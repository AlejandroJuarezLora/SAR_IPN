* SPICE3 file created from sarlogic.ext - technology: sky130B

.subckt sar_logic VGND VPWR cal clk clkc comp ctln[0] ctln[1] ctln[2] ctln[3] ctln[4]
+ ctln[5] ctln[6] ctln[7] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6]
+ ctlp[7] en result[0] result[1] result[2] result[3] result[4] result[5] result[6]
+ result[7] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1]
+ trimb[2] trimb[3] trimb[4] valid
* X0 VGND VPWR.t184 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=199 ps=2.08k w=0 l=0
* X1 VGND VPWR.t24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X2 VPWR VGND.t92 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=299 ps=2.85k w=0 l=0
* X3 VGND VPWR.t40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X4 VGND VPWR.t234 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X5 VGND VPWR.t167 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X6 VPWR VGND.t241 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X7 VGND VPWR.t9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X8 VPWR VGND.t32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X9 VPWR VGND.t38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X10 VPWR VGND.t168 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X11 VGND VPWR.t29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X12 VGND VPWR.t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X13 VPWR VGND.t9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X14 VPWR VGND.t117 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X15 VPWR VGND.t161 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X16 VGND VPWR.t155 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X17 VPWR VGND.t131 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X18 VGND VPWR.t194 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X19 VGND VPWR.t140 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X20 VPWR VGND.t94 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X21 VPWR VGND.t219 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X22 VPWR VGND.t190 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X23 VPWR VGND.t211 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X24 VGND VPWR.t241 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X25 VGND VPWR.t20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X26 VGND VPWR.t215 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X27 VPWR VGND.t235 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X28 VPWR VGND.t244 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X29 VPWR VGND.t74 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X30 VPWR VGND.t26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X31 VPWR VGND.t103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X32 VPWR VGND.t140 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X33 VPWR VGND.t10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X34 VPWR VGND.t192 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X35 VPWR VGND.t197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X36 VPWR VGND.t59 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X37 VGND VPWR.t57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X38 VPWR VGND.t107 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X39 VPWR VGND.t238 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X40 VGND VPWR.t8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X41 VGND VPWR.t137 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X42 VGND VPWR.t165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X43 VGND VPWR.t187 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X44 VPWR VGND.t57 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X45 VGND VPWR.t145 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X46 VPWR VGND.t172 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X47 VGND VPWR.t12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X48 VPWR VGND.t243 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X49 VGND VPWR.t10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X50 VPWR VGND.t16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X51 VGND VPWR.t192 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X52 VGND VPWR.t161 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X53 VGND VPWR.t242 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X54 VPWR VGND.t62 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X55 VPWR VGND.t12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X56 VGND VPWR.t49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X57 VGND VPWR.t235 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X58 VGND VPWR.t92 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X59 VPWR VGND.t159 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X60 VGND VPWR.t218 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X61 VPWR VGND.t242 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X62 VGND VPWR.t153 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X63 VPWR VGND.t49 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X64 VGND VPWR.t142 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X65 VPWR VGND.t226 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X66 VGND VPWR.t247 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X67 VPWR VGND.t2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X68 VPWR VGND.t164 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X69 VGND VPWR.t72 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X70 VPWR VGND.t143 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X71 VPWR VGND.t122 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X72 VPWR VGND.t142 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X73 VGND VPWR.t62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X74 VPWR VGND.t253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X75 VPWR VGND.t28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X76 VGND VPWR.t209 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X77 VPWR VGND.t213 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X78 VGND VPWR.t75 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X79 VPWR VGND.t163 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X80 VPWR VGND.t208 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X81 VPWR VGND.t175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X82 VPWR VGND.t118 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X83 clkbuf_0_clk/a_110_47# clk.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=0 l=0
* X84 VGND VPWR.t190 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X85 VPWR VGND.t202 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X86 VGND VPWR.t91 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X87 VGND VPWR.t46 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X88 VPWR VGND.t176 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X89 VPWR VGND.t101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X90 VPWR VGND.t75 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X91 VGND VPWR.t74 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X92 VGND VPWR.t96 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X93 VGND VPWR.t197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X94 VPWR VGND.t177 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X95 VGND VPWR.t162 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X96 VPWR VGND.t46 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X97 VGND VPWR.t47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X98 VGND VPWR.t135 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X99 VPWR VGND.t254 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X100 VGND VPWR.t128 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X101 VPWR VGND.t86 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X102 VPWR VGND.t135 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X103 VGND VPWR.t202 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X104 VPWR VGND.t171 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X105 VPWR VGND.t83 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X106 VGND VPWR.t65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X107 VPWR VGND.t236 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X108 VPWR VGND.t167 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X109 VPWR VGND.t109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X110 VGND VPWR.t156 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X111 VPWR VGND.t65 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X112 VPWR VGND.t40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X113 VGND VPWR.t79 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X114 VGND VPWR.t67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X115 VPWR VGND.t89 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X116 VPWR VGND.t19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X117 VGND VPWR.t2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X118 VPWR VGND.t127 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X119 VGND VPWR.t116 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X120 VPWR VGND.t20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X121 VGND VPWR.t252 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X122 VGND VPWR.t150 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X123 VPWR VGND.t24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X124 VGND VPWR.t31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X125 VGND VPWR.t90 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X126 VPWR VGND.t95 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X127 VGND VPWR.t233 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X128 VGND VPWR.t236 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X129 VGND VPWR.t163 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X130 VGND VPWR.t154 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X131 VPWR VGND.t71 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X132 VGND VPWR.t118 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X133 VGND VPWR.t97 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X134 VGND VPWR.t61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X135 VPWR VGND.t136 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X136 VPWR VGND.t31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X137 VPWR VGND.t137 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X138 VGND VPWR.t101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X139 VPWR VGND.t90 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X140 VGND VPWR.t195 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X141 VGND VPWR.t228 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X142 VGND VPWR.t180 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X143 VPWR VGND.t179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X144 VPWR VGND.t80 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X145 VGND VPWR.t81 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X146 VPWR VGND.t41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X147 VPWR VGND.t228 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X148 VPWR VGND.t120 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X149 VGND VPWR.t121 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X150 VGND VPWR.t86 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X151 VPWR VGND.t194 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X152 VPWR VGND.t214 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X153 VGND VPWR.t171 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X154 VGND VPWR.t83 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X155 VGND VPWR.t231 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X156 VGND VPWR.t43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X157 VGND VPWR.t206 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X158 VPWR VGND.t215 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X159 VPWR VGND.t199 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X160 VGND VPWR.t179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X161 VGND VPWR.t80 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X162 VPWR clk.t0 clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
* X163 VGND VPWR.t112 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X164 VPWR VGND.t206 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X165 VPWR VGND.t43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X166 VPWR VGND.t218 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X167 VPWR VGND.t239 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X168 VPWR VGND.t134 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X169 VGND VPWR.t39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X170 VGND VPWR.t129 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X171 VGND VPWR.t89 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X172 VGND VPWR.t205 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X173 VGND VPWR.t106 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X174 VPWR VGND.t209 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X175 VGND VPWR.t5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X176 VPWR VGND.t129 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X177 VPWR VGND.t70 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X178 VPWR VGND.t170 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X179 VGND VPWR.t220 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X180 VPWR VGND.t205 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X181 VPWR VGND.t104 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X182 VGND VPWR.t173 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X183 VGND VPWR.t125 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X184 VGND VPWR.t127 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X185 VGND VPWR.t27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X186 VPWR VGND.t247 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X187 VGND VPWR.t71 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X188 VPWR VGND.t4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X189 VPWR VGND.t88 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X190 VPWR VGND.t173 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X191 VGND VPWR.t30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X192 VGND VPWR.t151 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X193 VGND VPWR.t130 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X194 VPWR VGND.t72 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X195 VPWR VGND.t223 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X196 VGND VPWR.t44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X197 VGND VPWR.t70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X198 VPWR VGND.t147 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X199 VPWR VGND.t102 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X200 VPWR VGND.t30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X201 VGND VPWR.t66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X202 VGND VPWR.t182 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X203 VGND VPWR.t41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X204 VPWR VGND.t44 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X205 clkbuf_0_clk/a_110_47# clk.t3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
* X206 VGND VPWR.t68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X207 VGND VPWR.t183 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X208 VPWR VGND.t98 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X209 VPWR VGND.t96 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X210 VGND VPWR.t4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X211 VGND VPWR.t214 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X212 VGND VPWR.t166 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X213 VPWR VGND.t156 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X214 VPWR VGND.t232 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X215 VGND VPWR.t199 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X216 VGND VPWR.t157 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X217 VPWR VGND.t91 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X218 VPWR VGND.t162 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X219 VPWR VGND.t128 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X220 VGND VPWR.t6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X221 VPWR VGND.t53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X222 VGND VPWR.t239 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X223 VPWR VGND.t141 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X224 VPWR VGND.t47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X225 VPWR VGND.t150 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X226 VGND VPWR.t250 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X227 VPWR VGND.t111 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X228 VGND VPWR.t105 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X229 clkbuf_0_clk/a_110_47# clk.t6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0 l=0
* X230 VGND VPWR.t189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X231 VGND VPWR.t172 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X232 VGND VPWR.t170 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X233 VGND VPWR.t58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X234 VPWR VGND.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X235 VPWR VGND.t36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X236 VGND VPWR.t55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X237 VPWR VGND.t195 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X238 VPWR VGND.t189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X239 VGND VPWR.t77 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X240 VPWR VGND.t67 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X241 VGND VPWR.t232 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X242 VGND VPWR.t15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X243 VPWR VGND.t79 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X244 VGND VPWR.t45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X245 VPWR VGND.t196 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X246 VPWR VGND.t34 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X247 VPWR VGND.t55 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X248 VPWR clk.t7 clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
* X249 VGND VPWR.t88 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X250 VGND VPWR.t223 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X251 VPWR VGND.t132 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X252 VGND VPWR.t147 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X253 VGND VPWR.t102 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X254 VPWR VGND.t153 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X255 VGND VPWR.t139 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X256 VPWR VGND.t116 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X257 VGND VPWR.t144 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X258 VGND VPWR.t174 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X259 VGND VPWR.t138 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X260 VPWR VGND.t97 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X261 VPWR VGND.t8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X262 VPWR VGND.t152 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X263 VGND VPWR.t132 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X264 VGND VPWR.t69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X265 VPWR VGND.t231 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X266 VGND VPWR.t14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X267 VGND VPWR.t98 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X268 VPWR VGND.t165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X269 VPWR VGND.t154 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X270 VGND VPWR.t115 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X271 VGND VPWR.t169 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X272 VGND VPWR.t158 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X273 VPWR VGND.t61 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X274 VPWR VGND.t191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X275 VPWR VGND.t180 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X276 VPWR VGND.t69 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X277 VPWR VGND.t39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X278 VGND VPWR.t126 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X279 VGND VPWR.t23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X280 VGND VPWR.t133 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X281 VGND VPWR.t108 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X282 VPWR VGND.t121 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X283 VGND VPWR.t53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X284 VGND VPWR.t141 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X285 VPWR VGND.t81 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X286 VPWR VGND.t220 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X287 VGND VPWR.t100 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X288 VGND VPWR.t13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X289 VGND VPWR.t22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X290 VPWR VGND.t245 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X291 VGND VPWR.t111 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X292 VGND VPWR.t191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X293 VGND VPWR.t56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X294 VGND VPWR.t60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X295 VGND VPWR.t152 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X296 VGND VPWR.t1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X297 VGND VPWR.t36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X298 VGND VPWR.t99 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X299 VPWR VGND.t87 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X300 VPWR VGND.t56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X301 VPWR VGND.t66 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X302 VGND VPWR.t196 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X303 VPWR VGND.t182 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X304 VGND VPWR.t34 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X305 VGND VPWR.t64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X306 VPWR VGND.t76 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X307 VPWR VGND.t149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X308 VPWR VGND.t106 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X309 VPWR VGND.t35 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X310 VPWR VGND.t27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X311 VPWR VGND.t249 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X312 VGND clk.t5 clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
* X313 VPWR VGND.t157 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X314 VPWR VGND.t3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X315 VPWR VGND.t151 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X316 VGND VPWR.t225 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X317 VGND VPWR.t200 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X318 VGND VPWR.t110 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X319 VGND VPWR.t85 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X320 VGND VPWR.t211 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X321 VGND VPWR.t103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X322 VGND VPWR.t76 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X323 VPWR VGND.t130 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X324 VPWR VGND.t110 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X325 VPWR VGND.t105 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X326 VPWR VGND.t85 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X327 VPWR VGND.t6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X328 VPWR VGND.t84 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X329 VPWR VGND.t240 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X330 VGND VPWR.t160 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X331 VGND VPWR.t245 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X332 VPWR VGND.t188 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X333 VPWR VGND.t166 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X334 VPWR VGND.t123 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X335 VGND VPWR.t50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X336 VPWR VGND.t246 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X337 VPWR VGND.t183 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X338 VGND VPWR.t181 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X339 VPWR VGND.t45 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X340 VGND VPWR.t48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X341 VPWR VGND.t82 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X342 VGND VPWR.t87 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X343 VPWR VGND.t252 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X344 VGND VPWR.t124 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X345 VGND VPWR.t149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X346 clkbuf_0_clk/a_110_47# clk.t2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
* X347 VPWR VGND.t139 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X348 VPWR VGND.t233 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X349 VGND VPWR.t204 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X350 VGND VPWR.t119 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X351 VGND VPWR.t37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X352 VGND VPWR.t7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X353 VPWR VGND.t138 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X354 VPWR VGND.t250 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X355 VGND VPWR.t114 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X356 VPWR VGND.t146 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X357 VPWR VGND.t33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X358 VPWR VGND.t14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X359 VGND VPWR.t35 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X360 VPWR VGND.t119 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X361 VPWR VGND.t37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X362 VGND VPWR.t203 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X363 VGND VPWR.t136 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X364 VPWR VGND.t115 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X365 VPWR VGND.t11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X366 VPWR VGND.t15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X367 VPWR VGND.t58 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X368 VGND VPWR.t227 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X369 VGND VPWR.t246 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X370 VGND VPWR.t249 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X371 VPWR VGND.t93 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X372 VGND VPWR.t217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X373 VGND VPWR.t3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X374 VGND VPWR.t208 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X375 VPWR VGND.t77 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X376 VPWR VGND.t52 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X377 VGND VPWR.t175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X378 VPWR VGND.t108 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X379 VGND VPWR.t73 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X380 VPWR VGND.t230 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X381 VPWR VGND.t100 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X382 VPWR VGND.t22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X383 VGND VPWR.t33 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X384 VPWR VGND.t248 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X385 VGND VPWR.t11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X386 VGND VPWR.t84 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X387 VPWR VGND.t73 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X388 VPWR VGND.t112 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X389 VPWR VGND.t18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X390 VGND VPWR.t240 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X391 VPWR VGND.t51 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X392 VGND VPWR.t63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X393 VPWR comp.t0 input2/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=0 l=0
* X394 VGND VPWR.t146 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X395 VPWR VGND.t99 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X396 VPWR VGND.t169 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X397 VPWR VGND.t158 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X398 VGND VPWR.t123 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X399 VGND VPWR.t201 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X400 VGND VPWR.t188 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X401 VPWR VGND.t17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X402 VGND clk.t4 clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
* X403 VPWR VGND.t63 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X404 VGND VPWR.t148 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X405 VPWR VGND.t185 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X406 VPWR VGND.t5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X407 VGND VPWR.t82 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X408 VPWR VGND.t186 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X409 VPWR VGND.t174 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X410 VPWR VGND.t126 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X411 VPWR VGND.t23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X412 VPWR VGND.t148 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X413 VGND VPWR.t117 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X414 VGND VPWR.t18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X415 VPWR VGND.t13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X416 VGND VPWR.t51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X417 VGND VPWR.t237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X418 VGND VPWR.t198 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X419 VPWR VGND.t125 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X420 VGND VPWR.t143 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X421 VPWR VGND.t222 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X422 VPWR VGND.t237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X423 VGND VPWR.t42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X424 VGND VPWR.t21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X425 VGND VPWR.t244 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X426 VGND VPWR.t164 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X427 VGND VPWR.t26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X428 VPWR VGND.t200 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X429 VGND VPWR.t93 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X430 VPWR VGND.t42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X431 VPWR VGND.t64 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X432 VPWR VGND.t21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X433 VPWR VGND.t68 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X434 VGND VPWR.t185 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X435 VGND VPWR.t32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X436 VGND VPWR.t38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X437 VGND VPWR.t52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X438 VPWR VGND.t212 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X439 VGND VPWR.t168 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X440 VGND VPWR.t230 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X441 VGND VPWR.t16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X442 VGND VPWR.t229 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X443 VGND VPWR.t248 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X444 VPWR VGND.t181 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X445 VGND VPWR.t131 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X446 VGND VPWR.t94 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X447 VPWR VGND.t229 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X448 VPWR VGND.t216 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X449 VPWR VGND.t225 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X450 VPWR VGND.t50 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X451 VGND VPWR.t219 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X452 VGND VPWR.t120 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X453 VPWR VGND.t193 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X454 VGND VPWR.t17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X455 input1/a_75_212# cal.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0 l=0
* X456 VPWR VGND.t224 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X457 VGND VPWR.t159 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X458 VGND VPWR.t59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X459 VGND VPWR.t54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X460 VGND VPWR.t107 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X461 VPWR VGND.t78 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X462 VGND VPWR.t238 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X463 VGND VPWR.t122 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X464 VGND VPWR.t186 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X465 VPWR VGND.t160 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X466 VPWR VGND.t207 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X467 VGND VPWR.t226 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X468 VPWR VGND.t114 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X469 VGND VPWR.t28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X470 VPWR VGND.t54 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X471 VPWR rstn.t0 input4/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0 l=0
* X472 VGND VPWR.t216 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X473 input1/a_75_212# cal.t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0 l=0
* X474 VPWR VGND.t7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X475 VPWR VGND.t203 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X476 VPWR VGND.t184 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X477 VGND VPWR.t134 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X478 VGND VPWR.t221 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X479 VPWR VGND.t227 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X480 VGND VPWR.t243 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X481 VGND VPWR.t193 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X482 VGND VPWR.t222 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X483 VPWR VGND.t234 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X484 VPWR VGND.t210 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X485 VPWR VGND.t48 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X486 VPWR VGND.t221 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X487 VPWR VGND.t178 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X488 VPWR VGND.t29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X489 VGND VPWR.t104 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X490 VPWR VGND.t0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X491 VGND VPWR.t224 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X492 VPWR VGND.t251 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X493 VPWR VGND.t144 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X494 VPWR VGND.t124 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X495 VPWR VGND.t155 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X496 VGND VPWR.t212 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X497 VPWR VGND.t204 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X498 VGND VPWR.t210 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X499 VGND VPWR.t253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X500 VPWR VGND.t25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X501 VPWR VGND.t201 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X502 VGND VPWR.t178 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X503 VGND VPWR.t213 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X504 VPWR VGND.t133 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X505 VGND VPWR.t109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X506 input3/a_75_212# en.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0 l=0
* X507 VGND VPWR.t251 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X508 VPWR VGND.t217 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X509 VGND rstn.t1 input4/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0 l=0
* X510 VGND VPWR.t113 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X511 VGND VPWR.t176 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X512 VGND comp.t1 input2/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0 l=0
* X513 VGND VPWR.t19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X514 VPWR VGND.t187 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X515 VGND VPWR.t177 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X516 VPWR VGND.t145 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X517 VGND VPWR.t254 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X518 VPWR VGND.t113 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X519 VGND VPWR.t78 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X520 VGND VPWR.t25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X521 VPWR VGND.t60 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X522 VGND VPWR.t207 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X523 VPWR VGND.t198 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X524 input3/a_75_212# en.t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0 l=0
* X525 VGND VPWR.t95 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
C0 _109_ _332_/a_27_47# 4.37e-19
C1 trim_val\[0\] _108_ 0.37f
C2 trim_val\[0\] _332_/a_543_47# 1.9e-19
C3 net12 net26 0.102f
C4 _022_ _078_ 2.81e-20
C5 _304_/a_1283_21# _065_ 0.00232f
C6 _337_/a_1462_47# _049_ 4.02e-19
C7 net43 _314_/a_543_47# 0.157f
C8 clk _317_/a_1108_47# 0.00521f
C9 net34 net33 0.433f
C10 net5 net33 3.09e-19
C11 net22 mask\[0\] 0.297f
C12 _257_/a_27_297# net46 1.93e-20
C13 _315_/a_27_47# net14 0.0117f
C14 _290_/a_207_413# net40 1.78e-19
C15 trim_mask\[1\] net34 5.19e-20
C16 _189_/a_218_47# clknet_0_clk 0.0521f
C17 _340_/a_1602_47# _300_/a_47_47# 6.18e-20
C18 _290_/a_27_413# net34 0.0108f
C19 _306_/a_651_413# _101_ 7.37e-21
C20 output25/a_27_47# _310_/a_193_47# 2.18e-19
C21 _306_/a_1108_47# _063_ 9.17e-21
C22 _284_/a_68_297# _067_ 4.38e-19
C23 _222_/a_113_297# _222_/a_199_47# 2.42e-19
C24 clk _203_/a_59_75# 0.0113f
C25 _238_/a_75_212# _316_/a_27_47# 9.84e-19
C26 _270_/a_145_75# net16 4.09e-19
C27 VPWR _331_/a_1462_47# 7.03e-20
C28 net15 _090_ 7.61e-19
C29 _235_/a_79_21# _090_ 0.001f
C30 VPWR _260_/a_93_21# 0.142f
C31 _340_/a_1032_413# _132_ 6.76e-20
C32 _322_/a_651_413# mask\[3\] 0.0227f
C33 _032_ net19 1.11e-19
C34 _225_/a_109_297# net14 5.22e-19
C35 net4 _317_/a_1108_47# 0.0157f
C36 net44 net26 0.0747f
C37 _325_/a_27_47# _222_/a_113_297# 1.15e-19
C38 _232_/a_32_297# _098_ 6.57e-21
C39 VPWR _328_/a_448_47# 0.0795f
C40 _078_ _313_/a_1283_21# 3.27e-20
C41 _311_/a_1462_47# net19 5.5e-20
C42 cal_itt\[0\] _303_/a_639_47# 1.44e-19
C43 _071_ _303_/a_448_47# 6.22e-20
C44 _300_/a_377_297# cal_count\[3\] 3.69e-19
C45 _329_/a_1217_47# _026_ 7.86e-21
C46 output20/a_27_47# _312_/a_193_47# 0.00122f
C47 _337_/a_448_47# clknet_2_0__leaf_clk 0.00471f
C48 net28 _314_/a_805_47# 7.38e-19
C49 _108_ _279_/a_204_297# 0.0111f
C50 _239_/a_694_21# _003_ 3.62e-21
C51 output36/a_27_47# net16 3.37e-19
C52 _015_ _317_/a_27_47# 9.18e-22
C53 trim_mask\[3\] _330_/a_1283_21# 0.0628f
C54 _262_/a_109_297# cal_count\[3\] 2.87e-19
C55 _289_/a_68_297# net40 0.00492f
C56 result[3] _082_ 5.94e-19
C57 _058_ _092_ 9.34e-19
C58 VPWR _312_/a_1108_47# 0.302f
C59 _232_/a_32_297# clknet_0_clk 2.86e-21
C60 _110_ _113_ 0.255f
C61 clknet_2_0__leaf_clk net14 0.527f
C62 net45 _138_/a_27_47# 0.0027f
C63 _093_ fanout45/a_27_47# 2.06e-20
C64 VPWR _307_/a_27_47# 0.483f
C65 VPWR _323_/a_448_47# 0.0807f
C66 _253_/a_81_21# _086_ 3.17e-21
C67 _313_/a_761_289# _313_/a_639_47# 3.16e-19
C68 _313_/a_27_47# _313_/a_1217_47# 2.56e-19
C69 _336_/a_193_47# clknet_0_clk 7.24e-19
C70 _336_/a_1108_47# clkbuf_2_2__f_clk/a_110_47# 0.00155f
C71 _071_ _190_/a_655_47# 6.61e-21
C72 _051_ cal_itt\[3\] 3.84e-20
C73 clk _318_/a_1270_413# 3.55e-19
C74 _337_/a_1283_21# _065_ 5.5e-21
C75 _048_ _226_/a_303_47# 0.00242f
C76 trim_mask\[0\] _262_/a_193_297# 3.38e-19
C77 net46 trim_val\[4\] 0.00883f
C78 _326_/a_1108_47# net52 9.47e-19
C79 _323_/a_448_47# net53 1.6e-21
C80 ctln[2] trim_val\[2\] 1.8e-20
C81 net8 net48 0.0209f
C82 _110_ net2 1.31e-20
C83 _325_/a_1108_47# mask\[2\] 4.31e-20
C84 _060_ _092_ 0.0391f
C85 VPWR _341_/a_651_413# 0.133f
C86 _321_/a_761_289# clknet_2_1__leaf_clk 0.00609f
C87 _289_/a_68_297# _299_/a_215_297# 6.49e-20
C88 output33/a_27_47# net34 0.0216f
C89 _024_ _111_ 7.76e-21
C90 VPWR _333_/a_543_47# 0.216f
C91 _104_ _098_ 8.66e-21
C92 _063_ _203_/a_59_75# 3.84e-19
C93 _089_ _054_ 6.64e-21
C94 _090_ _049_ 0.385f
C95 _275_/a_81_21# _335_/a_27_47# 3.69e-19
C96 trim[1] _173_/a_27_47# 0.00392f
C97 output32/a_27_47# net32 0.237f
C98 _337_/a_27_47# _319_/a_1283_21# 1.4e-19
C99 _234_/a_109_297# _282_/a_68_297# 6.46e-21
C100 cal_count\[0\] _338_/a_27_47# 1.14e-19
C101 VPWR _265_/a_384_47# 2.76e-19
C102 _124_ _338_/a_652_21# 0.00466f
C103 net33 _133_ 5.06e-20
C104 ctln[2] net16 1.33e-20
C105 _208_/a_218_47# _077_ 2.88e-19
C106 _330_/a_193_47# _330_/a_651_413# 0.0346f
C107 _330_/a_543_47# _330_/a_1108_47# 7.99e-20
C108 _172_/a_68_297# _172_/a_150_297# 0.00477f
C109 _208_/a_439_47# _076_ 6.37e-19
C110 net31 net46 9.91e-19
C111 clk clknet_2_0__leaf_clk 0.0705f
C112 VPWR _308_/a_1108_47# 0.323f
C113 net27 _152_/a_150_297# 3.75e-19
C114 net55 _098_ 0.0966f
C115 _048_ _228_/a_79_21# 0.185f
C116 net47 net2 0.0188f
C117 _315_/a_1217_47# net14 2.37e-19
C118 _015_ _318_/a_543_47# 9.18e-19
C119 _167_/a_161_47# _243_/a_27_297# 0.0011f
C120 _104_ clknet_0_clk 0.0857f
C121 net24 result[2] 0.0288f
C122 _079_ mask\[0\] 0.111f
C123 VPWR _237_/a_76_199# 0.107f
C124 _319_/a_1270_413# clknet_0_clk 9.87e-20
C125 _242_/a_382_297# _049_ 3.21e-19
C126 _284_/a_68_297# _284_/a_150_297# 0.00477f
C127 mask\[1\] _208_/a_505_21# 5.76e-20
C128 net16 _298_/a_78_199# 1.26e-20
C129 net45 _331_/a_761_289# 0.169f
C130 net9 _304_/a_27_47# 0.00441f
C131 VPWR _320_/a_805_47# 4.48e-19
C132 _230_/a_59_75# _067_ 8.66e-19
C133 _091_ _194_/a_113_297# 3.02e-20
C134 clknet_0_clk net55 0.344f
C135 VPWR _339_/a_1032_413# 0.459f
C136 net43 _310_/a_805_47# 0.00368f
C137 net27 result[6] 9.45e-21
C138 mask\[1\] mask\[2\] 0.014f
C139 net4 clknet_2_0__leaf_clk 0.0188f
C140 net22 _121_ 7.52e-21
C141 _297_/a_377_297# _132_ 0.00372f
C142 _071_ _000_ 1.61e-20
C143 ctlp[6] _312_/a_448_47# 7.83e-20
C144 _324_/a_1270_413# net27 1.8e-20
C145 _047_ trim_val\[1\] 0.00257f
C146 _212_/a_113_297# _212_/a_199_47# 2.42e-19
C147 _253_/a_81_21# clknet_2_1__leaf_clk 6.49e-21
C148 net12 net2 0.00487f
C149 _305_/a_1108_47# clk 0.00238f
C150 _107_ _171_/a_27_47# 0.00468f
C151 _339_/a_193_47# _286_/a_76_199# 4.61e-20
C152 _339_/a_27_47# _286_/a_505_21# 0.033f
C153 net13 net41 0.00634f
C154 _325_/a_543_47# _325_/a_651_413# 0.0572f
C155 _325_/a_761_289# _325_/a_1270_413# 2.6e-19
C156 _325_/a_193_47# _325_/a_639_47# 2.28e-19
C157 _110_ trim_val\[1\] 8.48e-19
C158 cal_itt\[0\] _231_/a_161_47# 0.0693f
C159 net17 cal_count\[0\] 9.79e-21
C160 _189_/a_408_47# clk 0.00194f
C161 _110_ _336_/a_193_47# 0.0134f
C162 VPWR _324_/a_27_47# 0.454f
C163 _024_ _065_ 3.21e-19
C164 VPWR _307_/a_1217_47# 5.67e-20
C165 mask\[4\] _311_/a_1283_21# 0.0672f
C166 clknet_0_clk _067_ 0.00189f
C167 _226_/a_27_47# _075_ 0.0637f
C168 _226_/a_109_47# _062_ 0.00153f
C169 VPWR output6/a_27_47# 0.267f
C170 clknet_0_clk _070_ 0.00135f
C171 _023_ _011_ 0.00513f
C172 _313_/a_1108_47# _010_ 3.47e-19
C173 _334_/a_1283_21# _057_ 1.12e-19
C174 _305_/a_1108_47# net4 2.22e-21
C175 _324_/a_27_47# net53 0.0107f
C176 output8/a_27_47# _179_/a_27_47# 1.48e-19
C177 net2 net44 0.00953f
C178 _323_/a_193_47# _150_/a_27_47# 1.52e-19
C179 clknet_2_0__leaf_clk net52 0.139f
C180 net45 _101_ 0.349f
C181 output30/a_27_47# sample 0.338f
C182 VPWR _241_/a_388_297# 0.0139f
C183 _321_/a_639_47# _042_ 3.04e-19
C184 cal_itt\[0\] _001_ 0.0135f
C185 _278_/a_109_297# net40 0.0105f
C186 trim_mask\[4\] _049_ 0.161f
C187 _271_/a_75_212# _333_/a_27_47# 1.15e-19
C188 net47 _123_ 0.192f
C189 _316_/a_27_47# _316_/a_1108_47# 0.102f
C190 _316_/a_193_47# _316_/a_1283_21# 0.0424f
C191 _316_/a_761_289# _316_/a_543_47# 0.21f
C192 _189_/a_218_47# net44 2.22e-22
C193 _324_/a_27_47# _009_ 5.42e-21
C194 VPWR _303_/a_1108_47# 0.292f
C195 _340_/a_1140_413# _123_ 0.00163f
C196 VPWR output25/a_27_47# 0.3f
C197 net50 _335_/a_543_47# 0.00214f
C198 _168_/a_207_413# clknet_0_clk 2.23e-19
C199 trim_mask\[3\] _335_/a_1283_21# 0.0277f
C200 trim_val\[3\] _335_/a_1108_47# 0.00159f
C201 net28 net29 0.0207f
C202 _110_ _104_ 0.0117f
C203 _101_ _065_ 0.722f
C204 _008_ _311_/a_651_413# 2.01e-20
C205 _330_/a_761_289# _027_ 0.0431f
C206 _330_/a_193_47# net46 0.024f
C207 _301_/a_47_47# net2 0.00226f
C208 calibrate _260_/a_250_297# 0.0157f
C209 mask\[0\] clknet_0_clk 0.00866f
C210 _337_/a_651_413# net55 4.2e-19
C211 net15 _283_/a_75_212# 5.67e-19
C212 _231_/a_161_47# _108_ 2.1e-19
C213 state\[2\] _318_/a_805_47# 1.41e-19
C214 _341_/a_27_47# net2 1.15e-20
C215 _064_ _136_ 2.37e-19
C216 _158_/a_68_297# net29 0.105f
C217 _305_/a_1108_47# _063_ 2.71e-19
C218 _110_ net55 8.54e-21
C219 _146_/a_68_297# net52 0.00178f
C220 _320_/a_27_47# net45 1.04e-20
C221 _320_/a_761_289# clknet_2_0__leaf_clk 4.81e-19
C222 VPWR _309_/a_1270_413# 9.56e-19
C223 _061_ _301_/a_285_47# 2.07e-19
C224 VPWR _190_/a_465_47# 0.00182f
C225 _020_ _311_/a_1283_21# 6.17e-19
C226 net13 _094_ 0.0763f
C227 _113_ clknet_2_2__leaf_clk 0.174f
C228 trim_mask\[2\] _269_/a_81_21# 1.32e-20
C229 mask\[7\] _251_/a_109_297# 0.0111f
C230 _102_ _251_/a_27_297# 0.00446f
C231 clkbuf_2_1__f_clk/a_110_47# _016_ 0.0198f
C232 output32/a_27_47# clkc 4.89e-21
C233 _204_/a_75_212# _073_ 0.188f
C234 net9 _340_/a_476_47# 0.0153f
C235 _319_/a_27_47# _101_ 6.81e-20
C236 state\[2\] calibrate 0.62f
C237 net4 trim_mask\[1\] 2.12e-21
C238 _328_/a_27_47# _336_/a_27_47# 1.59e-21
C239 _327_/a_27_47# _267_/a_59_75# 5.67e-21
C240 state\[1\] _090_ 5.04e-20
C241 _307_/a_761_289# _074_ 0.00439f
C242 net4 _336_/a_761_289# 0.0085f
C243 _334_/a_27_47# _334_/a_193_47# 0.902f
C244 _329_/a_193_47# _258_/a_27_297# 3.43e-19
C245 _314_/a_27_47# _314_/a_761_289# 0.0701f
C246 _329_/a_1283_21# trim_mask\[0\] 5.88e-20
C247 trimb[1] cal_count\[0\] 4.96e-19
C248 output36/a_27_47# trimb[0] 0.339f
C249 VPWR _249_/a_109_47# 6.87e-19
C250 _324_/a_1283_21# net26 1.34e-21
C251 _326_/a_761_289# net28 9.18e-19
C252 VPWR _293_/a_299_297# 0.282f
C253 _228_/a_382_297# _228_/a_297_47# 8.13e-19
C254 _187_/a_212_413# trim_val\[0\] 1.02e-19
C255 net43 _306_/a_448_47# 5.43e-21
C256 _339_/a_193_47# cal_count\[0\] 0.498f
C257 _320_/a_27_47# _065_ 1.76e-20
C258 state\[2\] net45 0.0716f
C259 _169_/a_109_53# _050_ 3.88e-20
C260 _144_/a_27_47# _126_ 6.56e-22
C261 _064_ _119_ 0.0152f
C262 _216_/a_199_47# _082_ 0.00151f
C263 _110_ _114_ 0.103f
C264 _239_/a_694_21# _229_/a_27_297# 8.56e-21
C265 _227_/a_109_93# _092_ 4.21e-21
C266 _307_/a_543_47# clknet_2_0__leaf_clk 6.3e-19
C267 _307_/a_193_47# net45 0.0264f
C268 trim[3] _334_/a_761_289# 9.11e-20
C269 _110_ _336_/a_1462_47# 2.04e-19
C270 VPWR _324_/a_1217_47# 1.16e-19
C271 _336_/a_27_47# _266_/a_68_297# 5.87e-21
C272 _104_ net12 0.034f
C273 _060_ _226_/a_197_47# 1.78e-19
C274 _235_/a_297_47# _092_ 0.00256f
C275 _053_ _048_ 0.0572f
C276 _330_/a_1283_21# _108_ 4.09e-21
C277 _283_/a_75_212# _049_ 0.0032f
C278 net12 net55 0.00863f
C279 net47 _067_ 0.0716f
C280 _041_ _202_/a_79_21# 4.47e-20
C281 VPWR _322_/a_805_47# 2.57e-19
C282 _304_/a_27_47# _122_ 0.0101f
C283 net47 _070_ 0.00159f
C284 _053_ _330_/a_27_47# 9.79e-21
C285 _104_ _258_/a_373_47# 6.81e-19
C286 _083_ _311_/a_639_47# 2.45e-20
C287 clknet_2_1__leaf_clk net21 0.00953f
C288 _308_/a_651_413# _074_ 0.00538f
C289 fanout46/a_27_47# trim_mask\[4\] 0.00133f
C290 _273_/a_59_75# _272_/a_81_21# 0.00979f
C291 _030_ _333_/a_448_47# 0.158f
C292 ctln[7] _318_/a_651_413# 3.69e-20
C293 net13 _318_/a_639_47# 0.00132f
C294 _316_/a_1108_47# _316_/a_1217_47# 0.00742f
C295 _316_/a_1283_21# _316_/a_1462_47# 0.0074f
C296 _195_/a_218_47# _062_ 0.00222f
C297 _237_/a_505_21# calibrate 5.7e-20
C298 _237_/a_76_199# _093_ 4.41e-19
C299 _323_/a_193_47# _042_ 0.545f
C300 net43 _094_ 2.06e-20
C301 VPWR _281_/a_103_199# 0.455f
C302 _087_ _100_ 0.0124f
C303 clknet_2_1__leaf_clk _312_/a_1283_21# 3.11e-20
C304 net44 _319_/a_1270_413# 1.27e-20
C305 _078_ net14 0.304f
C306 _247_/a_109_47# mask\[2\] 8.74e-19
C307 _171_/a_27_47# _118_ 1.86e-20
C308 _326_/a_448_47# net43 2.56e-19
C309 _330_/a_1462_47# net46 0.00331f
C310 _134_ _135_ 0.259f
C311 _007_ _310_/a_193_47# 0.252f
C312 net2 _209_/a_27_47# 9.21e-20
C313 en_co_clk net51 1.77e-19
C314 _122_ _298_/a_292_297# 4.73e-19
C315 _323_/a_1108_47# clknet_2_1__leaf_clk 6.95e-20
C316 net44 net55 0.00485f
C317 _284_/a_68_297# clknet_2_3__leaf_clk 0.002f
C318 net13 _074_ 0.13f
C319 net4 _069_ 0.0991f
C320 _237_/a_218_374# _014_ 1.21e-19
C321 _074_ _155_/a_68_297# 0.0534f
C322 _181_/a_68_297# _108_ 0.0216f
C323 mask\[0\] _245_/a_27_297# 0.0739f
C324 _143_/a_68_297# _078_ 0.0426f
C325 _334_/a_543_47# net46 0.177f
C326 net15 _246_/a_373_47# 4.75e-19
C327 trim_val\[1\] clknet_2_2__leaf_clk 2.5e-20
C328 mask\[3\] _310_/a_193_47# 1.41e-20
C329 net25 _310_/a_761_289# 0.00128f
C330 _195_/a_76_199# _195_/a_218_47# 0.00783f
C331 _294_/a_150_297# _132_ 8.78e-19
C332 net9 _338_/a_193_47# 5.19e-20
C333 _327_/a_193_47# net46 0.0321f
C334 _336_/a_27_47# _028_ 1.05e-19
C335 _336_/a_193_47# clknet_2_2__leaf_clk 0.00584f
C336 cal_itt\[0\] _195_/a_218_374# 0.00697f
C337 cal_itt\[1\] _195_/a_505_21# 0.0052f
C338 _328_/a_639_47# trim_mask\[1\] 6.86e-21
C339 mask\[7\] _022_ 0.00132f
C340 cal_itt\[2\] cal_itt\[1\] 0.0472f
C341 result[1] _308_/a_193_47# 0.00876f
C342 net9 _340_/a_1224_47# 1.72e-20
C343 _319_/a_651_413# _016_ 6.95e-19
C344 _319_/a_639_47# net52 6.3e-20
C345 _304_/a_27_47# _304_/a_1283_21# 0.0436f
C346 _304_/a_193_47# _304_/a_543_47# 0.23f
C347 _121_ clknet_0_clk 0.0132f
C348 _230_/a_59_75# _230_/a_145_75# 0.00658f
C349 _221_/a_109_297# _084_ 0.00265f
C350 _092_ net30 0.0074f
C351 _329_/a_1283_21# _328_/a_1283_21# 1.06e-19
C352 _334_/a_543_47# _334_/a_639_47# 0.0138f
C353 _334_/a_193_47# _334_/a_1217_47# 2.36e-20
C354 _334_/a_761_289# _334_/a_805_47# 3.69e-19
C355 _329_/a_543_47# trim_mask\[2\] 2.01e-19
C356 _168_/a_297_47# clk 7.46e-19
C357 _314_/a_1108_47# _314_/a_1270_413# 0.00645f
C358 _314_/a_761_289# _314_/a_1217_47# 4.2e-19
C359 _314_/a_543_47# _314_/a_805_47# 0.00171f
C360 _034_ _192_/a_27_47# 3.76e-21
C361 _263_/a_79_21# net55 0.0508f
C362 net44 _070_ 0.00138f
C363 _058_ net46 0.0779f
C364 _327_/a_543_47# _327_/a_1108_47# 7.99e-20
C365 _327_/a_193_47# _327_/a_651_413# 0.0346f
C366 net17 net16 0.00167f
C367 _050_ net51 4.53e-21
C368 _336_/a_543_47# net19 0.00765f
C369 _335_/a_761_289# _027_ 1.21e-19
C370 _335_/a_193_47# net46 0.051f
C371 _322_/a_193_47# _074_ 0.0117f
C372 _069_ _063_ 0.0696f
C373 _307_/a_1462_47# net45 0.00342f
C374 _308_/a_1108_47# _319_/a_193_47# 9.39e-20
C375 _308_/a_27_47# _319_/a_448_47# 6.41e-22
C376 _168_/a_27_413# _331_/a_448_47# 2.27e-21
C377 _169_/a_215_311# _169_/a_373_53# 0.0026f
C378 _169_/a_109_53# _169_/a_301_53# 1.81e-19
C379 _169_/a_215_311# net54 6.47e-20
C380 VPWR _048_ 2.55f
C381 _262_/a_193_297# _190_/a_27_47# 8.1e-21
C382 _081_ net22 3.65e-20
C383 state\[2\] _239_/a_27_297# 3.98e-20
C384 _327_/a_651_413# _058_ 0.00331f
C385 net45 _241_/a_297_47# 1.02e-19
C386 _104_ clknet_2_2__leaf_clk 0.0678f
C387 VPWR _330_/a_27_47# 0.429f
C388 net15 _222_/a_113_297# 2.39e-19
C389 _257_/a_27_297# rebuffer3/a_75_212# 9.43e-22
C390 _332_/a_27_47# net46 0.331f
C391 _104_ _260_/a_584_47# 0.00332f
C392 _328_/a_543_47# net9 0.00272f
C393 _341_/a_27_47# _067_ 1.77e-19
C394 net3 net41 0.00983f
C395 _336_/a_543_47# _107_ 0.00213f
C396 net43 _074_ 0.0393f
C397 _002_ net19 1.69e-20
C398 _340_/a_476_47# _122_ 0.00178f
C399 trim_mask\[1\] _333_/a_448_47# 4.06e-19
C400 net49 _333_/a_1108_47# 0.00521f
C401 trim_val\[1\] _333_/a_651_413# 4.79e-19
C402 _274_/a_75_212# _114_ 0.00163f
C403 _304_/a_543_47# net18 0.00332f
C404 mask\[0\] net44 2.97e-19
C405 _051_ clone7/a_27_47# 1.21e-20
C406 clkbuf_2_1__f_clk/a_110_47# _040_ 0.00524f
C407 _301_/a_285_47# net16 0.00322f
C408 _092_ _072_ 4.89e-20
C409 _310_/a_27_47# _310_/a_1108_47# 0.102f
C410 _310_/a_193_47# _310_/a_1283_21# 0.0418f
C411 _310_/a_761_289# _310_/a_543_47# 0.21f
C412 net13 _243_/a_27_297# 0.00819f
C413 _276_/a_59_75# clkbuf_2_2__f_clk/a_110_47# 2.09e-21
C414 _327_/a_1283_21# _108_ 1.58e-19
C415 VPWR _325_/a_193_47# 0.591f
C416 _239_/a_694_21# _107_ 0.00576f
C417 VPWR _120_ 0.327f
C418 _046_ _313_/a_761_289# 0.00279f
C419 net21 _313_/a_27_47# 7.59e-19
C420 _335_/a_193_47# _335_/a_651_413# 0.0346f
C421 _335_/a_543_47# _335_/a_1108_47# 7.99e-20
C422 _005_ net45 8.46e-20
C423 _327_/a_27_47# _053_ 7.36e-20
C424 _097_ _090_ 7.45e-19
C425 result[4] _310_/a_193_47# 9.51e-19
C426 _305_/a_193_47# _092_ 1.07e-20
C427 _004_ net14 0.00343f
C428 _034_ clknet_2_0__leaf_clk 0.0621f
C429 _110_ net8 5.18e-21
C430 _230_/a_59_75# clknet_2_3__leaf_clk 0.00118f
C431 result[6] _011_ 0.0016f
C432 mask\[2\] net26 7.52e-20
C433 net35 _332_/a_1283_21# 0.019f
C434 _058_ _332_/a_448_47# 0.00217f
C435 _078_ net52 0.0217f
C436 _304_/a_543_47# _302_/a_27_297# 8.26e-20
C437 ctln[4] _057_ 1.27e-19
C438 net13 _232_/a_220_297# 9.18e-19
C439 VPWR _076_ 1.44f
C440 output35/a_27_47# net37 0.0127f
C441 net24 _041_ 0.0067f
C442 net2 _131_ 0.157f
C443 _135_ cal_count\[2\] 7.17e-20
C444 _327_/a_1462_47# net46 0.00407f
C445 net9 _341_/a_1283_21# 0.0146f
C446 _035_ net18 0.0212f
C447 net9 _333_/a_27_47# 2.54e-21
C448 _304_/a_448_47# _304_/a_639_47# 4.61e-19
C449 clkbuf_2_0__f_clk/a_110_47# _099_ 0.00122f
C450 trimb[1] net16 4.04e-20
C451 trim_mask\[2\] _033_ 0.00893f
C452 _339_/a_956_413# _123_ 0.00243f
C453 net43 _305_/a_448_47# 0.0148f
C454 net29 _085_ 1.86e-19
C455 trim[1] _047_ 0.122f
C456 _334_/a_448_47# _031_ 0.156f
C457 _076_ net53 0.0282f
C458 net16 _339_/a_193_47# 1.92e-21
C459 _214_/a_199_47# _078_ 2.65e-19
C460 _256_/a_27_297# net18 0.0106f
C461 clk _316_/a_1283_21# 5.68e-19
C462 _336_/a_761_289# _279_/a_396_47# 1.09e-19
C463 _336_/a_193_47# _279_/a_204_297# 7.53e-21
C464 ctlp[6] _156_/a_27_47# 0.001f
C465 _321_/a_27_47# _321_/a_1283_21# 0.0435f
C466 _321_/a_193_47# _321_/a_543_47# 0.22f
C467 net43 _146_/a_150_297# 3.43e-19
C468 _332_/a_543_47# _108_ 0.042f
C469 _332_/a_27_47# _332_/a_448_47# 0.0902f
C470 _332_/a_193_47# _332_/a_1108_47# 0.117f
C471 cal net1 0.0211f
C472 _110_ trim[1] 5.23e-20
C473 clknet_0_clk clknet_2_3__leaf_clk 0.00541f
C474 _106_ net19 0.159f
C475 _335_/a_1462_47# net46 0.00414f
C476 output14/a_27_47# _314_/a_193_47# 0.00632f
C477 _136_ net34 2.33e-20
C478 net23 clkbuf_2_1__f_clk/a_110_47# 0.00115f
C479 net5 _136_ 5.3e-20
C480 _049_ rebuffer5/a_161_47# 4.88e-19
C481 _125_ net37 0.00738f
C482 _168_/a_27_413# _028_ 4.62e-19
C483 _168_/a_207_413# clknet_2_2__leaf_clk 4.38e-20
C484 _094_ net3 0.0127f
C485 _053_ net54 1.84e-19
C486 state\[0\] _060_ 0.0791f
C487 _059_ _075_ 2.71e-19
C488 output7/a_27_47# clk 0.00341f
C489 fanout47/a_27_47# net4 0.229f
C490 _320_/a_761_289# _078_ 1.24e-19
C491 _320_/a_543_47# mask\[0\] 1.57e-20
C492 _304_/a_761_289# cal_count\[3\] 9.6e-21
C493 _337_/a_27_47# _337_/a_1283_21# 0.0435f
C494 _337_/a_193_47# _337_/a_543_47# 0.23f
C495 _304_/a_651_413# clknet_2_3__leaf_clk 6.03e-20
C496 _333_/a_761_289# net32 1.34e-19
C497 net4 _316_/a_1283_21# 0.00105f
C498 rebuffer4/a_27_47# rebuffer6/a_27_47# 1.62e-19
C499 _340_/a_1032_413# _298_/a_215_47# 1.11e-19
C500 _257_/a_109_47# trim_mask\[1\] 8.34e-19
C501 net9 _339_/a_652_21# 0.0048f
C502 _256_/a_27_297# _302_/a_27_297# 3.29e-21
C503 _250_/a_27_297# _249_/a_27_297# 8.82e-20
C504 VPWR _330_/a_1217_47# 8.79e-20
C505 trim_mask\[0\] clkbuf_2_2__f_clk/a_110_47# 4.42e-20
C506 _257_/a_27_297# _336_/a_1283_21# 1.8e-20
C507 cal_count\[1\] net2 0.914f
C508 _332_/a_1217_47# net46 2.95e-19
C509 _048_ _192_/a_548_47# 0.00535f
C510 _341_/a_193_47# _284_/a_68_297# 2.51e-20
C511 VPWR _007_ 0.791f
C512 _325_/a_1108_47# net26 7.08e-20
C513 _291_/a_35_297# cal_count\[0\] 0.103f
C514 _106_ _107_ 0.186f
C515 clknet_2_1__leaf_clk _045_ 0.0454f
C516 _340_/a_1224_47# _122_ 7.52e-20
C517 _104_ _279_/a_204_297# 5.82e-19
C518 net3 _192_/a_505_280# 0.0657f
C519 output7/a_27_47# net4 0.0341f
C520 _324_/a_27_47# mask\[6\] 4.25e-20
C521 clknet_2_1__leaf_clk _249_/a_109_297# 0.00341f
C522 _306_/a_761_289# rebuffer4/a_27_47# 2.69e-21
C523 VPWR _334_/a_761_289# 0.223f
C524 _053_ _068_ 0.00191f
C525 _310_/a_1108_47# _310_/a_1217_47# 0.00742f
C526 _310_/a_1283_21# _310_/a_1462_47# 0.0074f
C527 clkbuf_0_clk/a_110_47# clkbuf_2_3__f_clk/a_110_47# 0.00246f
C528 _314_/a_543_47# net29 0.00118f
C529 cal_count\[3\] clkbuf_2_3__f_clk/a_110_47# 0.0047f
C530 _048_ _262_/a_27_47# 0.101f
C531 _307_/a_543_47# _078_ 3.81e-19
C532 _307_/a_1108_47# net22 0.0601f
C533 VPWR _327_/a_27_47# 0.493f
C534 _307_/a_1283_21# mask\[0\] 0.00278f
C535 VPWR _325_/a_1462_47# 1.68e-19
C536 VPWR mask\[3\] 1.85f
C537 net31 _135_ 6.2e-21
C538 net21 _313_/a_1217_47# 5.32e-20
C539 _335_/a_761_289# _032_ 2.11e-19
C540 result[0] net22 0.00496f
C541 net16 _333_/a_805_47# 0.00127f
C542 _324_/a_805_47# clknet_2_1__leaf_clk 1.32e-19
C543 _302_/a_27_297# _302_/a_109_47# 0.00393f
C544 _340_/a_1602_47# _129_ 4.04e-19
C545 _123_ _131_ 2.67e-19
C546 result[4] _310_/a_1462_47# 2.78e-20
C547 net16 _109_ 0.0017f
C548 _311_/a_193_47# _311_/a_1270_413# 1.46e-19
C549 _311_/a_27_47# _311_/a_639_47# 3.82e-19
C550 _311_/a_543_47# _311_/a_448_47# 0.0498f
C551 _311_/a_761_289# _311_/a_651_413# 0.0977f
C552 _311_/a_1283_21# _311_/a_1108_47# 0.234f
C553 mask\[3\] net53 0.00181f
C554 net44 _121_ 2.33e-20
C555 _000_ _065_ 6.57e-20
C556 en_co_clk _192_/a_639_47# 1.02e-19
C557 output10/a_27_47# _335_/a_193_47# 2.95e-19
C558 _304_/a_761_289# _038_ 0.00102f
C559 _304_/a_448_47# _136_ 4.81e-19
C560 _104_ _257_/a_373_47# 6.81e-19
C561 VPWR _335_/a_27_47# 0.519f
C562 _071_ _306_/a_193_47# 6.82e-21
C563 cal_itt\[2\] _306_/a_1108_47# 1.91e-20
C564 _300_/a_377_297# en_co_clk 3.47e-21
C565 clknet_2_1__leaf_clk mask\[4\] 0.0601f
C566 trim[4] _332_/a_193_47# 1.01e-20
C567 _304_/a_1270_413# net47 4.46e-19
C568 net4 _287_/a_75_212# 1.58e-19
C569 _100_ _099_ 0.0406f
C570 _096_ _095_ 0.136f
C571 _326_/a_1108_47# _314_/a_27_47# 2.25e-20
C572 _326_/a_543_47# _314_/a_761_289# 3.17e-20
C573 _326_/a_761_289# _314_/a_543_47# 3.66e-20
C574 _326_/a_27_47# _314_/a_1108_47# 6.19e-20
C575 _048_ _093_ 0.153f
C576 net43 _002_ 0.311f
C577 en_co_clk _132_ 1.15e-19
C578 _256_/a_27_297# trim_mask\[0\] 0.177f
C579 _110_ clknet_2_3__leaf_clk 1.07e-20
C580 _340_/a_27_47# net47 0.0445f
C581 _336_/a_543_47# _118_ 0.0115f
C582 _336_/a_1283_21# trim_val\[4\] 0.063f
C583 VPWR _314_/a_1270_413# 7.89e-19
C584 _074_ net3 3.09e-20
C585 _106_ _279_/a_27_47# 0.00751f
C586 clknet_2_1__leaf_clk _220_/a_199_47# 2.53e-20
C587 _308_/a_1270_413# _078_ 1.46e-19
C588 VPWR rebuffer1/a_75_212# 0.231f
C589 _321_/a_448_47# _321_/a_639_47# 4.61e-19
C590 _074_ _080_ 0.235f
C591 _340_/a_652_21# _340_/a_562_413# 9.35e-20
C592 _340_/a_1182_261# _340_/a_1602_47# 0.144f
C593 _340_/a_476_47# _340_/a_381_47# 0.0356f
C594 _228_/a_382_297# _049_ 2.38e-19
C595 _088_ _170_/a_299_297# 0.0463f
C596 net2 _208_/a_505_21# 0.147f
C597 _052_ _170_/a_81_21# 0.00659f
C598 _302_/a_109_297# cal_count\[3\] 0.0172f
C599 _094_ fanout44/a_27_47# 5.81e-20
C600 _308_/a_1108_47# net24 3.38e-21
C601 _136_ _133_ 7.12e-19
C602 VPWR net54 0.751f
C603 VPWR _169_/a_373_53# 1.08e-19
C604 _038_ clkbuf_2_3__f_clk/a_110_47# 7.24e-21
C605 trim_mask\[0\] _162_/a_27_47# 0.00115f
C606 ctlp[0] _314_/a_448_47# 5.04e-19
C607 cal_count\[1\] _123_ 0.0248f
C608 net43 _319_/a_805_47# 0.00206f
C609 _090_ _240_/a_109_297# 3.4e-19
C610 _309_/a_27_47# _078_ 0.0158f
C611 _292_/a_493_297# net16 6.13e-20
C612 net3 _014_ 0.0126f
C613 _259_/a_27_297# trim_val\[3\] 7.23e-21
C614 trim[0] net33 0.00267f
C615 _326_/a_27_47# _310_/a_193_47# 2.81e-21
C616 _326_/a_193_47# _310_/a_27_47# 1.33e-20
C617 net47 _144_/a_27_47# 4.17e-20
C618 _048_ wire42/a_75_212# 0.0537f
C619 _337_/a_448_47# _337_/a_639_47# 4.61e-19
C620 _188_/a_27_47# _134_ 3.59e-21
C621 net31 _112_ 1.19e-20
C622 trim[0] trim_mask\[1\] 7.26e-19
C623 net47 clknet_2_3__leaf_clk 0.481f
C624 net2 _001_ 0.148f
C625 _062_ _203_/a_145_75# 6.54e-20
C626 net45 _330_/a_193_47# 5.82e-23
C627 VPWR _310_/a_1283_21# 0.392f
C628 _088_ _227_/a_368_53# 5.81e-20
C629 _066_ _092_ 0.0852f
C630 net9 _339_/a_1056_47# 2.24e-19
C631 _051_ _337_/a_1283_21# 7.17e-19
C632 _250_/a_109_47# mask\[5\] 0.00214f
C633 _333_/a_27_47# _055_ 3.54e-19
C634 net28 _022_ 8.53e-19
C635 _035_ _338_/a_652_21# 1.2e-19
C636 _329_/a_27_47# _025_ 1.44e-20
C637 net27 _224_/a_113_297# 0.0472f
C638 VPWR result[4] 0.264f
C639 _110_ _116_ 0.503f
C640 VPWR _068_ 0.958f
C641 _041_ net18 0.00946f
C642 net8 clknet_2_2__leaf_clk 0.0058f
C643 _321_/a_27_47# _101_ 0.457f
C644 _341_/a_193_47# _230_/a_59_75# 6.55e-21
C645 clknet_2_1__leaf_clk _020_ 0.349f
C646 _338_/a_1182_261# net18 0.00254f
C647 _320_/a_543_47# _121_ 5.22e-20
C648 output23/a_27_47# _080_ 0.00498f
C649 VPWR _327_/a_1217_47# 1.49e-19
C650 _041_ _129_ 0.00225f
C651 _094_ _137_/a_68_297# 5.3e-20
C652 ctlp[2] net39 0.0015f
C653 _313_/a_27_47# _045_ 9.7e-21
C654 _288_/a_59_75# trimb[4] 2.54e-20
C655 _302_/a_109_297# _038_ 0.0017f
C656 _169_/a_215_311# _318_/a_543_47# 4.71e-20
C657 _307_/a_543_47# _004_ 0.00161f
C658 _129_ _297_/a_129_47# 2.57e-19
C659 trim_val\[3\] trim_mask\[1\] 1.05e-21
C660 net28 _313_/a_1283_21# 0.15f
C661 _322_/a_761_289# _078_ 3.39e-21
C662 net50 _336_/a_27_47# 2.82e-21
C663 clknet_0_clk _016_ 7.76e-21
C664 _164_/a_161_47# _096_ 0.00593f
C665 output21/a_27_47# _078_ 1.82e-19
C666 VPWR fanout43/a_27_47# 0.456f
C667 net4 _261_/a_113_47# 1.27e-19
C668 VPWR _335_/a_1217_47# 6.15e-20
C669 net3 _243_/a_27_297# 0.00209f
C670 mask\[7\] net14 3.5e-19
C671 VPWR output35/a_27_47# 0.494f
C672 trimb[0] trimb[1] 0.0464f
C673 _245_/a_27_297# _245_/a_109_297# 0.171f
C674 VPWR _311_/a_448_47# 0.0796f
C675 VPWR net27 1.22f
C676 clknet_2_1__leaf_clk _222_/a_199_47# 4.52e-19
C677 net44 clknet_2_3__leaf_clk 0.00416f
C678 net46 net30 3.76e-21
C679 _042_ _084_ 6.34e-21
C680 _341_/a_448_47# _304_/a_761_289# 1.91e-20
C681 _340_/a_193_47# _063_ 3.52e-20
C682 _340_/a_1182_261# _041_ 4.68e-21
C683 _340_/a_586_47# net47 1.54e-19
C684 _325_/a_27_47# clknet_2_1__leaf_clk 0.253f
C685 _065_ _077_ 0.173f
C686 _106_ _118_ 0.00544f
C687 net27 net53 1.42e-19
C688 _311_/a_448_47# net53 0.00818f
C689 _123_ _001_ 0.0103f
C690 net23 net22 0.00148f
C691 _071_ net30 1.26e-19
C692 trim[0] output33/a_27_47# 9.86e-19
C693 output31/a_27_47# trim[2] 0.00245f
C694 VPWR _332_/a_805_47# 0.00186f
C695 input4/a_27_47# rstn 0.195f
C696 VPWR _186_/a_109_297# 0.00469f
C697 _028_ _098_ 1.39e-20
C698 _340_/a_193_47# _037_ 0.0834f
C699 _319_/a_193_47# _120_ 1.44e-20
C700 clknet_2_0__leaf_clk _075_ 0.00194f
C701 _038_ cal_count\[3\] 0.0219f
C702 _327_/a_193_47# _111_ 1.95e-19
C703 _277_/a_75_212# _117_ 0.212f
C704 en_co_clk _243_/a_373_47# 7.94e-20
C705 _337_/a_543_47# _090_ 8.11e-22
C706 VPWR _125_ 0.441f
C707 _134_ _298_/a_292_297# 6.3e-20
C708 _309_/a_1217_47# _078_ 0.0011f
C709 _309_/a_1462_47# mask\[0\] 2.34e-20
C710 _110_ _328_/a_27_47# 5.55e-20
C711 _301_/a_47_47# clknet_2_3__leaf_clk 0.117f
C712 _104_ trim_mask\[3\] 0.257f
C713 _323_/a_1108_47# _043_ 0.00275f
C714 _261_/a_113_47# _063_ 5.07e-19
C715 _309_/a_1270_413# net24 4.39e-19
C716 _337_/a_1270_413# net44 2.59e-19
C717 clknet_0_clk _028_ 8.37e-20
C718 clkbuf_2_2__f_clk/a_110_47# trim_mask\[4\] 2.14e-19
C719 output35/a_27_47# _161_/a_68_297# 0.00583f
C720 _341_/a_27_47# clknet_2_3__leaf_clk 0.8f
C721 output41/a_27_47# net41 0.223f
C722 net27 _009_ 3.17e-19
C723 net2 mask\[1\] 3.22e-20
C724 _233_/a_109_297# cal 0.00146f
C725 _233_/a_27_297# net1 0.0853f
C726 _058_ _111_ 0.0177f
C727 _074_ _082_ 0.102f
C728 _239_/a_277_297# _048_ 0.0172f
C729 _136_ net4 3e-20
C730 net12 net20 0.103f
C731 _291_/a_35_297# net16 0.00571f
C732 _081_ _245_/a_27_297# 1.53e-19
C733 VPWR _306_/a_27_47# 0.502f
C734 _247_/a_373_47# _018_ 2.47e-19
C735 clk _119_ 2.39e-20
C736 _110_ _266_/a_68_297# 0.106f
C737 _187_/a_27_413# _332_/a_1283_21# 1.11e-19
C738 _048_ _206_/a_27_93# 2.7e-20
C739 _338_/a_1296_47# net18 2.78e-19
C740 trim[1] trim_val\[0\] 0.00234f
C741 _326_/a_27_47# _224_/a_113_297# 2.65e-20
C742 _122_ _295_/a_113_47# 1.45e-19
C743 ctln[6] clk 1.18e-20
C744 _149_/a_68_297# _303_/a_193_47# 1.58e-19
C745 _189_/a_408_47# _075_ 1.97e-19
C746 _071_ _072_ 0.0822f
C747 _111_ _332_/a_27_47# 2.22e-19
C748 _231_/a_161_47# _067_ 0.0161f
C749 net51 _049_ 0.00338f
C750 _316_/a_761_289# _095_ 9.69e-20
C751 clk _331_/a_651_413# 0.00269f
C752 _323_/a_27_47# net47 0.296f
C753 clknet_2_2__leaf_clk clknet_2_3__leaf_clk 1.6e-20
C754 net44 net20 0.0362f
C755 _314_/a_1108_47# _011_ 1.26e-19
C756 cal_itt\[0\] net2 0.00936f
C757 ctln[6] _331_/a_1283_21# 1.83e-21
C758 _058_ rebuffer3/a_75_212# 0.0034f
C759 net4 _119_ 0.648f
C760 _104_ _330_/a_1283_21# 0.00112f
C761 _208_/a_505_21# _070_ 5.95e-22
C762 _327_/a_193_47# _065_ 1.61e-20
C763 cal_itt\[2\] _305_/a_1108_47# 0.00769f
C764 _306_/a_543_47# _306_/a_1108_47# 7.99e-20
C765 _306_/a_193_47# _306_/a_651_413# 0.0346f
C766 _076_ _202_/a_79_21# 9.14e-20
C767 cal_itt\[0\] _305_/a_1283_21# 1.59e-20
C768 _071_ _305_/a_193_47# 1.05e-19
C769 trim_val\[4\] _278_/a_27_47# 3.3e-19
C770 _118_ _278_/a_109_297# 5.24e-19
C771 net42 _226_/a_27_47# 4.92e-20
C772 _329_/a_639_47# trim_mask\[3\] 1.18e-19
C773 _326_/a_448_47# result[5] 2.53e-19
C774 _035_ _339_/a_476_47# 1.11e-21
C775 _331_/a_761_289# _331_/a_639_47# 3.16e-19
C776 _331_/a_27_47# _331_/a_1217_47# 2.56e-19
C777 _060_ calibrate 0.0293f
C778 net54 _093_ 0.0386f
C779 _037_ _136_ 0.00132f
C780 en_co_clk _206_/a_206_47# 2.33e-19
C781 _325_/a_193_47# mask\[6\] 0.0254f
C782 _245_/a_27_297# _016_ 0.11f
C783 _245_/a_109_47# net52 3.87e-21
C784 _001_ _067_ 9.01e-19
C785 _256_/a_27_297# trim_mask\[4\] 0.0098f
C786 _001_ _070_ 0.105f
C787 VPWR _235_/a_382_297# 0.00496f
C788 _325_/a_651_413# _042_ 4.99e-19
C789 _041_ _338_/a_652_21# 1.13e-19
C790 _308_/a_27_47# net14 0.00787f
C791 _185_/a_68_297# _232_/a_32_297# 1.12e-19
C792 _189_/a_218_47# _088_ 1.17e-19
C793 _338_/a_27_47# _338_/a_1602_47# 2.39e-19
C794 _338_/a_193_47# _338_/a_1032_413# 0.0573f
C795 VPWR _317_/a_27_47# 0.476f
C796 _058_ _065_ 8.88e-19
C797 VPWR _326_/a_27_47# 0.466f
C798 _086_ _310_/a_543_47# 2.06e-21
C799 _050_ _336_/a_448_47# 8.9e-21
C800 VPWR net10 0.359f
C801 _113_ _108_ 9.94e-20
C802 _058_ _135_ 1.25e-19
C803 mask\[7\] net52 0.195f
C804 _169_/a_109_53# state\[1\] 0.134f
C805 _292_/a_215_47# _122_ 0.107f
C806 _074_ _310_/a_448_47# 0.00248f
C807 _339_/a_1032_413# _129_ 6.61e-20
C808 _060_ net45 1.14e-19
C809 net25 clknet_2_1__leaf_clk 0.367f
C810 net4 _087_ 2.67e-20
C811 _229_/a_27_297# _089_ 0.113f
C812 ctlp[7] _313_/a_1462_47# 1.98e-20
C813 _327_/a_1462_47# _111_ 7.11e-19
C814 _170_/a_81_21# _170_/a_384_47# 0.00138f
C815 _092_ net40 1.05e-19
C816 _051_ _260_/a_250_297# 2.34e-19
C817 _297_/a_47_47# _297_/a_129_47# 0.00369f
C818 _116_ clknet_2_2__leaf_clk 2.26e-20
C819 output31/a_27_47# _055_ 0.224f
C820 _104_ _181_/a_68_297# 2.89e-19
C821 _078_ _208_/a_76_199# 9.44e-19
C822 _325_/a_27_47# _313_/a_27_47# 7.57e-19
C823 ctln[3] _057_ 0.0412f
C824 _259_/a_27_297# _335_/a_543_47# 0.00351f
C825 _341_/a_448_47# cal_count\[3\] 0.0163f
C826 clkbuf_2_1__f_clk/a_110_47# _141_/a_27_47# 4.1e-19
C827 mask\[0\] mask\[2\] 1.12e-19
C828 _341_/a_1217_47# clknet_2_3__leaf_clk 0.00112f
C829 net4 _266_/a_150_297# 1.65e-19
C830 net2 _108_ 4.09e-20
C831 net2 _332_/a_543_47# 1.14e-19
C832 _012_ cal 0.00363f
C833 _060_ _065_ 5.79e-21
C834 _323_/a_27_47# net44 0.00995f
C835 _092_ _003_ 4.53e-21
C836 state\[2\] _051_ 0.601f
C837 _116_ net11 5.63e-20
C838 _298_/a_292_297# cal_count\[2\] 7.38e-20
C839 _040_ clknet_0_clk 0.0218f
C840 VPWR _306_/a_1217_47# 7.1e-20
C841 _101_ _046_ 0.00309f
C842 net2 _288_/a_145_75# 0.00219f
C843 trim_val\[0\] clknet_2_3__leaf_clk 3.62e-22
C844 _321_/a_27_47# _248_/a_27_297# 1.74e-20
C845 trim_mask\[1\] _334_/a_1108_47# 9.68e-21
C846 _272_/a_299_297# _334_/a_543_47# 1.49e-19
C847 _053_ _262_/a_205_47# 1.72e-19
C848 _340_/a_1182_261# _339_/a_1032_413# 5.58e-20
C849 _340_/a_1032_413# _339_/a_1182_261# 7.12e-20
C850 _113_ _031_ 0.00248f
C851 _303_/a_543_47# _035_ 2.78e-21
C852 net15 _318_/a_193_47# 7.1e-21
C853 _336_/a_27_47# _052_ 3.51e-20
C854 cal_itt\[0\] _123_ 0.00309f
C855 mask\[1\] _319_/a_1270_413# 8.1e-21
C856 _329_/a_1283_21# _334_/a_27_47# 1.95e-20
C857 _095_ _098_ 2.5e-20
C858 trim_mask\[0\] _333_/a_543_47# 1.73e-19
C859 _294_/a_150_297# _130_ 0.00145f
C860 _303_/a_1108_47# net18 2.39e-19
C861 _029_ _332_/a_805_47# 9.23e-20
C862 VPWR _318_/a_543_47# 0.205f
C863 _315_/a_193_47# output41/a_27_47# 5.23e-20
C864 output18/a_27_47# net17 1.18e-20
C865 trim_mask\[0\] _265_/a_384_47# 0.0102f
C866 result[5] _074_ 2.8e-19
C867 net35 net33 0.415f
C868 _190_/a_215_47# clkbuf_2_3__f_clk/a_110_47# 3.87e-20
C869 net54 _243_/a_109_47# 1.14e-19
C870 _185_/a_68_297# net55 3.84e-19
C871 _181_/a_68_297# _067_ 3.4e-20
C872 _060_ _243_/a_109_297# 0.0101f
C873 _058_ _112_ 0.0036f
C874 _323_/a_1217_47# net47 6.03e-19
C875 _312_/a_639_47# net20 0.00117f
C876 net12 _028_ 0.00295f
C877 clknet_2_1__leaf_clk _310_/a_543_47# 0.0364f
C878 clknet_0_clk _095_ 0.161f
C879 _064_ _027_ 0.00142f
C880 _022_ _085_ 0.00128f
C881 output12/a_27_47# output13/a_27_47# 5.8e-21
C882 _336_/a_1108_47# _335_/a_27_47# 1.46e-19
C883 VPWR _233_/a_109_47# 1.28e-19
C884 net9 _267_/a_59_75# 3.47e-19
C885 output20/a_27_47# ctlp[6] 0.372f
C886 _341_/a_448_47# _038_ 0.186f
C887 _341_/a_805_47# _136_ 4.9e-19
C888 _301_/a_47_47# _301_/a_377_297# 0.00899f
C889 _326_/a_1283_21# net26 2.13e-20
C890 _331_/a_1108_47# _028_ 0.00379f
C891 _331_/a_448_47# clknet_2_2__leaf_clk 6.21e-19
C892 _331_/a_193_47# trim_mask\[4\] 5.49e-19
C893 net15 _317_/a_639_47# 0.00103f
C894 _281_/a_253_47# _316_/a_1283_21# 1.96e-20
C895 _317_/a_193_47# _317_/a_651_413# 0.0276f
C896 _317_/a_543_47# _317_/a_1108_47# 7.99e-20
C897 _325_/a_1462_47# mask\[6\] 0.00198f
C898 mask\[6\] mask\[3\] 8.02e-19
C899 _233_/a_109_47# valid 1.39e-19
C900 _328_/a_27_47# clknet_2_2__leaf_clk 0.862f
C901 _132_ output40/a_27_47# 7.25e-21
C902 _326_/a_543_47# _326_/a_1108_47# 7.99e-20
C903 _326_/a_193_47# _326_/a_651_413# 0.0346f
C904 _325_/a_1283_21# _078_ 1.76e-20
C905 _104_ _088_ 0.102f
C906 _263_/a_79_21# _263_/a_382_297# 0.00145f
C907 _074_ rebuffer6/a_27_47# 7.09e-21
C908 net49 _332_/a_193_47# 1.04e-19
C909 trim_val\[1\] _108_ 0.139f
C910 _112_ _332_/a_27_47# 6.36e-19
C911 _324_/a_1283_21# clknet_2_3__leaf_clk 5.51e-21
C912 VPWR _317_/a_1217_47# 2.84e-20
C913 _328_/a_543_47# _328_/a_651_413# 0.0572f
C914 _328_/a_761_289# _328_/a_1270_413# 2.6e-19
C915 _328_/a_193_47# _328_/a_639_47# 2.28e-19
C916 _328_/a_1108_47# trim_mask\[2\] 7.08e-20
C917 _341_/a_27_47# _341_/a_193_47# 0.64f
C918 VPWR _326_/a_1217_47# 1.17e-19
C919 VPWR _271_/a_75_212# 0.201f
C920 _050_ _033_ 9.69e-19
C921 _336_/a_193_47# _108_ 3.78e-19
C922 _320_/a_1283_21# net44 0.345f
C923 _291_/a_35_297# net40 2.3e-20
C924 _288_/a_59_75# net33 0.00892f
C925 net13 _337_/a_805_47# 4.26e-19
C926 _088_ net55 0.044f
C927 _309_/a_543_47# net14 0.0113f
C928 _106_ _062_ 0.0208f
C929 _293_/a_299_297# _129_ 0.00178f
C930 VPWR cal_itt\[3\] 0.557f
C931 _318_/a_193_47# _318_/a_761_289# 0.181f
C932 _318_/a_27_47# _318_/a_543_47# 0.115f
C933 _340_/a_476_47# cal_count\[2\] 2.99e-20
C934 cal_itt\[2\] _069_ 1.61e-19
C935 net42 _052_ 5.72e-21
C936 _103_ en_co_clk 1.3e-20
C937 _104_ _335_/a_1283_21# 8.76e-20
C938 _066_ net46 2.54e-19
C939 trim_val\[2\] net46 0.00547f
C940 net44 _312_/a_805_47# 0.00316f
C941 _110_ _279_/a_314_297# 0.004f
C942 VPWR _300_/a_285_47# 0.00701f
C943 _312_/a_193_47# _312_/a_651_413# 0.0346f
C944 _312_/a_543_47# _312_/a_1108_47# 7.99e-20
C945 _336_/a_639_47# net46 1.79e-19
C946 _312_/a_193_47# net19 4.79e-20
C947 _074_ net29 3.58e-19
C948 VPWR _305_/a_27_47# 0.48f
C949 _320_/a_1108_47# net52 2.33e-20
C950 _306_/a_543_47# clknet_2_0__leaf_clk 1.49e-19
C951 _306_/a_193_47# net45 4.54e-22
C952 clknet_2_1__leaf_clk _311_/a_1108_47# 0.00435f
C953 _015_ state\[2\] 8.91e-20
C954 _329_/a_448_47# net46 2.48e-19
C955 net28 net14 0.398f
C956 _078_ _314_/a_27_47# 9.87e-19
C957 _068_ _202_/a_79_21# 0.00218f
C958 cal_itt\[0\] _067_ 0.942f
C959 _043_ mask\[4\] 0.0799f
C960 VPWR _262_/a_205_47# 1.16e-19
C961 _323_/a_761_289# net19 0.00947f
C962 _041_ _339_/a_476_47# 0.043f
C963 mask\[1\] mask\[0\] 0.0883f
C964 trim[2] trim[3] 0.0486f
C965 cal_itt\[0\] _070_ 0.00994f
C966 net47 _339_/a_1140_413# 6.59e-19
C967 _305_/a_805_47# net51 1.55e-19
C968 _114_ _334_/a_448_47# 2.07e-19
C969 trim_val\[2\] _334_/a_639_47# 1.48e-19
C970 net16 net46 0.0561f
C971 _323_/a_543_47# _323_/a_651_413# 0.0572f
C972 _323_/a_761_289# _323_/a_1270_413# 2.6e-19
C973 _323_/a_193_47# _323_/a_639_47# 2.28e-19
C974 output24/a_27_47# mask\[1\] 2.25e-19
C975 _104_ _108_ 0.0175f
C976 _037_ _339_/a_27_47# 2.81e-20
C977 state\[2\] _242_/a_79_21# 0.00202f
C978 _140_/a_68_297# _101_ 0.00187f
C979 _040_ _245_/a_27_297# 1.86e-19
C980 VPWR _315_/a_448_47# 0.0865f
C981 _107_ _089_ 0.00335f
C982 _337_/a_1108_47# _092_ 2.64e-19
C983 net14 ctln[0] 0.00137f
C984 net3 _316_/a_1108_47# 9.66e-19
C985 trim_mask\[2\] _333_/a_761_289# 4.36e-20
C986 calibrate _227_/a_109_93# 3.13e-20
C987 _233_/a_27_297# _233_/a_109_297# 0.171f
C988 trim_mask\[2\] _115_ 0.0818f
C989 _292_/a_78_199# net47 0.00916f
C990 _306_/a_193_47# _065_ 1.17e-20
C991 _315_/a_448_47# valid 0.00102f
C992 _308_/a_651_413# _006_ 1.65e-21
C993 clkbuf_0_clk/a_110_47# _190_/a_215_47# 0.00413f
C994 en_co_clk clkc 0.00312f
C995 _103_ _050_ 0.0737f
C996 net34 _057_ 0.00351f
C997 net12 _205_/a_27_47# 0.00291f
C998 _306_/a_1108_47# _305_/a_543_47# 5.01e-19
C999 net31 net38 2.61e-20
C1000 _093_ _317_/a_27_47# 6.21e-22
C1001 calibrate _317_/a_193_47# 4.8e-21
C1002 net43 _321_/a_805_47# 0.00401f
C1003 _153_/a_27_47# _044_ 0.195f
C1004 VPWR _011_ 0.714f
C1005 _326_/a_761_289# _074_ 0.00387f
C1006 _320_/a_193_47# _320_/a_448_47# 0.0605f
C1007 _320_/a_761_289# _320_/a_1108_47# 0.0512f
C1008 _320_/a_27_47# _320_/a_651_413# 9.73e-19
C1009 _192_/a_639_47# _049_ 2.36e-20
C1010 _119_ _279_/a_396_47# 0.309f
C1011 _309_/a_193_47# _081_ 0.00817f
C1012 _168_/a_27_413# _052_ 0.00112f
C1013 net24 _007_ 3.43e-21
C1014 _189_/a_27_47# _306_/a_1108_47# 4.15e-22
C1015 _008_ _321_/a_1108_47# 1.37e-20
C1016 result[3] net14 8.01e-20
C1017 ctlp[0] _086_ 1.04e-19
C1018 net12 _040_ 1.15e-20
C1019 _331_/a_1462_47# trim_mask\[4\] 0.00102f
C1020 _228_/a_79_21# clone7/a_27_47# 2.84e-20
C1021 clknet_2_2__leaf_clk _028_ 0.00261f
C1022 net7 net45 1.3e-20
C1023 _237_/a_76_199# _090_ 0.192f
C1024 trim_mask\[4\] _260_/a_93_21# 0.0854f
C1025 cal_count\[1\] _144_/a_27_47# 0.0563f
C1026 _062_ _278_/a_109_297# 2.94e-21
C1027 _317_/a_761_289# _014_ 6.4e-19
C1028 _317_/a_543_47# clknet_2_0__leaf_clk 0.0306f
C1029 _317_/a_193_47# net45 0.0265f
C1030 _308_/a_193_47# _307_/a_761_289# 6.96e-20
C1031 _308_/a_27_47# _307_/a_543_47# 1.1e-20
C1032 _328_/a_1217_47# clknet_2_2__leaf_clk 1.2e-21
C1033 net27 output29/a_27_47# 1.35e-21
C1034 net17 _339_/a_381_47# 8.46e-20
C1035 VPWR _269_/a_384_47# 1.86e-19
C1036 _067_ _108_ 2.97e-19
C1037 _341_/a_761_289# _341_/a_805_47# 3.69e-19
C1038 _341_/a_193_47# _341_/a_1217_47# 2.36e-20
C1039 _341_/a_543_47# _341_/a_639_47# 0.0138f
C1040 net24 mask\[3\] 0.0026f
C1041 clk ctln[0] 0.0136f
C1042 _043_ _020_ 2.16e-21
C1043 net44 _205_/a_27_47# 0.00463f
C1044 _303_/a_27_47# _063_ 4.53e-21
C1045 _303_/a_543_47# _041_ 3.11e-20
C1046 net47 _303_/a_805_47# 0.00316f
C1047 _303_/a_27_47# _338_/a_381_47# 7.45e-21
C1048 cal_itt\[2\] _255_/a_27_47# 8.54e-20
C1049 _210_/a_113_297# _039_ 6.7e-20
C1050 net4 _279_/a_206_47# 3.06e-19
C1051 _146_/a_68_297# _018_ 0.00373f
C1052 _333_/a_193_47# _333_/a_543_47# 0.23f
C1053 _333_/a_27_47# _333_/a_1283_21# 0.0436f
C1054 _312_/a_193_47# _155_/a_68_297# 1.03e-20
C1055 net23 _245_/a_27_297# 0.0304f
C1056 net16 _332_/a_448_47# 4.27e-19
C1057 _040_ net44 0.279f
C1058 net12 _095_ 6.2e-21
C1059 net27 mask\[6\] 0.348f
C1060 net12 _322_/a_1283_21# 0.00904f
C1061 output8/a_27_47# trim[3] 6.33e-19
C1062 _265_/a_81_21# _265_/a_384_47# 0.00138f
C1063 net43 _102_ 0.00624f
C1064 _309_/a_1108_47# _101_ 0.00106f
C1065 net4 ctln[0] 0.0219f
C1066 _226_/a_27_47# _098_ 1.11e-20
C1067 _324_/a_1108_47# net44 0.248f
C1068 _312_/a_1462_47# net19 9.63e-20
C1069 _320_/a_1283_21# _209_/a_27_47# 0.0148f
C1070 calibrate _054_ 6.74e-19
C1071 VPWR _305_/a_1217_47# 9.49e-21
C1072 _048_ _337_/a_193_47# 1.59e-20
C1073 VPWR _250_/a_109_297# 0.204f
C1074 _026_ net46 0.0054f
C1075 calibrate net30 0.00261f
C1076 _308_/a_543_47# _308_/a_1108_47# 7.99e-20
C1077 _308_/a_193_47# _308_/a_651_413# 0.0346f
C1078 en_co_clk clkbuf_2_3__f_clk/a_110_47# 6.9e-19
C1079 _324_/a_1283_21# _323_/a_27_47# 0.00384f
C1080 clknet_2_1__leaf_clk net15 1.21f
C1081 _041_ _339_/a_1224_47# 0.00127f
C1082 _169_/a_215_311# clone7/a_27_47# 6.11e-19
C1083 net15 _319_/a_761_289# 0.00236f
C1084 _019_ _321_/a_1108_47# 4.75e-19
C1085 _114_ _031_ 0.00585f
C1086 _090_ _241_/a_388_297# 3.97e-19
C1087 _307_/a_1283_21# _307_/a_1108_47# 0.234f
C1088 _307_/a_761_289# _307_/a_651_413# 0.0977f
C1089 _307_/a_543_47# _307_/a_448_47# 0.0498f
C1090 _307_/a_27_47# _307_/a_639_47# 0.00188f
C1091 _307_/a_193_47# _307_/a_1270_413# 1.46e-19
C1092 _305_/a_543_47# _203_/a_59_75# 7.48e-19
C1093 _094_ clkbuf_2_0__f_clk/a_110_47# 0.00233f
C1094 clknet_0_clk _226_/a_27_47# 5.47e-20
C1095 result[0] _307_/a_1283_21# 1.48e-19
C1096 net9 _053_ 6.64e-20
C1097 _231_/a_161_47# clknet_2_3__leaf_clk 0.00105f
C1098 _250_/a_109_297# net53 0.0106f
C1099 VPWR _319_/a_1283_21# 0.368f
C1100 _322_/a_1283_21# net44 0.337f
C1101 _318_/a_193_47# state\[1\] 2.44e-21
C1102 _300_/a_47_47# _300_/a_285_47# 0.0175f
C1103 _318_/a_1283_21# net45 0.33f
C1104 net28 net52 0.00395f
C1105 _309_/a_27_47# _308_/a_27_47# 6.48e-21
C1106 _233_/a_373_47# calibrate 0.00153f
C1107 _233_/a_27_297# _012_ 0.152f
C1108 _340_/a_27_47# _001_ 1.09e-19
C1109 net45 net30 0.0259f
C1110 net30 rebuffer3/a_75_212# 2.94e-19
C1111 _036_ net47 0.0224f
C1112 _325_/a_193_47# _321_/a_193_47# 1.07e-20
C1113 net43 _006_ 0.00128f
C1114 _059_ _096_ 0.0162f
C1115 clone1/a_27_47# _170_/a_81_21# 8.07e-20
C1116 net52 _158_/a_68_297# 8.6e-20
C1117 net24 _310_/a_1283_21# 3.61e-22
C1118 _187_/a_212_413# net2 1.13e-20
C1119 en_co_clk _130_ 3.39e-20
C1120 _337_/a_193_47# _120_ 9.35e-20
C1121 _337_/a_761_289# en_co_clk 0.00551f
C1122 _100_ net41 0.0383f
C1123 _262_/a_27_47# _262_/a_205_47# 0.00762f
C1124 _262_/a_109_297# _262_/a_193_297# 0.0927f
C1125 _303_/a_193_47# net19 0.0168f
C1126 clkbuf_2_0__f_clk/a_110_47# _192_/a_505_280# 0.00268f
C1127 _001_ clknet_2_3__leaf_clk 0.381f
C1128 _065_ net30 0.634f
C1129 _339_/a_27_47# _339_/a_562_413# 6.02e-19
C1130 _339_/a_193_47# _339_/a_381_47# 0.149f
C1131 _339_/a_476_47# _339_/a_1032_413# 0.00329f
C1132 net37 _055_ 0.0027f
C1133 net13 _320_/a_448_47# 3.09e-19
C1134 _172_/a_150_297# _108_ 5.76e-19
C1135 _317_/a_639_47# state\[1\] 1.48e-19
C1136 _317_/a_1462_47# net45 0.00342f
C1137 output15/a_27_47# net15 0.191f
C1138 _320_/a_543_47# _040_ 0.0357f
C1139 input2/a_27_47# output5/a_27_47# 4.01e-20
C1140 _122_ net37 7.04e-21
C1141 _321_/a_1270_413# mask\[2\] 6e-20
C1142 _105_ net30 0.0135f
C1143 _315_/a_193_47# _315_/a_1270_413# 1.46e-19
C1144 _315_/a_27_47# _315_/a_639_47# 0.00188f
C1145 _315_/a_543_47# _315_/a_448_47# 0.0498f
C1146 _315_/a_761_289# _315_/a_651_413# 0.0977f
C1147 _315_/a_1283_21# _315_/a_1108_47# 0.234f
C1148 net21 _045_ 0.00973f
C1149 _337_/a_193_47# _076_ 3.9e-20
C1150 _104_ _170_/a_299_297# 0.021f
C1151 clknet_2_2__leaf_clk _279_/a_314_297# 6e-20
C1152 VPWR _336_/a_1270_413# 0.00122f
C1153 net19 _152_/a_68_297# 0.00139f
C1154 _218_/a_113_297# _101_ 2.38e-19
C1155 _110_ net50 0.0487f
C1156 _116_ trim_mask\[3\] 6.05e-19
C1157 _117_ trim_val\[3\] 0.00648f
C1158 _134_ _295_/a_113_47# 1.68e-19
C1159 clknet_2_1__leaf_clk _049_ 5.62e-19
C1160 VPWR _329_/a_1108_47# 0.307f
C1161 ctln[2] _334_/a_1283_21# 8.69e-19
C1162 net8 _334_/a_448_47# 0.00107f
C1163 _319_/a_761_289# _049_ 9.8e-19
C1164 _232_/a_32_297# _192_/a_174_21# 0.0237f
C1165 _323_/a_27_47# _044_ 4.75e-20
C1166 net46 net40 0.33f
C1167 _319_/a_27_47# net30 1.48e-19
C1168 _333_/a_448_47# _333_/a_639_47# 4.61e-19
C1169 output14/a_27_47# ctlp[1] 5.95e-22
C1170 net36 net34 0.206f
C1171 _136_ _193_/a_109_297# 4.88e-19
C1172 _243_/a_373_47# _049_ 1.84e-19
C1173 _286_/a_535_374# _123_ 0.00177f
C1174 trim_mask\[0\] _048_ 0.124f
C1175 _012_ _315_/a_1283_21# 4.1e-20
C1176 calibrate _315_/a_651_413# 0.0256f
C1177 _322_/a_543_47# _320_/a_1283_21# 1.58e-20
C1178 _326_/a_27_47# mask\[6\] 5.74e-21
C1179 en input4/a_27_47# 1.99e-20
C1180 _209_/a_27_47# _205_/a_27_47# 0.0152f
C1181 _334_/a_1270_413# net34 5.17e-20
C1182 _065_ _072_ 0.128f
C1183 clkbuf_0_clk/a_110_47# en_co_clk 3.63e-19
C1184 VPWR _021_ 0.367f
C1185 mask\[4\] net21 2.5e-19
C1186 state\[0\] _316_/a_27_47# 2.65e-19
C1187 _246_/a_27_297# net52 0.191f
C1188 _246_/a_109_47# _101_ 0.00183f
C1189 net12 _083_ 0.00879f
C1190 en_co_clk cal_count\[3\] 0.00244f
C1191 _308_/a_193_47# net43 0.0431f
C1192 _308_/a_761_289# _005_ 9.52e-19
C1193 _328_/a_761_289# _025_ 1.82e-19
C1194 _053_ clone7/a_27_47# 8.25e-20
C1195 VPWR net9 1.25f
C1196 clknet_2_0__leaf_clk _315_/a_639_47# 1.44e-19
C1197 net45 _315_/a_651_413# 0.0122f
C1198 clkbuf_2_1__f_clk/a_110_47# clknet_2_0__leaf_clk 0.0448f
C1199 cal_itt\[1\] _230_/a_59_75# 9.72e-19
C1200 _305_/a_651_413# _072_ 0.00299f
C1201 VPWR output16/a_27_47# 0.299f
C1202 _040_ _209_/a_27_47# 3.17e-19
C1203 _021_ net53 0.0551f
C1204 _194_/a_113_297# net30 7.16e-19
C1205 _305_/a_193_47# _065_ 7.67e-20
C1206 _107_ _279_/a_490_47# 5.99e-19
C1207 _092_ net19 0.00741f
C1208 _110_ _330_/a_1108_47# 0.0152f
C1209 _116_ _330_/a_1283_21# 1.78e-20
C1210 _181_/a_68_297# clknet_2_3__leaf_clk 3.62e-21
C1211 _327_/a_27_47# net18 0.0237f
C1212 net15 _313_/a_27_47# 0.00107f
C1213 _305_/a_1283_21# net2 1.58e-19
C1214 net8 _108_ 4.46e-19
C1215 _323_/a_1108_47# mask\[4\] 0.02f
C1216 _321_/a_193_47# mask\[3\] 2.82e-19
C1217 _321_/a_761_289# net25 4.62e-21
C1218 _305_/a_543_47# _305_/a_1108_47# 7.99e-20
C1219 _305_/a_193_47# _305_/a_651_413# 0.0346f
C1220 _281_/a_103_199# _090_ 0.139f
C1221 net12 _208_/a_218_374# 6.82e-19
C1222 net12 _207_/a_109_297# 4.37e-19
C1223 VPWR _313_/a_761_289# 0.225f
C1224 _239_/a_474_297# _049_ 0.00562f
C1225 _052_ _098_ 0.141f
C1226 _309_/a_27_47# _309_/a_543_47# 0.115f
C1227 _309_/a_193_47# _309_/a_761_289# 0.181f
C1228 _083_ net44 0.00381f
C1229 _061_ _135_ 5.21e-19
C1230 _262_/a_465_47# _105_ 0.00164f
C1231 _277_/a_75_212# _057_ 6.35e-20
C1232 VPWR trim[2] 0.606f
C1233 _021_ _009_ 2.08e-20
C1234 _106_ _227_/a_209_311# 5.89e-20
C1235 _332_/a_448_47# net40 6.16e-19
C1236 _323_/a_543_47# _000_ 1.96e-19
C1237 _192_/a_27_47# _096_ 4.47e-19
C1238 _322_/a_1283_21# _209_/a_27_47# 9.72e-19
C1239 cal_itt\[1\] clknet_0_clk 0.0151f
C1240 _335_/a_27_47# net18 2.82e-20
C1241 _206_/a_206_47# _049_ 2.08e-19
C1242 _269_/a_81_21# _269_/a_299_297# 0.0821f
C1243 _339_/a_1182_261# _339_/a_1296_47# 1.84e-19
C1244 _339_/a_1032_413# _339_/a_1224_47# 0.00536f
C1245 _081_ mask\[2\] 0.0816f
C1246 net34 _332_/a_1108_47# 4.6e-20
C1247 _189_/a_27_47# _189_/a_408_47# 0.0212f
C1248 clknet_0_clk _052_ 1.9e-20
C1249 _107_ _092_ 0.0107f
C1250 _126_ trimb[4] 0.00797f
C1251 _327_/a_27_47# _302_/a_27_297# 8.93e-19
C1252 net31 _333_/a_27_47# 1.1e-20
C1253 output31/a_27_47# _333_/a_1283_21# 0.00807f
C1254 trim[1] _108_ 3.27e-19
C1255 _038_ en_co_clk 2.04e-19
C1256 net12 _226_/a_27_47# 2.37e-20
C1257 _050_ _331_/a_27_47# 7.37e-19
C1258 net44 _207_/a_109_297# 2.44e-19
C1259 _053_ _122_ 0.203f
C1260 VPWR _234_/a_109_297# 0.00643f
C1261 _292_/a_215_47# _339_/a_1602_47# 9.75e-21
C1262 _276_/a_59_75# _335_/a_27_47# 0.00105f
C1263 net8 _031_ 0.00114f
C1264 cal_itt\[3\] _202_/a_79_21# 4.21e-22
C1265 net28 _155_/a_150_297# 8.39e-21
C1266 _078_ _018_ 0.00646f
C1267 clk _330_/a_448_47# 7.28e-19
C1268 _041_ rebuffer5/a_161_47# 4.56e-21
C1269 _279_/a_396_47# _279_/a_206_47# 0.00414f
C1270 _279_/a_204_297# _279_/a_314_297# 0.14f
C1271 _279_/a_27_47# _279_/a_490_47# 2.12e-19
C1272 _303_/a_543_47# _303_/a_1108_47# 7.99e-20
C1273 _303_/a_193_47# _303_/a_651_413# 0.0346f
C1274 _074_ _042_ 0.448f
C1275 _141_/a_27_47# clknet_0_clk 0.0326f
C1276 _253_/a_81_21# net25 8.35e-19
C1277 _290_/a_297_47# cal_count\[0\] 5.23e-19
C1278 mask\[5\] net19 0.033f
C1279 result[1] net45 3.22e-20
C1280 _341_/a_193_47# _231_/a_161_47# 3.72e-19
C1281 _237_/a_218_374# _092_ 5.89e-19
C1282 net54 _337_/a_193_47# 3.54e-19
C1283 _295_/a_113_47# cal_count\[2\] 5.18e-19
C1284 _006_ _080_ 9.8e-20
C1285 _048_ _090_ 0.549f
C1286 cal_itt\[0\] clknet_2_3__leaf_clk 0.042f
C1287 _322_/a_543_47# _205_/a_27_47# 0.00358f
C1288 net44 _226_/a_27_47# 4.7e-21
C1289 _314_/a_543_47# net14 0.00272f
C1290 _019_ _320_/a_193_47# 1.24e-19
C1291 _321_/a_193_47# _310_/a_1283_21# 3.21e-20
C1292 _321_/a_27_47# _310_/a_1108_47# 3.19e-20
C1293 net2 _123_ 0.0507f
C1294 _326_/a_543_47# _078_ 0.00326f
C1295 _324_/a_1283_21# _324_/a_1108_47# 0.234f
C1296 _324_/a_761_289# _324_/a_651_413# 0.0977f
C1297 _324_/a_543_47# _324_/a_448_47# 0.0498f
C1298 _324_/a_27_47# _324_/a_639_47# 0.00188f
C1299 _324_/a_193_47# _324_/a_1270_413# 1.46e-19
C1300 VPWR clone7/a_27_47# 0.24f
C1301 _306_/a_193_47# _204_/a_75_212# 5.35e-19
C1302 net13 _322_/a_448_47# 0.00788f
C1303 mask\[2\] _016_ 2.53e-20
C1304 net13 _092_ 0.0585f
C1305 _308_/a_1462_47# net43 0.00384f
C1306 _316_/a_193_47# net41 0.0258f
C1307 _097_ _233_/a_27_297# 7.99e-20
C1308 _319_/a_1108_47# net45 0.00151f
C1309 _319_/a_651_413# clknet_2_0__leaf_clk 0.00604f
C1310 mask\[1\] _245_/a_109_297# 0.0105f
C1311 _341_/a_193_47# _001_ 2.94e-19
C1312 _048_ _242_/a_382_297# 0.0158f
C1313 output21/a_27_47# net28 0.00665f
C1314 _189_/a_27_47# clone1/a_27_47# 4.91e-19
C1315 _309_/a_1283_21# net43 0.271f
C1316 _309_/a_193_47# net23 6.13e-20
C1317 clknet_2_0__leaf_clk _096_ 0.00191f
C1318 _325_/a_761_289# _046_ 0.00305f
C1319 _327_/a_27_47# trim_mask\[0\] 8.88e-19
C1320 _327_/a_1217_47# net18 5.39e-20
C1321 VPWR output8/a_27_47# 0.301f
C1322 mask\[7\] _314_/a_27_47# 1.54e-19
C1323 _263_/a_79_21# _226_/a_27_47# 2.58e-19
C1324 _305_/a_761_289# _002_ 0.0231f
C1325 _120_ _090_ 0.027f
C1326 net9 _300_/a_47_47# 0.00155f
C1327 net16 _111_ 7.22e-22
C1328 trim[4] net34 0.0953f
C1329 net5 trim[4] 2.79e-19
C1330 _319_/a_1108_47# _065_ 8.33e-19
C1331 net50 clknet_2_2__leaf_clk 0.0136f
C1332 _320_/a_1108_47# _208_/a_76_199# 6.13e-20
C1333 _030_ _173_/a_27_47# 1.16e-20
C1334 _292_/a_215_47# cal_count\[2\] 4.49e-19
C1335 _146_/a_150_297# _042_ 4.96e-19
C1336 _322_/a_193_47# _322_/a_448_47# 0.0594f
C1337 _322_/a_761_289# _322_/a_1108_47# 0.0512f
C1338 _322_/a_27_47# _322_/a_651_413# 9.73e-19
C1339 _056_ net33 0.0733f
C1340 _110_ _327_/a_1108_47# 0.00254f
C1341 _305_/a_805_47# clknet_2_1__leaf_clk 1.33e-20
C1342 _320_/a_193_47# _017_ 0.316f
C1343 _250_/a_27_297# clknet_2_1__leaf_clk 0.045f
C1344 clknet_2_3__leaf_clk _108_ 1.78e-19
C1345 net22 _315_/a_27_47# 2.45e-20
C1346 _259_/a_109_297# _064_ 0.0116f
C1347 VPWR _055_ 0.517f
C1348 _043_ _311_/a_1108_47# 2.32e-20
C1349 _327_/a_543_47# _136_ 0.00139f
C1350 _066_ rebuffer3/a_75_212# 1.04e-19
C1351 trim_mask\[1\] _336_/a_27_47# 4.07e-20
C1352 cal_itt\[1\] net47 0.00158f
C1353 _336_/a_27_47# _336_/a_761_289# 0.0532f
C1354 VPWR _122_ 1.1f
C1355 net9 _029_ 0.00231f
C1356 _081_ mask\[1\] 0.274f
C1357 clknet_2_1__leaf_clk _319_/a_543_47# 6.88e-19
C1358 _319_/a_27_47# _319_/a_1108_47# 0.102f
C1359 _319_/a_193_47# _319_/a_1283_21# 0.0424f
C1360 _319_/a_761_289# _319_/a_543_47# 0.21f
C1361 VPWR _073_ 0.396f
C1362 net13 mask\[5\] 9.08e-20
C1363 _083_ _209_/a_27_47# 1.29e-20
C1364 _308_/a_193_47# _080_ 6.57e-20
C1365 _249_/a_27_297# _249_/a_109_47# 0.00393f
C1366 _117_ _335_/a_543_47# 1.78e-19
C1367 _110_ _335_/a_1108_47# 1.75e-19
C1368 _280_/a_75_212# net46 0.00431f
C1369 net43 _092_ 2.25e-20
C1370 clk _027_ 0.00154f
C1371 _053_ _091_ 3.98e-19
C1372 _022_ _074_ 1.49e-19
C1373 net35 _136_ 4.2e-19
C1374 _066_ _065_ 0.107f
C1375 _303_/a_761_289# _000_ 3.71e-19
C1376 _097_ _315_/a_1283_21# 7.8e-21
C1377 _048_ trim_mask\[4\] 2.84e-20
C1378 VPWR _299_/a_27_413# 0.245f
C1379 _243_/a_27_297# _100_ 0.0743f
C1380 _103_ _049_ 0.0125f
C1381 _047_ _332_/a_1283_21# 1.23e-20
C1382 net2 _067_ 3.42e-19
C1383 _087_ _075_ 0.00266f
C1384 _089_ _062_ 5.29e-21
C1385 _324_/a_761_289# mask\[5\] 2.14e-19
C1386 net2 _070_ 0.38f
C1387 _059_ _098_ 1.04e-19
C1388 _034_ _099_ 1.39e-21
C1389 _317_/a_27_47# _316_/a_651_413# 2.78e-20
C1390 _282_/a_68_297# net30 1.63e-19
C1391 _110_ rebuffer2/a_75_212# 9.17e-19
C1392 _292_/a_78_199# cal_count\[1\] 0.00316f
C1393 _292_/a_215_47# _128_ 0.00844f
C1394 _305_/a_1283_21# _067_ 2.17e-19
C1395 _277_/a_75_212# _027_ 3.83e-21
C1396 _305_/a_1283_21# _070_ 0.00139f
C1397 trim_mask\[4\] _330_/a_27_47# 1.35e-21
C1398 clknet_2_2__leaf_clk _330_/a_1108_47# 0.0234f
C1399 _125_ _129_ 0.0064f
C1400 state\[0\] _167_/a_161_47# 0.00282f
C1401 _060_ _051_ 0.26f
C1402 net22 clknet_2_0__leaf_clk 0.0104f
C1403 net12 _052_ 0.00248f
C1404 net30 _278_/a_27_47# 0.00632f
C1405 _219_/a_109_297# _218_/a_113_297# 1.95e-20
C1406 net13 _019_ 0.105f
C1407 net4 _027_ 2.02e-19
C1408 _136_ _332_/a_761_289# 2.34e-20
C1409 _135_ net16 0.00779f
C1410 _104_ _336_/a_193_47# 0.287f
C1411 _059_ clknet_0_clk 0.0276f
C1412 _249_/a_109_297# mask\[4\] 0.0015f
C1413 _316_/a_1462_47# net41 0.00184f
C1414 _074_ _313_/a_1283_21# 3.85e-19
C1415 _053_ _302_/a_373_47# 0.00193f
C1416 _232_/a_32_297# net55 0.0307f
C1417 _329_/a_27_47# _064_ 3.82e-21
C1418 _092_ _118_ 9.2e-20
C1419 _331_/a_1108_47# _052_ 2.8e-19
C1420 net4 _195_/a_218_47# 7.62e-19
C1421 mask\[1\] _016_ 0.00155f
C1422 _330_/a_651_413# net19 0.00323f
C1423 VPWR ctln[1] 0.176f
C1424 trim_mask\[2\] _334_/a_193_47# 0.00989f
C1425 VPWR _304_/a_1283_21# 0.389f
C1426 _082_ _006_ 0.00503f
C1427 fanout46/a_27_47# _033_ 0.0622f
C1428 _335_/a_543_47# _119_ 1.05e-20
C1429 net14 _310_/a_805_47# 5.85e-19
C1430 _327_/a_1270_413# _024_ 4.33e-20
C1431 _327_/a_1217_47# trim_mask\[0\] 6.68e-21
C1432 net30 _204_/a_75_212# 0.0371f
C1433 mask\[7\] _314_/a_1217_47# 6.99e-20
C1434 output33/a_27_47# _056_ 0.171f
C1435 _130_ output40/a_27_47# 5.69e-21
C1436 _200_/a_80_21# net19 0.00424f
C1437 ctln[5] output12/a_27_47# 2.68e-20
C1438 _053_ _340_/a_381_47# 8.64e-20
C1439 mask\[6\] _250_/a_109_297# 0.0116f
C1440 net12 _311_/a_27_47# 7.12e-21
C1441 output31/a_27_47# net31 0.235f
C1442 state\[2\] _228_/a_79_21# 2.59e-20
C1443 _239_/a_694_21# _100_ 0.0016f
C1444 net43 mask\[5\] 2.36e-21
C1445 _306_/a_1108_47# clknet_0_clk 3.47e-19
C1446 _328_/a_543_47# _058_ 0.0026f
C1447 _322_/a_193_47# _019_ 0.253f
C1448 _019_ _248_/a_109_297# 0.00891f
C1449 mask\[2\] _205_/a_27_47# 3.88e-19
C1450 net48 net33 1.38e-20
C1451 _194_/a_113_297# _066_ 0.00936f
C1452 clkbuf_2_1__f_clk/a_110_47# _078_ 0.0012f
C1453 _121_ _192_/a_174_21# 7.67e-21
C1454 net48 trim_mask\[1\] 1.98e-20
C1455 trim_mask\[0\] output35/a_27_47# 9.4e-19
C1456 _272_/a_299_297# trim_val\[2\] 0.0171f
C1457 _202_/a_382_297# _202_/a_297_47# 8.13e-19
C1458 output37/a_27_47# net37 0.218f
C1459 _127_ net33 0.0235f
C1460 net13 _017_ 9.55e-19
C1461 _273_/a_59_75# net46 0.0121f
C1462 trim_mask\[1\] _336_/a_1217_47# 2.91e-21
C1463 _320_/a_1283_21# mask\[1\] 0.0914f
C1464 _200_/a_80_21# _107_ 9.99e-19
C1465 _336_/a_543_47# _336_/a_805_47# 0.00171f
C1466 _336_/a_761_289# _336_/a_1217_47# 4.2e-19
C1467 _336_/a_1108_47# _336_/a_1270_413# 0.00645f
C1468 _079_ _315_/a_27_47# 1.26e-20
C1469 cal_itt\[0\] _341_/a_193_47# 0.00165f
C1470 _336_/a_543_47# _264_/a_27_297# 8.17e-20
C1471 _040_ mask\[2\] 0.0363f
C1472 _123_ _067_ 5.69e-19
C1473 _281_/a_337_297# _092_ 0.00685f
C1474 _319_/a_1283_21# _319_/a_1462_47# 0.0074f
C1475 _319_/a_1108_47# _319_/a_1217_47# 0.00742f
C1476 net44 _311_/a_27_47# 0.304f
C1477 net10 net18 0.228f
C1478 _104_ net55 0.0665f
C1479 VPWR _091_ 0.348f
C1480 _290_/a_27_413# _127_ 6.21e-19
C1481 _048_ _283_/a_75_212# 8.48e-21
C1482 net16 _112_ 0.0667f
C1483 VPWR _256_/a_109_297# 0.184f
C1484 _272_/a_299_297# net16 0.00392f
C1485 _249_/a_109_297# _020_ 0.00169f
C1486 calibrate _316_/a_27_47# 2.84e-20
C1487 trim_mask\[0\] _332_/a_805_47# 8.96e-19
C1488 _329_/a_193_47# _329_/a_448_47# 0.0642f
C1489 _329_/a_761_289# _329_/a_1108_47# 0.0512f
C1490 _329_/a_27_47# _329_/a_651_413# 9.73e-19
C1491 VPWR _321_/a_1283_21# 0.39f
C1492 _115_ _334_/a_193_47# 0.00186f
C1493 net43 _019_ 6.48e-19
C1494 _093_ clone7/a_27_47# 3.26e-20
C1495 _204_/a_75_212# _072_ 2.13e-20
C1496 _024_ _053_ 5.87e-20
C1497 clknet_2_1__leaf_clk _313_/a_193_47# 0.597f
C1498 net54 _090_ 0.259f
C1499 VPWR _337_/a_1283_21# 0.36f
C1500 _327_/a_27_47# _265_/a_81_21# 1.9e-21
C1501 _300_/a_47_47# _122_ 3.83e-19
C1502 net50 _257_/a_373_47# 1.65e-19
C1503 clknet_2_0__leaf_clk _316_/a_761_289# 6.07e-21
C1504 _014_ _316_/a_193_47# 0.0222f
C1505 net45 _316_/a_27_47# 0.305f
C1506 _321_/a_1283_21# net53 0.00285f
C1507 cal_count\[1\] _036_ 2.79e-20
C1508 _341_/a_1283_21# _058_ 1.27e-20
C1509 state\[2\] _169_/a_215_311# 0.0739f
C1510 _015_ _060_ 0.0686f
C1511 _126_ net33 0.46f
C1512 _188_/a_27_47# _061_ 0.212f
C1513 _266_/a_68_297# _108_ 0.00179f
C1514 VPWR _138_/a_27_47# 0.257f
C1515 _111_ net40 0.0034f
C1516 _322_/a_1283_21# mask\[2\] 8.98e-21
C1517 _058_ _333_/a_27_47# 0.00266f
C1518 _101_ _311_/a_543_47# 3.18e-21
C1519 _128_ _291_/a_117_297# 2.33e-19
C1520 _290_/a_27_413# _126_ 0.0944f
C1521 net14 net41 0.0116f
C1522 net54 _242_/a_382_297# 1.17e-20
C1523 _020_ mask\[4\] 1.22e-19
C1524 _329_/a_761_289# net9 0.00805f
C1525 _064_ _106_ 0.00126f
C1526 _309_/a_193_47# _216_/a_113_297# 4.52e-20
C1527 _079_ clknet_2_0__leaf_clk 0.0308f
C1528 _134_ net37 1.79e-20
C1529 clknet_2_2__leaf_clk _052_ 2.54e-20
C1530 _052_ _260_/a_584_47# 0.00318f
C1531 _327_/a_1108_47# clknet_2_2__leaf_clk 3.11e-19
C1532 _327_/a_27_47# trim_mask\[4\] 0.00152f
C1533 clknet_0_clk _203_/a_59_75# 0.00228f
C1534 net46 net19 0.00497f
C1535 _341_/a_193_47# _108_ 1.06e-19
C1536 _325_/a_1270_413# net13 1.29e-19
C1537 VPWR _340_/a_381_47# 0.104f
C1538 clknet_0_clk _192_/a_27_47# 0.0127f
C1539 _041_ net51 4.43e-20
C1540 _175_/a_68_297# rebuffer1/a_75_212# 0.0215f
C1541 _333_/a_1283_21# net37 9e-19
C1542 _333_/a_193_47# rebuffer1/a_75_212# 1.72e-20
C1543 _333_/a_27_47# _332_/a_27_47# 5.12e-19
C1544 ctlp[1] _223_/a_109_297# 8.48e-19
C1545 VPWR _253_/a_384_47# 3.4e-19
C1546 net23 mask\[2\] 2.03e-20
C1547 _071_ net19 4.17e-19
C1548 net45 sample 4.04e-20
C1549 mask\[6\] _021_ 0.0173f
C1550 net26 clknet_2_3__leaf_clk 8.28e-19
C1551 net3 _092_ 0.0901f
C1552 _337_/a_761_289# _049_ 0.00926f
C1553 rebuffer3/a_75_212# net40 0.0347f
C1554 net33 _172_/a_68_297# 0.00219f
C1555 _210_/a_113_297# _210_/a_199_47# 2.42e-19
C1556 _277_/a_75_212# _032_ 0.109f
C1557 _125_ _297_/a_47_47# 0.001f
C1558 _337_/a_27_47# net30 2.09e-19
C1559 _335_/a_1108_47# clknet_2_2__leaf_clk 8.02e-20
C1560 _335_/a_27_47# trim_mask\[4\] 1.83e-22
C1561 trim_val\[1\] _172_/a_150_297# 0.00172f
C1562 trim_mask\[1\] _172_/a_68_297# 0.105f
C1563 _107_ net46 0.00233f
C1564 _341_/a_639_47# net46 0.00108f
C1565 _168_/a_207_413# net55 1.95e-21
C1566 _067_ _070_ 0.0808f
C1567 net12 _059_ 4.92e-20
C1568 net4 _032_ 3.38e-21
C1569 VPWR _198_/a_109_47# 1.68e-19
C1570 _333_/a_1108_47# net46 0.236f
C1571 result[2] clknet_2_1__leaf_clk 2.89e-20
C1572 clk net41 3.86e-20
C1573 _243_/a_109_47# clone7/a_27_47# 1.5e-19
C1574 mask\[1\] _205_/a_27_47# 9.85e-20
C1575 net45 _003_ 1.36e-21
C1576 _071_ _107_ 2.52e-19
C1577 VPWR _331_/a_761_289# 0.232f
C1578 _286_/a_535_374# clknet_2_3__leaf_clk 2.46e-19
C1579 _065_ net40 1.05e-19
C1580 VPWR _215_/a_109_297# 0.00533f
C1581 _332_/a_1283_21# clknet_2_2__leaf_clk 2.36e-21
C1582 _051_ _227_/a_109_93# 0.122f
C1583 _264_/a_27_297# _106_ 0.206f
C1584 mask\[6\] _313_/a_761_289# 1.34e-21
C1585 net44 _311_/a_1217_47# 4.56e-19
C1586 _135_ net40 7.13e-19
C1587 VPWR _258_/a_27_297# 0.205f
C1588 net27 _312_/a_543_47# 2.14e-19
C1589 _053_ _260_/a_250_297# 0.00772f
C1590 VPWR _024_ 0.523f
C1591 VPWR _147_/a_27_47# 0.286f
C1592 _233_/a_373_47# _013_ 5.79e-20
C1593 _329_/a_193_47# _026_ 0.228f
C1594 _094_ _337_/a_448_47# 0.025f
C1595 VPWR rstn 0.198f
C1596 mask\[1\] _040_ 0.41f
C1597 net28 _314_/a_27_47# 0.0118f
C1598 _051_ _235_/a_297_47# 1.85e-20
C1599 _036_ _001_ 0.00281f
C1600 _319_/a_1108_47# _282_/a_68_297# 4.85e-20
C1601 _102_ net29 2.32e-20
C1602 _306_/a_448_47# clk 7.3e-22
C1603 _262_/a_193_297# clkbuf_2_3__f_clk/a_110_47# 0.00178f
C1604 _064_ _278_/a_109_297# 5.72e-19
C1605 net4 net41 1.15e-19
C1606 _327_/a_1108_47# trim_val\[0\] 1.75e-21
C1607 _065_ _003_ 0.0016f
C1608 _059_ net44 0.00165f
C1609 net12 _306_/a_1108_47# 0.00227f
C1610 _317_/a_448_47# net14 1.74e-19
C1611 net45 _316_/a_1217_47# 4.56e-19
C1612 _314_/a_27_47# _158_/a_68_297# 2.64e-21
C1613 _187_/a_212_413# clknet_2_3__leaf_clk 0.00159f
C1614 _325_/a_1270_413# net43 2.06e-19
C1615 _255_/a_27_47# net42 5.16e-19
C1616 _103_ _254_/a_109_297# 0.0123f
C1617 _119_ _170_/a_81_21# 5.69e-21
C1618 state\[2\] _053_ 0.13f
C1619 clknet_2_0__leaf_clk clknet_0_clk 0.825f
C1620 _313_/a_27_47# _313_/a_193_47# 0.582f
C1621 _058_ _333_/a_1217_47# 1.11e-19
C1622 cal_count\[3\] _049_ 5.13e-20
C1623 clk _171_/a_27_47# 0.0124f
C1624 net46 _279_/a_27_47# 0.00143f
C1625 result[7] _078_ 2.78e-20
C1626 _308_/a_1283_21# _039_ 0.0101f
C1627 _309_/a_651_413# net25 1.1e-19
C1628 VPWR _101_ 1.68f
C1629 _185_/a_68_297# _095_ 5.79e-20
C1630 _331_/a_27_47# _049_ 2.8e-20
C1631 VPWR _338_/a_1032_413# 0.433f
C1632 _306_/a_1108_47# net44 0.249f
C1633 _059_ _263_/a_79_21# 0.0912f
C1634 _075_ _099_ 3.69e-19
C1635 input3/a_75_212# en 0.193f
C1636 _062_ _092_ 0.0592f
C1637 _333_/a_651_413# rebuffer2/a_75_212# 1.13e-19
C1638 _326_/a_193_47# _023_ 0.259f
C1639 _312_/a_193_47# _221_/a_109_297# 8.06e-20
C1640 _326_/a_543_47# mask\[7\] 0.00755f
C1641 _326_/a_761_289# _102_ 1.46e-19
C1642 _333_/a_1270_413# _108_ 2.09e-19
C1643 trim_mask\[3\] net50 0.158f
C1644 VPWR _297_/a_285_47# 9.42e-19
C1645 net4 _171_/a_27_47# 1.45e-20
C1646 _101_ net53 0.0933f
C1647 trim_val\[3\] _057_ 0.0206f
C1648 net37 cal_count\[2\] 1.17e-19
C1649 _286_/a_76_199# _338_/a_193_47# 0.00114f
C1650 _194_/a_113_297# net40 6.94e-19
C1651 _109_ _332_/a_193_47# 0.00209f
C1652 trim_val\[0\] _332_/a_1283_21# 0.0699f
C1653 _208_/a_76_199# _208_/a_535_374# 6.64e-19
C1654 _305_/a_1108_47# clknet_0_clk 1.24e-19
C1655 _066_ _278_/a_27_47# 3.47e-20
C1656 _304_/a_1108_47# _065_ 0.00918f
C1657 clk _317_/a_448_47# 0.00205f
C1658 net43 _314_/a_1283_21# 0.281f
C1659 _340_/a_476_47# cal_count\[0\] 7.26e-21
C1660 _336_/a_1283_21# net40 3.24e-21
C1661 net23 mask\[1\] 0.958f
C1662 net22 _078_ 0.0116f
C1663 _257_/a_109_297# net46 5.48e-21
C1664 _315_/a_193_47# net14 0.0145f
C1665 _051_ _054_ 0.0162f
C1666 _187_/a_27_413# _136_ 1.29e-19
C1667 _189_/a_408_47# clknet_0_clk 0.0319f
C1668 _051_ net30 0.705f
C1669 _340_/a_27_47# net2 1.21e-19
C1670 _290_/a_207_413# net34 0.0122f
C1671 _316_/a_1283_21# _096_ 6.93e-20
C1672 _101_ _009_ 5.33e-21
C1673 net15 net21 1.66e-20
C1674 VPWR output37/a_27_47# 0.457f
C1675 clk _203_/a_145_75# 9.6e-19
C1676 _136_ _268_/a_75_212# 0.0029f
C1677 VPWR _320_/a_27_47# 0.429f
C1678 _238_/a_75_212# _316_/a_193_47# 2.94e-19
C1679 net12 _203_/a_59_75# 2.86e-19
C1680 output16/a_27_47# output39/a_27_47# 8.52e-19
C1681 output27/a_27_47# output28/a_27_47# 0.00249f
C1682 _340_/a_1602_47# _132_ 6.93e-20
C1683 _167_/a_161_47# calibrate 1.95e-20
C1684 VPWR _260_/a_250_297# 0.332f
C1685 net43 _310_/a_27_47# 0.311f
C1686 _322_/a_1270_413# mask\[3\] 3.62e-19
C1687 _321_/a_651_413# clknet_2_0__leaf_clk 4.04e-20
C1688 _303_/a_543_47# _068_ 0.0027f
C1689 VPWR _328_/a_651_413# 0.133f
C1690 net2 _144_/a_27_47# 6.55e-20
C1691 cal_itt\[0\] _303_/a_805_47# 8.9e-20
C1692 _074_ net14 0.926f
C1693 _324_/a_27_47# _311_/a_1283_21# 2.45e-20
C1694 output20/a_27_47# _312_/a_761_289# 0.0034f
C1695 net2 clknet_2_3__leaf_clk 0.106f
C1696 net13 state\[0\] 0.143f
C1697 _337_/a_651_413# clknet_2_0__leaf_clk 1.08e-20
C1698 _108_ _279_/a_314_297# 0.0131f
C1699 net28 _314_/a_1217_47# 2.55e-20
C1700 result[6] _314_/a_639_47# 3.88e-19
C1701 _323_/a_27_47# net26 4.04e-19
C1702 _309_/a_1108_47# _310_/a_1108_47# 1.55e-20
C1703 _015_ _317_/a_193_47# 5.56e-20
C1704 trim_mask\[3\] _330_/a_1108_47# 0.00165f
C1705 _289_/a_150_297# net40 2.58e-19
C1706 _167_/a_161_47# net45 0.00532f
C1707 _262_/a_193_297# cal_count\[3\] 5.67e-19
C1708 _071_ net43 0.00629f
C1709 VPWR _312_/a_448_47# 0.0824f
C1710 state\[2\] VPWR 1.13f
C1711 _110_ _030_ 0.00981f
C1712 _014_ net14 3.31e-19
C1713 VPWR _323_/a_651_413# 0.134f
C1714 VPWR _307_/a_193_47# 0.581f
C1715 _074_ _143_/a_68_297# 2.68e-20
C1716 ctlp[3] ctlp[4] 0.00165f
C1717 clone1/a_27_47# _098_ 0.0229f
C1718 _010_ _223_/a_109_297# 0.0124f
C1719 net44 _203_/a_59_75# 1.65e-19
C1720 _068_ _190_/a_27_47# 0.00106f
C1721 _313_/a_543_47# _313_/a_639_47# 0.0138f
C1722 _313_/a_193_47# _313_/a_1217_47# 2.36e-20
C1723 _313_/a_761_289# _313_/a_805_47# 3.69e-19
C1724 _336_/a_448_47# clkbuf_2_2__f_clk/a_110_47# 9.38e-19
C1725 _312_/a_448_47# net53 7.79e-20
C1726 _051_ _072_ 8.19e-19
C1727 _337_/a_1108_47# _065_ 9.33e-19
C1728 net31 net37 0.249f
C1729 net46 _118_ 6.17e-20
C1730 _304_/a_27_47# _066_ 2.59e-21
C1731 clknet_0_clk clone1/a_27_47# 1.68e-20
C1732 VPWR _134_ 0.618f
C1733 _076_ rebuffer5/a_161_47# 0.0222f
C1734 net8 _114_ 3.77e-19
C1735 input2/a_27_47# _131_ 0.0115f
C1736 VPWR _341_/a_1270_413# 4.89e-19
C1737 _321_/a_543_47# clknet_2_1__leaf_clk 0.0142f
C1738 _312_/a_448_47# _009_ 0.158f
C1739 VPWR _333_/a_1283_21# 0.359f
C1740 _340_/a_27_47# _123_ 0.519f
C1741 _275_/a_299_297# _335_/a_27_47# 1.03e-19
C1742 _275_/a_81_21# _335_/a_193_47# 0.00133f
C1743 _294_/a_68_297# _125_ 6.58e-20
C1744 _337_/a_193_47# _319_/a_1283_21# 3.92e-20
C1745 _337_/a_27_47# _319_/a_1108_47# 3.29e-20
C1746 _050_ en_co_clk 0.112f
C1747 ctlp[1] _010_ 0.00232f
C1748 cal_count\[0\] _338_/a_193_47# 1.45e-19
C1749 _124_ _338_/a_476_47# 0.00285f
C1750 _330_/a_193_47# _330_/a_1270_413# 1.46e-19
C1751 _330_/a_27_47# _330_/a_639_47# 3.82e-19
C1752 _330_/a_543_47# _330_/a_448_47# 0.0498f
C1753 _330_/a_761_289# _330_/a_651_413# 0.0977f
C1754 _330_/a_1283_21# _330_/a_1108_47# 0.234f
C1755 clk _014_ 0.0041f
C1756 VPWR _308_/a_448_47# 0.0854f
C1757 _025_ net46 0.00717f
C1758 net12 clknet_2_0__leaf_clk 1.37e-19
C1759 _015_ _318_/a_1283_21# 4.1e-20
C1760 state\[2\] _318_/a_27_47# 6.3e-19
C1761 calibrate _229_/a_27_297# 0.0647f
C1762 _079_ _078_ 0.0139f
C1763 VPWR _237_/a_505_21# 0.224f
C1764 _123_ clknet_2_3__leaf_clk 0.156f
C1765 _004_ net22 0.00877f
C1766 mask\[1\] _208_/a_218_374# 1.34e-19
C1767 net45 _331_/a_543_47# 0.155f
C1768 net9 _304_/a_193_47# 0.0014f
C1769 _242_/a_297_47# _049_ 0.00675f
C1770 net27 _249_/a_27_297# 4e-20
C1771 VPWR _320_/a_1217_47# 2.71e-20
C1772 net10 trim_mask\[4\] 5.9e-22
C1773 VPWR _339_/a_1602_47# 0.199f
C1774 ctln[2] ctln[3] 0.00303f
C1775 net43 _310_/a_1217_47# 0.00157f
C1776 _208_/a_76_199# rebuffer4/a_27_47# 5.21e-19
C1777 _328_/a_1283_21# _271_/a_75_212# 2.79e-19
C1778 net4 _014_ 5.39e-20
C1779 _297_/a_129_47# _132_ 0.0018f
C1780 mask\[0\] _121_ 0.00291f
C1781 _047_ net33 0.0023f
C1782 ctlp[6] net19 1.79e-21
C1783 net44 clknet_2_0__leaf_clk 0.173f
C1784 _339_/a_193_47# _286_/a_505_21# 1.07e-19
C1785 _110_ net33 1.3e-20
C1786 _325_/a_27_47# _325_/a_1217_47# 2.56e-19
C1787 _325_/a_761_289# _325_/a_639_47# 3.16e-19
C1788 _110_ trim_mask\[1\] 0.0802f
C1789 cal_itt\[1\] _231_/a_161_47# 3.16e-19
C1790 VPWR _324_/a_193_47# 0.6f
C1791 mask\[3\] rebuffer5/a_161_47# 1.65e-21
C1792 _110_ _336_/a_761_289# 0.00634f
C1793 _104_ clknet_2_3__leaf_clk 1.02e-19
C1794 _074_ net52 0.0103f
C1795 _189_/a_408_47# net12 4.34e-22
C1796 VPWR _307_/a_1462_47# 2.57e-19
C1797 mask\[4\] _311_/a_1108_47# 0.0402f
C1798 _226_/a_197_47# _062_ 0.00623f
C1799 _226_/a_109_47# _075_ 1.72e-20
C1800 ctlp[7] net27 1.3e-20
C1801 net15 _241_/a_105_352# 0.00353f
C1802 _313_/a_448_47# _010_ 0.159f
C1803 _033_ clkbuf_2_2__f_clk/a_110_47# 0.065f
C1804 _334_/a_1108_47# _057_ 2.11e-20
C1805 _324_/a_193_47# net53 0.00258f
C1806 _304_/a_1270_413# _067_ 8.41e-20
C1807 VPWR _322_/a_27_47# 0.48f
C1808 VPWR _248_/a_27_297# 0.288f
C1809 VPWR _241_/a_297_47# 0.00555f
C1810 net9 net18 0.0456f
C1811 _321_/a_805_47# _042_ 2.51e-19
C1812 _337_/a_1283_21# _206_/a_27_93# 0.00185f
C1813 VPWR _257_/a_27_297# 0.22f
C1814 net27 _220_/a_113_297# 0.00977f
C1815 _305_/a_1108_47# net44 9.86e-21
C1816 _314_/a_27_47# _085_ 1.58e-21
C1817 net16 net38 0.0476f
C1818 cal_itt\[1\] _001_ 0.00103f
C1819 _278_/a_27_47# net40 0.039f
C1820 trim_mask\[2\] fanout46/a_27_47# 0.00289f
C1821 _181_/a_68_297# _181_/a_150_297# 0.00477f
C1822 output13/a_27_47# _318_/a_543_47# 1.95e-19
C1823 _316_/a_27_47# _316_/a_448_47# 0.0859f
C1824 _316_/a_193_47# _316_/a_1108_47# 0.125f
C1825 _189_/a_408_47# net44 1.14e-20
C1826 _248_/a_27_297# net53 0.221f
C1827 _322_/a_27_47# net53 2.38e-20
C1828 VPWR _303_/a_448_47# 0.0834f
C1829 _200_/a_80_21# _062_ 0.125f
C1830 net50 _335_/a_1283_21# 0.00823f
C1831 net4 _243_/a_27_297# 3.76e-21
C1832 trim_mask\[3\] _335_/a_1108_47# 0.00393f
C1833 VPWR cal_count\[2\] 0.615f
C1834 _116_ _104_ 1.8e-20
C1835 _171_/a_27_47# _279_/a_396_47# 2.25e-20
C1836 cal_count\[0\] _338_/a_796_47# 2.06e-20
C1837 _330_/a_543_47# _027_ 0.0336f
C1838 _330_/a_761_289# net46 0.159f
C1839 _134_ _300_/a_47_47# 7.21e-19
C1840 _301_/a_377_297# net2 7.35e-19
C1841 _336_/a_27_47# _119_ 0.0126f
C1842 clkbuf_0_clk/a_110_47# _202_/a_297_47# 6.77e-20
C1843 VPWR _005_ 0.428f
C1844 _067_ clknet_2_3__leaf_clk 0.0407f
C1845 _078_ clknet_0_clk 3.17e-20
C1846 clknet_2_3__leaf_clk _070_ 2.49e-20
C1847 _341_/a_193_47# net2 9.68e-20
C1848 _341_/a_1108_47# _300_/a_285_47# 8.66e-20
C1849 _158_/a_150_297# net29 2.03e-19
C1850 VPWR _219_/a_109_297# 0.00866f
C1851 net50 _108_ 0.13f
C1852 _320_/a_193_47# net45 4.53e-20
C1853 _320_/a_543_47# clknet_2_0__leaf_clk 0.0014f
C1854 output36/a_27_47# net34 0.0153f
C1855 output33/a_27_47# _047_ 4.2e-22
C1856 VPWR _309_/a_639_47# 4.66e-19
C1857 _162_/a_27_47# net32 5.19e-19
C1858 _020_ _311_/a_1108_47# 1.4e-20
C1859 VPWR _190_/a_655_47# 0.00379f
C1860 _030_ clknet_2_2__leaf_clk 0.179f
C1861 mask\[7\] _251_/a_109_47# 0.00419f
C1862 _102_ _251_/a_109_297# 6.74e-19
C1863 _238_/a_75_212# net14 2.88e-21
C1864 _204_/a_75_212# _003_ 0.109f
C1865 net9 _340_/a_1182_261# 9.58e-19
C1866 _319_/a_193_47# _101_ 0.00234f
C1867 _079_ _004_ 0.149f
C1868 _041_ clknet_2_1__leaf_clk 0.0101f
C1869 _255_/a_27_47# clknet_0_clk 9.47e-19
C1870 _102_ _042_ 1.59e-20
C1871 _219_/a_109_297# net53 8.05e-19
C1872 _307_/a_761_289# calibrate 3.2e-20
C1873 _307_/a_543_47# _074_ 0.0152f
C1874 output34/a_27_47# net46 8.6e-19
C1875 net4 _336_/a_543_47# 0.0072f
C1876 _334_/a_27_47# _334_/a_761_289# 0.0701f
C1877 _314_/a_193_47# _314_/a_761_289# 0.186f
C1878 _314_/a_27_47# _314_/a_543_47# 0.115f
C1879 VPWR _249_/a_373_47# 3.07e-19
C1880 _326_/a_543_47# net28 7.67e-20
C1881 _324_/a_1108_47# net26 1.04e-19
C1882 _002_ clk 5.38e-20
C1883 VPWR trim_val\[4\] 0.311f
C1884 _339_/a_652_21# cal_count\[0\] 0.0264f
C1885 _320_/a_193_47# _065_ 4.41e-20
C1886 _019_ _247_/a_27_297# 9.77e-21
C1887 VPWR _128_ 0.684f
C1888 _234_/a_109_297# _337_/a_193_47# 9.28e-20
C1889 _307_/a_761_289# net45 0.166f
C1890 _307_/a_1283_21# clknet_2_0__leaf_clk 3.93e-19
C1891 net47 _069_ 3.22e-19
C1892 _058_ _267_/a_59_75# 0.00906f
C1893 trim[3] _334_/a_543_47# 2.57e-20
C1894 VPWR _324_/a_1462_47# 3.61e-19
C1895 _185_/a_68_297# _185_/a_150_297# 0.00477f
C1896 _249_/a_373_47# net53 0.00204f
C1897 _336_/a_193_47# _266_/a_68_297# 2.02e-21
C1898 _060_ _226_/a_303_47# 0.00137f
C1899 calibrate _107_ 0.0534f
C1900 _322_/a_1283_21# net26 0.00125f
C1901 _251_/a_27_297# _046_ 5.07e-19
C1902 net27 _222_/a_113_297# 2.1e-19
C1903 _002_ net4 7.04e-21
C1904 _259_/a_27_297# clknet_2_2__leaf_clk 5.1e-19
C1905 state\[0\] net3 0.135f
C1906 _065_ net19 0.00893f
C1907 _330_/a_1108_47# _108_ 5.54e-22
C1908 VPWR net31 1.38f
C1909 clknet_2_0__leaf_clk _209_/a_27_47# 3.24e-21
C1910 ctln[2] net34 0.00136f
C1911 net17 _042_ 0.029f
C1912 net9 trim_mask\[0\] 0.0947f
C1913 _104_ _328_/a_27_47# 0.0099f
C1914 _304_/a_193_47# _122_ 0.00922f
C1915 VPWR _322_/a_1217_47# 7.57e-20
C1916 _053_ _330_/a_193_47# 1.33e-19
C1917 _083_ _311_/a_805_47# 1.62e-20
C1918 _336_/a_543_47# _063_ 2.94e-21
C1919 _274_/a_75_212# net33 7.24e-21
C1920 _267_/a_59_75# _332_/a_27_47# 0.00126f
C1921 _269_/a_299_297# _333_/a_761_289# 2.18e-19
C1922 _274_/a_75_212# trim_mask\[1\] 1.93e-19
C1923 _105_ net19 0.0167f
C1924 _182_/a_27_47# _058_ 0.196f
C1925 fanout47/a_27_47# clknet_0_clk 3.52e-21
C1926 net13 _318_/a_805_47# 5.87e-19
C1927 _316_/a_27_47# _013_ 0.218f
C1928 _195_/a_439_47# _062_ 0.00422f
C1929 _237_/a_505_21# _093_ 4.38e-19
C1930 VPWR _000_ 0.473f
C1931 _030_ trim_val\[0\] 0.00101f
C1932 _323_/a_761_289# _042_ 0.0184f
C1933 _071_ _062_ 2.92e-19
C1934 _192_/a_174_21# _095_ 0.0458f
C1935 trim_val\[3\] _032_ 2.72e-19
C1936 VPWR _281_/a_253_297# 0.00217f
C1937 clknet_2_1__leaf_clk _312_/a_1108_47# 1.32e-19
C1938 _309_/a_27_47# _074_ 0.0189f
C1939 cal_count\[1\] trimb[4] 5.25e-20
C1940 _087_ _096_ 3.13e-20
C1941 _089_ _100_ 0.243f
C1942 _308_/a_639_47# clknet_2_0__leaf_clk 1.44e-19
C1943 _326_/a_651_413# net43 0.0139f
C1944 _104_ _266_/a_68_297# 0.00161f
C1945 _007_ _310_/a_761_289# 0.00229f
C1946 _122_ _298_/a_493_297# 0.0108f
C1947 net42 _087_ 2.68e-20
C1948 _323_/a_448_47# clknet_2_1__leaf_clk 1.99e-19
C1949 _094_ _034_ 0.0183f
C1950 net13 calibrate 0.00629f
C1951 _000_ net53 0.00139f
C1952 clk _106_ 1.91e-20
C1953 _074_ _155_/a_150_297# 5.4e-19
C1954 _002_ net52 2.54e-20
C1955 _237_/a_218_374# net45 8.89e-20
C1956 _237_/a_535_374# _014_ 1.51e-20
C1957 net31 _161_/a_68_297# 4.7e-19
C1958 mask\[6\] _101_ 0.509f
C1959 net10 _275_/a_299_297# 4.27e-19
C1960 _058_ net37 3.24e-19
C1961 _181_/a_150_297# _108_ 5.77e-19
C1962 mask\[0\] _245_/a_109_297# 0.00641f
C1963 _078_ _245_/a_27_297# 6.43e-20
C1964 fanout43/a_27_47# _212_/a_113_297# 7.26e-19
C1965 _266_/a_68_297# net55 5.3e-21
C1966 _334_/a_1283_21# net46 0.278f
C1967 _143_/a_150_297# _078_ 0.00132f
C1968 _107_ _105_ 0.00862f
C1969 net25 _310_/a_543_47# 8.59e-19
C1970 _082_ _310_/a_27_47# 1.67e-19
C1971 trim_mask\[1\] clknet_2_2__leaf_clk 0.374f
C1972 _315_/a_1108_47# _241_/a_105_352# 5.06e-20
C1973 net9 _338_/a_652_21# 5.31e-20
C1974 _300_/a_47_47# cal_count\[2\] 8.29e-19
C1975 _327_/a_761_289# net46 0.17f
C1976 cal_itt\[0\] _195_/a_535_374# 0.00591f
C1977 cal_itt\[1\] _195_/a_218_374# 9.79e-19
C1978 _336_/a_193_47# _028_ 6.93e-20
C1979 _336_/a_761_289# clknet_2_2__leaf_clk 0.00214f
C1980 _328_/a_805_47# trim_mask\[1\] 4.53e-21
C1981 _102_ _022_ 1.9e-20
C1982 cal_itt\[0\] cal_itt\[1\] 0.944f
C1983 net13 net45 0.226f
C1984 net51 _076_ 0.092f
C1985 result[1] _308_/a_761_289# 0.00102f
C1986 _122_ net18 0.155f
C1987 _319_/a_1270_413# _016_ 1.55e-20
C1988 _304_/a_761_289# _304_/a_543_47# 0.21f
C1989 _304_/a_193_47# _304_/a_1283_21# 0.0424f
C1990 _304_/a_27_47# _304_/a_1108_47# 0.102f
C1991 _190_/a_27_47# cal_itt\[3\] 0.169f
C1992 _306_/a_27_47# rebuffer5/a_161_47# 0.0041f
C1993 _329_/a_1108_47# _328_/a_1283_21# 1.18e-19
C1994 _329_/a_1283_21# _328_/a_1108_47# 5.34e-20
C1995 output32/a_27_47# _162_/a_27_47# 4.49e-19
C1996 _334_/a_1108_47# _334_/a_1270_413# 0.00645f
C1997 _334_/a_761_289# _334_/a_1217_47# 4.2e-19
C1998 _334_/a_543_47# _334_/a_805_47# 0.00171f
C1999 _329_/a_1283_21# trim_mask\[2\] 0.0687f
C2000 net4 _106_ 0.0182f
C2001 _110_ _270_/a_59_75# 0.132f
C2002 _122_ _129_ 0.00432f
C2003 _263_/a_297_47# _096_ 1.97e-20
C2004 _263_/a_382_297# net55 0.00139f
C2005 _088_ _052_ 0.133f
C2006 _327_/a_1283_21# _327_/a_1108_47# 0.234f
C2007 _327_/a_761_289# _327_/a_651_413# 0.0977f
C2008 _327_/a_27_47# _327_/a_639_47# 0.00188f
C2009 _327_/a_193_47# _327_/a_1270_413# 1.46e-19
C2010 _327_/a_543_47# _327_/a_448_47# 0.0498f
C2011 _335_/a_543_47# _027_ 5.87e-19
C2012 _164_/a_161_47# _317_/a_1283_21# 7.1e-20
C2013 _335_/a_761_289# net46 0.189f
C2014 _074_ _248_/a_109_47# 4.39e-19
C2015 net12 _078_ 0.111f
C2016 _322_/a_761_289# _074_ 0.0107f
C2017 VPWR _156_/a_27_47# 0.277f
C2018 net13 _065_ 0.058f
C2019 _169_/a_109_53# net54 3.91e-19
C2020 _169_/a_215_311# _060_ 5.66e-19
C2021 output21/a_27_47# _074_ 0.0289f
C2022 _299_/a_27_413# _129_ 0.0652f
C2023 _136_ _284_/a_68_297# 0.00218f
C2024 VPWR en 0.243f
C2025 net2 _040_ 1.61e-21
C2026 _081_ mask\[0\] 1.69e-19
C2027 _327_/a_1270_413# _058_ 1.09e-19
C2028 _078_ _159_/a_27_47# 0.0319f
C2029 _322_/a_193_47# net45 5.96e-21
C2030 VPWR _330_/a_193_47# 0.589f
C2031 _104_ _028_ 4.91e-20
C2032 _332_/a_193_47# net46 0.595f
C2033 _292_/a_78_199# net2 0.0528f
C2034 _328_/a_1283_21# net9 0.0067f
C2035 trimb[0] net38 0.00705f
C2036 _194_/a_113_297# _107_ 5.69e-20
C2037 en valid 0.00147f
C2038 _341_/a_193_47# _067_ 2.28e-20
C2039 _164_/a_161_47# _192_/a_174_21# 1.47e-20
C2040 _083_ net26 0.256f
C2041 _336_/a_1283_21# _107_ 3.14e-19
C2042 _106_ _063_ 0.0377f
C2043 mask\[6\] _312_/a_448_47# 2.83e-21
C2044 net13 _319_/a_27_47# 1.88e-21
C2045 trim_mask\[1\] _333_/a_651_413# 0.00123f
C2046 trim_val\[1\] _333_/a_1270_413# 1.87e-19
C2047 _021_ _312_/a_543_47# 2.75e-20
C2048 _340_/a_1182_261# _122_ 0.00579f
C2049 _325_/a_27_47# net15 8.47e-19
C2050 _078_ net44 0.0366f
C2051 net15 en_co_clk 0.00947f
C2052 _235_/a_79_21# en_co_clk 0.00618f
C2053 trim_val\[0\] net33 0.0273f
C2054 _298_/a_78_199# _133_ 0.243f
C2055 _310_/a_27_47# _310_/a_448_47# 0.0931f
C2056 _310_/a_193_47# _310_/a_1108_47# 0.117f
C2057 net13 _243_/a_109_297# 0.00326f
C2058 _156_/a_27_47# _009_ 1.44e-19
C2059 _307_/a_27_47# _210_/a_113_297# 7.96e-20
C2060 _327_/a_1108_47# _108_ 1.55e-19
C2061 VPWR _325_/a_761_289# 0.207f
C2062 _341_/a_1283_21# net16 2.94e-20
C2063 _239_/a_27_297# _107_ 0.00349f
C2064 _159_/a_27_47# _313_/a_651_413# 8.84e-19
C2065 net21 _313_/a_193_47# 8.73e-19
C2066 _046_ _313_/a_543_47# 2.94e-19
C2067 net43 net45 0.392f
C2068 _335_/a_193_47# _335_/a_1270_413# 1.46e-19
C2069 _335_/a_27_47# _335_/a_639_47# 4.78e-19
C2070 _335_/a_543_47# _335_/a_448_47# 0.0498f
C2071 _335_/a_761_289# _335_/a_651_413# 0.0977f
C2072 _335_/a_1283_21# _335_/a_1108_47# 0.234f
C2073 net16 _333_/a_27_47# 0.0152f
C2074 _324_/a_27_47# clknet_2_1__leaf_clk 0.248f
C2075 mask\[3\] net51 4.53e-21
C2076 net47 fanout47/a_27_47# 0.19f
C2077 net26 _208_/a_218_374# 6.87e-20
C2078 result[4] _310_/a_761_289# 2.56e-19
C2079 _313_/a_1283_21# _312_/a_193_47# 9.64e-21
C2080 _313_/a_1108_47# _312_/a_27_47# 1.26e-20
C2081 _058_ _332_/a_651_413# 9.61e-19
C2082 net35 _332_/a_1108_47# 0.00429f
C2083 mask\[0\] _016_ 0.0328f
C2084 net13 _232_/a_304_297# 9e-19
C2085 VPWR _077_ 0.279f
C2086 net24 _101_ 0.00937f
C2087 _053_ _058_ 0.00145f
C2088 net9 _341_/a_1108_47# 0.00738f
C2089 net43 _065_ 0.0751f
C2090 _303_/a_193_47# _042_ 2.78e-21
C2091 _050_ net15 3.54e-20
C2092 _235_/a_79_21# _050_ 2.2e-19
C2093 _304_/a_1283_21# _304_/a_1462_47# 0.0074f
C2094 _304_/a_1108_47# _304_/a_1217_47# 0.00742f
C2095 clkbuf_2_0__f_clk/a_110_47# _092_ 0.0808f
C2096 _339_/a_1140_413# _123_ 0.00177f
C2097 net43 _305_/a_651_413# 0.0135f
C2098 _256_/a_109_297# net18 0.00587f
C2099 _336_/a_543_47# _279_/a_396_47# 0.00228f
C2100 _336_/a_1283_21# _279_/a_27_47# 0.00531f
C2101 rebuffer3/a_75_212# _118_ 1.4e-20
C2102 clk _316_/a_1108_47# 5.5e-19
C2103 _108_ rebuffer2/a_75_212# 0.196f
C2104 _308_/a_27_47# net22 1.73e-19
C2105 output25/a_27_47# clknet_2_1__leaf_clk 0.0196f
C2106 _321_/a_761_289# _321_/a_543_47# 0.21f
C2107 _321_/a_193_47# _321_/a_1283_21# 0.0424f
C2108 _321_/a_27_47# _321_/a_1108_47# 0.102f
C2109 _332_/a_27_47# _332_/a_651_413# 9.73e-19
C2110 _332_/a_761_289# _332_/a_1108_47# 0.0512f
C2111 _332_/a_193_47# _332_/a_448_47# 0.0564f
C2112 output14/a_27_47# _314_/a_761_289# 0.00321f
C2113 _292_/a_78_199# _123_ 0.0968f
C2114 en_co_clk _049_ 0.459f
C2115 _168_/a_207_413# _028_ 0.00369f
C2116 net43 _319_/a_27_47# 0.298f
C2117 _042_ _152_/a_68_297# 1.02e-20
C2118 _320_/a_543_47# _078_ 7.94e-20
C2119 _337_/a_761_289# _337_/a_543_47# 0.21f
C2120 _337_/a_193_47# _337_/a_1283_21# 0.0418f
C2121 _337_/a_27_47# _337_/a_1108_47# 0.102f
C2122 _304_/a_543_47# cal_count\[3\] 3.03e-21
C2123 _232_/a_32_297# _095_ 4.99e-19
C2124 clkbuf_2_2__f_clk/a_110_47# _331_/a_27_47# 3.93e-19
C2125 _216_/a_199_47# _018_ 3.21e-20
C2126 _333_/a_543_47# net32 1.22e-19
C2127 net24 _320_/a_27_47# 1.18e-19
C2128 _340_/a_1602_47# _298_/a_215_47# 3.17e-21
C2129 net4 _316_/a_1108_47# 0.00387f
C2130 net9 _339_/a_476_47# 0.0108f
C2131 _126_ _339_/a_27_47# 1.75e-20
C2132 _319_/a_1283_21# _283_/a_75_212# 8.51e-19
C2133 net9 trim_mask\[4\] 2.61e-20
C2134 _257_/a_373_47# trim_mask\[1\] 0.00366f
C2135 _340_/a_27_47# clknet_2_3__leaf_clk 0.24f
C2136 _256_/a_109_297# _302_/a_27_297# 4.61e-21
C2137 _250_/a_27_297# _249_/a_109_297# 1.58e-19
C2138 _302_/a_373_47# net18 5.13e-19
C2139 VPWR _330_/a_1462_47# 0.00178f
C2140 _090_ clone7/a_27_47# 6.18e-19
C2141 _257_/a_27_297# _336_/a_1108_47# 3.7e-19
C2142 _332_/a_1462_47# net46 0.00196f
C2143 _036_ net2 0.152f
C2144 net47 _287_/a_75_212# 0.0126f
C2145 clkbuf_2_1__f_clk/a_110_47# _246_/a_27_297# 0.0105f
C2146 _105_ _118_ 0.00226f
C2147 _048_ _192_/a_639_47# 0.00353f
C2148 _291_/a_117_297# cal_count\[0\] 0.00146f
C2149 _015_ _316_/a_27_47# 3.05e-21
C2150 _340_/a_1296_47# _122_ 6.42e-19
C2151 _104_ _279_/a_314_297# 6.76e-19
C2152 net3 _192_/a_476_47# 9.36e-19
C2153 net25 net15 4.23e-21
C2154 _324_/a_193_47# mask\[6\] 6.26e-20
C2155 net33 _131_ 0.00541f
C2156 _306_/a_543_47# rebuffer4/a_27_47# 1.06e-19
C2157 VPWR _334_/a_543_47# 0.226f
C2158 _255_/a_27_47# clknet_2_2__leaf_clk 4.21e-20
C2159 _103_ _260_/a_93_21# 1.08e-20
C2160 _314_/a_1283_21# net29 0.0966f
C2161 _048_ _262_/a_109_297# 0.0145f
C2162 _307_/a_448_47# net22 1.88e-19
C2163 VPWR _327_/a_193_47# 0.555f
C2164 _307_/a_1108_47# mask\[0\] 8.21e-19
C2165 _307_/a_1283_21# _078_ 0.0109f
C2166 _059_ _088_ 7.29e-21
C2167 _050_ _049_ 0.4f
C2168 trim[4] net35 0.0161f
C2169 net21 _313_/a_1462_47# 1.36e-19
C2170 _335_/a_543_47# _032_ 0.00164f
C2171 _302_/a_27_297# _302_/a_373_47# 0.0134f
C2172 _299_/a_27_413# _297_/a_47_47# 3.62e-19
C2173 _250_/a_27_297# mask\[4\] 2.19e-19
C2174 output35/a_27_47# comp 3.98e-20
C2175 _311_/a_193_47# _311_/a_639_47# 2.28e-19
C2176 _311_/a_761_289# _311_/a_1270_413# 2.6e-19
C2177 _311_/a_543_47# _311_/a_651_413# 0.0572f
C2178 output27/a_27_47# result[5] 0.158f
C2179 net27 _311_/a_1283_21# 2.42e-19
C2180 _270_/a_59_75# clknet_2_2__leaf_clk 0.0016f
C2181 _322_/a_448_47# _042_ 2.87e-20
C2182 _256_/a_27_297# cal_count\[3\] 3.52e-20
C2183 _078_ _209_/a_27_47# 0.223f
C2184 VPWR _058_ 1.27f
C2185 _304_/a_651_413# _136_ 3.08e-19
C2186 _304_/a_543_47# _038_ 2.52e-20
C2187 _064_ _092_ 0.00523f
C2188 VPWR _335_/a_193_47# 0.627f
C2189 clknet_2_0__leaf_clk mask\[2\] 8.35e-19
C2190 trim[4] _332_/a_761_289# 1.68e-19
C2191 _305_/a_27_47# rebuffer5/a_161_47# 5.84e-21
C2192 _304_/a_639_47# net47 9.54e-19
C2193 _326_/a_543_47# _314_/a_543_47# 0.00139f
C2194 _326_/a_1108_47# _314_/a_193_47# 5.19e-20
C2195 _326_/a_193_47# _314_/a_1108_47# 3.21e-21
C2196 _096_ _099_ 0.28f
C2197 _100_ _092_ 9.61e-20
C2198 _194_/a_113_297# _118_ 3.83e-19
C2199 net55 _095_ 0.0478f
C2200 cal_count\[1\] net33 0.0109f
C2201 trim_mask\[0\] _091_ 7.39e-20
C2202 _258_/a_27_297# net18 0.00591f
C2203 _024_ net18 0.029f
C2204 _340_/a_193_47# net47 0.203f
C2205 _256_/a_109_297# trim_mask\[0\] 0.0828f
C2206 _336_/a_1283_21# _118_ 1.64e-20
C2207 _336_/a_1108_47# trim_val\[4\] 0.00135f
C2208 _147_/a_27_47# net18 0.00164f
C2209 VPWR _314_/a_639_47# 4.68e-19
C2210 _097_ _241_/a_105_352# 8.1e-19
C2211 calibrate net3 0.00995f
C2212 _106_ _279_/a_396_47# 0.00425f
C2213 clknet_0_clk _119_ 0.0394f
C2214 VPWR _332_/a_27_47# 0.484f
C2215 _094_ _075_ 1.22e-19
C2216 _321_/a_1283_21# _321_/a_1462_47# 0.0074f
C2217 _321_/a_1108_47# _321_/a_1217_47# 0.00742f
C2218 _340_/a_652_21# _340_/a_956_413# 3.11e-19
C2219 _340_/a_1032_413# _340_/a_1602_47# 0.111f
C2220 _340_/a_476_47# _340_/a_562_413# 0.00972f
C2221 output8/a_27_47# _175_/a_68_297# 8.9e-21
C2222 _228_/a_79_21# _054_ 1.26e-20
C2223 _228_/a_297_47# _049_ 0.0486f
C2224 _052_ _170_/a_299_297# 0.0718f
C2225 _308_/a_448_47# net24 9.84e-21
C2226 VPWR _060_ 0.535f
C2227 net28 result[7] 0.11f
C2228 _036_ _123_ 0.012f
C2229 _253_/a_81_21# _253_/a_299_297# 0.0821f
C2230 _008_ _042_ 6.43e-21
C2231 net43 _319_/a_1217_47# 4.13e-19
C2232 _087_ _098_ 0.105f
C2233 _309_/a_193_47# _078_ 0.0278f
C2234 net3 net45 0.264f
C2235 _107_ _278_/a_27_47# 9.64e-19
C2236 _292_/a_215_47# net16 0.00111f
C2237 _259_/a_109_297# trim_val\[3\] 1.23e-20
C2238 _259_/a_27_297# trim_mask\[3\] 0.172f
C2239 _326_/a_761_289# _310_/a_27_47# 3.13e-20
C2240 _326_/a_193_47# _310_/a_193_47# 3.85e-21
C2241 _341_/a_1283_21# net40 1.69e-20
C2242 _337_/a_1283_21# _337_/a_1462_47# 0.0074f
C2243 _337_/a_1108_47# _337_/a_1217_47# 0.00742f
C2244 _080_ net45 0.00397f
C2245 trim[0] net49 1.66e-19
C2246 output26/a_27_47# net26 0.18f
C2247 VPWR _310_/a_1108_47# 0.286f
C2248 _037_ _298_/a_78_199# 0.106f
C2249 _051_ _337_/a_1108_47# 1.6e-19
C2250 ctln[4] net46 1.77e-19
C2251 output36/a_27_47# output38/a_27_47# 0.00249f
C2252 _325_/a_1283_21# _074_ 0.00417f
C2253 trim_mask\[2\] clkbuf_2_2__f_clk/a_110_47# 1.07e-19
C2254 _250_/a_373_47# mask\[5\] 2.82e-19
C2255 _021_ _249_/a_27_297# 7.91e-20
C2256 _175_/a_68_297# _055_ 3.39e-19
C2257 _025_ _336_/a_1283_21# 6.6e-21
C2258 _333_/a_193_47# _055_ 1.23e-19
C2259 _167_/a_161_47# _051_ 0.311f
C2260 _042_ mask\[5\] 0.00943f
C2261 _035_ _338_/a_476_47# 0.0103f
C2262 _329_/a_193_47# _025_ 9.52e-21
C2263 net27 _224_/a_199_47# 6.1e-21
C2264 output27/a_27_47# net29 5.41e-20
C2265 _341_/a_1108_47# _122_ 9.16e-20
C2266 _091_ _191_/a_27_297# 1.14e-19
C2267 _270_/a_59_75# trim_val\[0\] 1.89e-21
C2268 _110_ _117_ 0.0389f
C2269 _161_/a_68_297# _332_/a_27_47# 5.68e-21
C2270 _306_/a_27_47# net51 0.00529f
C2271 net3 _065_ 0.0566f
C2272 _321_/a_193_47# _101_ 0.493f
C2273 _338_/a_1032_413# net18 0.00919f
C2274 _324_/a_639_47# _021_ 1.9e-19
C2275 state\[1\] en_co_clk 6.36e-19
C2276 _110_ _136_ 5.58e-19
C2277 VPWR _327_/a_1462_47# 2.34e-19
C2278 clkbuf_0_clk/a_110_47# _198_/a_27_47# 0.0095f
C2279 _263_/a_297_47# _098_ 1.51e-19
C2280 net15 _039_ 8.96e-21
C2281 _313_/a_193_47# _045_ 1.48e-20
C2282 _129_ _297_/a_285_47# 0.0619f
C2283 _307_/a_1283_21# _004_ 1.29e-20
C2284 trimb[1] net34 0.0785f
C2285 _321_/a_27_47# _214_/a_113_297# 8.73e-21
C2286 trim_mask\[3\] trim_mask\[1\] 1.44e-19
C2287 _057_ _056_ 8.97e-20
C2288 net28 _313_/a_1108_47# 0.044f
C2289 _311_/a_27_47# net26 0.0437f
C2290 _322_/a_543_47# _078_ 7.59e-21
C2291 _259_/a_27_297# _330_/a_1283_21# 0.00828f
C2292 mask\[0\] _095_ 0.00186f
C2293 net50 _336_/a_193_47# 1.03e-20
C2294 _019_ _042_ 7.08e-19
C2295 _074_ _314_/a_27_47# 0.00141f
C2296 _164_/a_161_47# net55 8.54e-19
C2297 net47 _136_ 0.00242f
C2298 _329_/a_27_47# trim_val\[3\] 8.78e-20
C2299 VPWR _335_/a_1462_47# 7.25e-20
C2300 _102_ net14 1.21e-20
C2301 _331_/a_27_47# _331_/a_193_47# 0.725f
C2302 _053_ _227_/a_109_93# 8.89e-20
C2303 VPWR _311_/a_651_413# 0.133f
C2304 _245_/a_27_297# _245_/a_109_47# 0.00393f
C2305 calibrate _062_ 3.45e-19
C2306 _110_ _119_ 0.00786f
C2307 mask\[1\] clknet_2_0__leaf_clk 7.16e-19
C2308 _050_ state\[1\] 4.82e-20
C2309 _258_/a_27_297# trim_mask\[0\] 6.41e-20
C2310 trim_mask\[2\] _256_/a_27_297# 5.93e-21
C2311 _340_/a_796_47# net47 0.00187f
C2312 trim_mask\[0\] _024_ 0.123f
C2313 _323_/a_27_47# clknet_2_3__leaf_clk 1.16e-20
C2314 _340_/a_1032_413# _041_ 9.24e-22
C2315 _266_/a_68_297# clknet_2_3__leaf_clk 3.57e-20
C2316 _325_/a_193_47# clknet_2_1__leaf_clk 0.00758f
C2317 _311_/a_651_413# net53 0.00167f
C2318 net23 mask\[0\] 0.241f
C2319 VPWR _332_/a_1217_47# 1.35e-19
C2320 clknet_2_1__leaf_clk _120_ 8.85e-21
C2321 _340_/a_652_21# _037_ 7.99e-19
C2322 _319_/a_761_289# _120_ 2.43e-20
C2323 _005_ net24 0.00456f
C2324 net23 output24/a_27_47# 0.0138f
C2325 _062_ rebuffer3/a_75_212# 9.39e-20
C2326 _051_ _331_/a_543_47# 0.00194f
C2327 _327_/a_761_289# _111_ 2.55e-19
C2328 fanout44/a_27_47# net45 0.165f
C2329 cal_count\[0\] net37 2.9e-19
C2330 _134_ _298_/a_493_297# 8.56e-20
C2331 _006_ net14 0.0111f
C2332 _309_/a_1462_47# _078_ 0.00213f
C2333 _110_ _328_/a_193_47# 4.66e-20
C2334 _104_ net50 0.363f
C2335 _323_/a_448_47# _043_ 7.3e-22
C2336 clkbuf_0_clk/a_110_47# _041_ 6.5e-21
C2337 net9 _178_/a_68_297# 2.97e-19
C2338 _051_ _229_/a_27_297# 6.43e-21
C2339 _337_/a_639_47# net44 1.79e-19
C2340 _053_ _286_/a_76_199# 1.01e-19
C2341 _039_ _049_ 1.46e-19
C2342 _341_/a_193_47# clknet_2_3__leaf_clk 0.526f
C2343 _233_/a_109_47# cal 1.54e-19
C2344 _233_/a_109_297# net1 0.00511f
C2345 clknet_2_1__leaf_clk _076_ 0.0855f
C2346 net43 _282_/a_68_297# 6.96e-20
C2347 _236_/a_109_297# _096_ 0.0114f
C2348 _058_ _029_ 0.00671f
C2349 _239_/a_474_297# _048_ 0.0991f
C2350 net43 _313_/a_639_47# 2.48e-19
C2351 _065_ _062_ 1.86e-19
C2352 _015_ _167_/a_161_47# 0.0131f
C2353 _291_/a_117_297# net16 7.79e-19
C2354 fanout44/a_27_47# _065_ 0.024f
C2355 VPWR _306_/a_193_47# 0.602f
C2356 _146_/a_68_297# mask\[1\] 1.08e-21
C2357 _269_/a_299_297# _334_/a_193_47# 2.19e-21
C2358 _061_ net37 0.00617f
C2359 mask\[6\] _156_/a_27_47# 7.31e-22
C2360 _110_ _266_/a_150_297# 4.96e-19
C2361 _187_/a_27_413# _332_/a_1108_47# 0.00112f
C2362 _187_/a_212_413# _332_/a_1283_21# 4.47e-19
C2363 _105_ _062_ 2.74e-19
C2364 _326_/a_193_47# _224_/a_113_297# 4.52e-20
C2365 _134_ _129_ 0.0297f
C2366 _149_/a_68_297# _303_/a_761_289# 5.23e-19
C2367 _306_/a_651_413# rebuffer6/a_27_47# 6.28e-21
C2368 _294_/a_68_297# _299_/a_27_413# 0.00519f
C2369 net12 ctln[6] 0.02f
C2370 _029_ _332_/a_27_47# 0.285f
C2371 _195_/a_76_199# _065_ 8.83e-20
C2372 _053_ _054_ 0.339f
C2373 _316_/a_543_47# _095_ 4.5e-19
C2374 net45 _137_/a_68_297# 0.00161f
C2375 VPWR ctlp[3] 0.283f
C2376 _040_ _121_ 2.96e-20
C2377 clk _331_/a_1270_413# 5.04e-20
C2378 fanout44/a_27_47# _319_/a_27_47# 6.12e-21
C2379 _254_/a_109_297# _050_ 1.84e-20
C2380 _053_ net30 0.173f
C2381 _323_/a_193_47# net47 0.0258f
C2382 _170_/a_81_21# net41 1.75e-22
C2383 _001_ _069_ 0.216f
C2384 _314_/a_448_47# _011_ 0.16f
C2385 output7/a_27_47# net6 3.17e-21
C2386 ctln[6] _331_/a_1108_47# 3.54e-20
C2387 net55 _226_/a_27_47# 5.75e-19
C2388 cal_itt\[1\] net2 5.03e-19
C2389 _136_ _301_/a_47_47# 0.144f
C2390 _104_ _330_/a_1108_47# 5.9e-20
C2391 _306_/a_1283_21# _306_/a_1108_47# 0.234f
C2392 _306_/a_761_289# _306_/a_651_413# 0.0977f
C2393 _306_/a_543_47# _306_/a_448_47# 0.0498f
C2394 _306_/a_27_47# _306_/a_639_47# 0.00188f
C2395 _306_/a_193_47# _306_/a_1270_413# 1.46e-19
C2396 cal_itt\[0\] _305_/a_1108_47# 7.11e-20
C2397 VPWR _227_/a_109_93# 0.165f
C2398 _118_ _278_/a_27_47# 0.068f
C2399 _329_/a_805_47# trim_mask\[3\] 4.63e-20
C2400 _341_/a_27_47# _136_ 0.0151f
C2401 net12 _087_ 0.00185f
C2402 _331_/a_543_47# _331_/a_639_47# 0.0138f
C2403 _331_/a_193_47# _331_/a_1217_47# 2.36e-20
C2404 _331_/a_761_289# _331_/a_805_47# 3.69e-19
C2405 _331_/a_27_47# _260_/a_93_21# 4.97e-21
C2406 _060_ _093_ 0.00231f
C2407 _325_/a_761_289# mask\[6\] 0.0219f
C2408 _007_ clknet_2_1__leaf_clk 0.233f
C2409 _245_/a_109_297# _016_ 0.00452f
C2410 _245_/a_373_47# net52 0.00236f
C2411 VPWR output20/a_27_47# 0.41f
C2412 _256_/a_109_297# trim_mask\[4\] 0.00264f
C2413 VPWR _235_/a_297_47# 0.00571f
C2414 VPWR net7 0.521f
C2415 net12 _312_/a_27_47# 1.3e-19
C2416 _041_ _338_/a_476_47# 3.12e-19
C2417 _308_/a_193_47# net14 0.0121f
C2418 _189_/a_408_47# _088_ 6.59e-20
C2419 _338_/a_27_47# _338_/a_381_47# 0.0685f
C2420 _338_/a_193_47# _338_/a_1602_47# 4.3e-19
C2421 _338_/a_652_21# _338_/a_1032_413# 0.00971f
C2422 VPWR _317_/a_193_47# 0.273f
C2423 _113_ rebuffer2/a_75_212# 3.36e-21
C2424 VPWR _326_/a_193_47# 0.589f
C2425 output10/a_27_47# ctln[4] 0.159f
C2426 net13 _321_/a_27_47# 4.31e-21
C2427 _030_ _108_ 1.99e-20
C2428 _121_ _095_ 7.97e-19
C2429 cal _315_/a_448_47# 0.00123f
C2430 _102_ net52 0.17f
C2431 clknet_2_0__leaf_clk _244_/a_27_297# 0.0417f
C2432 mask\[3\] clknet_2_1__leaf_clk 0.737f
C2433 _074_ _310_/a_651_413# 0.00464f
C2434 _194_/a_113_297# _062_ 4.43e-19
C2435 _304_/a_193_47# cal_count\[2\] 1.23e-21
C2436 net13 _337_/a_27_47# 0.0153f
C2437 _336_/a_1283_21# _062_ 3.55e-19
C2438 _170_/a_299_297# _170_/a_384_47# 1.48e-19
C2439 net2 input2/a_27_47# 0.178f
C2440 _297_/a_47_47# _297_/a_285_47# 0.0175f
C2441 _117_ clknet_2_2__leaf_clk 8.95e-22
C2442 _048_ _033_ 3.33e-21
C2443 state\[2\] trim_mask\[0\] 0.00126f
C2444 VPWR _286_/a_76_199# 0.105f
C2445 _325_/a_193_47# _313_/a_27_47# 7.04e-19
C2446 _313_/a_1108_47# _084_ 1.37e-20
C2447 _259_/a_27_297# _335_/a_1283_21# 3.08e-19
C2448 _097_ en_co_clk 0.00288f
C2449 _136_ clknet_2_2__leaf_clk 0.00225f
C2450 net44 _312_/a_27_47# 0.299f
C2451 output35/a_27_47# _132_ 4.05e-20
C2452 _341_/a_651_413# cal_count\[3\] 0.0265f
C2453 _078_ mask\[2\] 0.208f
C2454 _341_/a_1462_47# clknet_2_3__leaf_clk 0.00219f
C2455 _033_ _330_/a_27_47# 6.44e-20
C2456 _012_ net1 0.0346f
C2457 _323_/a_193_47# net44 0.00488f
C2458 _051_ net19 7.23e-20
C2459 _320_/a_448_47# _143_/a_68_297# 9.86e-19
C2460 _117_ net11 1.72e-19
C2461 _298_/a_493_297# cal_count\[2\] 1.79e-19
C2462 net47 _339_/a_27_47# 0.0527f
C2463 _257_/a_27_297# net18 0.00956f
C2464 VPWR _306_/a_1462_47# 1.48e-19
C2465 _305_/a_27_47# net51 0.0281f
C2466 trim_mask\[0\] _134_ 1.05e-19
C2467 _321_/a_193_47# _248_/a_27_297# 1.67e-19
C2468 _053_ _262_/a_465_47# 0.00116f
C2469 _340_/a_1032_413# _339_/a_1032_413# 7.46e-19
C2470 _235_/a_79_21# _049_ 0.00169f
C2471 _327_/a_1283_21# trim_mask\[1\] 5.11e-23
C2472 net15 _049_ 0.0163f
C2473 _030_ _031_ 2.09e-19
C2474 _307_/a_651_413# net14 9.07e-20
C2475 result[7] _085_ 1.61e-21
C2476 _303_/a_1283_21# _035_ 0.00101f
C2477 _336_/a_193_47# _052_ 1.27e-20
C2478 cal_itt\[1\] _123_ 4.01e-20
C2479 _263_/a_79_21# _087_ 0.00945f
C2480 _326_/a_651_413# net29 1.1e-19
C2481 _306_/a_1283_21# _203_/a_59_75# 0.00131f
C2482 _099_ _098_ 0.0998f
C2483 trim_mask\[0\] _333_/a_1283_21# 2.4e-20
C2484 _125_ _132_ 0.00249f
C2485 net39 net38 0.067f
C2486 VPWR _054_ 0.243f
C2487 net27 _086_ 0.193f
C2488 VPWR _318_/a_1283_21# 0.405f
C2489 _029_ _332_/a_1217_47# 2.47e-21
C2490 trim[3] trim_val\[2\] 8.5e-19
C2491 _088_ clone1/a_27_47# 0.00314f
C2492 VPWR net30 4.34f
C2493 _119_ clknet_2_2__leaf_clk 0.358f
C2494 _042_ _310_/a_27_47# 1.81e-20
C2495 _190_/a_465_47# clkbuf_2_3__f_clk/a_110_47# 1.07e-20
C2496 _051_ _107_ 0.156f
C2497 _060_ _243_/a_109_47# 0.00527f
C2498 net12 _320_/a_1108_47# 7.6e-22
C2499 _323_/a_1462_47# net47 0.00223f
C2500 _312_/a_805_47# net20 4.97e-19
C2501 net43 _321_/a_27_47# 0.446f
C2502 trim_mask\[1\] _335_/a_1283_21# 1.15e-20
C2503 _129_ cal_count\[2\] 0.127f
C2504 clknet_0_clk _099_ 2.05e-20
C2505 clknet_2_1__leaf_clk _310_/a_1283_21# 0.0376f
C2506 _064_ net46 0.0173f
C2507 cal_itt\[2\] _002_ 0.0339f
C2508 _336_/a_1108_47# _335_/a_193_47# 3.03e-19
C2509 VPWR _233_/a_373_47# 4.86e-19
C2510 net43 _337_/a_27_47# 5.87e-20
C2511 _341_/a_1217_47# _136_ 1.18e-19
C2512 _103_ _048_ 0.481f
C2513 _301_/a_47_47# _301_/a_129_47# 0.00369f
C2514 _331_/a_761_289# trim_mask\[4\] 5.6e-19
C2515 _331_/a_448_47# _028_ 0.17f
C2516 net15 _317_/a_805_47# 5.85e-19
C2517 _182_/a_27_47# net16 7.97e-19
C2518 net9 _334_/a_27_47# 0.00213f
C2519 _317_/a_193_47# _317_/a_1270_413# 1.46e-19
C2520 _317_/a_27_47# _317_/a_639_47# 0.00188f
C2521 _317_/a_543_47# _317_/a_448_47# 0.0498f
C2522 _317_/a_761_289# _317_/a_651_413# 0.0977f
C2523 _317_/a_1283_21# _317_/a_1108_47# 0.234f
C2524 result[4] clknet_2_1__leaf_clk 0.0505f
C2525 _233_/a_373_47# valid 1.33e-19
C2526 _258_/a_27_297# trim_mask\[4\] 0.0102f
C2527 _326_/a_1283_21# _326_/a_1108_47# 0.234f
C2528 _326_/a_761_289# _326_/a_651_413# 0.0977f
C2529 _326_/a_543_47# _326_/a_448_47# 0.0498f
C2530 _326_/a_27_47# _326_/a_639_47# 0.00188f
C2531 _326_/a_193_47# _326_/a_1270_413# 1.46e-19
C2532 _328_/a_193_47# clknet_2_2__leaf_clk 0.596f
C2533 trim_val\[1\] rebuffer2/a_75_212# 1.75e-20
C2534 net33 _108_ 0.34f
C2535 _024_ trim_mask\[4\] 4.44e-19
C2536 trim_mask\[1\] _108_ 0.0105f
C2537 _112_ _332_/a_193_47# 0.00101f
C2538 _263_/a_79_21# _263_/a_297_47# 0.0326f
C2539 _104_ _052_ 0.434f
C2540 ctln[6] net11 6.71e-19
C2541 VPWR _317_/a_1462_47# 7.03e-20
C2542 _338_/a_1032_413# _338_/a_1056_47# 0.0016f
C2543 _338_/a_381_47# _338_/a_586_47# 3.7e-19
C2544 _324_/a_1108_47# clknet_2_3__leaf_clk 2.62e-19
C2545 _328_/a_27_47# _328_/a_1217_47# 2.56e-19
C2546 _328_/a_761_289# _328_/a_639_47# 3.16e-19
C2547 _341_/a_27_47# _341_/a_761_289# 0.0531f
C2548 VPWR _326_/a_1462_47# 0.00178f
C2549 _336_/a_761_289# _108_ 0.00893f
C2550 _320_/a_1108_47# net44 0.234f
C2551 _288_/a_145_75# net33 6.02e-19
C2552 net47 _303_/a_27_47# 0.304f
C2553 result[7] _314_/a_543_47# 3.7e-20
C2554 net18 trim_val\[4\] 1.73e-21
C2555 _052_ net55 0.0806f
C2556 net16 net37 2.55e-20
C2557 net13 _051_ 0.0111f
C2558 cal_itt\[0\] _069_ 0.257f
C2559 _318_/a_193_47# _318_/a_543_47# 0.217f
C2560 _318_/a_27_47# _318_/a_1283_21# 0.0436f
C2561 VPWR _072_ 1.06f
C2562 _290_/a_207_413# _288_/a_59_75# 1.16e-19
C2563 _340_/a_1182_261# cal_count\[2\] 0.00355f
C2564 VPWR cal_count\[0\] 1.12f
C2565 state\[2\] _090_ 3.14e-19
C2566 output18/a_27_47# ctlp[4] 0.168f
C2567 _128_ _129_ 4.32e-20
C2568 _104_ _335_/a_1108_47# 7.7e-20
C2569 net44 _312_/a_1217_47# 6.03e-19
C2570 _110_ _279_/a_206_47# 0.00264f
C2571 _312_/a_193_47# _312_/a_1270_413# 1.46e-19
C2572 _312_/a_27_47# _312_/a_639_47# 0.00188f
C2573 _312_/a_543_47# _312_/a_448_47# 0.0498f
C2574 _312_/a_761_289# _312_/a_651_413# 0.0977f
C2575 _312_/a_1283_21# _312_/a_1108_47# 0.234f
C2576 _336_/a_805_47# net46 0.0019f
C2577 _264_/a_27_297# net46 4.18e-20
C2578 VPWR _305_/a_193_47# 0.524f
C2579 _320_/a_448_47# net52 5.81e-19
C2580 _306_/a_1283_21# clknet_2_0__leaf_clk 1.09e-20
C2581 clknet_2_1__leaf_clk _311_/a_448_47# 1.68e-20
C2582 net27 clknet_2_1__leaf_clk 0.0557f
C2583 _329_/a_651_413# net46 0.0122f
C2584 _078_ _314_/a_193_47# 0.00266f
C2585 _068_ _202_/a_382_297# 4e-19
C2586 _323_/a_543_47# net19 0.00603f
C2587 cal_itt\[1\] _067_ 0.258f
C2588 _060_ _206_/a_27_93# 0.00643f
C2589 _031_ net33 2.32e-21
C2590 mask\[1\] _078_ 0.975f
C2591 VPWR _262_/a_465_47# 3.05e-19
C2592 _041_ _339_/a_1182_261# 0.0204f
C2593 _065_ rebuffer6/a_27_47# 3.73e-19
C2594 net47 _339_/a_586_47# 1.16e-19
C2595 cal_itt\[1\] _070_ 1.5e-19
C2596 _257_/a_27_297# trim_mask\[0\] 6.95e-19
C2597 _192_/a_174_21# _192_/a_27_47# 0.267f
C2598 trim_mask\[1\] _031_ 2.04e-20
C2599 _309_/a_27_47# _102_ 4.1e-21
C2600 trim_val\[2\] _334_/a_805_47# 9.25e-20
C2601 _323_/a_27_47# _323_/a_1217_47# 2.56e-19
C2602 _323_/a_761_289# _323_/a_639_47# 3.16e-19
C2603 _037_ _339_/a_193_47# 2.07e-20
C2604 cal_itt\[2\] _106_ 1.12e-20
C2605 net31 _129_ 1.41e-20
C2606 VPWR _061_ 0.248f
C2607 state\[2\] _242_/a_382_297# 2.81e-19
C2608 output22/a_27_47# _307_/a_27_47# 0.0112f
C2609 output34/a_27_47# _179_/a_27_47# 4.2e-19
C2610 VPWR _315_/a_651_413# 0.138f
C2611 _306_/a_639_47# cal_itt\[3\] 2.69e-19
C2612 _337_/a_448_47# _092_ 0.00126f
C2613 _233_/a_27_297# _233_/a_109_47# 0.00393f
C2614 trim_mask\[2\] _333_/a_543_47# 2.97e-20
C2615 calibrate _227_/a_209_311# 2.51e-19
C2616 _289_/a_68_297# _288_/a_59_75# 0.00852f
C2617 _292_/a_292_297# net47 4.05e-19
C2618 _306_/a_761_289# _065_ 1.3e-21
C2619 clkbuf_0_clk/a_110_47# _190_/a_465_47# 0.00282f
C2620 _315_/a_651_413# valid 7.82e-19
C2621 _036_ _340_/a_27_47# 0.00113f
C2622 _128_ _340_/a_1182_261# 3.45e-20
C2623 _326_/a_27_47# _086_ 2.59e-20
C2624 net36 _126_ 6.86e-20
C2625 _303_/a_27_47# net44 0.00597f
C2626 _093_ _317_/a_193_47# 3.73e-21
C2627 ctln[3] net46 4.12e-20
C2628 net43 _321_/a_1217_47# 0.00134f
C2629 _326_/a_543_47# _074_ 0.0147f
C2630 output33/a_27_47# _108_ 6.33e-19
C2631 net2 trimb[4] 1.08e-19
C2632 _320_/a_543_47# _320_/a_1108_47# 7.99e-20
C2633 _320_/a_193_47# _320_/a_651_413# 0.0276f
C2634 _119_ _279_/a_204_297# 3.48e-19
C2635 ctln[6] ctln[7] 0.00465f
C2636 _309_/a_27_47# _006_ 0.169f
C2637 _309_/a_761_289# _081_ 1.59e-19
C2638 _033_ _335_/a_27_47# 5.24e-22
C2639 _107_ _242_/a_79_21# 0.0112f
C2640 _168_/a_207_413# _052_ 0.0801f
C2641 _036_ _144_/a_27_47# 6.61e-21
C2642 _306_/a_27_47# clknet_2_1__leaf_clk 5.04e-20
C2643 net15 state\[1\] 1.16e-19
C2644 _235_/a_79_21# state\[1\] 1.16e-21
C2645 _237_/a_505_21# _090_ 0.147f
C2646 trim_mask\[4\] _260_/a_250_297# 0.11f
C2647 _061_ _161_/a_68_297# 2.27e-20
C2648 _062_ _278_/a_27_47# 0.0522f
C2649 _187_/a_212_413# _187_/a_297_47# 0.00539f
C2650 _317_/a_1283_21# clknet_2_0__leaf_clk 0.0495f
C2651 _317_/a_543_47# _014_ 0.00234f
C2652 _317_/a_761_289# net45 0.166f
C2653 _036_ clknet_2_3__leaf_clk 0.0321f
C2654 _059_ _232_/a_32_297# 4.28e-19
C2655 _308_/a_193_47# _307_/a_543_47# 1.91e-19
C2656 _328_/a_1462_47# clknet_2_2__leaf_clk 2.16e-19
C2657 net13 _046_ 7.78e-20
C2658 _262_/a_27_47# net30 0.00193f
C2659 _341_/a_543_47# _341_/a_805_47# 0.00171f
C2660 _341_/a_761_289# _341_/a_1217_47# 4.2e-19
C2661 _341_/a_1108_47# _341_/a_1270_413# 0.00645f
C2662 _081_ _040_ 0.165f
C2663 _048_ clkbuf_2_3__f_clk/a_110_47# 0.00413f
C2664 _053_ _066_ 0.0928f
C2665 _303_/a_193_47# _063_ 8.5e-21
C2666 net47 _303_/a_1217_47# 8.66e-19
C2667 net28 _159_/a_27_47# 1.04e-20
C2668 trim_mask\[0\] trim_val\[4\] 0.0422f
C2669 _304_/a_543_47# en_co_clk 2.76e-20
C2670 _315_/a_543_47# net30 4.91e-21
C2671 net4 _279_/a_490_47# 0.00201f
C2672 _333_/a_1283_21# _175_/a_68_297# 1.68e-20
C2673 state\[2\] trim_mask\[4\] 0.168f
C2674 _333_/a_27_47# _333_/a_1108_47# 0.102f
C2675 _333_/a_193_47# _333_/a_1283_21# 0.0424f
C2676 _333_/a_761_289# _333_/a_543_47# 0.21f
C2677 _255_/a_27_47# _088_ 2.94e-20
C2678 net16 _332_/a_651_413# 0.00193f
C2679 net23 _245_/a_109_297# 0.00553f
C2680 clk _092_ 0.034f
C2681 _015_ net13 0.171f
C2682 _267_/a_59_75# net40 2.5e-20
C2683 clknet_2_0__leaf_clk _192_/a_174_21# 8.64e-21
C2684 _318_/a_448_47# _318_/a_639_47# 4.61e-19
C2685 net12 _322_/a_1108_47# 0.00241f
C2686 _297_/a_47_47# cal_count\[2\] 8.68e-19
C2687 _097_ net1 3.15e-20
C2688 net12 _099_ 0.00188f
C2689 _051_ _118_ 2.39e-21
C2690 _265_/a_299_297# _265_/a_384_47# 1.48e-19
C2691 _146_/a_68_297# net26 8.47e-20
C2692 VPWR result[1] 0.361f
C2693 net43 _023_ 0.00545f
C2694 _324_/a_448_47# net44 0.00198f
C2695 _324_/a_27_47# _312_/a_1283_21# 1.2e-19
C2696 _320_/a_1108_47# _209_/a_27_47# 2.12e-19
C2697 VPWR _305_/a_1462_47# 3.12e-19
C2698 net31 trim_mask\[0\] 3.14e-19
C2699 VPWR _250_/a_109_47# 6.5e-19
C2700 VPWR _251_/a_27_297# 0.259f
C2701 _093_ net30 9.79e-21
C2702 _308_/a_1283_21# _308_/a_1108_47# 0.234f
C2703 _308_/a_761_289# _308_/a_651_413# 0.0977f
C2704 _308_/a_543_47# _308_/a_448_47# 0.0498f
C2705 _308_/a_27_47# _308_/a_639_47# 0.00188f
C2706 _308_/a_193_47# _308_/a_1270_413# 1.46e-19
C2707 _041_ _339_/a_1296_47# 0.00205f
C2708 _094_ clkbuf_2_1__f_clk/a_110_47# 2.84e-21
C2709 net2 _203_/a_59_75# 7.02e-22
C2710 _324_/a_1283_21# _323_/a_193_47# 0.00889f
C2711 _324_/a_1108_47# _323_/a_27_47# 2.06e-19
C2712 net3 _337_/a_27_47# 6.19e-19
C2713 net15 _319_/a_543_47# 0.00861f
C2714 _307_/a_543_47# _307_/a_651_413# 0.0572f
C2715 _307_/a_761_289# _307_/a_1270_413# 2.6e-19
C2716 _307_/a_193_47# _307_/a_639_47# 2.28e-19
C2717 net4 _092_ 0.0098f
C2718 _326_/a_27_47# clknet_2_1__leaf_clk 0.371f
C2719 _078_ _244_/a_27_297# 4.42e-20
C2720 _249_/a_27_297# _101_ 0.103f
C2721 result[0] _307_/a_1108_47# 3.43e-19
C2722 _293_/a_81_21# _041_ 0.00233f
C2723 state\[1\] _049_ 6.95e-20
C2724 _309_/a_1108_47# _214_/a_113_297# 6.28e-19
C2725 VPWR _319_/a_1108_47# 0.297f
C2726 _322_/a_1108_47# net44 0.255f
C2727 _318_/a_1108_47# net45 0.242f
C2728 net27 _313_/a_27_47# 3.51e-20
C2729 _309_/a_27_47# _308_/a_193_47# 1.51e-19
C2730 _309_/a_193_47# _308_/a_27_47# 4.17e-21
C2731 _233_/a_373_47# _093_ 0.00193f
C2732 _233_/a_109_297# _012_ 0.0526f
C2733 net3 _013_ 1.05e-19
C2734 _340_/a_193_47# _001_ 5.65e-20
C2735 net50 clknet_2_3__leaf_clk 3.78e-21
C2736 output35/a_27_47# net32 0.00105f
C2737 wire42/a_75_212# net30 1.1e-19
C2738 _059_ net55 0.186f
C2739 _078_ _310_/a_1270_413# 1.98e-19
C2740 net23 _081_ 0.0986f
C2741 clone1/a_27_47# _170_/a_299_297# 4.68e-19
C2742 net43 _046_ 0.0109f
C2743 cal_itt\[0\] fanout47/a_27_47# 0.00255f
C2744 _128_ _297_/a_47_47# 1.51e-21
C2745 _061_ _300_/a_47_47# 2.52e-20
C2746 _096_ net41 1.83e-20
C2747 _303_/a_761_289# net19 0.00894f
C2748 _337_/a_543_47# en_co_clk 0.003f
C2749 _262_/a_27_47# _262_/a_465_47# 0.013f
C2750 net37 net40 0.016f
C2751 _323_/a_1108_47# _303_/a_1108_47# 1.46e-20
C2752 _323_/a_543_47# _303_/a_651_413# 4.92e-20
C2753 _339_/a_652_21# _339_/a_381_47# 7.79e-20
C2754 _339_/a_193_47# _339_/a_562_413# 4.45e-20
C2755 _339_/a_1182_261# _339_/a_1032_413# 0.344f
C2756 _339_/a_27_47# _339_/a_956_413# 0.00159f
C2757 _322_/a_1270_413# _101_ 1.37e-19
C2758 _063_ _092_ 0.367f
C2759 _041_ mask\[4\] 1.8e-20
C2760 net13 _320_/a_651_413# 0.00125f
C2761 _270_/a_59_75# _108_ 1.9e-19
C2762 _263_/a_79_21# _099_ 0.0441f
C2763 _317_/a_805_47# state\[1\] 9.25e-20
C2764 _320_/a_1283_21# _040_ 0.00251f
C2765 VPWR _066_ 0.621f
C2766 VPWR trim_val\[2\] 0.557f
C2767 _113_ _030_ 0.0189f
C2768 _315_/a_193_47# _315_/a_639_47# 2.28e-19
C2769 _315_/a_761_289# _315_/a_1270_413# 2.6e-19
C2770 _315_/a_543_47# _315_/a_651_413# 0.0572f
C2771 _337_/a_761_289# _076_ 1.76e-19
C2772 _048_ cal_count\[3\] 0.0554f
C2773 _104_ _170_/a_384_47# 3.55e-19
C2774 VPWR _336_/a_639_47# 5.1e-19
C2775 net19 _152_/a_150_297# 1.13e-19
C2776 _116_ net50 0.00151f
C2777 _117_ trim_mask\[3\] 6.22e-19
C2778 _101_ _220_/a_113_297# 1.76e-20
C2779 net4 _199_/a_109_297# 7.7e-19
C2780 VPWR _329_/a_448_47# 0.0853f
C2781 net44 _246_/a_27_297# 2.21e-20
C2782 ctln[2] _334_/a_1108_47# 1.72e-20
C2783 net8 _334_/a_651_413# 0.00203f
C2784 _110_ _057_ 0.0685f
C2785 _319_/a_543_47# _049_ 8.73e-19
C2786 _232_/a_32_297# _192_/a_27_47# 8.26e-19
C2787 _323_/a_193_47# _044_ 1.39e-21
C2788 _319_/a_193_47# net30 9.05e-20
C2789 _333_/a_1108_47# _333_/a_1217_47# 0.00742f
C2790 _333_/a_1283_21# _333_/a_1462_47# 0.0074f
C2791 VPWR net16 2.18f
C2792 _312_/a_1108_47# _045_ 9.55e-21
C2793 _340_/a_1602_47# en_co_clk 5.5e-22
C2794 net23 _016_ 0.0433f
C2795 net34 net46 0.00589f
C2796 _050_ _337_/a_543_47# 5.57e-20
C2797 _093_ _315_/a_651_413# 8.82e-19
C2798 _012_ _315_/a_1108_47# 1.26e-19
C2799 calibrate _315_/a_1270_413# 4.47e-19
C2800 _074_ _315_/a_639_47# 0.00164f
C2801 _331_/a_27_47# _330_/a_27_47# 0.0967f
C2802 _326_/a_193_47# mask\[6\] 4.14e-20
C2803 fanout44/a_27_47# _337_/a_27_47# 8.93e-21
C2804 _257_/a_27_297# trim_mask\[4\] 0.0106f
C2805 _324_/a_1270_413# net19 3.32e-20
C2806 _187_/a_212_413# net33 0.0027f
C2807 clkbuf_2_0__f_clk/a_110_47# calibrate 7e-21
C2808 _136_ _001_ 0.00119f
C2809 state\[0\] _316_/a_193_47# 5.34e-19
C2810 _246_/a_109_297# net52 0.0143f
C2811 net12 _084_ 0.00227f
C2812 _308_/a_761_289# net43 0.175f
C2813 _308_/a_543_47# _005_ 0.00362f
C2814 cal_itt\[0\] _287_/a_75_212# 0.00199f
C2815 _328_/a_543_47# _025_ 6.4e-19
C2816 _143_/a_68_297# _017_ 3.47e-19
C2817 _086_ _011_ 0.184f
C2818 net45 _315_/a_1270_413# 1.7e-19
C2819 _305_/a_1270_413# _072_ 5.67e-19
C2820 _198_/a_27_47# en_co_clk 1.18e-19
C2821 _051_ net3 0.0124f
C2822 _094_ _096_ 2.17e-19
C2823 trim_mask\[3\] _119_ 0.0315f
C2824 clkbuf_2_0__f_clk/a_110_47# net45 9.16e-19
C2825 _116_ _330_/a_1108_47# 1.53e-20
C2826 _097_ net15 0.211f
C2827 _327_/a_193_47# net18 0.00863f
C2828 net15 _313_/a_193_47# 1.11e-19
C2829 _305_/a_1108_47# net2 1.43e-20
C2830 net43 _320_/a_651_413# 2.97e-20
C2831 _323_/a_448_47# mask\[4\] 1.8e-19
C2832 _321_/a_543_47# net25 2.89e-20
C2833 _321_/a_761_289# mask\[3\] 5.12e-21
C2834 _305_/a_1283_21# _305_/a_1108_47# 0.234f
C2835 _305_/a_761_289# _305_/a_651_413# 0.0977f
C2836 _305_/a_543_47# _305_/a_448_47# 0.0498f
C2837 _305_/a_27_47# _305_/a_639_47# 3.82e-19
C2838 _305_/a_193_47# _305_/a_1270_413# 1.46e-19
C2839 _309_/a_27_47# _309_/a_1283_21# 0.0436f
C2840 _309_/a_193_47# _309_/a_543_47# 0.217f
C2841 VPWR _313_/a_543_47# 0.227f
C2842 net44 _084_ 1.46e-19
C2843 output32/a_27_47# output35/a_27_47# 0.003f
C2844 net43 _140_/a_68_297# 3.96e-19
C2845 clkbuf_2_0__f_clk/a_110_47# _065_ 0.0331f
C2846 _058_ net18 0.0388f
C2847 _328_/a_27_47# net50 5.21e-21
C2848 _332_/a_651_413# net40 6.24e-19
C2849 _192_/a_505_280# _096_ 3.38e-20
C2850 _305_/a_27_47# clknet_2_1__leaf_clk 0.26f
C2851 _322_/a_1108_47# _209_/a_27_47# 1.04e-19
C2852 net1 _316_/a_639_47# 7.19e-21
C2853 _335_/a_193_47# net18 1.54e-19
C2854 _053_ net40 0.00149f
C2855 _019_ net52 9.79e-21
C2856 _339_/a_1032_413# _339_/a_1296_47# 0.00384f
C2857 _269_/a_81_21# _269_/a_384_47# 0.00138f
C2858 _168_/a_27_413# _171_/a_27_47# 0.00107f
C2859 _113_ net33 4.06e-22
C2860 trim[1] rebuffer2/a_75_212# 2.73e-19
C2861 _189_/a_218_47# _189_/a_408_47# 0.097f
C2862 _327_/a_193_47# _302_/a_27_297# 5.93e-20
C2863 _113_ trim_mask\[1\] 0.0392f
C2864 _030_ trim_val\[1\] 1.15e-19
C2865 net31 _333_/a_193_47# 9.64e-20
C2866 trim[4] output5/a_27_47# 0.00118f
C2867 _275_/a_81_21# net19 2.46e-21
C2868 _293_/a_81_21# _339_/a_1032_413# 1.08e-19
C2869 _050_ _331_/a_193_47# 0.00139f
C2870 trim_mask\[4\] trim_val\[4\] 0.336f
C2871 comp _299_/a_27_413# 4.35e-19
C2872 cal_count\[1\] _339_/a_27_47# 1.09e-19
C2873 _276_/a_59_75# _335_/a_193_47# 1.13e-21
C2874 _119_ _330_/a_1283_21# 4.21e-20
C2875 VPWR _026_ 0.389f
C2876 net51 _073_ 2.67e-20
C2877 _101_ rebuffer5/a_161_47# 0.0034f
C2878 clkbuf_2_0__f_clk/a_110_47# _319_/a_27_47# 4.99e-19
C2879 _294_/a_68_297# cal_count\[2\] 0.101f
C2880 _072_ _202_/a_79_21# 0.171f
C2881 _166_/a_161_47# _087_ 1.03e-19
C2882 _058_ _302_/a_27_297# 0.00216f
C2883 _279_/a_204_297# _279_/a_206_47# 1.91e-19
C2884 _279_/a_396_47# _279_/a_490_47# 0.0245f
C2885 _303_/a_1283_21# _303_/a_1108_47# 0.234f
C2886 _303_/a_761_289# _303_/a_651_413# 0.0977f
C2887 _303_/a_27_47# _303_/a_639_47# 0.00188f
C2888 _303_/a_193_47# _303_/a_1270_413# 1.46e-19
C2889 _303_/a_543_47# _303_/a_448_47# 0.0498f
C2890 net2 net33 0.612f
C2891 output28/a_27_47# result[6] 0.332f
C2892 _020_ _312_/a_1108_47# 6.99e-22
C2893 _253_/a_299_297# net25 5.91e-19
C2894 clknet_2_1__leaf_clk _011_ 0.185f
C2895 _237_/a_218_47# _099_ 0.00187f
C2896 _068_ clkbuf_2_3__f_clk/a_110_47# 2.29e-19
C2897 net54 _337_/a_761_289# 1.02e-19
C2898 _078_ net26 0.062f
C2899 _323_/a_448_47# _020_ 0.158f
C2900 cal_itt\[1\] clknet_2_3__leaf_clk 0.00118f
C2901 _305_/a_193_47# _202_/a_79_21# 2.48e-19
C2902 _290_/a_27_413# net2 5.47e-21
C2903 _322_/a_1283_21# _205_/a_27_47# 0.00472f
C2904 _019_ _320_/a_761_289# 1.17e-19
C2905 _169_/a_215_311# _167_/a_161_47# 7.46e-19
C2906 _314_/a_1283_21# net14 0.00117f
C2907 _094_ net22 0.00156f
C2908 VPWR _316_/a_27_47# 0.522f
C2909 _321_/a_193_47# _310_/a_1108_47# 2.49e-20
C2910 _321_/a_448_47# _310_/a_27_47# 6.41e-22
C2911 _051_ _062_ 0.0941f
C2912 _256_/a_373_47# net46 5.19e-20
C2913 calibrate _100_ 0.631f
C2914 _324_/a_543_47# _324_/a_651_413# 0.0572f
C2915 _324_/a_761_289# _324_/a_1270_413# 2.6e-19
C2916 _324_/a_193_47# _324_/a_639_47# 2.28e-19
C2917 net13 _322_/a_651_413# 0.00105f
C2918 _300_/a_47_47# net16 2.14e-19
C2919 _017_ net52 0.0168f
C2920 _064_ rebuffer3/a_75_212# 0.00294f
C2921 _316_/a_761_289# net41 0.0219f
C2922 _319_/a_1270_413# clknet_2_0__leaf_clk 4.01e-19
C2923 _015_ net3 0.0538f
C2924 mask\[1\] _245_/a_109_47# 0.00256f
C2925 _200_/a_80_21# net4 0.00116f
C2926 _048_ _242_/a_297_47# 0.0482f
C2927 _014_ _096_ 7.19e-19
C2928 _309_/a_1108_47# net43 0.221f
C2929 net6 ctln[0] 0.0657f
C2930 _325_/a_651_413# _159_/a_27_47# 1.26e-19
C2931 _325_/a_543_47# _046_ 1.31e-19
C2932 clknet_2_0__leaf_clk net55 3.53e-19
C2933 net14 _310_/a_27_47# 0.00725f
C2934 _110_ _027_ 0.00725f
C2935 _327_/a_1462_47# net18 5.71e-20
C2936 _327_/a_193_47# trim_mask\[0\] 0.00497f
C2937 _324_/a_27_47# mask\[4\] 9.76e-21
C2938 _229_/a_27_297# _228_/a_79_21# 5.4e-20
C2939 _053_ _304_/a_1108_47# 7.74e-19
C2940 mask\[7\] _314_/a_193_47# 5.51e-19
C2941 _305_/a_543_47# _002_ 0.0364f
C2942 net31 trimb[2] 3.03e-20
C2943 net9 _300_/a_377_297# 5.89e-20
C2944 net16 _029_ 4.6e-19
C2945 _309_/a_448_47# _309_/a_639_47# 4.61e-19
C2946 _232_/a_32_297# _232_/a_114_297# 0.0139f
C2947 _320_/a_1108_47# _208_/a_505_21# 5.98e-21
C2948 VPWR sample 0.531f
C2949 net23 _040_ 0.0546f
C2950 _190_/a_215_47# _190_/a_465_47# 0.089f
C2951 _321_/a_27_47# _247_/a_27_297# 0.00133f
C2952 _057_ clknet_2_2__leaf_clk 2.3e-19
C2953 VPWR net40 2.22f
C2954 trim_mask\[0\] _058_ 0.142f
C2955 _322_/a_543_47# _322_/a_1108_47# 7.99e-20
C2956 _322_/a_193_47# _322_/a_651_413# 0.0306f
C2957 net43 result[6] 7.22e-20
C2958 _064_ _105_ 3.99e-19
C2959 _250_/a_109_297# clknet_2_1__leaf_clk 9.25e-19
C2960 _320_/a_761_289# _017_ 7.03e-19
C2961 _320_/a_1108_47# mask\[2\] 5.22e-21
C2962 trim_val\[1\] net33 0.127f
C2963 _272_/a_81_21# _056_ 2.92e-20
C2964 result[7] _074_ 1.76e-20
C2965 _335_/a_1462_47# net18 3.94e-19
C2966 _332_/a_1283_21# clknet_2_3__leaf_clk 1.26e-21
C2967 valid sample 0.0379f
C2968 mask\[0\] _315_/a_27_47# 1.54e-19
C2969 net22 _315_/a_193_47# 0.00108f
C2970 trim_val\[1\] trim_mask\[1\] 0.32f
C2971 _259_/a_109_47# _064_ 0.00153f
C2972 _259_/a_27_297# _104_ 0.201f
C2973 _253_/a_81_21# _310_/a_1283_21# 6.89e-19
C2974 _327_/a_1283_21# _136_ 0.00212f
C2975 _327_/a_27_47# _038_ 2.98e-20
C2976 trim_mask\[1\] _336_/a_193_47# 0.00141f
C2977 _200_/a_80_21# _063_ 0.0782f
C2978 _123_ net33 4.06e-22
C2979 _336_/a_27_47# _336_/a_543_47# 0.109f
C2980 _336_/a_193_47# _336_/a_761_289# 0.175f
C2981 net2 _069_ 0.0612f
C2982 output35/a_27_47# _130_ 0.00105f
C2983 clknet_2_1__leaf_clk _319_/a_1283_21# 0.0013f
C2984 _050_ _260_/a_93_21# 0.0243f
C2985 _319_/a_27_47# _319_/a_448_47# 0.0867f
C2986 VPWR _003_ 0.418f
C2987 _319_/a_193_47# _319_/a_1108_47# 0.125f
C2988 _308_/a_761_289# _080_ 4.22e-19
C2989 result[4] _253_/a_81_21# 9.76e-20
C2990 _305_/a_1283_21# _069_ 5.34e-20
C2991 VPWR _149_/a_68_297# 0.179f
C2992 _128_ _339_/a_1224_47# 1.82e-19
C2993 _110_ _335_/a_448_47# 0.00206f
C2994 trim_mask\[0\] _332_/a_27_47# 0.00555f
C2995 VPWR trimb[0] 0.581f
C2996 _249_/a_27_297# _249_/a_373_47# 0.0134f
C2997 _293_/a_81_21# _293_/a_299_297# 0.0821f
C2998 _303_/a_543_47# _000_ 0.00213f
C2999 _074_ net22 0.191f
C3000 _097_ _315_/a_1108_47# 2.42e-20
C3001 VPWR _299_/a_215_297# 0.207f
C3002 _243_/a_109_297# _100_ 0.00161f
C3003 _243_/a_27_297# _096_ 0.0924f
C3004 _089_ _075_ 5.41e-22
C3005 _047_ _332_/a_1108_47# 1.66e-19
C3006 clkbuf_0_clk/a_110_47# _068_ 0.0139f
C3007 _324_/a_543_47# mask\[5\] 2.57e-19
C3008 _324_/a_27_47# _020_ 6.39e-20
C3009 _034_ _092_ 0.00377f
C3010 _071_ clk 6.42e-20
C3011 _317_/a_193_47# _316_/a_651_413# 5.3e-20
C3012 _317_/a_448_47# _316_/a_761_289# 1.99e-20
C3013 _317_/a_1283_21# _316_/a_1283_21# 1.13e-19
C3014 _292_/a_78_199# _036_ 0.106f
C3015 _337_/a_1283_21# net51 9.5e-20
C3016 _277_/a_75_212# net46 0.00127f
C3017 _305_/a_1108_47# _067_ 7.47e-19
C3018 _305_/a_1108_47# _070_ 0.00102f
C3019 clknet_2_2__leaf_clk _330_/a_448_47# 0.0254f
C3020 net44 rebuffer4/a_27_47# 0.00187f
C3021 _125_ _130_ 4.49e-21
C3022 VPWR _316_/a_1217_47# 3.62e-20
C3023 net22 _014_ 5.06e-20
C3024 mask\[0\] clknet_2_0__leaf_clk 0.0635f
C3025 _064_ _194_/a_113_297# 0.0518f
C3026 _104_ trim_mask\[1\] 0.212f
C3027 net4 net46 0.0382f
C3028 _136_ _332_/a_543_47# 8.86e-19
C3029 _136_ _108_ 0.008f
C3030 _064_ _336_/a_1283_21# 2.96e-19
C3031 _104_ _336_/a_761_289# 0.0473f
C3032 _249_/a_109_47# mask\[4\] 0.00134f
C3033 _237_/a_76_199# en_co_clk 4.52e-20
C3034 _013_ output41/a_27_47# 2.01e-20
C3035 _097_ _012_ 7.01e-20
C3036 _074_ _313_/a_1108_47# 6.62e-20
C3037 _232_/a_114_297# net55 0.00257f
C3038 _329_/a_193_47# _064_ 5.56e-20
C3039 net4 _195_/a_439_47# 4.03e-19
C3040 _071_ net4 1.18e-21
C3041 trim_mask\[2\] _334_/a_761_289# 1.47e-20
C3042 VPWR _304_/a_1108_47# 0.307f
C3043 _104_ clone1/a_27_47# 1.3e-19
C3044 mask\[3\] net21 9.79e-21
C3045 _327_/a_1462_47# trim_mask\[0\] 5.41e-21
C3046 _087_ _088_ 4.44e-20
C3047 _164_/a_161_47# _095_ 5.12e-19
C3048 output23/a_27_47# net22 6.71e-20
C3049 net2 _078_ 6.06e-20
C3050 _200_/a_209_297# net19 0.00228f
C3051 _251_/a_27_297# mask\[6\] 0.132f
C3052 mask\[6\] _250_/a_109_47# 0.00348f
C3053 clone1/a_27_47# net55 0.181f
C3054 net12 _311_/a_193_47# 1.11e-19
C3055 state\[2\] _228_/a_382_297# 1.95e-19
C3056 net52 _310_/a_27_47# 5.43e-22
C3057 _308_/a_27_47# mask\[1\] 3.15e-20
C3058 cal_itt\[1\] _266_/a_68_297# 8.13e-20
C3059 _240_/a_109_297# _049_ 5.97e-22
C3060 _123_ _069_ 5.86e-20
C3061 _119_ _108_ 0.00869f
C3062 _328_/a_1283_21# _058_ 0.0034f
C3063 _239_/a_694_21# net42 1.79e-19
C3064 net46 _063_ 1.01e-21
C3065 _113_ _270_/a_59_75# 0.11f
C3066 _021_ clknet_2_1__leaf_clk 0.143f
C3067 trim_mask\[2\] _335_/a_27_47# 3.11e-19
C3068 state\[0\] clk 2.86e-19
C3069 net48 net49 0.00261f
C3070 _272_/a_384_47# trim_val\[2\] 3.41e-19
C3071 _272_/a_81_21# net48 0.00566f
C3072 _023_ _310_/a_448_47# 4.05e-19
C3073 _037_ net46 1.3e-20
C3074 trim_mask\[1\] _336_/a_1462_47# 1.97e-21
C3075 _273_/a_145_75# net46 3.61e-19
C3076 _320_/a_1108_47# mask\[1\] 0.0542f
C3077 _071_ _063_ 0.0685f
C3078 clknet_0_clk _171_/a_27_47# 0.00186f
C3079 _200_/a_209_297# _107_ 4.95e-20
C3080 _322_/a_1283_21# _083_ 4.82e-19
C3081 _321_/a_543_47# net15 0.00541f
C3082 cal_itt\[0\] _341_/a_761_289# 1.25e-20
C3083 _336_/a_1283_21# _264_/a_27_297# 1.04e-19
C3084 _079_ _315_/a_193_47# 7.45e-20
C3085 _336_/a_27_47# _106_ 0.0015f
C3086 _281_/a_253_47# _092_ 0.0386f
C3087 trim[4] _047_ 0.0025f
C3088 _005_ _213_/a_109_297# 0.0125f
C3089 net44 _311_/a_193_47# 0.0334f
C3090 _107_ _228_/a_79_21# 0.00492f
C3091 _300_/a_47_47# net40 0.00196f
C3092 _290_/a_207_413# _127_ 0.0902f
C3093 _053_ _331_/a_543_47# 1.42e-21
C3094 trim_mask\[2\] rebuffer1/a_75_212# 0.053f
C3095 VPWR _256_/a_109_47# 6.98e-20
C3096 _110_ _032_ 0.111f
C3097 calibrate _316_/a_193_47# 4.87e-20
C3098 _093_ _316_/a_27_47# 2.78e-20
C3099 _235_/a_79_21# _337_/a_543_47# 1.39e-19
C3100 trim_mask\[0\] _332_/a_1217_47# 0.00108f
C3101 _329_/a_543_47# _329_/a_1108_47# 7.99e-20
C3102 _329_/a_193_47# _329_/a_651_413# 0.0346f
C3103 _249_/a_109_47# _020_ 6.05e-20
C3104 _235_/a_297_47# _337_/a_193_47# 6.67e-21
C3105 VPWR _321_/a_1108_47# 0.304f
C3106 state\[0\] net4 0.0129f
C3107 clknet_2_1__leaf_clk _313_/a_761_289# 0.0433f
C3108 _060_ _090_ 0.00512f
C3109 _306_/a_27_47# clkbuf_0_clk/a_110_47# 1.17e-20
C3110 VPWR _337_/a_1108_47# 0.288f
C3111 _286_/a_76_199# net18 0.0103f
C3112 clkbuf_2_0__f_clk/a_110_47# _282_/a_68_297# 0.0126f
C3113 VPWR _167_/a_161_47# 0.611f
C3114 _321_/a_1108_47# net53 4.72e-19
C3115 _006_ _310_/a_651_413# 1.1e-20
C3116 _014_ _316_/a_761_289# 0.00576f
C3117 clknet_2_0__leaf_clk _316_/a_543_47# 2.38e-19
C3118 net45 _316_/a_193_47# 0.0342f
C3119 _144_/a_27_47# trimb[4] 4.07e-21
C3120 _074_ _079_ 0.0789f
C3121 clknet_2_2__leaf_clk _027_ 0.0294f
C3122 _094_ clknet_0_clk 0.0166f
C3123 state\[2\] _169_/a_109_53# 0.0798f
C3124 _029_ net40 0.0203f
C3125 _322_/a_1108_47# mask\[2\] 8.23e-21
C3126 _058_ _333_/a_193_47# 0.00218f
C3127 _328_/a_639_47# net46 0.00181f
C3128 _122_ _132_ 7.95e-21
C3129 fanout45/a_27_47# net15 0.00307f
C3130 _058_ _265_/a_81_21# 0.0124f
C3131 _290_/a_207_413# _126_ 0.194f
C3132 _128_ _291_/a_285_297# 0.072f
C3133 _329_/a_543_47# net9 0.00535f
C3134 _301_/a_285_47# _332_/a_761_289# 8.57e-20
C3135 _028_ _052_ 0.207f
C3136 net2 fanout47/a_27_47# 5.94e-20
C3137 _023_ result[5] 8.38e-19
C3138 _327_/a_193_47# trim_mask\[4\] 0.00205f
C3139 _327_/a_448_47# clknet_2_2__leaf_clk 0.00253f
C3140 _226_/a_27_47# _095_ 3.66e-19
C3141 _299_/a_27_413# _132_ 0.0119f
C3142 _101_ net51 0.426f
C3143 _326_/a_27_47# _253_/a_81_21# 1.02e-19
C3144 VPWR _340_/a_562_413# 0.00334f
C3145 clknet_0_clk _192_/a_505_280# 0.0117f
C3146 _175_/a_150_297# rebuffer1/a_75_212# 1e-19
C3147 _121_ clknet_2_0__leaf_clk 0.0275f
C3148 ctlp[7] _156_/a_27_47# 3.27e-19
C3149 _333_/a_761_289# rebuffer1/a_75_212# 2.09e-20
C3150 _333_/a_27_47# _332_/a_193_47# 7.12e-22
C3151 _115_ rebuffer1/a_75_212# 9.01e-19
C3152 net30 net18 5.08e-20
C3153 _069_ _067_ 0.0468f
C3154 _069_ _070_ 0.13f
C3155 _304_/a_193_47# cal_count\[0\] 7.48e-20
C3156 _304_/a_543_47# _124_ 8.48e-20
C3157 net42 _106_ 2.06e-19
C3158 _265_/a_81_21# _332_/a_27_47# 3.01e-20
C3159 _058_ trim_mask\[4\] 0.134f
C3160 _337_/a_543_47# _049_ 0.0111f
C3161 net52 _310_/a_1217_47# 9.61e-21
C3162 _005_ _212_/a_113_297# 6.78e-19
C3163 _337_/a_193_47# net30 7.21e-20
C3164 _335_/a_448_47# clknet_2_2__leaf_clk 2.28e-19
C3165 VPWR _280_/a_75_212# 0.209f
C3166 trim_mask\[1\] _172_/a_150_297# 5.26e-20
C3167 net49 _172_/a_68_297# 0.00295f
C3168 _289_/a_68_297# _126_ 0.106f
C3169 trim_mask\[0\] _227_/a_109_93# 0.0225f
C3170 output9/a_27_47# ctln[3] 0.159f
C3171 _341_/a_805_47# net46 0.00322f
C3172 _246_/a_27_297# mask\[2\] 0.112f
C3173 net27 net21 0.448f
C3174 mask\[0\] _319_/a_639_47# 0.00449f
C3175 VPWR _198_/a_181_47# 2.14e-19
C3176 _333_/a_448_47# net46 0.0181f
C3177 fanout46/a_27_47# clkbuf_2_2__f_clk/a_110_47# 0.0029f
C3178 _307_/a_27_47# _039_ 7.99e-19
C3179 net12 net41 5.07e-20
C3180 VPWR _331_/a_543_47# 0.216f
C3181 _286_/a_218_47# clknet_2_3__leaf_clk 2.48e-19
C3182 _332_/a_1108_47# clknet_2_2__leaf_clk 2.43e-21
C3183 _051_ _227_/a_209_311# 0.00701f
C3184 mask\[6\] _313_/a_543_47# 8.25e-21
C3185 net44 _311_/a_1462_47# 0.00222f
C3186 VPWR _258_/a_109_297# 0.191f
C3187 net27 _312_/a_1283_21# 0.0716f
C3188 cal_itt\[0\] _303_/a_27_47# 1.43e-19
C3189 _053_ _260_/a_256_47# 0.00107f
C3190 _329_/a_761_289# _026_ 7.06e-19
C3191 _094_ _337_/a_651_413# 8.78e-22
C3192 _104_ _255_/a_27_47# 0.096f
C3193 net13 _169_/a_215_311# 0.0132f
C3194 VPWR _229_/a_27_297# 0.362f
C3195 _135_ net34 1.32e-20
C3196 _035_ _124_ 0.00385f
C3197 net28 _314_/a_193_47# 0.0133f
C3198 net5 _135_ 1.05e-19
C3199 _309_/a_27_47# _310_/a_27_47# 2.63e-19
C3200 _023_ net29 1.43e-21
C3201 output25/a_27_47# net25 0.179f
C3202 _064_ _278_/a_27_47# 0.00201f
C3203 cal_count\[0\] net18 0.00559f
C3204 _281_/a_103_199# en_co_clk 0.171f
C3205 net12 _306_/a_448_47# 0.00883f
C3206 _255_/a_27_47# net55 0.00894f
C3207 _317_/a_651_413# net14 2.17e-19
C3208 net45 _316_/a_1462_47# 0.00196f
C3209 _326_/a_651_413# net14 0.00477f
C3210 _325_/a_639_47# net43 0.00118f
C3211 _053_ net19 0.0347f
C3212 cal_count\[0\] _129_ 0.0507f
C3213 _134_ comp 1.07e-19
C3214 _313_/a_27_47# _313_/a_761_289# 0.0535f
C3215 net46 _279_/a_396_47# 7.7e-19
C3216 net35 _109_ 3.95e-20
C3217 _308_/a_1108_47# _039_ 0.00137f
C3218 net8 net33 1.21e-19
C3219 mask\[7\] net26 0.0661f
C3220 trim[2] net32 6.26e-20
C3221 _308_/a_1283_21# fanout43/a_27_47# 0.00444f
C3222 _331_/a_193_47# _049_ 1.54e-19
C3223 _185_/a_68_297# _099_ 7.19e-21
C3224 VPWR _338_/a_1602_47# 0.184f
C3225 _306_/a_448_47# net44 6.13e-19
C3226 _168_/a_207_413# _168_/a_297_47# 0.00476f
C3227 _046_ net29 0.00419f
C3228 _059_ _263_/a_382_297# 0.016f
C3229 _075_ _092_ 0.0268f
C3230 input3/a_75_212# net3 0.108f
C3231 _326_/a_1283_21# mask\[7\] 0.0788f
C3232 _326_/a_543_47# _102_ 1.05e-19
C3233 _326_/a_761_289# _023_ 8.7e-19
C3234 trim_mask\[0\] _054_ 5.81e-20
C3235 _053_ _107_ 0.0484f
C3236 VPWR _273_/a_59_75# 0.226f
C3237 trim_mask\[0\] net30 0.0433f
C3238 _050_ _281_/a_103_199# 0.018f
C3239 trim_mask\[3\] _057_ 0.00172f
C3240 output39/a_27_47# net16 0.00133f
C3241 VPWR output18/a_27_47# 0.291f
C3242 _286_/a_76_199# _338_/a_652_21# 1.79e-19
C3243 _208_/a_76_199# _208_/a_218_47# 0.00783f
C3244 trim_val\[0\] _332_/a_1108_47# 0.0019f
C3245 VPWR _214_/a_113_297# 0.235f
C3246 net43 _314_/a_1108_47# 0.242f
C3247 clk _317_/a_651_413# 0.00154f
C3248 _340_/a_1182_261# cal_count\[0\] 1.02e-20
C3249 net12 _094_ 1.21e-20
C3250 mask\[0\] _078_ 0.177f
C3251 _257_/a_109_47# net46 1.94e-21
C3252 _032_ clknet_2_2__leaf_clk 0.0022f
C3253 _315_/a_761_289# net14 0.0127f
C3254 trim[1] net33 0.00648f
C3255 _051_ _318_/a_1108_47# 2.53e-19
C3256 _187_/a_212_413# _136_ 1.66e-19
C3257 _340_/a_193_47# net2 1.9e-19
C3258 _048_ en_co_clk 0.0131f
C3259 _290_/a_297_47# net34 1.65e-19
C3260 _141_/a_27_47# _040_ 0.193f
C3261 cal_itt\[2\] _092_ 0.0943f
C3262 clkbuf_0_clk/a_110_47# cal_itt\[3\] 0.01f
C3263 VPWR _320_/a_193_47# 0.358f
C3264 mask\[1\] _246_/a_27_297# 0.06f
C3265 _325_/a_1283_21# _019_ 9.46e-20
C3266 _167_/a_161_47# _093_ 2.98e-20
C3267 VPWR _260_/a_256_47# 1.63e-19
C3268 net43 _310_/a_193_47# 0.0404f
C3269 mask\[3\] mask\[4\] 0.0432f
C3270 _287_/a_75_212# _123_ 2.48e-19
C3271 _322_/a_639_47# mask\[3\] 2.74e-19
C3272 _032_ net11 1.11e-19
C3273 VPWR _328_/a_1270_413# 4.98e-19
C3274 cal_itt\[0\] _303_/a_1217_47# 1.13e-19
C3275 calibrate net14 0.0958f
C3276 _300_/a_285_47# cal_count\[3\] 0.0353f
C3277 output20/a_27_47# _312_/a_543_47# 0.0111f
C3278 _324_/a_193_47# _311_/a_1283_21# 4.08e-19
C3279 _324_/a_27_47# _311_/a_1108_47# 2.8e-21
C3280 _094_ net44 0.14f
C3281 _191_/a_27_297# net30 0.00331f
C3282 net13 _053_ 5.12e-19
C3283 net22 output30/a_27_47# 0.00146f
C3284 _305_/a_27_47# clkbuf_0_clk/a_110_47# 7.19e-20
C3285 _125_ _339_/a_1182_261# 9.71e-21
C3286 net28 _314_/a_1462_47# 7.77e-20
C3287 _323_/a_193_47# net26 0.00549f
C3288 _108_ _279_/a_206_47# 0.0318f
C3289 fanout47/a_27_47# _067_ 5.48e-19
C3290 net50 _330_/a_1108_47# 1.17e-20
C3291 _325_/a_27_47# _325_/a_193_47# 0.854f
C3292 fanout47/a_27_47# _070_ 1.46e-19
C3293 VPWR _312_/a_651_413# 0.142f
C3294 VPWR net19 1.54f
C3295 en_co_clk _120_ 0.129f
C3296 net45 net14 0.0278f
C3297 VPWR _307_/a_761_289# 0.207f
C3298 VPWR _323_/a_1270_413# 5.68e-19
C3299 _050_ _048_ 0.175f
C3300 _239_/a_694_21# _098_ 0.127f
C3301 _068_ _190_/a_215_47# 0.00289f
C3302 _313_/a_1108_47# _313_/a_1270_413# 0.00645f
C3303 _313_/a_761_289# _313_/a_1217_47# 4.2e-19
C3304 _313_/a_543_47# _313_/a_805_47# 0.00171f
C3305 _336_/a_651_413# clkbuf_2_2__f_clk/a_110_47# 0.00129f
C3306 _337_/a_448_47# _065_ 1.52e-19
C3307 trim_mask\[0\] _262_/a_465_47# 4.46e-19
C3308 net12 _318_/a_639_47# 2.31e-19
C3309 _326_/a_651_413# net52 1.99e-20
C3310 output36/a_27_47# _126_ 2.66e-19
C3311 fanout45/a_27_47# state\[1\] 0.0119f
C3312 _321_/a_27_47# _042_ 0.106f
C3313 _339_/a_1032_413# output40/a_27_47# 1.1e-20
C3314 en_co_clk _076_ 0.129f
C3315 _077_ rebuffer5/a_161_47# 0.0119f
C3316 _061_ trim_mask\[0\] 5.78e-19
C3317 trim[4] trim_val\[0\] 1.61e-19
C3318 comp cal_count\[2\] 8.28e-20
C3319 _322_/a_27_47# net51 3.21e-20
C3320 _260_/a_93_21# _049_ 0.11f
C3321 VPWR _107_ 1.04f
C3322 _321_/a_1283_21# clknet_2_1__leaf_clk 0.0101f
C3323 clk calibrate 6.08e-20
C3324 VPWR _333_/a_1108_47# 0.293f
C3325 net32 _055_ 0.0157f
C3326 net12 _074_ 4.02e-19
C3327 trim[1] output33/a_27_47# 7.46e-20
C3328 _340_/a_193_47# _123_ 0.0182f
C3329 _136_ net2 0.0141f
C3330 _275_/a_81_21# _335_/a_761_289# 0.00132f
C3331 _275_/a_299_297# _335_/a_193_47# 6.67e-20
C3332 _294_/a_150_297# _125_ 2.38e-20
C3333 _050_ _120_ 0.0965f
C3334 _090_ net30 9.79e-21
C3335 _041_ _124_ 0.112f
C3336 cal_count\[0\] _338_/a_652_21# 2.2e-20
C3337 _330_/a_193_47# _330_/a_639_47# 2.28e-19
C3338 _330_/a_761_289# _330_/a_1270_413# 2.6e-19
C3339 _330_/a_543_47# _330_/a_651_413# 0.0572f
C3340 _143_/a_68_297# _065_ 8.62e-20
C3341 calibrate _331_/a_1283_21# 1.23e-19
C3342 clk net45 0.323f
C3343 trim_mask\[4\] _227_/a_109_93# 3.9e-21
C3344 VPWR _308_/a_651_413# 0.144f
C3345 _237_/a_76_199# net15 0.00477f
C3346 _048_ _228_/a_297_47# 0.00637f
C3347 _074_ _159_/a_27_47# 1.62e-19
C3348 cal_count\[0\] _297_/a_47_47# 4.49e-21
C3349 _015_ _318_/a_1108_47# 1.26e-19
C3350 state\[2\] _318_/a_193_47# 0.00416f
C3351 calibrate net4 2.6e-19
C3352 mask\[4\] _068_ 3.07e-20
C3353 _004_ mask\[0\] 8.96e-20
C3354 VPWR _237_/a_218_374# 0.00203f
C3355 net27 _045_ 6.13e-19
C3356 mask\[1\] _208_/a_535_374# 2.87e-20
C3357 net16 _298_/a_493_297# 3.42e-20
C3358 net45 _331_/a_1283_21# 0.338f
C3359 _081_ clknet_2_0__leaf_clk 2.17e-20
C3360 _074_ net44 0.137f
C3361 VPWR _320_/a_1462_47# 6.24e-19
C3362 _066_ net18 0.0344f
C3363 VPWR _339_/a_381_47# 0.104f
C3364 net43 _310_/a_1462_47# 0.00413f
C3365 ctlp[2] trimb[3] 0.00996f
C3366 result[5] result[6] 0.035f
C3367 _208_/a_505_21# rebuffer4/a_27_47# 0.00391f
C3368 _328_/a_193_47# _113_ 8.33e-20
C3369 _328_/a_27_47# _030_ 2.88e-20
C3370 _328_/a_1108_47# _271_/a_75_212# 4.38e-19
C3371 clk _065_ 2.07e-20
C3372 trim_mask\[2\] _271_/a_75_212# 8.82e-19
C3373 net4 net45 0.179f
C3374 _297_/a_285_47# _132_ 0.067f
C3375 VPWR net13 1.38f
C3376 VPWR _155_/a_68_297# 0.169f
C3377 _078_ _010_ 8.71e-19
C3378 _047_ net49 4.23e-21
C3379 VPWR _279_/a_27_47# 0.238f
C3380 _125_ _339_/a_1296_47# 7.89e-21
C3381 _339_/a_27_47# _286_/a_535_374# 7e-20
C3382 VPWR output28/a_27_47# 0.402f
C3383 net12 _305_/a_448_47# 2.34e-19
C3384 trim_mask\[3\] _027_ 0.0622f
C3385 trim_val\[3\] net46 0.075f
C3386 _193_/a_109_297# net46 1.51e-19
C3387 _325_/a_761_289# _325_/a_805_47# 3.69e-19
C3388 _325_/a_193_47# _325_/a_1217_47# 2.36e-20
C3389 _325_/a_543_47# _325_/a_639_47# 0.0138f
C3390 _307_/a_1283_21# _094_ 8.61e-21
C3391 _053_ _118_ 1.98e-19
C3392 net13 net53 0.0143f
C3393 _110_ _272_/a_81_21# 4.04e-19
C3394 _110_ net49 8.81e-19
C3395 net9 _298_/a_215_47# 2.06e-20
C3396 _079_ output30/a_27_47# 0.00107f
C3397 _293_/a_81_21# _125_ 0.206f
C3398 _110_ _336_/a_543_47# 0.00179f
C3399 VPWR _324_/a_761_289# 0.22f
C3400 output14/a_27_47# net28 0.0464f
C3401 net31 comp 0.149f
C3402 net16 _129_ 0.791f
C3403 VPWR net39 0.307f
C3404 _302_/a_27_297# _066_ 0.278f
C3405 net43 _224_/a_113_297# 0.0107f
C3406 net4 _065_ 0.0126f
C3407 _329_/a_27_47# _110_ 1.2e-19
C3408 mask\[4\] _311_/a_448_47# 0.0249f
C3409 net27 mask\[4\] 9.99e-19
C3410 _226_/a_197_47# _075_ 0.00123f
C3411 net15 _241_/a_388_297# 0.00192f
C3412 _146_/a_68_297# _081_ 1.07e-20
C3413 clknet_0_clk _106_ 5.55e-20
C3414 _324_/a_761_289# net53 5.65e-19
C3415 _321_/a_27_47# _022_ 7.92e-21
C3416 _169_/a_215_311# net3 5.43e-20
C3417 output34/a_27_47# trim[3] 0.337f
C3418 _136_ _123_ 5.71e-19
C3419 _237_/a_76_199# _049_ 2.74e-19
C3420 _155_/a_68_297# _009_ 2.08e-21
C3421 net45 net52 0.356f
C3422 clknet_2_0__leaf_clk _016_ 0.0814f
C3423 net4 _105_ 0.00345f
C3424 VPWR _322_/a_193_47# 0.407f
C3425 VPWR _248_/a_109_297# 0.199f
C3426 _337_/a_1108_47# _206_/a_27_93# 0.00254f
C3427 _321_/a_1217_47# _042_ 1.61e-19
C3428 _063_ rebuffer3/a_75_212# 6.07e-20
C3429 VPWR _257_/a_109_297# 0.196f
C3430 _083_ _311_/a_27_47# 0.0291f
C3431 _303_/a_27_47# net26 6.75e-20
C3432 _305_/a_448_47# net44 0.00192f
C3433 net27 _220_/a_199_47# 0.00142f
C3434 _059_ _095_ 7.45e-19
C3435 trim[4] _131_ 3.48e-21
C3436 trim_mask\[4\] _054_ 1.48e-20
C3437 _069_ clknet_2_3__leaf_clk 4.01e-20
C3438 _322_/a_1217_47# net51 1.93e-20
C3439 trim_mask\[4\] net30 1.57e-19
C3440 _262_/a_27_47# net19 0.00233f
C3441 net13 _318_/a_27_47# 0.0199f
C3442 _316_/a_27_47# _316_/a_651_413# 9.73e-19
C3443 _316_/a_761_289# _316_/a_1108_47# 0.0512f
C3444 _316_/a_193_47# _316_/a_448_47# 0.0642f
C3445 _248_/a_109_297# net53 0.00625f
C3446 _322_/a_193_47# net53 2.02e-19
C3447 VPWR _303_/a_651_413# 0.143f
C3448 _200_/a_209_297# _062_ 0.0075f
C3449 _064_ _051_ 0.00148f
C3450 net50 _335_/a_1108_47# 0.0118f
C3451 result[6] net29 5.77e-20
C3452 cal_count\[0\] _338_/a_1056_47# 4.68e-20
C3453 _340_/a_1182_261# net16 7.99e-19
C3454 _117_ _104_ 8.64e-20
C3455 _179_/a_27_47# net34 0.12f
C3456 net52 _065_ 0.00701f
C3457 _330_/a_1283_21# _027_ 0.0413f
C3458 _330_/a_543_47# net46 0.152f
C3459 _065_ _063_ 4.66e-19
C3460 _188_/a_27_47# net34 0.00426f
C3461 _188_/a_27_47# net5 0.11f
C3462 _336_/a_193_47# _119_ 0.00802f
C3463 net54 en_co_clk 0.012f
C3464 _307_/a_1108_47# _315_/a_27_47# 4.72e-21
C3465 _307_/a_761_289# _315_/a_543_47# 5.13e-21
C3466 trim[1] _270_/a_59_75# 2.55e-20
C3467 _307_/a_543_47# _315_/a_761_289# 5.13e-21
C3468 _307_/a_27_47# _315_/a_1108_47# 4.72e-21
C3469 output32/a_27_47# _055_ 6.66e-22
C3470 VPWR net43 4.66f
C3471 calibrate _260_/a_346_47# 0.00602f
C3472 _015_ clkbuf_2_0__f_clk/a_110_47# 3.35e-20
C3473 _037_ _065_ 1.04e-20
C3474 _341_/a_761_289# net2 1.57e-22
C3475 _051_ _100_ 0.00624f
C3476 cal en 0.0365f
C3477 _105_ _063_ 0.127f
C3478 _320_/a_1283_21# clknet_2_0__leaf_clk 2.89e-20
C3479 _107_ _262_/a_27_47# 0.00775f
C3480 net43 net53 0.0152f
C3481 VPWR _309_/a_805_47# 2.95e-19
C3482 _057_ _108_ 2.53e-21
C3483 net27 _020_ 2.32e-20
C3484 _074_ _312_/a_639_47# 5.75e-21
C3485 mask\[7\] _251_/a_373_47# 9.47e-19
C3486 _328_/a_27_47# trim_mask\[1\] 0.0506f
C3487 _200_/a_80_21# cal_itt\[2\] 0.137f
C3488 trim_mask\[0\] _066_ 0.0715f
C3489 clknet_2_1__leaf_clk _101_ 1.01f
C3490 net12 _239_/a_694_21# 0.0098f
C3491 net9 _340_/a_1032_413# 0.00332f
C3492 net28 net26 1.3e-20
C3493 _319_/a_27_47# net52 5.23e-20
C3494 _092_ _170_/a_81_21# 6.21e-19
C3495 _007_ net25 0.0825f
C3496 net4 _336_/a_1283_21# 5.48e-19
C3497 _334_/a_193_47# _334_/a_761_289# 0.186f
C3498 _334_/a_27_47# _334_/a_543_47# 0.107f
C3499 _314_/a_193_47# _314_/a_543_47# 0.23f
C3500 _314_/a_27_47# _314_/a_1283_21# 0.0436f
C3501 en_co_clk _068_ 0.0292f
C3502 VPWR _118_ 0.292f
C3503 _339_/a_476_47# cal_count\[0\] 0.0503f
C3504 _320_/a_761_289# _065_ 7.65e-21
C3505 trim_mask\[0\] net16 0.0753f
C3506 _019_ _247_/a_109_297# 6.51e-21
C3507 _097_ fanout45/a_27_47# 2.22e-19
C3508 net12 _002_ 4.08e-19
C3509 net54 _050_ 2.65e-19
C3510 _104_ _119_ 0.103f
C3511 net25 mask\[3\] 0.199f
C3512 ctln[5] _330_/a_193_47# 1.07e-20
C3513 _307_/a_543_47# net45 0.153f
C3514 mask\[1\] rebuffer4/a_27_47# 2.18e-20
C3515 net9 cal_count\[3\] 0.129f
C3516 _307_/a_1108_47# clknet_2_0__leaf_clk 3.1e-19
C3517 wire42/a_75_212# net19 4.1e-22
C3518 trim[3] _334_/a_1283_21# 2.13e-19
C3519 _051_ _264_/a_27_297# 1.79e-20
C3520 _058_ _267_/a_145_75# 2.95e-19
C3521 net2 _339_/a_27_47# 1.57e-19
C3522 _074_ _209_/a_27_47# 0.00126f
C3523 _110_ _106_ 0.0828f
C3524 _336_/a_761_289# _266_/a_68_297# 4.53e-19
C3525 result[0] clknet_2_0__leaf_clk 0.152f
C3526 _093_ _107_ 1.73e-19
C3527 _136_ _067_ 8.31e-19
C3528 _251_/a_109_297# _046_ 1.51e-19
C3529 _237_/a_76_199# _315_/a_1108_47# 7.92e-21
C3530 net27 _222_/a_199_47# 0.00143f
C3531 _031_ _057_ 6.44e-20
C3532 ctlp[6] output21/a_27_47# 4.08e-19
C3533 _259_/a_109_297# clknet_2_2__leaf_clk 6.37e-21
C3534 _320_/a_27_47# clknet_2_1__leaf_clk 0.00248f
C3535 _320_/a_448_47# clkbuf_2_1__f_clk/a_110_47# 9.72e-19
C3536 _053_ net3 1.05e-20
C3537 VPWR _322_/a_1462_47# 0.00178f
C3538 _304_/a_761_289# _122_ 0.00631f
C3539 input3/a_75_212# output41/a_27_47# 0.0101f
C3540 _104_ _328_/a_193_47# 2.53e-20
C3541 _283_/a_75_212# net30 0.0273f
C3542 VPWR _025_ 0.333f
C3543 _336_/a_1283_21# _063_ 4.46e-19
C3544 _325_/a_27_47# net27 1.97e-20
C3545 _002_ net44 0.0123f
C3546 _308_/a_639_47# _074_ 0.00194f
C3547 _190_/a_27_47# net30 0.00291f
C3548 _107_ wire42/a_75_212# 0.00449f
C3549 net15 _281_/a_103_199# 0.0132f
C3550 ctln[7] _318_/a_639_47# 6.41e-20
C3551 net13 _318_/a_1217_47# 1.14e-19
C3552 _334_/a_193_47# rebuffer1/a_75_212# 1.5e-19
C3553 _316_/a_193_47# _013_ 0.223f
C3554 ctlp[1] mask\[7\] 5.33e-20
C3555 _329_/a_27_47# _274_/a_75_212# 8.25e-21
C3556 _237_/a_218_374# _093_ 1.07e-19
C3557 _323_/a_543_47# _042_ 0.0296f
C3558 trim_mask\[3\] _032_ 0.00318f
C3559 _192_/a_174_21# _099_ 4.16e-20
C3560 _192_/a_27_47# _095_ 0.149f
C3561 VPWR _281_/a_337_297# 0.00302f
C3562 clknet_2_1__leaf_clk _312_/a_448_47# 4.56e-19
C3563 _309_/a_193_47# _074_ 0.0142f
C3564 _087_ net55 0.0879f
C3565 _308_/a_1270_413# net45 1.41e-19
C3566 _186_/a_109_297# en_co_clk 9.86e-20
C3567 _326_/a_1270_413# net43 2.06e-19
C3568 net16 _297_/a_47_47# 1.68e-20
C3569 _007_ _310_/a_543_47# 5.1e-19
C3570 _122_ _298_/a_215_47# 0.0601f
C3571 net9 _038_ 1.21e-20
C3572 net13 _093_ 5.91e-20
C3573 net18 net40 0.0116f
C3574 _015_ _100_ 3.26e-20
C3575 net31 _161_/a_150_297# 2.19e-20
C3576 output10/a_27_47# trim_val\[3\] 0.0101f
C3577 ctln[4] _275_/a_81_21# 8.88e-19
C3578 _309_/a_27_47# net45 2.73e-20
C3579 mask\[0\] _245_/a_109_47# 0.0011f
C3580 _078_ _245_/a_109_297# 1.34e-20
C3581 _334_/a_1108_47# net46 0.237f
C3582 net49 clknet_2_2__leaf_clk 3.7e-21
C3583 net25 _310_/a_1283_21# 0.129f
C3584 _082_ _310_/a_193_47# 0.00178f
C3585 _129_ net40 0.083f
C3586 _315_/a_27_47# _095_ 5.58e-22
C3587 output27/a_27_47# _314_/a_27_47# 3.9e-19
C3588 net9 _338_/a_476_47# 7.29e-20
C3589 _300_/a_377_297# cal_count\[2\] 2.46e-19
C3590 _327_/a_543_47# net46 0.156f
C3591 _100_ _242_/a_79_21# 0.109f
C3592 _336_/a_543_47# clknet_2_2__leaf_clk 0.00149f
C3593 cal_itt\[1\] _195_/a_535_374# 1.1e-19
C3594 cal_itt\[0\] _195_/a_218_47# 2.23e-19
C3595 cal_itt\[2\] _071_ 0.447f
C3596 net51 _077_ 1.67e-19
C3597 result[1] _308_/a_543_47# 2.56e-19
C3598 _078_ net20 1.54e-19
C3599 _329_/a_27_47# clknet_2_2__leaf_clk 0.266f
C3600 _304_/a_193_47# _304_/a_1108_47# 0.125f
C3601 _304_/a_27_47# _304_/a_448_47# 0.0826f
C3602 _258_/a_27_297# _033_ 9.34e-20
C3603 _339_/a_27_47# _123_ 0.522f
C3604 fanout47/a_27_47# clknet_2_3__leaf_clk 1.9e-20
C3605 _040_ clknet_2_0__leaf_clk 0.0704f
C3606 _190_/a_215_47# cal_itt\[3\] 0.00223f
C3607 result[4] net25 1.25e-20
C3608 _190_/a_27_47# _072_ 3.88e-19
C3609 _329_/a_1108_47# _328_/a_1108_47# 4.15e-21
C3610 _329_/a_1108_47# trim_mask\[2\] 0.00264f
C3611 _314_/a_448_47# _314_/a_639_47# 4.61e-19
C3612 _026_ trim_mask\[0\] 1.75e-20
C3613 _132_ cal_count\[2\] 0.00622f
C3614 _110_ _270_/a_145_75# 0.00123f
C3615 _263_/a_297_47# net55 0.00256f
C3616 _302_/a_27_297# net40 1.71e-19
C3617 net35 net46 0.00522f
C3618 _327_/a_193_47# _327_/a_639_47# 2.28e-19
C3619 _327_/a_761_289# _327_/a_1270_413# 2.6e-19
C3620 _327_/a_543_47# _327_/a_651_413# 0.0572f
C3621 _048_ net15 0.0177f
C3622 _235_/a_79_21# _048_ 0.0273f
C3623 _032_ _330_/a_1283_21# 4.72e-19
C3624 _335_/a_543_47# net46 0.187f
C3625 _281_/a_103_199# _049_ 0.00104f
C3626 _164_/a_161_47# _317_/a_1108_47# 8.6e-20
C3627 _322_/a_543_47# _074_ 0.00617f
C3628 net34 net38 0.481f
C3629 _169_/a_109_53# _060_ 0.00124f
C3630 _059_ _226_/a_27_47# 0.00764f
C3631 _299_/a_215_297# _129_ 0.12f
C3632 _299_/a_27_413# _130_ 0.0431f
C3633 _053_ _062_ 0.162f
C3634 mask\[7\] _313_/a_448_47# 4.96e-21
C3635 _304_/a_27_47# _133_ 0.00172f
C3636 _136_ _284_/a_150_297# 1.5e-19
C3637 _006_ net22 7.26e-21
C3638 VPWR net3 2.8f
C3639 _081_ _078_ 0.0714f
C3640 _327_/a_639_47# _058_ 9.54e-19
C3641 VPWR _080_ 0.292f
C3642 clknet_2_0__leaf_clk _095_ 0.0837f
C3643 VPWR _330_/a_761_289# 0.209f
C3644 _027_ _108_ 8.23e-22
C3645 _332_/a_761_289# net46 0.181f
C3646 trim_mask\[2\] net9 0.0102f
C3647 _328_/a_1108_47# net9 0.0101f
C3648 _105_ _279_/a_396_47# 9.38e-20
C3649 _146_/a_68_297# _040_ 1.18e-21
C3650 _306_/a_27_47# _050_ 3.23e-20
C3651 _336_/a_1108_47# _107_ 0.00111f
C3652 trim_val\[2\] _175_/a_68_297# 0.202f
C3653 _340_/a_1032_413# _122_ 0.0353f
C3654 net13 _319_/a_193_47# 1.73e-20
C3655 trim_mask\[1\] _333_/a_1270_413# 1.17e-20
C3656 _112_ _333_/a_448_47# 0.00367f
C3657 net49 _333_/a_651_413# 0.00301f
C3658 _304_/a_1108_47# net18 6.42e-19
C3659 _324_/a_27_47# _250_/a_27_297# 1.46e-20
C3660 _235_/a_382_297# en_co_clk 3.21e-19
C3661 net15 _120_ 0.0591f
C3662 _298_/a_292_297# _133_ 0.00556f
C3663 _053_ _195_/a_76_199# 0.00262f
C3664 _310_/a_27_47# _310_/a_651_413# 9.73e-19
C3665 _310_/a_761_289# _310_/a_1108_47# 0.0512f
C3666 _310_/a_193_47# _310_/a_448_47# 0.0594f
C3667 net49 trim_val\[0\] 4.74e-20
C3668 net13 _243_/a_109_47# 0.00167f
C3669 _307_/a_193_47# _210_/a_113_297# 1.15e-19
C3670 _329_/a_1108_47# _115_ 5.13e-21
C3671 VPWR _325_/a_543_47# 0.202f
C3672 _327_/a_448_47# _108_ 9.48e-19
C3673 _239_/a_277_297# _107_ 5.69e-19
C3674 net21 _313_/a_761_289# 9.46e-19
C3675 net16 _175_/a_68_297# 0.00422f
C3676 _335_/a_193_47# _335_/a_639_47# 2.28e-19
C3677 _335_/a_761_289# _335_/a_1270_413# 2.6e-19
C3678 _335_/a_543_47# _335_/a_651_413# 0.0572f
C3679 net23 clknet_2_0__leaf_clk 7.41e-19
C3680 _324_/a_193_47# clknet_2_1__leaf_clk 0.0064f
C3681 net16 _333_/a_193_47# 0.0161f
C3682 result[4] _310_/a_543_47# 0.00118f
C3683 _122_ cal_count\[3\] 4.88e-19
C3684 trim_mask\[2\] trim[2] 1.25e-19
C3685 VPWR output34/a_27_47# 0.421f
C3686 _287_/a_75_212# clknet_2_3__leaf_clk 4.39e-22
C3687 clk _204_/a_75_212# 4.17e-19
C3688 net16 _265_/a_81_21# 0.0035f
C3689 trim_mask\[0\] net40 0.00625f
C3690 _107_ _206_/a_27_93# 1.04e-19
C3691 net31 _132_ 0.00487f
C3692 _048_ _049_ 0.598f
C3693 _091_ clkbuf_2_3__f_clk/a_110_47# 0.00418f
C3694 _313_/a_1108_47# _312_/a_193_47# 9.89e-22
C3695 _058_ _332_/a_1270_413# 3.02e-20
C3696 _078_ _016_ 3.68e-20
C3697 _189_/a_27_47# _092_ 0.018f
C3698 _066_ trim_mask\[4\] 2.16e-20
C3699 clknet_2_1__leaf_clk _248_/a_27_297# 2.24e-20
C3700 _322_/a_27_47# clknet_2_1__leaf_clk 0.243f
C3701 _127_ trimb[1] 6.52e-19
C3702 _336_/a_639_47# trim_mask\[4\] 0.00435f
C3703 _106_ clknet_2_2__leaf_clk 1.18e-19
C3704 net9 _115_ 2.05e-20
C3705 net43 _305_/a_1270_413# 2.53e-19
C3706 _256_/a_109_47# net18 4.58e-20
C3707 clk _316_/a_448_47# 2.08e-19
C3708 _336_/a_543_47# _279_/a_204_297# 4.32e-20
C3709 _336_/a_1108_47# _279_/a_27_47# 7.96e-19
C3710 _034_ _065_ 0.148f
C3711 _308_/a_27_47# mask\[0\] 6.38e-21
C3712 _308_/a_193_47# net22 8.85e-20
C3713 net24 _214_/a_113_297# 0.0111f
C3714 _321_/a_193_47# _321_/a_1108_47# 0.125f
C3715 _321_/a_27_47# _321_/a_448_47# 0.0859f
C3716 _332_/a_1108_47# _108_ 8.3e-20
C3717 _340_/a_27_47# _340_/a_193_47# 0.779f
C3718 _332_/a_193_47# _332_/a_651_413# 0.0276f
C3719 _332_/a_543_47# _332_/a_1108_47# 7.99e-20
C3720 _308_/a_27_47# output24/a_27_47# 3.92e-20
C3721 output14/a_27_47# _314_/a_543_47# 0.00343f
C3722 net27 _310_/a_543_47# 1.76e-21
C3723 _120_ _049_ 0.0916f
C3724 _164_/a_161_47# clknet_2_0__leaf_clk 4.38e-20
C3725 _292_/a_292_297# _123_ 0.00337f
C3726 VPWR _062_ 3.68f
C3727 _286_/a_439_47# _001_ 4.44e-20
C3728 _005_ clknet_2_1__leaf_clk 1.3e-21
C3729 net43 _319_/a_193_47# 0.0243f
C3730 _063_ _278_/a_27_47# 3.44e-19
C3731 _191_/a_27_297# net40 1.45e-19
C3732 VPWR fanout44/a_27_47# 0.305f
C3733 clkbuf_0_clk/a_110_47# _304_/a_1283_21# 1.75e-20
C3734 _185_/a_68_297# net41 0.0201f
C3735 net47 _298_/a_78_199# 8.16e-19
C3736 _232_/a_32_297# _099_ 0.0651f
C3737 mask\[7\] _010_ 0.00329f
C3738 _320_/a_1283_21# _078_ 4.8e-19
C3739 _337_/a_193_47# _337_/a_1108_47# 0.123f
C3740 _337_/a_27_47# _337_/a_448_47# 0.0897f
C3741 trimb[1] _126_ 4.36e-19
C3742 _038_ _122_ 0.00538f
C3743 _304_/a_639_47# clknet_2_3__leaf_clk 2.64e-19
C3744 _333_/a_1283_21# net32 0.00146f
C3745 net13 mask\[6\] 0.015f
C3746 net24 _320_/a_193_47# 9.63e-20
C3747 net26 _085_ 1.3e-20
C3748 _297_/a_47_47# net40 0.015f
C3749 _319_/a_1108_47# _283_/a_75_212# 0.00442f
C3750 mask\[6\] _155_/a_68_297# 0.193f
C3751 _340_/a_193_47# clknet_2_3__leaf_clk 0.0106f
C3752 _257_/a_109_297# _336_/a_1108_47# 1.54e-19
C3753 _076_ _049_ 0.143f
C3754 clkbuf_2_1__f_clk/a_110_47# _246_/a_109_297# 2.46e-19
C3755 trimb[2] net16 3.94e-19
C3756 _306_/a_1217_47# _050_ 3.14e-20
C3757 _291_/a_285_297# cal_count\[0\] 0.0075f
C3758 _015_ _316_/a_193_47# 7.75e-21
C3759 VPWR _195_/a_76_199# 0.103f
C3760 net3 _192_/a_548_47# 0.00123f
C3761 _097_ _237_/a_76_199# 0.0806f
C3762 _303_/a_27_47# _067_ 1.31e-22
C3763 mask\[3\] net15 0.00596f
C3764 clknet_2_1__leaf_clk _249_/a_373_47# 0.00105f
C3765 _303_/a_27_47# _070_ 8.05e-20
C3766 fanout43/a_27_47# _039_ 2.5e-19
C3767 _304_/a_27_47# net4 1.42e-21
C3768 VPWR _334_/a_1283_21# 0.379f
C3769 _326_/a_27_47# net25 2.09e-19
C3770 _013_ net14 3.23e-20
C3771 output8/a_27_47# trim_mask\[2\] 3e-19
C3772 _314_/a_1108_47# net29 0.0124f
C3773 _294_/a_68_297# net16 2.83e-19
C3774 _048_ _262_/a_193_297# 0.0224f
C3775 _307_/a_651_413# net22 0.00352f
C3776 VPWR _327_/a_761_289# 0.221f
C3777 _307_/a_1108_47# _078_ 0.0138f
C3778 VPWR _082_ 0.403f
C3779 net43 _202_/a_79_21# 0.00122f
C3780 result[0] _078_ 4.11e-20
C3781 _335_/a_1283_21# _032_ 1.97e-20
C3782 _088_ net41 1.32e-20
C3783 _074_ mask\[2\] 0.00154f
C3784 _299_/a_215_297# _297_/a_47_47# 4.73e-20
C3785 _322_/a_193_47# mask\[6\] 5.57e-22
C3786 _250_/a_109_297# mask\[4\] 3.11e-19
C3787 en_co_clk cal_itt\[3\] 1.08e-19
C3788 _280_/a_75_212# net18 6.73e-20
C3789 _328_/a_1283_21# net40 1.77e-21
C3790 _311_/a_761_289# _311_/a_639_47# 3.16e-19
C3791 _311_/a_27_47# _311_/a_1217_47# 2.56e-19
C3792 VPWR _137_/a_68_297# 0.186f
C3793 net43 output29/a_27_47# 4.29e-20
C3794 _072_ rebuffer5/a_161_47# 4.08e-21
C3795 _091_ cal_count\[3\] 2.04e-19
C3796 _322_/a_651_413# _042_ 2.18e-20
C3797 state\[2\] _103_ 0.00629f
C3798 _304_/a_1270_413# _136_ 1.97e-21
C3799 _310_/a_193_47# net29 9.97e-20
C3800 VPWR _335_/a_761_289# 0.212f
C3801 trim[4] _332_/a_543_47# 7.31e-20
C3802 _305_/a_27_47# en_co_clk 3.78e-21
C3803 _026_ trim_mask\[4\] 1.16e-19
C3804 _304_/a_805_47# net47 0.00316f
C3805 _194_/a_199_47# _118_ 9.57e-20
C3806 _096_ _092_ 0.276f
C3807 net55 _099_ 0.103f
C3808 _018_ _310_/a_27_47# 2.75e-21
C3809 _258_/a_109_297# net18 0.00283f
C3810 net43 mask\[6\] 0.414f
C3811 net54 _235_/a_79_21# 0.201f
C3812 _340_/a_652_21# net47 0.159f
C3813 _037_ _304_/a_27_47# 0.00269f
C3814 clk _013_ 1.58e-19
C3815 _336_/a_1108_47# _118_ 8.28e-20
C3816 VPWR _314_/a_805_47# 2.69e-19
C3817 _093_ net3 0.0565f
C3818 _065_ _208_/a_76_199# 0.158f
C3819 _097_ _241_/a_388_297# 0.0012f
C3820 _106_ _279_/a_204_297# 0.00183f
C3821 net42 _092_ 0.0793f
C3822 VPWR _332_/a_193_47# 0.275f
C3823 ctlp[1] net28 3.32e-19
C3824 _340_/a_193_47# _340_/a_586_47# 0.00206f
C3825 _302_/a_373_47# cal_count\[3\] 0.00137f
C3826 _136_ clknet_2_3__leaf_clk 0.181f
C3827 _088_ _171_/a_27_47# 5.46e-19
C3828 _048_ state\[1\] 6.16e-19
C3829 _253_/a_81_21# _253_/a_384_47# 0.00138f
C3830 net43 _319_/a_1462_47# 0.00223f
C3831 ctlp[1] _158_/a_68_297# 3.63e-19
C3832 _309_/a_761_289# _078_ 0.0257f
C3833 _064_ _275_/a_81_21# 1.27e-19
C3834 _259_/a_27_297# net50 0.0102f
C3835 _259_/a_109_297# trim_mask\[3\] 0.0193f
C3836 _323_/a_1283_21# _149_/a_68_297# 0.00781f
C3837 _326_/a_761_289# _310_/a_193_47# 6.88e-21
C3838 _326_/a_27_47# _310_/a_543_47# 6.4e-21
C3839 _326_/a_543_47# _310_/a_27_47# 9.08e-19
C3840 _078_ _205_/a_27_47# 0.0386f
C3841 trim[0] _112_ 1.79e-20
C3842 VPWR _310_/a_448_47# 0.08f
C3843 _037_ _298_/a_292_297# 0.00106f
C3844 _038_ _091_ 1.84e-20
C3845 _325_/a_1108_47# _074_ 7.48e-19
C3846 _025_ _336_/a_1108_47# 6.48e-20
C3847 _265_/a_81_21# net40 1.62e-20
C3848 input2/a_27_47# trimb[4] 0.00219f
C3849 _333_/a_761_289# _055_ 2.51e-21
C3850 net24 net13 2.64e-19
C3851 clknet_0_clk _089_ 2.95e-21
C3852 _041_ _035_ 0.126f
C3853 _035_ _338_/a_1182_261# 1.83e-21
C3854 clkbuf_2_1__f_clk/a_110_47# _017_ 0.0101f
C3855 _078_ _040_ 0.00184f
C3856 output32/a_27_47# _333_/a_1283_21# 9.15e-19
C3857 _338_/a_1224_47# _122_ 1.73e-19
C3858 _341_/a_448_47# _122_ 3.67e-19
C3859 _116_ _117_ 0.224f
C3860 _321_/a_761_289# _101_ 0.0432f
C3861 _321_/a_27_47# net52 0.0211f
C3862 _306_/a_193_47# net51 0.00189f
C3863 _134_ clkc 2.48e-19
C3864 _338_/a_1602_47# net18 7.99e-19
C3865 cal_count\[1\] _289_/a_68_297# 0.145f
C3866 _324_/a_805_47# _021_ 7.78e-20
C3867 _303_/a_1217_47# _070_ 6.83e-20
C3868 _262_/a_27_47# _062_ 3.41e-21
C3869 cal_itt\[1\] _203_/a_59_75# 5.31e-20
C3870 output18/a_27_47# net18 0.172f
C3871 clknet_2_1__leaf_clk _156_/a_27_47# 5.37e-20
C3872 _171_/a_27_47# _108_ 1.1e-19
C3873 _125_ output40/a_27_47# 0.0129f
C3874 net54 _049_ 0.392f
C3875 _302_/a_373_47# _038_ 1.97e-19
C3876 trim_mask\[4\] net40 0.00108f
C3877 _060_ _318_/a_193_47# 9.79e-21
C3878 _307_/a_1108_47# _004_ 5.47e-21
C3879 _307_/a_651_413# _079_ 4.5e-20
C3880 net50 trim_mask\[1\] 0.191f
C3881 _311_/a_193_47# net26 0.555f
C3882 net28 _313_/a_448_47# 0.0249f
C3883 output39/a_27_47# net39 0.203f
C3884 VPWR _247_/a_27_297# 0.26f
C3885 result[0] _004_ 0.00119f
C3886 _322_/a_1283_21# _078_ 0.0128f
C3887 _259_/a_27_297# _330_/a_1108_47# 3.98e-19
C3888 _074_ _314_/a_193_47# 0.00484f
C3889 _187_/a_27_413# net46 3.5e-19
C3890 clk input4/a_27_47# 0.00296f
C3891 net27 net15 0.008f
C3892 _074_ mask\[1\] 0.0263f
C3893 _329_/a_27_47# trim_mask\[3\] 0.00556f
C3894 net3 _243_/a_109_47# 8.21e-21
C3895 _331_/a_27_47# _331_/a_761_289# 0.0623f
C3896 _339_/a_1182_261# _122_ 2.09e-19
C3897 _023_ net14 0.0179f
C3898 _254_/a_109_297# _048_ 0.0011f
C3899 _053_ _227_/a_209_311# 6.7e-20
C3900 _245_/a_27_297# _245_/a_373_47# 0.0134f
C3901 VPWR _311_/a_1270_413# 4.91e-19
C3902 _268_/a_75_212# net46 0.0145f
C3903 VPWR result[5] 0.317f
C3904 _325_/a_193_47# _250_/a_27_297# 5.85e-20
C3905 calibrate _075_ 1.61e-20
C3906 _051_ clk 0.357f
C3907 net47 _338_/a_27_47# 0.101f
C3908 output24/a_27_47# result[3] 0.00182f
C3909 _258_/a_109_297# trim_mask\[0\] 3.49e-20
C3910 input1/a_75_212# _315_/a_27_47# 1.03e-21
C3911 _340_/a_1056_47# net47 0.00215f
C3912 _033_ trim_val\[4\] 5.22e-21
C3913 _325_/a_761_289# clknet_2_1__leaf_clk 6.93e-20
C3914 _311_/a_1270_413# net53 4.26e-20
C3915 net23 _078_ 0.0113f
C3916 input4/a_27_47# net4 0.109f
C3917 _319_/a_1283_21# en_co_clk 2.97e-21
C3918 _340_/a_476_47# _037_ 0.00265f
C3919 _319_/a_543_47# _120_ 1.27e-19
C3920 net31 net32 0.0992f
C3921 net43 net24 0.07f
C3922 _224_/a_113_297# net29 0.00958f
C3923 _340_/a_1032_413# _297_/a_285_47# 4.99e-20
C3924 _327_/a_543_47# _111_ 2.05e-19
C3925 wire42/a_75_212# _062_ 4.31e-19
C3926 VPWR output41/a_27_47# 0.437f
C3927 net19 net18 3.97e-19
C3928 _134_ _298_/a_215_47# 0.00196f
C3929 VPWR rebuffer6/a_27_47# 0.261f
C3930 _294_/a_68_297# net40 0.0078f
C3931 _301_/a_129_47# clknet_2_3__leaf_clk 0.0029f
C3932 _110_ _328_/a_761_289# 5.43e-20
C3933 net9 _178_/a_150_297# 6.58e-20
C3934 _167_/a_161_47# _090_ 8.23e-21
C3935 _051_ net4 0.324f
C3936 _097_ _281_/a_103_199# 3.28e-19
C3937 _337_/a_805_47# net44 0.0019f
C3938 _338_/a_1140_413# clknet_2_3__leaf_clk 9.56e-19
C3939 _291_/a_35_297# _127_ 0.37f
C3940 output41/a_27_47# valid 0.336f
C3941 _341_/a_761_289# clknet_2_3__leaf_clk 0.0701f
C3942 clknet_2_1__leaf_clk _077_ 2.07e-20
C3943 _233_/a_109_47# net1 0.00521f
C3944 _002_ _001_ 2.75e-20
C3945 trimb[0] trimb[2] 0.0503f
C3946 _024_ _038_ 0.00259f
C3947 net43 _313_/a_805_47# 0.00191f
C3948 rebuffer6/a_27_47# net53 0.12f
C3949 fanout46/a_27_47# _335_/a_27_47# 7.43e-20
C3950 _291_/a_285_297# net16 0.00445f
C3951 _276_/a_59_75# net19 5.08e-21
C3952 net2 rebuffer4/a_27_47# 0.0326f
C3953 VPWR _306_/a_761_289# 0.219f
C3954 _269_/a_81_21# _334_/a_543_47# 1.89e-20
C3955 VPWR _221_/a_109_297# 0.00572f
C3956 _034_ _282_/a_68_297# 1.49e-19
C3957 _340_/a_27_47# _339_/a_27_47# 3.88e-20
C3958 _187_/a_212_413# _332_/a_1108_47# 4.77e-20
C3959 net47 net17 1.8e-20
C3960 input1/a_75_212# clknet_2_0__leaf_clk 6.32e-20
C3961 _107_ net18 2.1e-20
C3962 _134_ _130_ 0.00574f
C3963 output22/a_27_47# _138_/a_27_47# 1.07e-20
C3964 _149_/a_68_297# _303_/a_543_47# 0.00374f
C3965 VPWR net29 1.12f
C3966 _294_/a_150_297# _299_/a_27_413# 1.95e-19
C3967 _029_ _332_/a_193_47# 0.218f
C3968 _195_/a_505_21# _065_ 2.68e-19
C3969 _051_ _063_ 7.4e-20
C3970 _316_/a_1283_21# _095_ 4.44e-20
C3971 net45 _137_/a_150_297# 1.59e-19
C3972 output38/a_27_47# net38 0.215f
C3973 _291_/a_35_297# _126_ 0.00393f
C3974 _144_/a_27_47# _339_/a_27_47# 1.08e-19
C3975 cal_itt\[2\] _065_ 0.00575f
C3976 fanout44/a_27_47# _319_/a_193_47# 1.05e-19
C3977 clk _331_/a_639_47# 0.00121f
C3978 _185_/a_68_297# _243_/a_27_297# 8.18e-19
C3979 net51 net30 8.47e-20
C3980 _058_ _269_/a_81_21# 3.09e-19
C3981 _323_/a_761_289# net47 0.166f
C3982 _339_/a_27_47# clknet_2_3__leaf_clk 0.22f
C3983 _314_/a_651_413# _011_ 0.00105f
C3984 _312_/a_27_47# net20 0.0263f
C3985 net28 _010_ 0.0643f
C3986 _136_ _301_/a_377_297# 0.00188f
C3987 _141_/a_27_47# clknet_2_0__leaf_clk 3.11e-19
C3988 _306_/a_543_47# _306_/a_651_413# 0.0572f
C3989 _306_/a_761_289# _306_/a_1270_413# 2.6e-19
C3990 _306_/a_193_47# _306_/a_639_47# 2.28e-19
C3991 cal_itt\[1\] _305_/a_1108_47# 3.79e-21
C3992 _076_ _202_/a_297_47# 6.01e-21
C3993 VPWR _227_/a_209_311# 0.2f
C3994 _221_/a_109_297# _009_ 0.0113f
C3995 _341_/a_193_47# _136_ 0.0113f
C3996 _235_/a_79_21# _235_/a_382_297# 0.00145f
C3997 cal_itt\[2\] _105_ 9.08e-20
C3998 net12 _089_ 0.0146f
C3999 _331_/a_1108_47# _331_/a_1270_413# 0.00645f
C4000 _331_/a_761_289# _331_/a_1217_47# 4.2e-19
C4001 _331_/a_543_47# _331_/a_805_47# 0.00171f
C4002 _339_/a_1296_47# _122_ 9.69e-20
C4003 net15 _317_/a_27_47# 0.0147f
C4004 _331_/a_193_47# _260_/a_93_21# 5.77e-21
C4005 _097_ _048_ 0.0686f
C4006 _010_ _158_/a_68_297# 2.42e-19
C4007 _326_/a_27_47# net15 6.55e-22
C4008 _325_/a_543_47# mask\[6\] 0.0357f
C4009 _083_ _078_ 0.147f
C4010 _015_ clk 0.0298f
C4011 _256_/a_109_47# trim_mask\[4\] 2.05e-19
C4012 net12 _312_/a_193_47# 8.37e-19
C4013 _325_/a_639_47# _042_ 1.01e-19
C4014 _306_/a_27_47# _049_ 8.61e-19
C4015 _041_ _338_/a_1182_261# 8.03e-20
C4016 net47 _338_/a_586_47# 0.00227f
C4017 _308_/a_1283_21# _138_/a_27_47# 5.15e-19
C4018 _308_/a_761_289# net14 0.0137f
C4019 _338_/a_27_47# _338_/a_562_413# 0.0018f
C4020 _338_/a_193_47# _338_/a_381_47# 0.152f
C4021 _338_/a_476_47# _338_/a_1032_413# 0.00329f
C4022 VPWR _317_/a_761_289# 0.216f
C4023 VPWR _326_/a_761_289# 0.217f
C4024 _328_/a_27_47# _328_/a_193_47# 0.578f
C4025 net9 en_co_clk 0.0171f
C4026 _258_/a_27_297# trim_mask\[2\] 0.172f
C4027 trim_mask\[2\] _024_ 3e-21
C4028 VPWR ctln[4] 0.193f
C4029 net13 _321_/a_193_47# 1.73e-20
C4030 cal _315_/a_651_413# 5.19e-19
C4031 _023_ net52 6.2e-21
C4032 net54 state\[1\] 0.201f
C4033 _229_/a_27_297# _090_ 0.159f
C4034 state\[2\] _331_/a_27_47# 1.55e-21
C4035 net13 _337_/a_193_47# 0.0177f
C4036 _228_/a_79_21# _100_ 0.0112f
C4037 _293_/a_81_21# _299_/a_27_413# 9.18e-21
C4038 trim_mask\[0\] net19 0.287f
C4039 output31/a_27_47# net34 0.0251f
C4040 VPWR _286_/a_505_21# 0.149f
C4041 _078_ _208_/a_218_374# 4.08e-19
C4042 _134_ cal_count\[3\] 0.0058f
C4043 _015_ net4 0.0171f
C4044 net31 output32/a_27_47# 0.00233f
C4045 _056_ net46 4.84e-20
C4046 _325_/a_193_47# _313_/a_193_47# 1.55e-20
C4047 _325_/a_27_47# _313_/a_761_289# 4.52e-22
C4048 net51 _072_ 2.5e-20
C4049 _259_/a_27_297# _335_/a_1108_47# 0.00164f
C4050 _259_/a_109_297# _335_/a_1283_21# 3.4e-19
C4051 _341_/a_1270_413# cal_count\[3\] 4.21e-19
C4052 net44 _312_/a_193_47# 0.0322f
C4053 _237_/a_76_199# fanout45/a_27_47# 2.12e-21
C4054 _033_ _330_/a_193_47# 4.32e-20
C4055 _135_ _332_/a_761_289# 3.35e-21
C4056 _336_/a_27_47# net46 0.296f
C4057 _192_/a_174_21# net41 2.35e-21
C4058 _303_/a_27_47# clknet_2_3__leaf_clk 0.851f
C4059 _323_/a_761_289# net44 0.00124f
C4060 _298_/a_215_47# cal_count\[2\] 0.072f
C4061 _298_/a_78_199# _131_ 0.00179f
C4062 _230_/a_59_75# _092_ 0.0421f
C4063 net47 _339_/a_193_47# 0.207f
C4064 net31 clkc 0.146f
C4065 _305_/a_193_47# net51 0.00359f
C4066 _257_/a_109_297# net18 0.0056f
C4067 _101_ net21 3.33e-21
C4068 net52 _046_ 1.65e-19
C4069 _321_/a_193_47# _248_/a_109_297# 2.5e-19
C4070 _062_ _206_/a_27_93# 0.00558f
C4071 trim_val\[2\] _334_/a_27_47# 2.46e-19
C4072 VPWR _296_/a_113_47# 4.45e-20
C4073 ctlp[1] _085_ 0.0037f
C4074 _323_/a_27_47# _323_/a_193_47# 0.9f
C4075 _340_/a_1602_47# _339_/a_1032_413# 1.29e-19
C4076 trim_mask\[0\] _107_ 0.0667f
C4077 _303_/a_1108_47# _035_ 7.31e-20
C4078 _266_/a_68_297# _266_/a_150_297# 0.00477f
C4079 _092_ _098_ 0.0892f
C4080 trim_mask\[0\] _333_/a_1108_47# 3.4e-19
C4081 _029_ _332_/a_1462_47# 6.53e-22
C4082 VPWR _318_/a_1108_47# 0.309f
C4083 _052_ clone1/a_27_47# 4.47e-19
C4084 _119_ _028_ 2.08e-20
C4085 _280_/a_75_212# trim_mask\[4\] 2.45e-20
C4086 _042_ _310_/a_193_47# 2.53e-20
C4087 _190_/a_655_47# clkbuf_2_3__f_clk/a_110_47# 2.98e-21
C4088 _169_/a_215_311# _100_ 3.01e-21
C4089 _060_ _243_/a_373_47# 0.0045f
C4090 net43 _321_/a_193_47# 0.0461f
C4091 _312_/a_1217_47# net20 8.49e-20
C4092 net24 _080_ 0.0117f
C4093 trim_mask\[1\] _335_/a_1108_47# 3.39e-21
C4094 _130_ cal_count\[2\] 0.15f
C4095 clknet_0_clk _092_ 0.206f
C4096 clknet_2_1__leaf_clk _310_/a_1108_47# 0.0679f
C4097 _047_ _109_ 6.2e-21
C4098 _104_ _027_ 0.146f
C4099 net43 _337_/a_193_47# 3.14e-20
C4100 _341_/a_1462_47# _136_ 1.99e-19
C4101 _301_/a_47_47# _301_/a_285_47# 0.0175f
C4102 _331_/a_651_413# _028_ 0.00136f
C4103 _331_/a_543_47# trim_mask\[4\] 3.65e-19
C4104 _110_ _109_ 0.126f
C4105 net15 _317_/a_1217_47# 2.97e-20
C4106 _292_/a_215_47# _133_ 1.3e-20
C4107 net33 rebuffer2/a_75_212# 1.19e-19
C4108 _317_/a_193_47# _317_/a_639_47# 2.28e-19
C4109 _317_/a_761_289# _317_/a_1270_413# 2.6e-19
C4110 _317_/a_543_47# _317_/a_651_413# 0.0572f
C4111 net9 _334_/a_193_47# 0.00121f
C4112 _328_/a_761_289# clknet_2_2__leaf_clk 0.0443f
C4113 en_co_clk clone7/a_27_47# 0.00156f
C4114 output14/a_27_47# _074_ 1.54e-19
C4115 _258_/a_109_297# trim_mask\[4\] 0.00592f
C4116 trim_mask\[1\] rebuffer2/a_75_212# 1.16e-20
C4117 _332_/a_1283_21# net33 5.11e-20
C4118 _326_/a_543_47# _326_/a_651_413# 0.0572f
C4119 _326_/a_761_289# _326_/a_1270_413# 2.6e-19
C4120 _326_/a_193_47# _326_/a_639_47# 2.28e-19
C4121 _216_/a_113_297# _078_ 0.0784f
C4122 _107_ _191_/a_27_297# 9.44e-19
C4123 _337_/a_27_47# _034_ 0.139f
C4124 _263_/a_382_297# _263_/a_297_47# 8.13e-19
C4125 net49 _108_ 0.119f
C4126 _338_/a_1182_261# _338_/a_1296_47# 1.84e-19
C4127 _338_/a_1032_413# _338_/a_1224_47# 0.00536f
C4128 _341_/a_27_47# _341_/a_543_47# 0.111f
C4129 _341_/a_193_47# _341_/a_761_289# 0.169f
C4130 _328_/a_761_289# _328_/a_805_47# 3.69e-19
C4131 _328_/a_193_47# _328_/a_1217_47# 2.36e-20
C4132 _328_/a_543_47# _328_/a_639_47# 0.0138f
C4133 _059_ clknet_2_0__leaf_clk 2.05e-19
C4134 _336_/a_543_47# _108_ 4.04e-19
C4135 _320_/a_448_47# net44 5.91e-20
C4136 net13 _321_/a_1462_47# 2.3e-19
C4137 _341_/a_1283_21# _037_ 9.46e-20
C4138 net47 _303_/a_193_47# 0.032f
C4139 net18 _118_ 1.71e-19
C4140 trim_mask\[0\] _279_/a_27_47# 0.028f
C4141 rebuffer4/a_27_47# _070_ 5.08e-20
C4142 net46 _173_/a_27_47# 5.03e-19
C4143 _313_/a_448_47# _085_ 1.78e-19
C4144 _094_ _192_/a_174_21# 4.06e-19
C4145 _308_/a_27_47# _016_ 2.75e-21
C4146 _340_/a_1032_413# cal_count\[2\] 0.0129f
C4147 cal_itt\[1\] _069_ 0.208f
C4148 _318_/a_27_47# _318_/a_1108_47# 0.102f
C4149 _318_/a_193_47# _318_/a_1283_21# 0.0424f
C4150 _318_/a_761_289# _318_/a_543_47# 0.21f
C4151 VPWR _150_/a_27_47# 0.246f
C4152 net27 _250_/a_27_297# 8.68e-19
C4153 _064_ _335_/a_1270_413# 6.72e-20
C4154 net48 net46 9.52e-19
C4155 net44 _312_/a_1462_47# 0.00288f
C4156 _110_ _279_/a_490_47# 1.61e-20
C4157 _312_/a_193_47# _312_/a_639_47# 2.28e-19
C4158 _312_/a_761_289# _312_/a_1270_413# 2.6e-19
C4159 _312_/a_543_47# _312_/a_651_413# 0.0572f
C4160 _309_/a_1283_21# _245_/a_27_297# 1.68e-20
C4161 _336_/a_1217_47# net46 2.95e-19
C4162 _309_/a_1108_47# _143_/a_68_297# 1.04e-20
C4163 calibrate _170_/a_81_21# 0.0066f
C4164 VPWR _305_/a_761_289# 0.22f
C4165 _320_/a_651_413# net52 1.67e-19
C4166 _306_/a_1108_47# clknet_2_0__leaf_clk 6.95e-20
C4167 _306_/a_543_47# net45 1e-21
C4168 result[6] net14 4.91e-20
C4169 _329_/a_1270_413# net46 3.67e-19
C4170 _195_/a_218_47# _067_ 1.53e-20
C4171 _050_ clone7/a_27_47# 5.91e-21
C4172 _048_ _240_/a_109_297# 3.92e-19
C4173 _078_ _314_/a_761_289# 0.00156f
C4174 _068_ _202_/a_297_47# 2.69e-19
C4175 net8 _057_ 0.159f
C4176 _323_/a_1283_21# net19 0.00502f
C4177 _041_ _339_/a_1032_413# 0.044f
C4178 net47 _339_/a_796_47# 7.37e-19
C4179 _025_ net18 0.00262f
C4180 _303_/a_1108_47# _198_/a_27_47# 5.29e-21
C4181 _192_/a_174_21# _192_/a_505_280# 0.145f
C4182 trim_val\[2\] _334_/a_1217_47# 1.34e-19
C4183 _309_/a_27_47# _023_ 1.73e-22
C4184 _323_/a_761_289# _323_/a_805_47# 3.69e-19
C4185 _323_/a_193_47# _323_/a_1217_47# 2.36e-20
C4186 _323_/a_543_47# _323_/a_639_47# 0.0138f
C4187 net31 _130_ 0.00142f
C4188 state\[2\] _242_/a_297_47# 0.00228f
C4189 output22/a_27_47# _307_/a_193_47# 2.18e-19
C4190 VPWR _315_/a_1270_413# 5.74e-19
C4191 _058_ net32 0.00353f
C4192 _306_/a_805_47# cal_itt\[3\] 1.57e-19
C4193 _107_ _090_ 0.00633f
C4194 _106_ _088_ 3.91e-20
C4195 _122_ en_co_clk 0.465f
C4196 _064_ _053_ 0.0826f
C4197 _329_/a_27_47# _031_ 8.51e-20
C4198 _233_/a_27_297# _233_/a_373_47# 0.0134f
C4199 _048_ clkbuf_2_2__f_clk/a_110_47# 3.38e-21
C4200 VPWR clkbuf_2_0__f_clk/a_110_47# 1.3f
C4201 _003_ rebuffer5/a_161_47# 2.29e-19
C4202 _306_/a_543_47# _065_ 2.85e-21
C4203 net16 _334_/a_1217_47# 6.83e-21
C4204 _315_/a_1270_413# valid 2.99e-20
C4205 _308_/a_639_47# _006_ 1.56e-20
C4206 clkbuf_0_clk/a_110_47# _190_/a_655_47# 0.00389f
C4207 _074_ net26 1.16f
C4208 net12 _152_/a_68_297# 4.73e-20
C4209 _128_ _340_/a_1032_413# 0.0117f
C4210 _036_ _340_/a_193_47# 1.63e-19
C4211 state\[0\] _096_ 2.01e-19
C4212 _326_/a_193_47# _086_ 0.00579f
C4213 clkbuf_2_2__f_clk/a_110_47# _330_/a_27_47# 0.0293f
C4214 _303_/a_193_47# net44 0.00334f
C4215 _306_/a_1283_21# _305_/a_448_47# 3.74e-19
C4216 _049_ cal_itt\[3\] 2.9e-21
C4217 en_co_clk _299_/a_27_413# 1.69e-19
C4218 net43 _321_/a_1462_47# 0.00288f
C4219 _326_/a_1283_21# _074_ 5.88e-20
C4220 _320_/a_1283_21# _320_/a_1108_47# 0.234f
C4221 _320_/a_761_289# _320_/a_651_413# 0.0977f
C4222 _320_/a_543_47# _320_/a_448_47# 0.0498f
C4223 _320_/a_27_47# _320_/a_639_47# 3.82e-19
C4224 _320_/a_193_47# _320_/a_1270_413# 1.46e-19
C4225 _119_ _279_/a_314_297# 0.0111f
C4226 _001_ _298_/a_78_199# 9.76e-20
C4227 _107_ _242_/a_382_297# 3.55e-19
C4228 _309_/a_193_47# _006_ 0.252f
C4229 _323_/a_27_47# _303_/a_27_47# 1.62e-20
C4230 _309_/a_543_47# _081_ 6.06e-19
C4231 _033_ _335_/a_193_47# 6.71e-22
C4232 _227_/a_209_311# wire42/a_75_212# 7.99e-20
C4233 _168_/a_297_47# _052_ 0.00101f
C4234 result[2] _007_ 4.52e-19
C4235 cal_count\[3\] trim_val\[4\] 1.44e-20
C4236 ctlp[0] _011_ 4.62e-19
C4237 _228_/a_297_47# clone7/a_27_47# 3.22e-20
C4238 trim_mask\[4\] _260_/a_256_47# 4.14e-20
C4239 _237_/a_218_374# _090_ 1.53e-19
C4240 _306_/a_193_47# clknet_2_1__leaf_clk 1.45e-19
C4241 net47 _092_ 0.0024f
C4242 _305_/a_27_47# _049_ 5.51e-20
C4243 _317_/a_1283_21# _014_ 1.29e-20
C4244 _317_/a_1108_47# clknet_2_0__leaf_clk 0.0701f
C4245 _317_/a_27_47# state\[1\] 1.28e-19
C4246 _317_/a_543_47# net45 0.153f
C4247 _308_/a_761_289# _307_/a_543_47# 7.82e-20
C4248 _308_/a_27_47# _307_/a_1108_47# 4.25e-21
C4249 _308_/a_543_47# _307_/a_761_289# 2.14e-20
C4250 _308_/a_1108_47# _307_/a_27_47# 3.02e-20
C4251 output27/a_27_47# result[7] 0.00234f
C4252 _262_/a_109_297# net30 1.47e-19
C4253 result[0] _308_/a_27_47# 0.00211f
C4254 net16 comp 3e-20
C4255 net44 _152_/a_68_297# 0.00258f
C4256 _232_/a_32_297# net41 4.77e-21
C4257 _050_ _073_ 3.44e-20
C4258 net13 _090_ 0.0117f
C4259 _303_/a_761_289# _063_ 7.96e-20
C4260 _106_ _108_ 0.174f
C4261 mask\[6\] _247_/a_27_297# 1.11e-20
C4262 _303_/a_1108_47# _041_ 4.03e-20
C4263 net47 _303_/a_1462_47# 0.00392f
C4264 _134_ _265_/a_299_297# 7.39e-21
C4265 _304_/a_1283_21# en_co_clk 6.54e-20
C4266 trim_mask\[0\] _118_ 0.202f
C4267 trim_mask\[4\] net19 0.00699f
C4268 _010_ _085_ 0.19f
C4269 _333_/a_27_47# _333_/a_448_47# 0.0864f
C4270 _333_/a_193_47# _333_/a_1108_47# 0.125f
C4271 _268_/a_75_212# _111_ 0.19f
C4272 net23 _245_/a_109_47# 0.00378f
C4273 net16 _332_/a_1270_413# 1.39e-19
C4274 net46 _172_/a_68_297# 0.00178f
C4275 _318_/a_1108_47# _318_/a_1217_47# 0.00742f
C4276 _318_/a_1283_21# _318_/a_1462_47# 0.0074f
C4277 clknet_2_0__leaf_clk _192_/a_27_47# 3.69e-20
C4278 net12 _092_ 0.00962f
C4279 _297_/a_377_297# cal_count\[2\] 5.95e-20
C4280 _078_ _311_/a_27_47# 2.01e-19
C4281 _104_ _032_ 3.44e-21
C4282 _309_/a_651_413# _101_ 1.95e-20
C4283 _324_/a_651_413# net44 0.0154f
C4284 _324_/a_27_47# _312_/a_1108_47# 7.23e-19
C4285 _324_/a_193_47# _312_/a_1283_21# 1.08e-19
C4286 _048_ _337_/a_543_47# 5.1e-21
C4287 VPWR _251_/a_109_297# 0.181f
C4288 VPWR _250_/a_373_47# 7.67e-19
C4289 _248_/a_27_297# net21 8.05e-21
C4290 _185_/a_68_297# _316_/a_1108_47# 3.02e-20
C4291 _308_/a_543_47# _308_/a_651_413# 0.0572f
C4292 _308_/a_761_289# _308_/a_1270_413# 2.6e-19
C4293 _308_/a_193_47# _308_/a_639_47# 2.28e-19
C4294 net33 trimb[4] 3.24e-19
C4295 trim_mask\[2\] _257_/a_27_297# 0.0648f
C4296 _324_/a_1108_47# _323_/a_193_47# 7.71e-20
C4297 _025_ trim_mask\[0\] 0.00129f
C4298 _107_ trim_mask\[4\] 0.0049f
C4299 VPWR _042_ 6.5f
C4300 net3 _337_/a_193_47# 6.11e-19
C4301 net15 _319_/a_1283_21# 8.76e-19
C4302 _087_ _095_ 3.83e-20
C4303 _307_/a_27_47# _307_/a_1217_47# 2.56e-19
C4304 _307_/a_761_289# _307_/a_639_47# 3.16e-19
C4305 _326_/a_193_47# clknet_2_1__leaf_clk 0.0253f
C4306 clknet_2_0__leaf_clk _315_/a_27_47# 0.271f
C4307 _101_ _045_ 7.28e-21
C4308 VPWR _064_ 0.74f
C4309 _200_/a_80_21# _230_/a_59_75# 0.0212f
C4310 _249_/a_109_297# _101_ 0.0106f
C4311 result[0] _307_/a_448_47# 6.73e-19
C4312 _290_/a_27_413# trimb[4] 9.58e-19
C4313 _191_/a_27_297# _118_ 7.13e-19
C4314 VPWR _319_/a_448_47# 0.0846f
C4315 _250_/a_373_47# net53 0.00193f
C4316 _322_/a_448_47# net44 7.6e-19
C4317 trim[3] net34 0.0749f
C4318 _318_/a_448_47# net45 2.45e-19
C4319 net27 _313_/a_193_47# 5.06e-22
C4320 net44 _092_ 7.09e-20
C4321 _309_/a_27_47# _308_/a_761_289# 3.48e-21
C4322 _309_/a_193_47# _308_/a_193_47# 1.43e-21
C4323 input3/a_75_212# net14 0.00162f
C4324 _233_/a_109_47# _012_ 3.65e-20
C4325 _109_ clknet_2_2__leaf_clk 0.00148f
C4326 _042_ net53 0.369f
C4327 _104_ net41 1.28e-20
C4328 cal_count\[0\] _132_ 8.08e-21
C4329 _091_ en_co_clk 0.00219f
C4330 _182_/a_27_47# net34 3.82e-22
C4331 net12 _008_ 0.00728f
C4332 output29/a_27_47# net29 0.173f
C4333 VPWR _100_ 0.397f
C4334 _325_/a_193_47# _321_/a_543_47# 8.89e-21
C4335 _188_/a_27_47# net35 1.73e-19
C4336 output32/a_27_47# _058_ 0.0029f
C4337 net24 _310_/a_448_47# 2.92e-21
C4338 _306_/a_1283_21# _002_ 2.36e-19
C4339 _320_/a_193_47# _283_/a_75_212# 5.64e-21
C4340 _187_/a_27_413# _135_ 0.00107f
C4341 _103_ _060_ 8.17e-21
C4342 _337_/a_1283_21# en_co_clk 0.125f
C4343 net55 net41 9.56e-19
C4344 _303_/a_543_47# net19 0.0109f
C4345 _291_/a_35_297# net47 8.66e-20
C4346 _094_ _232_/a_32_297# 1.95e-21
C4347 _108_ _278_/a_109_297# 1.2e-19
C4348 _042_ _009_ 5.83e-21
C4349 _192_/a_174_21# _243_/a_27_297# 4.67e-19
C4350 cal _316_/a_27_47# 8.2e-19
C4351 _200_/a_80_21# clknet_0_clk 4.96e-19
C4352 _270_/a_59_75# rebuffer2/a_75_212# 3.49e-20
C4353 net12 mask\[5\] 0.318f
C4354 mask\[4\] _101_ 0.366f
C4355 _339_/a_652_21# _339_/a_562_413# 9.35e-20
C4356 _339_/a_1182_261# _339_/a_1602_47# 0.144f
C4357 _339_/a_476_47# _339_/a_381_47# 0.0356f
C4358 net34 net37 2.05f
C4359 net13 _320_/a_1270_413# 1.5e-19
C4360 _081_ _246_/a_27_297# 2.76e-19
C4361 net5 net37 0.00267f
C4362 _263_/a_79_21# _092_ 0.00326f
C4363 mask\[6\] net29 6.37e-19
C4364 _341_/a_27_47# _092_ 0.00324f
C4365 _317_/a_1217_47# state\[1\] 1.2e-19
C4366 _008_ net44 0.00112f
C4367 _320_/a_1108_47# _040_ 0.0346f
C4368 output13/a_27_47# net13 0.241f
C4369 _315_/a_761_289# _315_/a_639_47# 3.16e-19
C4370 _315_/a_27_47# _315_/a_1217_47# 2.56e-19
C4371 output22/a_27_47# _005_ 1.31e-20
C4372 _337_/a_543_47# _076_ 1.22e-19
C4373 trim_mask\[4\] _279_/a_27_47# 0.0227f
C4374 VPWR _336_/a_805_47# 2.92e-19
C4375 VPWR _264_/a_27_297# 0.651f
C4376 clk input3/a_75_212# 0.00131f
C4377 _117_ net50 9.65e-19
C4378 _104_ _171_/a_27_47# 0.0483f
C4379 VPWR _329_/a_651_413# 0.145f
C4380 net4 _199_/a_193_297# 4.24e-19
C4381 net8 _334_/a_1270_413# 1.46e-19
C4382 trim_mask\[2\] trim_val\[4\] 0.00455f
C4383 _319_/a_1283_21# _049_ 0.00262f
C4384 _116_ _057_ 6.5e-20
C4385 _078_ _247_/a_373_47# 1.2e-20
C4386 clknet_2_1__leaf_clk net30 2.02e-20
C4387 net24 _247_/a_27_297# 5.06e-20
C4388 net50 _136_ 0.00145f
C4389 _312_/a_448_47# _045_ 2.21e-19
C4390 net44 mask\[5\] 0.0328f
C4391 _062_ net18 2.2e-19
C4392 net20 _084_ 0.00131f
C4393 _335_/a_27_47# clkbuf_2_2__f_clk/a_110_47# 9.57e-20
C4394 _050_ _337_/a_1283_21# 0.00416f
C4395 _002_ net26 4.53e-21
C4396 net55 _171_/a_27_47# 4.04e-19
C4397 _286_/a_439_47# _123_ 0.00504f
C4398 _331_/a_193_47# _330_/a_27_47# 0.00133f
C4399 _331_/a_27_47# _330_/a_193_47# 0.00133f
C4400 _074_ _315_/a_805_47# 6.43e-19
C4401 calibrate _315_/a_639_47# 2.29e-19
C4402 net54 _240_/a_109_297# 1.28e-21
C4403 trim_val\[0\] _109_ 0.00388f
C4404 _012_ _315_/a_448_47# 0.16f
C4405 _326_/a_761_289# mask\[6\] 2.18e-21
C4406 fanout44/a_27_47# _337_/a_193_47# 4.94e-20
C4407 _257_/a_109_297# trim_mask\[4\] 0.0018f
C4408 clkbuf_2_0__f_clk/a_110_47# _093_ 2.69e-21
C4409 VPWR _022_ 0.439f
C4410 state\[0\] _316_/a_761_289# 2.3e-19
C4411 _308_/a_543_47# net43 0.156f
C4412 _308_/a_27_47# net23 2.87e-19
C4413 _308_/a_1283_21# _005_ 4.73e-20
C4414 _328_/a_1283_21# _025_ 6.78e-21
C4415 clknet_2_0__leaf_clk _315_/a_1217_47# 2.56e-19
C4416 VPWR ctln[3] 0.189f
C4417 net45 _315_/a_639_47# 9.54e-19
C4418 clkbuf_2_1__f_clk/a_110_47# net45 0.158f
C4419 _020_ _101_ 0.00744f
C4420 _094_ net55 0.323f
C4421 net50 _119_ 0.00107f
C4422 _019_ net44 5.55e-19
C4423 trimb[2] net39 0.00735f
C4424 _305_/a_543_47# _065_ 3.64e-20
C4425 _327_/a_761_289# net18 7.42e-19
C4426 _327_/a_27_47# _256_/a_27_297# 5.24e-19
C4427 ctln[2] _108_ 1.05e-19
C4428 comp net40 2.43e-19
C4429 _097_ _317_/a_27_47# 4.22e-21
C4430 _321_/a_543_47# mask\[3\] 2.36e-20
C4431 clknet_2_1__leaf_clk _072_ 1.55e-20
C4432 _305_/a_543_47# _305_/a_651_413# 0.0572f
C4433 _305_/a_761_289# _305_/a_1270_413# 2.6e-19
C4434 _305_/a_193_47# _305_/a_639_47# 2.28e-19
C4435 net12 _208_/a_218_47# 1.76e-19
C4436 VPWR _313_/a_1283_21# 0.374f
C4437 _309_/a_761_289# _309_/a_543_47# 0.21f
C4438 _309_/a_193_47# _309_/a_1283_21# 0.0424f
C4439 _309_/a_27_47# _309_/a_1108_47# 0.102f
C4440 clkbuf_2_1__f_clk/a_110_47# _065_ 6.09e-19
C4441 _324_/a_1108_47# _303_/a_27_47# 1.54e-20
C4442 net37 _133_ 2.9e-20
C4443 _305_/a_193_47# clknet_2_1__leaf_clk 9.3e-19
C4444 _241_/a_105_352# _241_/a_297_47# 0.00424f
C4445 _232_/a_32_297# _014_ 1.2e-20
C4446 _071_ clknet_0_clk 0.0306f
C4447 _269_/a_299_297# _269_/a_384_47# 1.48e-19
C4448 _030_ net33 1.44e-20
C4449 _030_ trim_mask\[1\] 0.104f
C4450 _113_ net49 0.0029f
C4451 _234_/a_109_297# net15 0.00108f
C4452 _293_/a_299_297# _339_/a_1032_413# 4.14e-20
C4453 cal_itt\[1\] _304_/a_639_47# 1.4e-19
C4454 _210_/a_113_297# net30 0.0281f
C4455 _050_ _331_/a_761_289# 0.00234f
C4456 clkbuf_2_1__f_clk/a_110_47# _319_/a_27_47# 0.0219f
C4457 trim_mask\[4\] _118_ 0.0192f
C4458 comp _299_/a_215_297# 3.56e-19
C4459 _324_/a_1283_21# _152_/a_68_297# 0.00189f
C4460 _325_/a_27_47# _101_ 0.00168f
C4461 cal_count\[1\] _339_/a_193_47# 6.28e-20
C4462 _036_ _339_/a_27_47# 0.145f
C4463 _128_ _339_/a_1182_261# 0.0153f
C4464 en_co_clk _101_ 0.00249f
C4465 _119_ _330_/a_1108_47# 7.31e-20
C4466 net44 _017_ 2.51e-19
C4467 clkbuf_2_0__f_clk/a_110_47# _319_/a_193_47# 5.02e-20
C4468 net51 _003_ 0.00476f
C4469 cal_itt\[3\] _202_/a_297_47# 1.98e-21
C4470 _058_ _302_/a_109_297# 0.00122f
C4471 _279_/a_314_297# _279_/a_206_47# 5.08e-20
C4472 net21 _156_/a_27_47# 1.65e-19
C4473 _303_/a_193_47# _303_/a_639_47# 2.28e-19
C4474 _303_/a_761_289# _303_/a_1270_413# 2.6e-19
C4475 _303_/a_543_47# _303_/a_651_413# 0.0572f
C4476 _048_ _260_/a_93_21# 4.7e-21
C4477 trim_mask\[0\] _062_ 0.245f
C4478 _325_/a_448_47# mask\[7\] 5.89e-20
C4479 mask\[7\] _216_/a_113_297# 1.54e-19
C4480 _253_/a_299_297# mask\[3\] 1.23e-21
C4481 _087_ _226_/a_27_47# 0.0764f
C4482 _237_/a_218_47# _092_ 9.49e-19
C4483 _237_/a_439_47# _099_ 0.00174f
C4484 _292_/a_78_199# _292_/a_292_297# 0.013f
C4485 net54 _337_/a_543_47# 1.26e-21
C4486 cal_itt\[1\] _261_/a_113_47# 2.8e-20
C4487 _290_/a_207_413# net2 1.2e-19
C4488 _094_ mask\[0\] 0.0519f
C4489 _314_/a_1108_47# net14 0.00242f
C4490 _322_/a_1108_47# _205_/a_27_47# 0.00157f
C4491 _169_/a_109_53# _167_/a_161_47# 3.05e-19
C4492 VPWR _316_/a_193_47# 0.613f
C4493 _041_ _076_ 0.0928f
C4494 net3 _090_ 0.0948f
C4495 _025_ trim_mask\[4\] 0.016f
C4496 _326_/a_1108_47# _078_ 0.00364f
C4497 _051_ _075_ 0.15f
C4498 _324_/a_27_47# _324_/a_1217_47# 2.56e-19
C4499 _324_/a_761_289# _324_/a_639_47# 3.16e-19
C4500 _259_/a_27_297# trim_mask\[1\] 6.42e-20
C4501 calibrate _096_ 0.00876f
C4502 _306_/a_543_47# _204_/a_75_212# 3.36e-19
C4503 _103_ _227_/a_109_93# 0.0392f
C4504 _316_/a_193_47# valid 8.33e-20
C4505 _316_/a_543_47# net41 0.0356f
C4506 _237_/a_76_199# _281_/a_103_199# 4.52e-20
C4507 ctlp[7] _155_/a_68_297# 0.00111f
C4508 _232_/a_32_297# _243_/a_27_297# 0.0115f
C4509 net42 calibrate 3.11e-19
C4510 _047_ net46 6.63e-19
C4511 mask\[1\] _245_/a_373_47# 9.32e-19
C4512 _341_/a_543_47# _001_ 2.66e-19
C4513 net43 _283_/a_75_212# 0.0336f
C4514 net16 _132_ 4.18e-20
C4515 net45 _096_ 1.24e-19
C4516 _189_/a_408_47# clone1/a_27_47# 1.76e-20
C4517 _309_/a_448_47# net43 2.79e-19
C4518 net14 _310_/a_193_47# 0.0102f
C4519 _058_ cal_count\[3\] 0.00167f
C4520 _116_ _027_ 1.29e-20
C4521 _110_ net46 0.393f
C4522 _324_/a_193_47# mask\[4\] 1.34e-20
C4523 _327_/a_761_289# trim_mask\[0\] 7.95e-19
C4524 _033_ net30 2.25e-21
C4525 _002_ net2 0.0574f
C4526 mask\[7\] _314_/a_761_289# 2.25e-19
C4527 _191_/a_27_297# _062_ 0.125f
C4528 _305_/a_1283_21# _002_ 0.00336f
C4529 net2 _289_/a_68_297# 0.183f
C4530 _250_/a_27_297# _250_/a_109_297# 0.171f
C4531 net9 _300_/a_129_47# 4.46e-19
C4532 _309_/a_1283_21# _309_/a_1462_47# 0.0074f
C4533 _309_/a_1108_47# _309_/a_1217_47# 0.00742f
C4534 _152_/a_68_297# _044_ 0.109f
C4535 _232_/a_32_297# _232_/a_220_297# 0.00132f
C4536 trim[1] trim[4] 0.0419f
C4537 _190_/a_215_47# _190_/a_655_47# 0.0234f
C4538 _321_/a_193_47# _247_/a_27_297# 1.24e-19
C4539 _321_/a_27_47# _247_/a_109_297# 3.77e-20
C4540 ctlp[1] _074_ 5.89e-19
C4541 _322_/a_1283_21# _322_/a_1108_47# 0.234f
C4542 _322_/a_761_289# _322_/a_651_413# 0.0977f
C4543 _322_/a_543_47# _322_/a_448_47# 0.0498f
C4544 _322_/a_27_47# _322_/a_639_47# 0.00188f
C4545 _322_/a_193_47# _322_/a_1270_413# 1.46e-19
C4546 _248_/a_27_297# mask\[4\] 0.0892f
C4547 _322_/a_27_47# mask\[4\] 5.48e-19
C4548 _110_ _327_/a_651_413# 6.5e-21
C4549 _095_ _099_ 0.0338f
C4550 _065_ _096_ 2.11e-19
C4551 _251_/a_27_297# clknet_2_1__leaf_clk 0.0348f
C4552 trim_mask\[1\] net33 2.41e-19
C4553 _320_/a_543_47# _017_ 5.03e-19
C4554 _320_/a_448_47# mask\[2\] 1.38e-19
C4555 _272_/a_299_297# _056_ 9.9e-20
C4556 _332_/a_1108_47# clknet_2_3__leaf_clk 1.88e-21
C4557 _169_/a_215_311# clk 2.62e-20
C4558 trim_val\[1\] net49 0.115f
C4559 net22 _315_/a_761_289# 9.38e-20
C4560 _078_ _315_/a_27_47# 6.64e-20
C4561 VPWR net34 1.22f
C4562 _259_/a_373_47# _064_ 8.77e-19
C4563 _259_/a_109_297# _104_ 0.0106f
C4564 _253_/a_299_297# _310_/a_1283_21# 2.28e-19
C4565 _253_/a_81_21# _310_/a_1108_47# 4.33e-19
C4566 VPWR net5 0.48f
C4567 _327_/a_1108_47# _136_ 0.00119f
C4568 trim_mask\[1\] _336_/a_761_289# 4.87e-20
C4569 _200_/a_209_297# _063_ 0.0069f
C4570 _336_/a_27_47# _336_/a_1283_21# 0.0436f
C4571 _336_/a_193_47# _336_/a_543_47# 0.224f
C4572 cal_itt\[0\] _338_/a_27_47# 0.00494f
C4573 _040_ _246_/a_27_297# 0.0849f
C4574 _050_ _260_/a_250_297# 0.00209f
C4575 _314_/a_27_47# _046_ 6.7e-21
C4576 _006_ mask\[1\] 3.35e-19
C4577 _319_/a_761_289# _319_/a_1108_47# 0.0512f
C4578 _319_/a_27_47# _319_/a_651_413# 9.73e-19
C4579 _319_/a_193_47# _319_/a_448_47# 0.0612f
C4580 _138_/a_27_47# _039_ 0.194f
C4581 _305_/a_1108_47# _069_ 3.66e-20
C4582 _134_ en_co_clk 0.0584f
C4583 net25 _101_ 1.56e-20
C4584 net16 _269_/a_81_21# 0.00875f
C4585 VPWR _149_/a_150_297# 0.00228f
C4586 net42 _105_ 0.00141f
C4587 _237_/a_76_199# _048_ 0.0676f
C4588 _128_ _339_/a_1296_47# 3.98e-19
C4589 mask\[3\] _041_ 8.1e-20
C4590 _110_ _335_/a_651_413# 7.89e-21
C4591 trim_mask\[0\] _332_/a_193_47# 0.00645f
C4592 _293_/a_81_21# _293_/a_384_47# 0.00138f
C4593 _273_/a_59_75# _334_/a_27_47# 0.00722f
C4594 _058_ _038_ 0.00111f
C4595 ctlp[7] net43 1.17e-19
C4596 calibrate net22 1.75e-20
C4597 _169_/a_215_311# net4 0.0528f
C4598 _303_/a_1283_21# _000_ 9.79e-21
C4599 _074_ mask\[0\] 1.13e-20
C4600 _293_/a_81_21# _128_ 3.86e-19
C4601 VPWR _299_/a_298_297# 0.195f
C4602 _243_/a_109_297# _096_ 0.016f
C4603 _243_/a_27_297# net55 0.149f
C4604 _243_/a_109_47# _100_ 4.58e-19
C4605 _103_ _054_ 5.3e-21
C4606 _219_/a_109_297# mask\[4\] 4.12e-19
C4607 output24/a_27_47# _074_ 0.0126f
C4608 _324_/a_1283_21# mask\[5\] 0.0652f
C4609 _324_/a_193_47# _020_ 3.29e-20
C4610 _103_ net30 0.102f
C4611 state\[2\] _050_ 0.711f
C4612 _317_/a_1108_47# _316_/a_1283_21# 3.54e-22
C4613 _292_/a_493_297# cal_count\[1\] 0.00124f
C4614 _292_/a_292_297# _036_ 0.00106f
C4615 _337_/a_1108_47# net51 5.9e-20
C4616 _119_ _052_ 2.32e-21
C4617 _028_ _330_/a_448_47# 1.13e-20
C4618 clknet_2_2__leaf_clk _330_/a_651_413# 0.00252f
C4619 _331_/a_448_47# _027_ 9.25e-21
C4620 _161_/a_68_297# net34 0.0078f
C4621 VPWR _316_/a_1462_47# 6.13e-20
C4622 net22 net45 0.156f
C4623 output15/a_27_47# _251_/a_27_297# 7.82e-21
C4624 _078_ clknet_2_0__leaf_clk 0.006f
C4625 _017_ _209_/a_27_47# 7.14e-22
C4626 ctln[1] net15 0.00218f
C4627 _064_ _336_/a_1108_47# 1.31e-19
C4628 _104_ _336_/a_543_47# 0.0247f
C4629 _237_/a_505_21# en_co_clk 5.93e-19
C4630 _232_/a_304_297# _096_ 3.87e-19
C4631 _232_/a_220_297# net55 7.38e-19
C4632 _289_/a_68_297# _123_ 6.19e-21
C4633 _329_/a_27_47# _104_ 1.59e-19
C4634 _330_/a_639_47# net19 8.45e-19
C4635 trim_mask\[2\] _334_/a_543_47# 2.23e-19
C4636 VPWR _304_/a_448_47# 0.0846f
C4637 _049_ _073_ 6.44e-20
C4638 _335_/a_1108_47# _119_ 1.34e-21
C4639 _328_/a_27_47# _327_/a_448_47# 9.89e-21
C4640 _094_ _121_ 0.0342f
C4641 _087_ _052_ 3.07e-19
C4642 _089_ _088_ 5.01e-19
C4643 net22 _065_ 8.97e-21
C4644 _071_ net44 2.38e-20
C4645 trim[2] _176_/a_27_47# 8.02e-19
C4646 _164_/a_161_47# _099_ 6.81e-20
C4647 output33/a_27_47# net33 0.251f
C4648 net23 _246_/a_27_297# 5.34e-20
C4649 _200_/a_209_47# net19 6.7e-19
C4650 _304_/a_761_289# _286_/a_76_199# 9.16e-22
C4651 _251_/a_109_297# mask\[6\] 0.00335f
C4652 mask\[6\] _250_/a_373_47# 0.00163f
C4653 _250_/a_27_297# _021_ 0.119f
C4654 output23/a_27_47# output24/a_27_47# 0.0217f
C4655 output31/a_27_47# trim[0] 0.337f
C4656 state\[2\] _228_/a_297_47# 3.69e-19
C4657 _239_/a_694_21# net55 1.38e-19
C4658 mask\[6\] _042_ 1.95e-19
C4659 _308_/a_193_47# mask\[1\] 6.5e-20
C4660 _146_/a_68_297# _078_ 5.82e-19
C4661 _321_/a_27_47# _018_ 0.285f
C4662 _301_/a_47_47# net46 3.11e-20
C4663 _328_/a_1108_47# _058_ 0.00215f
C4664 trim_mask\[2\] _058_ 0.00127f
C4665 _309_/a_1283_21# mask\[2\] 1.21e-20
C4666 _322_/a_543_47# _019_ 3.53e-19
C4667 _019_ _248_/a_373_47# 1.97e-19
C4668 _239_/a_27_297# net42 0.00125f
C4669 VPWR _133_ 1.11f
C4670 _030_ _270_/a_59_75# 3.44e-19
C4671 _113_ _270_/a_145_75# 0.00141f
C4672 trim_mask\[2\] _335_/a_193_47# 1.44e-20
C4673 _341_/a_27_47# net46 0.296f
C4674 net14 _224_/a_113_297# 5.51e-19
C4675 _078_ _315_/a_1217_47# 6.12e-20
C4676 _121_ _192_/a_505_280# 9.37e-20
C4677 _053_ clk 0.00574f
C4678 _237_/a_505_21# _050_ 0.00133f
C4679 _272_/a_299_297# net48 0.0911f
C4680 _272_/a_81_21# _114_ 0.118f
C4681 mask\[5\] _044_ 0.162f
C4682 _274_/a_75_212# net46 0.0272f
C4683 net12 state\[0\] 1.7e-20
C4684 _284_/a_68_297# rebuffer3/a_75_212# 2.15e-21
C4685 _041_ _068_ 0.0507f
C4686 _320_/a_448_47# mask\[1\] 0.0111f
C4687 _200_/a_209_47# _107_ 1.42e-19
C4688 _336_/a_448_47# _336_/a_639_47# 4.61e-19
C4689 _322_/a_1108_47# _083_ 0.00198f
C4690 _000_ mask\[4\] 3.63e-20
C4691 _004_ _315_/a_27_47# 1.61e-20
C4692 cal_itt\[0\] _341_/a_543_47# 5.19e-21
C4693 _336_/a_1108_47# _264_/a_27_297# 1.59e-20
C4694 _336_/a_193_47# _106_ 7.03e-20
C4695 ctln[4] net18 0.00336f
C4696 net44 _311_/a_761_289# 0.165f
C4697 _107_ _228_/a_382_297# 2.25e-19
C4698 _290_/a_297_47# _127_ 8.17e-20
C4699 VPWR _256_/a_373_47# 1.35e-19
C4700 _249_/a_373_47# _020_ 0.00133f
C4701 _116_ _032_ 0.0668f
C4702 _093_ _316_/a_193_47# 6.32e-20
C4703 calibrate _316_/a_761_289# 6.54e-20
C4704 trim_mask\[0\] _332_/a_1462_47# 0.00222f
C4705 _329_/a_1283_21# _329_/a_1108_47# 0.234f
C4706 _329_/a_761_289# _329_/a_651_413# 0.0977f
C4707 _329_/a_543_47# _329_/a_448_47# 0.0498f
C4708 _329_/a_27_47# _329_/a_639_47# 0.00188f
C4709 _329_/a_193_47# _329_/a_1270_413# 1.46e-19
C4710 VPWR _321_/a_448_47# 0.0842f
C4711 trim_mask\[4\] _062_ 1.19e-20
C4712 _231_/a_161_47# _092_ 0.368f
C4713 _124_ _122_ 0.00765f
C4714 clkbuf_2_1__f_clk/a_110_47# _282_/a_68_297# 1.45e-21
C4715 net5 _300_/a_47_47# 7.07e-21
C4716 clknet_2_1__leaf_clk _313_/a_543_47# 0.0347f
C4717 net43 _222_/a_113_297# 1.63e-19
C4718 _053_ net4 1.21f
C4719 _156_/a_27_47# _045_ 0.197f
C4720 _306_/a_193_47# clkbuf_0_clk/a_110_47# 2.77e-19
C4721 _284_/a_68_297# _065_ 0.164f
C4722 VPWR _337_/a_448_47# 0.083f
C4723 _236_/a_109_297# _095_ 5.38e-19
C4724 _132_ net40 0.201f
C4725 _286_/a_505_21# net18 4.43e-19
C4726 en_co_clk cal_count\[2\] 1.66e-19
C4727 _110_ output10/a_27_47# 4.1e-20
C4728 clknet_2_0__leaf_clk _316_/a_1283_21# 3.04e-21
C4729 _014_ _316_/a_543_47# 0.0124f
C4730 net45 _316_/a_761_289# 0.165f
C4731 _002_ _067_ 1.66e-21
C4732 _002_ _070_ 9.91e-19
C4733 _028_ _027_ 0.00438f
C4734 clknet_2_2__leaf_clk net46 0.838f
C4735 state\[1\] clone7/a_27_47# 0.214f
C4736 state\[2\] _169_/a_301_53# 1.57e-21
C4737 VPWR net14 1.38f
C4738 _322_/a_448_47# mask\[2\] 0.00264f
C4739 net43 rebuffer5/a_161_47# 0.0504f
C4740 _058_ _333_/a_761_289# 6.41e-19
C4741 _328_/a_805_47# net46 0.00371f
C4742 _128_ _291_/a_285_47# 0.00206f
C4743 cal_count\[1\] _291_/a_35_297# 4.78e-21
C4744 clkbuf_2_3__f_clk/a_110_47# net30 0.00182f
C4745 _058_ _265_/a_299_297# 0.00973f
C4746 _290_/a_297_47# _126_ 1.43e-19
C4747 net14 valid 0.00598f
C4748 fanout45/a_27_47# _317_/a_27_47# 9.76e-20
C4749 _329_/a_1283_21# net9 3.47e-19
C4750 _104_ _106_ 0.00183f
C4751 _309_/a_543_47# _216_/a_113_297# 2.12e-19
C4752 _079_ net45 0.004f
C4753 _004_ clknet_2_0__leaf_clk 0.107f
C4754 _074_ _010_ 0.0801f
C4755 _327_/a_651_413# clknet_2_2__leaf_clk 9.04e-19
C4756 VPWR _143_/a_68_297# 0.168f
C4757 _061_ clkc 4.9e-19
C4758 _226_/a_27_47# _099_ 2.83e-19
C4759 _325_/a_805_47# net13 1.81e-19
C4760 _299_/a_215_297# _132_ 0.00272f
C4761 _326_/a_193_47# _253_/a_81_21# 2.09e-19
C4762 _326_/a_27_47# _253_/a_299_297# 9.57e-19
C4763 _053_ _063_ 0.696f
C4764 VPWR _340_/a_956_413# 0.00403f
C4765 _106_ net55 0.00408f
C4766 _333_/a_543_47# rebuffer1/a_75_212# 3.33e-19
C4767 _333_/a_193_47# _332_/a_193_47# 5.9e-22
C4768 _275_/a_81_21# trim_val\[3\] 0.185f
C4769 _041_ _125_ 0.0167f
C4770 _053_ _037_ 0.00216f
C4771 mask\[6\] _022_ 0.0576f
C4772 _265_/a_81_21# _332_/a_193_47# 0.00351f
C4773 _320_/a_1108_47# _141_/a_27_47# 2e-19
C4774 _337_/a_1283_21# _049_ 0.0176f
C4775 _179_/a_27_47# _056_ 6.48e-19
C4776 _176_/a_27_47# _055_ 3.12e-22
C4777 net52 _310_/a_1462_47# 5.5e-20
C4778 net43 _212_/a_113_297# 0.00838f
C4779 net49 _172_/a_150_297# 3.05e-19
C4780 _289_/a_150_297# _126_ 4.96e-19
C4781 VPWR clk 4.31f
C4782 trim_mask\[0\] _227_/a_209_311# 0.228f
C4783 net24 _042_ 1.88e-19
C4784 _048_ _281_/a_103_199# 0.017f
C4785 _341_/a_1217_47# net46 4.13e-19
C4786 _246_/a_109_297# mask\[2\] 0.0456f
C4787 net16 net32 1.21e-20
C4788 mask\[0\] _319_/a_805_47# 0.00218f
C4789 _309_/a_1283_21# mask\[1\] 0.00327f
C4790 _333_/a_651_413# net46 0.0122f
C4791 clk valid 5.35e-20
C4792 calibrate _098_ 0.382f
C4793 VPWR _277_/a_75_212# 0.261f
C4794 net31 en_co_clk 2.05e-20
C4795 _307_/a_193_47# _039_ 0.00143f
C4796 VPWR _331_/a_1283_21# 0.391f
C4797 _286_/a_439_47# clknet_2_3__leaf_clk 3.34e-19
C4798 trim_val\[0\] net46 0.00414f
C4799 _051_ _227_/a_296_53# 1.93e-20
C4800 _332_/a_448_47# clknet_2_2__leaf_clk 0.00155f
C4801 mask\[6\] _313_/a_1283_21# 1.6e-20
C4802 output25/a_27_47# _007_ 0.0163f
C4803 ctln[5] net19 0.00146f
C4804 _062_ _190_/a_27_47# 2.48e-19
C4805 _199_/a_109_297# _001_ 0.0121f
C4806 net27 _312_/a_1108_47# 0.00276f
C4807 _053_ _260_/a_346_47# 8.87e-19
C4808 cal_itt\[0\] _303_/a_193_47# 3.26e-19
C4809 _311_/a_1283_21# net19 0.00189f
C4810 _300_/a_47_47# _133_ 4.7e-21
C4811 _329_/a_543_47# _026_ 0.00195f
C4812 VPWR net4 4.23f
C4813 net13 _169_/a_109_53# 0.00396f
C4814 net28 _314_/a_761_289# 0.00719f
C4815 result[6] _314_/a_27_47# 0.00742f
C4816 _059_ _087_ 6.38e-19
C4817 _309_/a_193_47# _310_/a_27_47# 6.43e-21
C4818 _309_/a_27_47# _310_/a_193_47# 0.00127f
C4819 calibrate clknet_0_clk 1.42e-19
C4820 _281_/a_253_297# en_co_clk 0.00324f
C4821 _327_/a_1283_21# _109_ 1.29e-19
C4822 _281_/a_103_199# _120_ 0.0845f
C4823 net18 _150_/a_27_47# 0.111f
C4824 net12 _306_/a_651_413# 0.00178f
C4825 _325_/a_805_47# net43 0.00192f
C4826 cal_count\[0\] _130_ 7.12e-22
C4827 net45 clknet_0_clk 0.0745f
C4828 _313_/a_193_47# _313_/a_761_289# 0.176f
C4829 _313_/a_27_47# _313_/a_543_47# 0.106f
C4830 _019_ mask\[2\] 0.3f
C4831 clk _318_/a_27_47# 0.0539f
C4832 clkbuf_0_clk/a_110_47# net30 0.00164f
C4833 cal_count\[3\] net30 0.00416f
C4834 net15 _101_ 0.749f
C4835 output37/a_27_47# output40/a_27_47# 0.00222f
C4836 _309_/a_448_47# _082_ 1.16e-19
C4837 clknet_2_1__leaf_clk _003_ 3.91e-19
C4838 _102_ net26 0.408f
C4839 VPWR net52 1.43f
C4840 _308_/a_1108_47# fanout43/a_27_47# 0.00423f
C4841 net8 _272_/a_81_21# 0.00281f
C4842 VPWR _063_ 2.18f
C4843 _185_/a_68_297# _092_ 5.9e-22
C4844 VPWR _338_/a_381_47# 0.104f
C4845 _306_/a_651_413# net44 0.013f
C4846 _059_ _263_/a_297_47# 0.0535f
C4847 _326_/a_1108_47# mask\[7\] 0.0223f
C4848 _326_/a_543_47# _023_ 0.00115f
C4849 _326_/a_1283_21# _102_ 0.00375f
C4850 VPWR _037_ 1.06f
C4851 clknet_0_clk _065_ 0.288f
C4852 VPWR _273_/a_145_75# 5.67e-19
C4853 _325_/a_1108_47# mask\[5\] 1.74e-20
C4854 net4 _318_/a_27_47# 5.02e-19
C4855 _213_/a_109_297# _080_ 0.00379f
C4856 net50 _057_ 8.88e-20
C4857 _050_ _281_/a_253_297# 3.07e-19
C4858 _286_/a_76_199# _338_/a_476_47# 0.00437f
C4859 _109_ _108_ 0.00222f
C4860 _304_/a_651_413# _065_ 9.08e-20
C4861 clk _317_/a_1270_413# 8.78e-20
C4862 net43 _314_/a_448_47# 2.56e-19
C4863 _340_/a_1032_413# cal_count\[0\] 2.03e-20
C4864 clknet_0_clk _105_ 0.0125f
C4865 _315_/a_543_47# net14 0.00521f
C4866 _187_/a_297_47# _136_ 1.17e-19
C4867 trim[1] net49 1.86e-19
C4868 _110_ _111_ 0.00413f
C4869 _320_/a_27_47# net15 4.44e-21
C4870 _048_ _120_ 0.0423f
C4871 _123_ _298_/a_78_199# 0.094f
C4872 mask\[2\] _017_ 0.0217f
C4873 _319_/a_27_47# clknet_0_clk 0.00149f
C4874 cal_itt\[0\] _092_ 0.0807f
C4875 output20/a_27_47# net21 4.43e-21
C4876 fanout47/a_27_47# _069_ 0.0024f
C4877 clkbuf_0_clk/a_110_47# _072_ 0.0135f
C4878 VPWR _320_/a_761_289# 0.206f
C4879 _052_ _099_ 1.41e-19
C4880 _088_ _092_ 6.57e-20
C4881 mask\[1\] _246_/a_109_297# 0.00164f
C4882 VPWR _260_/a_346_47# 1.94e-19
C4883 net43 _310_/a_761_289# 0.174f
C4884 _325_/a_1108_47# _019_ 2.67e-19
C4885 _322_/a_805_47# mask\[3\] 4.33e-20
C4886 net4 _317_/a_1270_413# 1.46e-19
C4887 net22 _282_/a_68_297# 1.48e-20
C4888 output25/a_27_47# result[4] 0.0022f
C4889 result[3] output26/a_27_47# 1.88e-20
C4890 VPWR _328_/a_639_47# 3.07e-19
C4891 _101_ _049_ 0.00159f
C4892 _078_ _313_/a_651_413# 4.99e-19
C4893 cal_itt\[0\] _303_/a_1462_47# 5.1e-19
C4894 _093_ net14 0.0132f
C4895 ctlp[6] net44 2.53e-19
C4896 _324_/a_193_47# _311_/a_1108_47# 7.02e-21
C4897 _324_/a_761_289# _311_/a_1283_21# 5.29e-20
C4898 _048_ _076_ 1.71e-19
C4899 _324_/a_27_47# net27 2.02e-19
C4900 _210_/a_113_297# sample 3.8e-19
C4901 mask\[0\] output30/a_27_47# 2.42e-21
C4902 net13 net51 4.16e-20
C4903 _305_/a_193_47# clkbuf_0_clk/a_110_47# 0.00157f
C4904 _125_ _339_/a_1032_413# 1.43e-20
C4905 _337_/a_651_413# net45 6.88e-20
C4906 _108_ _279_/a_490_47# 0.0194f
C4907 _323_/a_761_289# net26 3.76e-20
C4908 _239_/a_474_297# _003_ 7.81e-21
C4909 _325_/a_27_47# _325_/a_761_289# 0.0701f
C4910 _053_ _279_/a_396_47# 0.00233f
C4911 net16 clkc 3e-20
C4912 VPWR _312_/a_1270_413# 7.19e-19
C4913 _061_ cal_count\[3\] 5.28e-20
C4914 VPWR _307_/a_543_47# 0.207f
C4915 VPWR _323_/a_639_47# 7.45e-19
C4916 _226_/a_27_47# _226_/a_109_47# 0.00578f
C4917 _239_/a_27_297# _098_ 0.00811f
C4918 _068_ _190_/a_465_47# 0.00437f
C4919 _080_ _212_/a_113_297# 0.0993f
C4920 VPWR output38/a_27_47# 0.445f
C4921 _074_ net20 0.00949f
C4922 net12 _318_/a_805_47# 1.31e-19
C4923 _042_ net18 0.169f
C4924 net45 _245_/a_27_297# 0.0631f
C4925 _326_/a_1270_413# net52 5.26e-21
C4926 _019_ mask\[1\] 2.67e-20
C4927 _321_/a_193_47# _042_ 0.00809f
C4928 _092_ _108_ 7.49e-20
C4929 _064_ net18 0.0288f
C4930 cal_itt\[0\] _199_/a_109_297# 4.74e-19
C4931 _260_/a_250_297# _049_ 0.033f
C4932 _321_/a_1108_47# clknet_2_1__leaf_clk 0.00232f
C4933 _028_ _171_/a_27_47# 4.32e-20
C4934 _258_/a_27_297# fanout46/a_27_47# 2.53e-20
C4935 VPWR _333_/a_448_47# 0.1f
C4936 net12 calibrate 0.0079f
C4937 _340_/a_652_21# _123_ 0.0316f
C4938 _275_/a_81_21# _335_/a_543_47# 0.0059f
C4939 _189_/a_27_47# _051_ 0.114f
C4940 cal_count\[0\] _338_/a_476_47# 0.00994f
C4941 _330_/a_761_289# _330_/a_639_47# 3.16e-19
C4942 _330_/a_27_47# _330_/a_1217_47# 2.56e-19
C4943 _143_/a_150_297# _065_ 8.49e-22
C4944 net47 _065_ 0.453f
C4945 calibrate _331_/a_1108_47# 7.33e-19
C4946 trim_mask\[4\] _227_/a_209_311# 8.9e-21
C4947 _074_ _081_ 0.0746f
C4948 VPWR _308_/a_1270_413# 8.34e-19
C4949 _066_ clkbuf_2_3__f_clk/a_110_47# 5.74e-19
C4950 _337_/a_27_47# _096_ 0.00163f
C4951 state\[2\] _049_ 0.00628f
C4952 net12 net45 0.0673f
C4953 state\[2\] _318_/a_761_289# 0.00114f
C4954 _064_ _302_/a_27_297# 3.11e-19
C4955 _015_ _318_/a_448_47# 0.16f
C4956 clk wire42/a_75_212# 0.00295f
C4957 _305_/a_27_47# _041_ 1.2e-20
C4958 net43 net51 0.382f
C4959 _093_ net4 2.32e-20
C4960 _262_/a_27_47# _063_ 0.171f
C4961 _004_ _078_ 1.57e-20
C4962 VPWR _237_/a_535_374# 8.37e-19
C4963 VPWR _309_/a_27_47# 0.486f
C4964 net45 _331_/a_1108_47# 0.255f
C4965 VPWR _339_/a_562_413# 0.00343f
C4966 mask\[1\] _017_ 0.00371f
C4967 _328_/a_193_47# _030_ 0.0025f
C4968 mask\[7\] _146_/a_68_297# 2.69e-19
C4969 VPWR _155_/a_150_297# 0.00138f
C4970 net12 _065_ 0.0165f
C4971 net44 net45 0.00514f
C4972 VPWR _279_/a_396_47# 0.277f
C4973 net12 _305_/a_651_413# 3.15e-19
C4974 net50 _027_ 0.002f
C4975 _307_/a_1108_47# _094_ 3.31e-23
C4976 _325_/a_543_47# _325_/a_805_47# 0.00171f
C4977 _325_/a_761_289# _325_/a_1217_47# 4.2e-19
C4978 _325_/a_1108_47# _325_/a_1270_413# 0.00645f
C4979 trim_mask\[3\] net46 0.0635f
C4980 _259_/a_27_297# _119_ 4.94e-19
C4981 _216_/a_113_297# _216_/a_199_47# 2.42e-19
C4982 _335_/a_27_47# _330_/a_27_47# 9.7e-19
C4983 _110_ _112_ 0.251f
C4984 _110_ _272_/a_299_297# 1.47e-19
C4985 _051_ _336_/a_27_47# 5.67e-19
C4986 _293_/a_299_297# _125_ 0.00884f
C4987 output34/a_27_47# _334_/a_27_47# 4.36e-20
C4988 _110_ _336_/a_1283_21# 0.00565f
C4989 VPWR _324_/a_543_47# 0.214f
C4990 _136_ net33 3.56e-20
C4991 net16 _130_ 0.0061f
C4992 net43 _224_/a_199_47# 1.59e-19
C4993 _329_/a_193_47# _110_ 2.48e-19
C4994 calibrate _263_/a_79_21# 3.97e-19
C4995 _302_/a_109_297# _066_ 0.0697f
C4996 _226_/a_303_47# _075_ 0.00549f
C4997 _322_/a_27_47# net15 6.81e-20
C4998 net15 _241_/a_297_47# 0.00587f
C4999 net54 _048_ 0.0101f
C5000 VPWR _201_/a_113_47# 1.33e-19
C5001 output29/a_27_47# net14 0.0211f
C5002 net44 _065_ 0.752f
C5003 output39/a_27_47# net34 4.68e-19
C5004 _324_/a_543_47# net53 8.7e-19
C5005 _321_/a_193_47# _022_ 7.1e-19
C5006 _058_ en_co_clk 9.63e-19
C5007 _169_/a_109_53# net3 4.79e-20
C5008 _237_/a_505_21# _049_ 8.24e-19
C5009 _323_/a_1283_21# _150_/a_27_47# 2.18e-19
C5010 ctln[3] net18 2.83e-20
C5011 VPWR _322_/a_761_289# 0.214f
C5012 VPWR _248_/a_109_47# 4.34e-19
C5013 mask\[3\] _076_ 7.04e-19
C5014 _304_/a_27_47# _284_/a_68_297# 1.21e-20
C5015 VPWR _257_/a_109_47# 7.06e-20
C5016 _064_ trim_mask\[0\] 0.46f
C5017 _303_/a_193_47# net26 4.16e-20
C5018 _083_ _311_/a_193_47# 5.05e-19
C5019 _059_ _099_ 0.0305f
C5020 _305_/a_651_413# net44 0.00382f
C5021 VPWR output21/a_27_47# 0.455f
C5022 _341_/a_27_47# rebuffer3/a_75_212# 2.11e-19
C5023 _063_ wire42/a_75_212# 1.25e-20
C5024 _111_ clknet_2_2__leaf_clk 0.0731f
C5025 _095_ net41 4.84e-20
C5026 _338_/a_27_47# _123_ 0.0015f
C5027 net13 _318_/a_193_47# 0.0212f
C5028 _316_/a_193_47# _316_/a_651_413# 0.0346f
C5029 _316_/a_543_47# _316_/a_1108_47# 7.99e-20
C5030 _248_/a_109_47# net53 0.00321f
C5031 _322_/a_761_289# net53 4.45e-21
C5032 trim_mask\[0\] _100_ 1.03e-20
C5033 VPWR _303_/a_1270_413# 7.9e-19
C5034 mask\[6\] net14 4.06e-22
C5035 clkbuf_2_0__f_clk/a_110_47# _090_ 0.00855f
C5036 net50 _335_/a_448_47# 7.97e-20
C5037 net44 _319_/a_27_47# 3.16e-20
C5038 _308_/a_27_47# clknet_2_0__leaf_clk 0.266f
C5039 _340_/a_1032_413# net16 8.39e-19
C5040 _330_/a_1108_47# _027_ 0.0566f
C5041 _330_/a_1283_21# net46 0.336f
C5042 _301_/a_47_47# _135_ 0.398f
C5043 _301_/a_285_47# net2 3.31e-19
C5044 _060_ en_co_clk 0.00965f
C5045 _066_ cal_count\[3\] 0.139f
C5046 clk _202_/a_79_21# 1.37e-19
C5047 _307_/a_1108_47# _315_/a_193_47# 5.53e-21
C5048 _307_/a_193_47# _315_/a_1108_47# 5.53e-21
C5049 _341_/a_27_47# _065_ 0.0135f
C5050 _341_/a_27_47# _135_ 1.04e-20
C5051 _051_ _096_ 4.33e-21
C5052 _106_ clknet_2_3__leaf_clk 4.29e-19
C5053 _250_/a_27_297# _101_ 0.0912f
C5054 _306_/a_1283_21# _092_ 1.19e-19
C5055 clkc net40 1.65e-19
C5056 cal net3 0.00534f
C5057 _320_/a_543_47# net45 4.02e-20
C5058 _320_/a_1108_47# clknet_2_0__leaf_clk 1.96e-19
C5059 _107_ _262_/a_109_297# 0.00217f
C5060 VPWR _034_ 0.596f
C5061 net31 output40/a_27_47# 0.00659f
C5062 net42 _051_ 0.00681f
C5063 VPWR _309_/a_1217_47# 5.34e-19
C5064 net45 clknet_2_2__leaf_clk 0.00335f
C5065 net16 cal_count\[3\] 2.33e-19
C5066 clknet_2_2__leaf_clk rebuffer3/a_75_212# 9.57e-19
C5067 _064_ _191_/a_27_297# 0.195f
C5068 output20/a_27_47# _045_ 6.23e-19
C5069 _053_ _193_/a_109_297# 1.93e-19
C5070 _328_/a_193_47# trim_mask\[1\] 0.554f
C5071 _074_ _312_/a_805_47# 2.48e-21
C5072 _200_/a_80_21# cal_itt\[0\] 0.066f
C5073 _200_/a_209_297# cal_itt\[2\] 0.0327f
C5074 net12 _239_/a_27_297# 0.00146f
C5075 _319_/a_193_47# net52 8.1e-20
C5076 net4 _194_/a_199_47# 2.28e-19
C5077 _007_ mask\[3\] 1.14e-19
C5078 trim_mask\[0\] _264_/a_27_297# 5.26e-21
C5079 net4 _336_/a_1108_47# 0.00131f
C5080 _329_/a_27_47# _328_/a_27_47# 2.08e-20
C5081 _334_/a_193_47# _334_/a_543_47# 0.23f
C5082 _334_/a_27_47# _334_/a_1283_21# 0.0436f
C5083 _314_/a_27_47# _314_/a_1108_47# 0.102f
C5084 _314_/a_193_47# _314_/a_1283_21# 0.0424f
C5085 _314_/a_761_289# _314_/a_543_47# 0.21f
C5086 result[0] _074_ 0.0228f
C5087 _339_/a_1182_261# cal_count\[0\] 0.065f
C5088 _320_/a_543_47# _065_ 8.11e-20
C5089 _181_/a_68_297# net46 2.99e-19
C5090 net8 ctln[2] 0.00686f
C5091 fanout47/a_27_47# _287_/a_75_212# 1.92e-20
C5092 state\[0\] _166_/a_161_47# 2.4e-19
C5093 state\[2\] state\[1\] 0.204f
C5094 clknet_2_2__leaf_clk _065_ 0.00202f
C5095 _214_/a_113_297# clknet_2_1__leaf_clk 2.91e-20
C5096 _060_ _050_ 2.31e-19
C5097 _335_/a_448_47# _330_/a_1108_47# 2.39e-19
C5098 _197_/a_113_297# _063_ 0.0474f
C5099 _307_/a_448_47# clknet_2_0__leaf_clk 0.00107f
C5100 _307_/a_1283_21# net45 0.291f
C5101 net2 _339_/a_193_47# 4.56e-20
C5102 trim[3] _334_/a_1108_47# 4.32e-19
C5103 _111_ trim_val\[0\] 4.54e-20
C5104 _336_/a_543_47# _266_/a_68_297# 1.1e-20
C5105 _038_ _066_ 0.257f
C5106 _105_ clknet_2_2__leaf_clk 4.87e-20
C5107 _094_ _095_ 0.0016f
C5108 _259_/a_109_47# clknet_2_2__leaf_clk 3.13e-21
C5109 _164_/a_161_47# net41 1.53e-19
C5110 _320_/a_193_47# clknet_2_1__leaf_clk 1.11e-20
C5111 VPWR trim[0] 0.554f
C5112 _338_/a_27_47# _067_ 1.25e-19
C5113 _304_/a_543_47# _122_ 0.0129f
C5114 _333_/a_1283_21# _176_/a_27_47# 1.3e-19
C5115 _325_/a_193_47# net27 9.9e-20
C5116 _168_/a_27_413# _051_ 0.13f
C5117 _308_/a_805_47# _074_ 6.63e-19
C5118 _104_ _089_ 0.00112f
C5119 _274_/a_75_212# _112_ 4.98e-19
C5120 _182_/a_27_47# net35 0.11f
C5121 output22/a_27_47# result[1] 0.00288f
C5122 result[0] output23/a_27_47# 1.11e-20
C5123 ctln[7] _318_/a_805_47# 2.48e-20
C5124 net13 _318_/a_1462_47# 1.57e-19
C5125 _316_/a_761_289# _013_ 3.21e-20
C5126 _329_/a_193_47# _274_/a_75_212# 1.35e-19
C5127 _237_/a_535_374# _093_ 7.79e-20
C5128 _113_ _109_ 3.58e-19
C5129 _192_/a_174_21# _092_ 0.00143f
C5130 _192_/a_27_47# _099_ 3.79e-20
C5131 _323_/a_1283_21# _042_ 0.0354f
C5132 _192_/a_505_280# _095_ 0.0569f
C5133 net50 _032_ 0.0063f
C5134 VPWR _281_/a_253_47# 0.00365f
C5135 _089_ net55 3.16e-19
C5136 _090_ _100_ 0.179f
C5137 clknet_2_1__leaf_clk net19 5.46e-19
C5138 _065_ _209_/a_27_47# 0.0703f
C5139 _326_/a_639_47# net43 9.54e-19
C5140 _074_ _205_/a_27_47# 0.334f
C5141 _008_ net26 0.317f
C5142 net24 net14 0.00633f
C5143 _033_ _280_/a_75_212# 0.109f
C5144 _015_ _096_ 2.48e-19
C5145 _237_/a_505_21# state\[1\] 3.95e-20
C5146 mask\[6\] net52 0.201f
C5147 ctln[4] _275_/a_299_297# 0.00151f
C5148 output10/a_27_47# trim_mask\[3\] 0.0104f
C5149 net35 net37 0.0143f
C5150 net28 _225_/a_109_297# 3.5e-19
C5151 _309_/a_193_47# net45 2.05e-19
C5152 _059_ _236_/a_109_297# 4.7e-21
C5153 VPWR trim_val\[3\] 0.258f
C5154 _074_ _040_ 4.02e-21
C5155 VPWR _193_/a_109_297# 0.00563f
C5156 _303_/a_193_47# net2 1.18e-20
C5157 _304_/a_27_47# clknet_0_clk 1.69e-20
C5158 result[4] _007_ 7.64e-20
C5159 _334_/a_448_47# net46 0.0181f
C5160 net25 _310_/a_1108_47# 0.0523f
C5161 mask\[3\] _310_/a_1283_21# 0.00292f
C5162 _082_ _310_/a_761_289# 0.00213f
C5163 _112_ clknet_2_2__leaf_clk 0.00632f
C5164 VPWR _208_/a_76_199# 0.117f
C5165 _035_ _122_ 3.09e-20
C5166 _130_ net40 0.0102f
C5167 _315_/a_1108_47# _241_/a_297_47# 2e-20
C5168 _315_/a_27_47# _099_ 1.82e-20
C5169 net9 _041_ 0.00973f
C5170 net24 _143_/a_68_297# 0.105f
C5171 mask\[5\] net26 0.00797f
C5172 net9 _338_/a_1182_261# 0.0012f
C5173 _327_/a_1283_21# net46 0.294f
C5174 cal_itt\[1\] _195_/a_218_47# 1.04e-19
C5175 cal_itt\[0\] _195_/a_439_47# 7.96e-19
C5176 _336_/a_543_47# _028_ 4.82e-20
C5177 _336_/a_1283_21# clknet_2_2__leaf_clk 0.00137f
C5178 ctln[7] net45 3.98e-19
C5179 trim_mask\[2\] trim_val\[2\] 0.319f
C5180 cal_itt\[0\] _071_ 9.45e-19
C5181 result[1] _308_/a_1283_21# 1.68e-19
C5182 net34 _129_ 9.43e-20
C5183 _304_/a_193_47# _304_/a_448_47# 0.0604f
C5184 _304_/a_761_289# _304_/a_1108_47# 0.0512f
C5185 _304_/a_27_47# _304_/a_651_413# 9.73e-19
C5186 _329_/a_193_47# clknet_2_2__leaf_clk 0.00202f
C5187 mask\[7\] _078_ 0.362f
C5188 _258_/a_109_297# _033_ 6.44e-20
C5189 _162_/a_27_47# _055_ 1.54e-20
C5190 _339_/a_193_47# _123_ 0.017f
C5191 _190_/a_465_47# cal_itt\[3\] 8.18e-20
C5192 _149_/a_68_297# _043_ 0.105f
C5193 _334_/a_448_47# _334_/a_639_47# 4.61e-19
C5194 _314_/a_1108_47# _314_/a_1217_47# 0.00742f
C5195 _314_/a_1283_21# _314_/a_1462_47# 0.0074f
C5196 _329_/a_448_47# trim_mask\[2\] 8.76e-20
C5197 trim_mask\[2\] net16 0.0178f
C5198 _327_/a_761_289# _327_/a_639_47# 3.16e-19
C5199 _327_/a_27_47# _327_/a_1217_47# 2.56e-19
C5200 _336_/a_448_47# net19 0.00617f
C5201 _032_ _330_/a_1108_47# 0.00731f
C5202 _335_/a_1283_21# net46 0.367f
C5203 _281_/a_253_297# _049_ 3.38e-21
C5204 _322_/a_1283_21# _074_ 0.00292f
C5205 _288_/a_59_75# net37 0.00414f
C5206 _059_ _226_/a_109_47# 8.6e-21
C5207 state\[0\] _185_/a_68_297# 0.167f
C5208 _293_/a_81_21# cal_count\[0\] 0.115f
C5209 _306_/a_27_47# _076_ 0.0196f
C5210 net51 _062_ 7.83e-21
C5211 _299_/a_298_297# _129_ 0.0763f
C5212 _299_/a_215_297# _130_ 0.135f
C5213 _304_/a_193_47# _133_ 0.0012f
C5214 _019_ net26 6.44e-20
C5215 _266_/a_68_297# _106_ 0.149f
C5216 net27 _007_ 2.83e-20
C5217 _340_/a_1032_413# net40 8.48e-21
C5218 _333_/a_27_47# _173_/a_27_47# 1.35e-20
C5219 _327_/a_805_47# _058_ 4.69e-19
C5220 _322_/a_543_47# net45 4.28e-20
C5221 clknet_2_0__leaf_clk _099_ 3.7e-20
C5222 _014_ _095_ 0.123f
C5223 _064_ trim_mask\[4\] 0.254f
C5224 VPWR _330_/a_543_47# 0.21f
C5225 output24/a_27_47# _006_ 0.00974f
C5226 en_co_clk _227_/a_109_93# 2.05e-21
C5227 net46 _108_ 0.0945f
C5228 _332_/a_543_47# net46 0.183f
C5229 _328_/a_448_47# net9 5.07e-19
C5230 clkbuf_2_0__f_clk/a_110_47# _283_/a_75_212# 3.13e-21
C5231 net43 _086_ 0.011f
C5232 _304_/a_1283_21# _035_ 1.83e-21
C5233 _164_/a_161_47# _192_/a_505_280# 1.86e-20
C5234 _306_/a_193_47# _050_ 1.23e-21
C5235 net27 mask\[3\] 1.52e-20
C5236 net13 clknet_2_1__leaf_clk 7.95e-20
C5237 _336_/a_448_47# _107_ 5.02e-19
C5238 trim_val\[2\] _175_/a_150_297# 7.85e-19
C5239 net23 _074_ 0.211f
C5240 _112_ _333_/a_651_413# 8.3e-19
C5241 net49 _333_/a_1270_413# 1.1e-19
C5242 clknet_2_1__leaf_clk _155_/a_68_297# 0.0393f
C5243 _340_/a_1602_47# _122_ 0.00134f
C5244 _337_/a_27_47# clknet_0_clk 0.0239f
C5245 _115_ trim_val\[2\] 0.0012f
C5246 _235_/a_297_47# en_co_clk 0.00145f
C5247 _324_/a_193_47# _250_/a_27_297# 2.84e-19
C5248 cal_count\[3\] net40 0.412f
C5249 _298_/a_493_297# _133_ 9.81e-19
C5250 _310_/a_193_47# _310_/a_651_413# 0.0276f
C5251 _310_/a_543_47# _310_/a_1108_47# 7.99e-20
C5252 net13 _243_/a_373_47# 1.99e-19
C5253 output28/a_27_47# clknet_2_1__leaf_clk 0.0131f
C5254 clknet_2_3__leaf_clk _298_/a_78_199# 1.63e-19
C5255 _314_/a_27_47# _224_/a_113_297# 0.00106f
C5256 cal_itt\[2\] _053_ 3.35e-19
C5257 _093_ _034_ 1.2e-21
C5258 VPWR _325_/a_1283_21# 0.382f
C5259 fanout46/a_27_47# trim_val\[4\] 0.00159f
C5260 _239_/a_474_297# _107_ 0.00144f
C5261 net21 _313_/a_543_47# 0.00136f
C5262 _046_ _313_/a_1108_47# 6.99e-20
C5263 net16 _175_/a_150_297# 3.12e-19
C5264 _335_/a_761_289# _335_/a_639_47# 3.16e-19
C5265 _335_/a_27_47# _335_/a_1217_47# 2.56e-19
C5266 net16 _333_/a_761_289# 0.00842f
C5267 _324_/a_761_289# clknet_2_1__leaf_clk 4.73e-19
C5268 _115_ net16 0.013f
C5269 result[4] _310_/a_1283_21# 3.24e-19
C5270 net16 _265_/a_299_297# 0.00719f
C5271 _311_/a_27_47# _311_/a_193_47# 0.855f
C5272 net12 _204_/a_75_212# 0.00856f
C5273 _050_ _227_/a_109_93# 1.83e-20
C5274 _058_ _332_/a_639_47# 8.33e-19
C5275 _189_/a_218_47# _092_ 0.00259f
C5276 _031_ net46 0.438f
C5277 net24 net52 0.0116f
C5278 _322_/a_193_47# clknet_2_1__leaf_clk 0.00174f
C5279 clknet_2_1__leaf_clk _248_/a_109_297# 6.27e-22
C5280 _315_/a_1462_47# _095_ 1.1e-19
C5281 _315_/a_1217_47# _099_ 2.14e-20
C5282 clknet_2_0__leaf_clk _246_/a_27_297# 0.0312f
C5283 _129_ _133_ 0.108f
C5284 net9 _341_/a_651_413# 3.15e-19
C5285 _336_/a_805_47# trim_mask\[4\] 0.00213f
C5286 _264_/a_27_297# trim_mask\[4\] 5.68e-19
C5287 output23/a_27_47# net23 0.181f
C5288 _329_/a_1462_47# clknet_2_2__leaf_clk 4.85e-19
C5289 _304_/a_27_47# net47 0.301f
C5290 _243_/a_27_297# _095_ 8.62e-21
C5291 net43 _305_/a_639_47# 1.79e-19
C5292 _256_/a_27_297# _256_/a_109_297# 0.171f
C5293 _336_/a_543_47# _279_/a_314_297# 5.26e-20
C5294 _026_ trim_mask\[2\] 0.0595f
C5295 net16 _339_/a_1182_261# 8.18e-19
C5296 clk _316_/a_651_413# 1.11e-19
C5297 VPWR _314_/a_27_47# 0.459f
C5298 _308_/a_761_289# net22 1.74e-19
C5299 _308_/a_193_47# mask\[0\] 3.45e-20
C5300 _308_/a_27_47# _078_ 0.00772f
C5301 _332_/a_448_47# _108_ 0.0154f
C5302 _321_/a_193_47# _321_/a_448_47# 0.0604f
C5303 _321_/a_761_289# _321_/a_1108_47# 0.0512f
C5304 _321_/a_27_47# _321_/a_651_413# 9.73e-19
C5305 _332_/a_193_47# _332_/a_1270_413# 1.46e-19
C5306 _332_/a_27_47# _332_/a_639_47# 0.00188f
C5307 _332_/a_543_47# _332_/a_448_47# 0.0498f
C5308 _332_/a_761_289# _332_/a_651_413# 0.0977f
C5309 _332_/a_1283_21# _332_/a_1108_47# 0.234f
C5310 net24 _214_/a_199_47# 4.81e-19
C5311 _038_ net40 2.03e-19
C5312 _340_/a_27_47# _340_/a_652_21# 0.185f
C5313 _308_/a_193_47# output24/a_27_47# 1.55e-19
C5314 net44 _204_/a_75_212# 1.06e-20
C5315 _033_ net19 0.00928f
C5316 _186_/a_109_297# net54 1.18e-20
C5317 net43 clknet_2_1__leaf_clk 0.305f
C5318 VPWR _075_ 0.573f
C5319 _292_/a_493_297# _123_ 4.54e-20
C5320 en_co_clk net30 0.00826f
C5321 net43 _319_/a_761_289# 0.16f
C5322 output31/a_27_47# _056_ 1.1e-19
C5323 net31 _176_/a_27_47# 5.31e-19
C5324 clkbuf_0_clk/a_110_47# _304_/a_1108_47# 4.44e-19
C5325 _320_/a_1108_47# _078_ 8.98e-19
C5326 _337_/a_193_47# _337_/a_448_47# 0.0642f
C5327 _337_/a_761_289# _337_/a_1108_47# 0.0512f
C5328 _337_/a_27_47# _337_/a_651_413# 9.73e-19
C5329 _232_/a_32_297# _092_ 0.113f
C5330 _333_/a_1108_47# net32 5.89e-19
C5331 _340_/a_1182_261# _133_ 9.84e-20
C5332 mask\[6\] _155_/a_150_297# 2.29e-19
C5333 net9 _339_/a_1032_413# 7.41e-19
C5334 _083_ _074_ 0.0735f
C5335 _340_/a_652_21# clknet_2_3__leaf_clk 9.5e-21
C5336 _051_ _098_ 0.00409f
C5337 _048_ cal_itt\[3\] 2.38e-19
C5338 _326_/a_27_47# _007_ 0.00105f
C5339 _333_/a_27_47# _172_/a_68_297# 3.35e-19
C5340 _042_ _249_/a_27_297# 0.0295f
C5341 _041_ _122_ 0.0417f
C5342 _338_/a_1182_261# _122_ 0.00536f
C5343 _291_/a_285_47# cal_count\[0\] 0.00164f
C5344 _033_ _107_ 0.00183f
C5345 VPWR _195_/a_505_21# 0.21f
C5346 _097_ _237_/a_505_21# 2.46e-19
C5347 _104_ _279_/a_490_47# 0.00142f
C5348 VPWR cal_itt\[2\] 0.738f
C5349 net3 _192_/a_639_47# 0.00452f
C5350 _303_/a_193_47# _067_ 9.32e-21
C5351 _324_/a_543_47# mask\[6\] 7.79e-22
C5352 _324_/a_27_47# _021_ 0.279f
C5353 _303_/a_193_47# _070_ 1.44e-19
C5354 _304_/a_193_47# net4 8.89e-21
C5355 _239_/a_694_21# _095_ 1.94e-20
C5356 VPWR _334_/a_1108_47# 0.303f
C5357 _326_/a_193_47# net25 1.29e-19
C5358 _291_/a_35_297# net2 5.01e-19
C5359 _051_ clknet_0_clk 1.46f
C5360 _314_/a_448_47# net29 8.96e-20
C5361 _048_ _262_/a_205_47# 3.16e-19
C5362 VPWR _327_/a_543_47# 0.22f
C5363 _307_/a_651_413# mask\[0\] 1.44e-20
C5364 _307_/a_1270_413# net22 2.15e-19
C5365 _050_ _054_ 0.0156f
C5366 _335_/a_1108_47# _032_ 1.92e-19
C5367 _050_ net30 4.74e-19
C5368 _313_/a_27_47# _155_/a_68_297# 3.73e-21
C5369 _052_ net41 0.00169f
C5370 cal output41/a_27_47# 0.0251f
C5371 input1/a_75_212# net41 0.0639f
C5372 _299_/a_298_297# _297_/a_47_47# 5.42e-19
C5373 _236_/a_109_297# clknet_2_0__leaf_clk 1.15e-20
C5374 en_co_clk _072_ 1.19e-19
C5375 _311_/a_543_47# _311_/a_639_47# 0.0138f
C5376 _311_/a_193_47# _311_/a_1217_47# 2.36e-20
C5377 _311_/a_761_289# _311_/a_805_47# 3.69e-19
C5378 VPWR _137_/a_150_297# 0.00231f
C5379 output21/a_27_47# mask\[6\] 0.00634f
C5380 VPWR net35 0.519f
C5381 output10/a_27_47# _335_/a_1283_21# 1.15e-19
C5382 _304_/a_639_47# _136_ 2.96e-19
C5383 _104_ _092_ 1.49e-20
C5384 output38/a_27_47# output39/a_27_47# 0.0523f
C5385 VPWR _335_/a_543_47# 0.212f
C5386 VPWR output11/a_27_47# 0.276f
C5387 net45 mask\[2\] 6.57e-20
C5388 trim[4] _332_/a_1283_21# 4.74e-19
C5389 _305_/a_193_47# en_co_clk 3.91e-21
C5390 _277_/a_75_212# net18 8.68e-19
C5391 _304_/a_193_47# _063_ 0.00209f
C5392 net12 _337_/a_27_47# 1.79e-21
C5393 _304_/a_1217_47# net47 8.02e-19
C5394 _076_ cal_itt\[3\] 1.53e-20
C5395 _341_/a_27_47# _304_/a_27_47# 4.05e-20
C5396 net55 _092_ 0.222f
C5397 output22/a_27_47# sample 4.4e-21
C5398 result[0] output30/a_27_47# 0.00176f
C5399 _258_/a_109_47# net18 2.46e-19
C5400 _258_/a_27_297# _256_/a_27_297# 1.26e-20
C5401 _060_ _235_/a_79_21# 7.13e-20
C5402 _340_/a_476_47# net47 0.205f
C5403 _256_/a_373_47# trim_mask\[0\] 0.00145f
C5404 _256_/a_27_297# _024_ 0.121f
C5405 _037_ _304_/a_193_47# 8.53e-19
C5406 _061_ en_co_clk 0.0379f
C5407 VPWR _314_/a_1217_47# 1.22e-19
C5408 net4 net18 4.59e-22
C5409 _097_ _241_/a_297_47# 0.0499f
C5410 _106_ _279_/a_314_297# 3.92e-19
C5411 _065_ _208_/a_505_21# 0.0772f
C5412 _308_/a_1462_47# mask\[0\] 4.24e-19
C5413 _308_/a_1217_47# _078_ 3.07e-19
C5414 net43 _210_/a_113_297# 1.58e-19
C5415 VPWR _332_/a_761_289# 0.221f
C5416 _340_/a_27_47# _340_/a_1056_47# 0.00248f
C5417 _228_/a_297_47# _054_ 7.75e-20
C5418 output31/a_27_47# _173_/a_27_47# 0.00944f
C5419 _103_ _107_ 0.0467f
C5420 _052_ _171_/a_27_47# 4.28e-20
C5421 result[6] result[7] 0.0507f
C5422 _293_/a_81_21# net16 0.00959f
C5423 _277_/a_75_212# _276_/a_59_75# 0.0157f
C5424 net26 _310_/a_27_47# 1.7e-19
C5425 mask\[2\] _065_ 1.79e-20
C5426 ctlp[0] _314_/a_639_47# 3.92e-20
C5427 _305_/a_27_47# _076_ 0.0104f
C5428 _308_/a_27_47# _004_ 2.88e-20
C5429 VPWR _288_/a_59_75# 0.212f
C5430 _253_/a_299_297# _253_/a_384_47# 1.48e-19
C5431 _217_/a_109_297# _074_ 0.00223f
C5432 net35 _161_/a_68_297# 2.12e-19
C5433 _309_/a_543_47# _078_ 0.00886f
C5434 _309_/a_1283_21# mask\[0\] 1.94e-19
C5435 _001_ _065_ 0.437f
C5436 _259_/a_109_297# net50 0.00887f
C5437 _259_/a_109_47# trim_mask\[3\] 0.00453f
C5438 _064_ _275_/a_299_297# 1.87e-19
C5439 _326_/a_27_47# _310_/a_1283_21# 3.63e-19
C5440 _326_/a_193_47# _310_/a_543_47# 1.44e-20
C5441 _326_/a_543_47# _310_/a_193_47# 5.84e-21
C5442 _337_/a_27_47# net44 0.298f
C5443 _309_/a_27_47# net24 0.0466f
C5444 _276_/a_59_75# net4 7.64e-22
C5445 _338_/a_27_47# clknet_2_3__leaf_clk 0.781f
C5446 net51 rebuffer6/a_27_47# 3.53e-19
C5447 VPWR _310_/a_651_413# 0.134f
C5448 _067_ _092_ 0.0862f
C5449 _133_ _297_/a_47_47# 0.148f
C5450 net43 _313_/a_27_47# 0.306f
C5451 net34 _175_/a_68_297# 0.00256f
C5452 net34 _333_/a_193_47# 2.12e-20
C5453 _333_/a_543_47# _055_ 1.88e-20
C5454 _035_ _338_/a_1032_413# 4.03e-20
C5455 _110_ _051_ 3.65e-20
C5456 _319_/a_27_47# mask\[2\] 7.21e-21
C5457 result[5] _224_/a_199_47# 5.81e-21
C5458 net28 _078_ 0.0029f
C5459 _242_/a_79_21# _098_ 0.0614f
C5460 _188_/a_27_47# trim_val\[0\] 1.76e-19
C5461 _306_/a_761_289# net51 2.89e-19
C5462 _063_ net18 2.7e-19
C5463 _321_/a_543_47# _101_ 0.0338f
C5464 _321_/a_193_47# net52 0.0131f
C5465 _338_/a_381_47# net18 0.00126f
C5466 _324_/a_1217_47# _021_ 2.14e-20
C5467 _321_/a_1283_21# _041_ 9.15e-20
C5468 cal_count\[1\] _289_/a_150_297# 0.00101f
C5469 _015_ clknet_0_clk 2e-20
C5470 _037_ net18 1.21e-20
C5471 _231_/a_161_47# _194_/a_113_297# 3.63e-19
C5472 _053_ _170_/a_81_21# 0.186f
C5473 _339_/a_1182_261# net40 4.04e-20
C5474 _060_ _049_ 0.00176f
C5475 _307_/a_448_47# _004_ 0.16f
C5476 _198_/a_27_47# _198_/a_109_47# 0.00517f
C5477 _057_ net33 4.43e-21
C5478 VPWR _247_/a_109_297# 0.177f
C5479 _311_/a_761_289# net26 0.0191f
C5480 _322_/a_1108_47# _078_ 0.0161f
C5481 output27/a_27_47# net26 5.05e-21
C5482 mask\[0\] _092_ 2e-19
C5483 trim_mask\[0\] clk 0.00535f
C5484 _259_/a_109_297# _330_/a_1108_47# 1.52e-19
C5485 _080_ clknet_2_1__leaf_clk 5.41e-19
C5486 _329_/a_193_47# trim_mask\[3\] 0.003f
C5487 cal_itt\[2\] _262_/a_27_47# 1.31e-19
C5488 _326_/a_27_47# net27 0.00215f
C5489 _287_/a_75_212# _339_/a_27_47# 2.52e-21
C5490 net3 _243_/a_373_47# 1.2e-19
C5491 _331_/a_193_47# _331_/a_761_289# 0.18f
C5492 _331_/a_27_47# _331_/a_543_47# 0.112f
C5493 _339_/a_1032_413# _122_ 0.00357f
C5494 _185_/a_68_297# calibrate 5.21e-20
C5495 VPWR _311_/a_639_47# 2.33e-19
C5496 _325_/a_27_47# _251_/a_27_297# 0.00122f
C5497 _325_/a_193_47# _250_/a_109_297# 6.47e-20
C5498 result[3] _078_ 3.52e-19
C5499 _199_/a_109_297# _070_ 1.38e-19
C5500 clkbuf_2_3__f_clk/a_110_47# net19 0.018f
C5501 net47 _338_/a_193_47# 0.509f
C5502 mask\[1\] net45 0.124f
C5503 net12 _051_ 0.23f
C5504 _340_/a_1224_47# net47 8.78e-19
C5505 _185_/a_68_297# net45 3.5e-20
C5506 _325_/a_543_47# clknet_2_1__leaf_clk 0.00214f
C5507 _311_/a_639_47# net53 6.89e-19
C5508 trim_mask\[0\] net4 0.0222f
C5509 _319_/a_1108_47# en_co_clk 3.26e-22
C5510 ctlp[7] _313_/a_1283_21# 0.00107f
C5511 _340_/a_1182_261# _037_ 0.00151f
C5512 _005_ result[2] 4.79e-21
C5513 _224_/a_199_47# net29 5.38e-19
C5514 _327_/a_1283_21# _111_ 0.0362f
C5515 trimb[2] net34 0.0773f
C5516 _043_ net19 0.0119f
C5517 output31/a_27_47# _172_/a_68_297# 0.001f
C5518 _059_ net41 0.174f
C5519 output26/a_27_47# _074_ 1.55e-19
C5520 _294_/a_150_297# net40 4.26e-19
C5521 _301_/a_285_47# clknet_2_3__leaf_clk 0.0449f
C5522 _320_/a_651_413# clknet_0_clk 4.43e-19
C5523 mask\[1\] _065_ 0.00925f
C5524 _337_/a_1217_47# net44 6.03e-19
C5525 _239_/a_694_21# _226_/a_27_47# 0.00111f
C5526 _107_ clkbuf_2_3__f_clk/a_110_47# 0.0141f
C5527 _291_/a_117_297# _127_ 0.00787f
C5528 _294_/a_68_297# net34 3.27e-20
C5529 _341_/a_543_47# clknet_2_3__leaf_clk 0.0431f
C5530 calibrate _088_ 0.218f
C5531 _336_/a_1283_21# _330_/a_1283_21# 7.1e-20
C5532 state\[0\] _192_/a_174_21# 1.68e-21
C5533 _233_/a_373_47# net1 0.00105f
C5534 _074_ input1/a_75_212# 0.00827f
C5535 _058_ fanout46/a_27_47# 1.08e-19
C5536 _113_ net46 0.14f
C5537 output20/a_27_47# ctlp[5] 5.22e-20
C5538 _051_ net44 0.00365f
C5539 net30 _039_ 9.56e-19
C5540 net43 _313_/a_1217_47# 2.95e-19
C5541 _329_/a_27_47# _330_/a_1108_47# 2.73e-20
C5542 fanout46/a_27_47# _335_/a_193_47# 1.22e-19
C5543 _291_/a_285_47# net16 5.96e-19
C5544 VPWR _306_/a_543_47# 0.221f
C5545 _340_/a_193_47# _339_/a_27_47# 0.00126f
C5546 _340_/a_27_47# _339_/a_193_47# 0.00117f
C5547 _188_/a_27_47# _131_ 7.53e-22
C5548 trim_mask\[0\] _063_ 0.271f
C5549 _307_/a_27_47# _138_/a_27_47# 0.0025f
C5550 trim[1] _109_ 6.11e-20
C5551 net4 _191_/a_27_297# 8.17e-19
C5552 en_co_clk _066_ 2.69e-21
C5553 _326_/a_543_47# _224_/a_113_297# 2.12e-19
C5554 _050_ _319_/a_1108_47# 3.91e-20
C5555 _068_ cal_itt\[3\] 3.49e-19
C5556 VPWR _170_/a_81_21# 0.205f
C5557 net2 net46 1.9e-19
C5558 _029_ _332_/a_761_289# 9.46e-20
C5559 _111_ _108_ 0.0474f
C5560 state\[2\] fanout45/a_27_47# 2.77e-20
C5561 _316_/a_1283_21# _099_ 5.48e-21
C5562 _316_/a_1108_47# _095_ 9.99e-20
C5563 _291_/a_117_297# _126_ 7.6e-19
C5564 _144_/a_27_47# _339_/a_193_47# 3.33e-21
C5565 _051_ _263_/a_79_21# 0.0135f
C5566 clk _331_/a_805_47# 5.18e-19
C5567 _185_/a_68_297# _243_/a_109_297# 7.35e-20
C5568 cal_itt\[0\] _065_ 0.0235f
C5569 _162_/a_27_47# _333_/a_1283_21# 0.00139f
C5570 _058_ _269_/a_299_297# 6.04e-19
C5571 _323_/a_543_47# net47 0.153f
C5572 net16 en_co_clk 0.045f
C5573 _170_/a_384_47# net41 4.96e-22
C5574 _339_/a_193_47# clknet_2_3__leaf_clk 0.00203f
C5575 trim_mask\[2\] _280_/a_75_212# 0.0345f
C5576 _071_ net2 1.4e-19
C5577 _312_/a_193_47# net20 0.0347f
C5578 VPWR _018_ 0.477f
C5579 _181_/a_68_297# _336_/a_1283_21# 0.00107f
C5580 _136_ _301_/a_129_47# 4.21e-19
C5581 _104_ _330_/a_651_413# 6.03e-20
C5582 _259_/a_27_297# _027_ 0.118f
C5583 _306_/a_27_47# _306_/a_1217_47# 2.56e-19
C5584 _306_/a_761_289# _306_/a_639_47# 3.16e-19
C5585 _293_/a_81_21# net40 0.00278f
C5586 _110_ _333_/a_27_47# 6.35e-19
C5587 cal_itt\[2\] _305_/a_1270_413# 9.87e-20
C5588 _071_ _305_/a_1283_21# 0.0266f
C5589 net50 _106_ 2.39e-21
C5590 VPWR _227_/a_296_53# 4.83e-20
C5591 _341_/a_761_289# _136_ 0.00384f
C5592 net15 net7 0.109f
C5593 _235_/a_79_21# _235_/a_297_47# 0.0326f
C5594 net15 _317_/a_193_47# 0.0174f
C5595 _331_/a_761_289# _260_/a_93_21# 7.97e-21
C5596 _081_ _006_ 0.117f
C5597 _292_/a_78_199# _298_/a_78_199# 8.87e-19
C5598 _325_/a_1283_21# mask\[6\] 0.129f
C5599 _245_/a_373_47# _016_ 1.97e-19
C5600 _041_ _101_ 0.0098f
C5601 _191_/a_27_297# _063_ 0.045f
C5602 clkbuf_0_clk/a_110_47# net19 0.0206f
C5603 cal_count\[3\] net19 0.00666f
C5604 _256_/a_373_47# trim_mask\[4\] 2.84e-19
C5605 _159_/a_27_47# _046_ 0.198f
C5606 _078_ _084_ 0.00638f
C5607 _306_/a_193_47# _049_ 4.22e-19
C5608 _041_ _338_/a_1032_413# 3.51e-19
C5609 _308_/a_543_47# net14 0.00542f
C5610 _338_/a_652_21# _338_/a_381_47# 7.79e-20
C5611 _338_/a_193_47# _338_/a_562_413# 4.45e-20
C5612 _338_/a_1182_261# _338_/a_1032_413# 0.344f
C5613 _338_/a_27_47# _338_/a_956_413# 0.00294f
C5614 net47 _338_/a_796_47# 0.00291f
C5615 VPWR _317_/a_543_47# 0.205f
C5616 _308_/a_1108_47# _138_/a_27_47# 1.9e-19
C5617 _059_ _094_ 0.0451f
C5618 _328_/a_27_47# _328_/a_761_289# 0.0535f
C5619 VPWR _326_/a_543_47# 0.212f
C5620 _258_/a_109_297# trim_mask\[2\] 0.0116f
C5621 _311_/a_1108_47# _072_ 2.67e-20
C5622 _108_ rebuffer3/a_75_212# 0.221f
C5623 _121_ _092_ 1.03e-21
C5624 _060_ state\[1\] 0.0926f
C5625 _074_ _310_/a_639_47# 0.00204f
C5626 _082_ clknet_2_1__leaf_clk 0.00131f
C5627 net45 _244_/a_27_297# 6.53e-19
C5628 output29/a_27_47# _314_/a_27_47# 0.0106f
C5629 net4 _090_ 3.3e-20
C5630 _317_/a_1108_47# net41 3.16e-21
C5631 _331_/a_27_47# net19 0.00294f
C5632 _326_/a_651_413# output14/a_27_47# 1.35e-20
C5633 net13 _337_/a_761_289# 0.00672f
C5634 state\[2\] _331_/a_193_47# 1.43e-20
C5635 _228_/a_382_297# _100_ 6.54e-20
C5636 net12 _242_/a_79_21# 0.00775f
C5637 _051_ clknet_2_2__leaf_clk 5.36e-19
C5638 VPWR _286_/a_218_374# 0.00203f
C5639 net36 net33 0.157f
C5640 _325_/a_27_47# _313_/a_543_47# 3.71e-21
C5641 _325_/a_543_47# _313_/a_27_47# 8.17e-21
C5642 _065_ _108_ 8.54e-20
C5643 _107_ cal_count\[3\] 0.00455f
C5644 trim_val\[1\] net46 0.0319f
C5645 _323_/a_1283_21# net4 5.5e-20
C5646 net44 _312_/a_761_289# 0.17f
C5647 net2 _332_/a_448_47# 1.91e-19
C5648 _336_/a_193_47# net46 0.0247f
C5649 _065_ _244_/a_27_297# 0.0937f
C5650 _227_/a_109_93# _049_ 0.00546f
C5651 _323_/a_543_47# net44 0.00197f
C5652 _192_/a_27_47# net41 2.68e-21
C5653 _303_/a_193_47# clknet_2_3__leaf_clk 0.588f
C5654 _320_/a_27_47# _041_ 7.84e-19
C5655 cal_itt\[0\] _194_/a_113_297# 3.46e-19
C5656 _230_/a_145_75# _092_ 0.00232f
C5657 _149_/a_68_297# mask\[4\] 0.195f
C5658 net47 _339_/a_652_21# 0.158f
C5659 cal_itt\[2\] _202_/a_79_21# 0.00349f
C5660 clkbuf_2_2__f_clk/a_110_47# trim_val\[4\] 1.41e-19
C5661 _257_/a_27_297# _256_/a_27_297# 8.33e-19
C5662 _305_/a_761_289# net51 4.95e-19
C5663 _075_ _206_/a_27_93# 0.159f
C5664 _272_/a_81_21# _334_/a_651_413# 5.04e-20
C5665 trim_val\[2\] _334_/a_193_47# 4.18e-19
C5666 _231_/a_161_47# _278_/a_27_47# 3.92e-20
C5667 _323_/a_27_47# _323_/a_761_289# 0.0701f
C5668 _340_/a_1602_47# _339_/a_1602_47# 1.04e-20
C5669 VPWR _187_/a_27_413# 0.217f
C5670 _140_/a_68_297# _245_/a_27_297# 7.94e-19
C5671 _336_/a_543_47# _052_ 1.55e-20
C5672 net15 net30 0.429f
C5673 _306_/a_27_47# cal_itt\[3\] 1.84e-19
C5674 _189_/a_27_47# _053_ 2.5e-19
C5675 _048_ clone7/a_27_47# 2.01e-20
C5676 trim_mask\[2\] _273_/a_59_75# 0.0537f
C5677 VPWR _268_/a_75_212# 0.257f
C5678 net27 _011_ 0.0592f
C5679 result[5] _086_ 3.98e-19
C5680 net16 _334_/a_193_47# 3.08e-20
C5681 VPWR _318_/a_448_47# 0.0829f
C5682 _315_/a_27_47# net41 1.9e-20
C5683 _308_/a_193_47# _081_ 1.5e-21
C5684 _042_ _310_/a_761_289# 2.1e-20
C5685 cal_count\[0\] output40/a_27_47# 3.06e-19
C5686 clk trim_mask\[4\] 0.00945f
C5687 _169_/a_215_311# _096_ 6.38e-21
C5688 net43 _321_/a_761_289# 0.182f
C5689 _312_/a_1462_47# net20 1.27e-19
C5690 clknet_2_1__leaf_clk _310_/a_448_47# 0.0289f
C5691 _104_ net46 0.688f
C5692 _078_ _085_ 0.00491f
C5693 net43 _337_/a_761_289# 6.51e-20
C5694 _341_/a_639_47# _038_ 0.00196f
C5695 _331_/a_639_47# clknet_2_2__leaf_clk 2.44e-19
C5696 _331_/a_1283_21# trim_mask\[4\] 0.0893f
C5697 clkbuf_2_3__f_clk/a_110_47# _118_ 2.47e-19
C5698 _260_/a_93_21# _260_/a_250_297# 0.188f
C5699 _317_/a_761_289# _317_/a_639_47# 3.16e-19
C5700 _317_/a_27_47# _317_/a_1217_47# 2.56e-19
C5701 net9 _334_/a_761_289# 3.21e-19
C5702 _258_/a_109_47# trim_mask\[4\] 1.17e-19
C5703 _328_/a_543_47# clknet_2_2__leaf_clk 0.0363f
C5704 _332_/a_1108_47# net33 1.36e-19
C5705 _326_/a_27_47# _326_/a_1217_47# 2.56e-19
C5706 _326_/a_761_289# _326_/a_639_47# 3.16e-19
C5707 net49 rebuffer2/a_75_212# 0.111f
C5708 _325_/a_651_413# _078_ 2.26e-19
C5709 _216_/a_199_47# _078_ 0.00136f
C5710 state\[0\] _232_/a_32_297# 8.12e-19
C5711 _337_/a_193_47# _034_ 0.293f
C5712 _194_/a_113_297# _108_ 5.02e-19
C5713 _327_/a_27_47# net9 5.13e-22
C5714 net4 trim_mask\[4\] 0.0156f
C5715 net49 _332_/a_1283_21# 1.28e-21
C5716 _112_ _108_ 0.00294f
C5717 _112_ _332_/a_543_47# 1.87e-20
C5718 _338_/a_1032_413# _338_/a_1296_47# 0.00384f
C5719 _328_/a_543_47# _328_/a_805_47# 0.00171f
C5720 _328_/a_761_289# _328_/a_1217_47# 4.2e-19
C5721 _328_/a_1108_47# _328_/a_1270_413# 0.00645f
C5722 _341_/a_27_47# _341_/a_1283_21# 0.0436f
C5723 _341_/a_193_47# _341_/a_543_47# 0.206f
C5724 _336_/a_1283_21# _108_ 0.00369f
C5725 _320_/a_651_413# net44 0.0122f
C5726 _127_ net37 0.00111f
C5727 _341_/a_1108_47# _037_ 2.26e-19
C5728 net47 _303_/a_761_289# 0.171f
C5729 _329_/a_1108_47# rebuffer1/a_75_212# 2.03e-20
C5730 trim_mask\[0\] _279_/a_396_47# 0.0296f
C5731 _256_/a_27_297# trim_val\[4\] 5.6e-20
C5732 _053_ _336_/a_27_47# 0.00136f
C5733 clknet_2_0__leaf_clk net41 0.123f
C5734 _309_/a_448_47# net14 0.00314f
C5735 _049_ _054_ 0.243f
C5736 state\[2\] _260_/a_93_21# 0.00652f
C5737 _094_ _192_/a_27_47# 3.55e-19
C5738 _273_/a_59_75# _115_ 0.119f
C5739 net30 _049_ 0.0182f
C5740 _340_/a_1602_47# cal_count\[2\] 0.132f
C5741 _318_/a_27_47# _318_/a_448_47# 0.0931f
C5742 _318_/a_193_47# _318_/a_1108_47# 0.119f
C5743 _048_ _073_ 7.12e-19
C5744 clknet_2_1__leaf_clk _247_/a_27_297# 0.0724f
C5745 clknet_2_3__leaf_clk _092_ 0.0956f
C5746 net27 _250_/a_109_297# 6.97e-20
C5747 _104_ _335_/a_651_413# 1.87e-19
C5748 _042_ _311_/a_1283_21# 7.31e-20
C5749 _203_/a_59_75# _203_/a_145_75# 0.00658f
C5750 _114_ net46 0.0171f
C5751 _086_ net29 0.162f
C5752 _312_/a_761_289# _312_/a_639_47# 3.16e-19
C5753 _312_/a_27_47# _312_/a_1217_47# 2.56e-19
C5754 net43 _253_/a_81_21# 0.0109f
C5755 _309_/a_1283_21# _245_/a_109_297# 7.64e-22
C5756 _309_/a_1108_47# _245_/a_27_297# 3.74e-22
C5757 rstn output6/a_27_47# 4.51e-19
C5758 input4/a_27_47# net6 0.00163f
C5759 _312_/a_1283_21# net19 0.00166f
C5760 _336_/a_1462_47# net46 0.00196f
C5761 calibrate _170_/a_299_297# 0.0408f
C5762 _286_/a_76_199# _124_ 0.0999f
C5763 _306_/a_448_47# clknet_2_0__leaf_clk 1.99e-19
C5764 en_co_clk net40 0.084f
C5765 VPWR _305_/a_543_47# 0.214f
C5766 _195_/a_439_47# _067_ 0.0061f
C5767 result[5] clknet_2_1__leaf_clk 0.0773f
C5768 _329_/a_639_47# net46 9.54e-19
C5769 _078_ _314_/a_543_47# 6.41e-19
C5770 _071_ _067_ 0.0665f
C5771 _323_/a_1108_47# net19 0.0132f
C5772 trim_mask\[4\] _063_ 1.61e-20
C5773 net47 _339_/a_1056_47# 7.28e-19
C5774 _041_ _339_/a_1602_47# 0.0475f
C5775 _071_ _070_ 1.97e-19
C5776 _126_ net37 0.458f
C5777 _192_/a_27_47# _192_/a_505_280# 0.103f
C5778 _192_/a_174_21# _192_/a_476_47# 0.00228f
C5779 _307_/a_27_47# _307_/a_193_47# 0.806f
C5780 net20 _152_/a_68_297# 1.58e-20
C5781 _321_/a_1108_47# mask\[4\] 1.5e-19
C5782 _309_/a_543_47# mask\[7\] 8.38e-21
C5783 trim_val\[2\] _334_/a_1462_47# 6.42e-19
C5784 _323_/a_543_47# _323_/a_805_47# 0.00171f
C5785 _323_/a_761_289# _323_/a_1217_47# 4.2e-19
C5786 _323_/a_1108_47# _323_/a_1270_413# 0.00645f
C5787 net43 clkbuf_0_clk/a_110_47# 4.46e-19
C5788 VPWR _189_/a_27_47# 0.327f
C5789 cal_itt\[1\] _106_ 8.72e-20
C5790 _333_/a_27_47# clknet_2_2__leaf_clk 0.235f
C5791 output31/a_27_47# _047_ 2.51e-19
C5792 net31 _162_/a_27_47# 0.149f
C5793 _304_/a_27_47# _001_ 0.323f
C5794 VPWR clkbuf_2_1__f_clk/a_110_47# 1.22f
C5795 VPWR _315_/a_639_47# 8.62e-19
C5796 _306_/a_1217_47# cal_itt\[3\] 1.52e-19
C5797 _329_/a_193_47# _031_ 1.39e-19
C5798 en_co_clk _003_ 9.3e-20
C5799 _292_/a_215_47# net47 1.11e-19
C5800 _324_/a_27_47# _101_ 2.95e-20
C5801 clk _190_/a_27_47# 1.17e-19
C5802 _128_ _340_/a_1602_47# 7.48e-19
C5803 clknet_2_1__leaf_clk rebuffer6/a_27_47# 0.0024f
C5804 mask\[7\] net28 0.0586f
C5805 _326_/a_761_289# _086_ 6.54e-20
C5806 _326_/a_27_47# _011_ 1.73e-19
C5807 clkbuf_2_2__f_clk/a_110_47# _330_/a_193_47# 0.0169f
C5808 state\[0\] net55 0.00109f
C5809 _049_ _072_ 1.81e-20
C5810 _303_/a_761_289# net44 2.45e-19
C5811 _306_/a_1283_21# _305_/a_651_413# 8.82e-19
C5812 trim[4] net33 3.24e-19
C5813 _103_ _062_ 2.33e-19
C5814 _053_ net42 0.0279f
C5815 _320_/a_543_47# _320_/a_651_413# 0.0572f
C5816 _320_/a_761_289# _320_/a_1270_413# 2.6e-19
C5817 _320_/a_193_47# _320_/a_639_47# 2.28e-19
C5818 _309_/a_1283_21# _081_ 0.00119f
C5819 _309_/a_761_289# _006_ 6.55e-19
C5820 _107_ _242_/a_297_47# 0.00311f
C5821 _323_/a_27_47# _303_/a_193_47# 9.08e-21
C5822 _323_/a_193_47# _303_/a_27_47# 4.37e-21
C5823 _076_ _073_ 7.03e-20
C5824 trim_val\[3\] net18 0.00706f
C5825 mask\[7\] _158_/a_68_297# 0.188f
C5826 _193_/a_109_297# net18 6.37e-19
C5827 cal_count\[3\] _118_ 0.0221f
C5828 _296_/a_113_47# _132_ 0.00948f
C5829 _322_/a_27_47# _041_ 7.15e-20
C5830 _306_/a_761_289# clknet_2_1__leaf_clk 1.63e-19
C5831 _235_/a_297_47# state\[1\] 4.89e-22
C5832 trim_mask\[4\] _260_/a_346_47# 3.96e-19
C5833 _237_/a_535_374# _090_ 0.00106f
C5834 _094_ clknet_2_0__leaf_clk 0.0325f
C5835 clknet_2_1__leaf_clk _221_/a_109_297# 0.00422f
C5836 _317_/a_1108_47# _014_ 5.47e-21
C5837 _317_/a_448_47# clknet_2_0__leaf_clk 0.017f
C5838 _317_/a_1283_21# net45 0.337f
C5839 _317_/a_193_47# state\[1\] 1.92e-19
C5840 mask\[5\] _153_/a_27_47# 0.00284f
C5841 _308_/a_1108_47# _307_/a_193_47# 5.24e-20
C5842 VPWR _056_ 0.517f
C5843 _308_/a_193_47# _307_/a_1108_47# 6.41e-22
C5844 _308_/a_543_47# _307_/a_543_47# 8.87e-19
C5845 net13 net21 0.13f
C5846 _262_/a_193_297# net30 6.47e-19
C5847 _321_/a_27_47# mask\[2\] 9e-19
C5848 _315_/a_27_47# _315_/a_193_47# 0.888f
C5849 net21 _155_/a_68_297# 0.00231f
C5850 calibrate _192_/a_174_21# 4.35e-21
C5851 _006_ _040_ 1e-19
C5852 _341_/a_448_47# _341_/a_639_47# 4.61e-19
C5853 VPWR _336_/a_27_47# 0.513f
C5854 _050_ _003_ 3.51e-20
C5855 _110_ _275_/a_81_21# 0.0625f
C5856 _276_/a_59_75# trim_val\[3\] 2.68e-19
C5857 clknet_2_1__leaf_clk net29 0.00238f
C5858 mask\[6\] _247_/a_109_297# 5.16e-21
C5859 _065_ net26 2.68e-20
C5860 net37 output5/a_27_47# 6.9e-20
C5861 _333_/a_27_47# _333_/a_651_413# 9.73e-19
C5862 _333_/a_761_289# _333_/a_1108_47# 0.0512f
C5863 _333_/a_193_47# _333_/a_448_47# 0.0642f
C5864 _268_/a_75_212# _029_ 0.116f
C5865 net23 _245_/a_373_47# 0.00101f
C5866 clknet_2_0__leaf_clk _192_/a_505_280# 1.98e-21
C5867 trim_val\[0\] _333_/a_27_47# 2.17e-20
C5868 cal_itt\[0\] _278_/a_27_47# 6.48e-20
C5869 _078_ _311_/a_193_47# 5.67e-20
C5870 _251_/a_27_297# net15 0.0133f
C5871 _074_ _315_/a_27_47# 0.0275f
C5872 _324_/a_1270_413# net44 3.33e-19
C5873 _324_/a_193_47# _312_/a_1108_47# 1.89e-19
C5874 _324_/a_761_289# _312_/a_1283_21# 9.96e-21
C5875 _334_/a_27_47# net34 2.68e-20
C5876 _124_ cal_count\[0\] 0.0173f
C5877 _063_ _190_/a_27_47# 0.0985f
C5878 VPWR _251_/a_109_47# 4.28e-19
C5879 _053_ _168_/a_27_413# 1.27e-19
C5880 _248_/a_109_297# net21 2.6e-21
C5881 net12 _218_/a_113_297# 0.00206f
C5882 _308_/a_27_47# _308_/a_1217_47# 2.56e-19
C5883 _308_/a_761_289# _308_/a_639_47# 3.16e-19
C5884 _008_ net20 7.12e-22
C5885 trim_mask\[2\] _257_/a_109_297# 0.00203f
C5886 _324_/a_1283_21# _323_/a_543_47# 3.32e-19
C5887 net15 _319_/a_1108_47# 9.63e-19
C5888 _192_/a_174_21# _065_ 0.122f
C5889 _014_ _315_/a_27_47# 1.2e-20
C5890 _307_/a_761_289# _307_/a_805_47# 3.69e-19
C5891 _307_/a_193_47# _307_/a_1217_47# 2.36e-20
C5892 _307_/a_543_47# _307_/a_639_47# 0.0138f
C5893 clknet_2_0__leaf_clk _315_/a_193_47# 0.0103f
C5894 net54 clone7/a_27_47# 0.179f
C5895 _087_ _099_ 0.153f
C5896 _326_/a_761_289# clknet_2_1__leaf_clk 4.07e-20
C5897 _249_/a_109_47# _101_ 0.00599f
C5898 _074_ _225_/a_109_297# 0.00107f
C5899 result[0] _307_/a_651_413# 5.48e-19
C5900 VPWR _319_/a_651_413# 0.143f
C5901 _322_/a_651_413# net44 0.0122f
C5902 _318_/a_651_413# net45 0.0122f
C5903 net27 _313_/a_761_289# 2.51e-21
C5904 _309_/a_27_47# _308_/a_543_47# 3.47e-19
C5905 _309_/a_193_47# _308_/a_761_289# 2.21e-21
C5906 _233_/a_373_47# _012_ 1.97e-19
C5907 output15/a_27_47# net29 8.41e-19
C5908 _128_ _041_ 0.012f
C5909 VPWR _096_ 0.938f
C5910 mask\[5\] net20 0.0649f
C5911 _325_/a_27_47# _321_/a_1108_47# 8.37e-21
C5912 output38/a_27_47# trimb[2] 0.337f
C5913 net23 _006_ 0.00178f
C5914 net43 net21 0.0413f
C5915 VPWR net42 0.687f
C5916 _306_/a_1108_47# _002_ 8.81e-19
C5917 _187_/a_212_413# _135_ 4.37e-19
C5918 _337_/a_1108_47# en_co_clk 0.05f
C5919 _074_ clknet_2_0__leaf_clk 0.167f
C5920 _303_/a_1283_21# net19 1.08e-19
C5921 VPWR _173_/a_27_47# 0.221f
C5922 _108_ _278_/a_27_47# 3.51e-19
C5923 cal _316_/a_193_47# 2.27e-19
C5924 net1 _316_/a_27_47# 3.65e-20
C5925 _339_/a_652_21# _339_/a_956_413# 3.11e-19
C5926 _339_/a_1032_413# _339_/a_1602_47# 0.111f
C5927 _339_/a_476_47# _339_/a_562_413# 0.00972f
C5928 _263_/a_297_47# _099_ 0.0373f
C5929 net8 net46 0.041f
C5930 _289_/a_68_297# trimb[4] 1.71e-19
C5931 _341_/a_193_47# _092_ 7.25e-19
C5932 _317_/a_1462_47# state\[1\] 6.42e-19
C5933 clknet_2_0__leaf_clk _014_ 0.0967f
C5934 _005_ _307_/a_27_47# 1.8e-20
C5935 _320_/a_448_47# _040_ 0.0214f
C5936 _062_ clkbuf_2_3__f_clk/a_110_47# 0.159f
C5937 cal_itt\[0\] _304_/a_27_47# 2.9e-21
C5938 VPWR net48 0.412f
C5939 _315_/a_543_47# _315_/a_639_47# 0.0138f
C5940 _315_/a_193_47# _315_/a_1217_47# 2.36e-20
C5941 _315_/a_761_289# _315_/a_805_47# 3.69e-19
C5942 _337_/a_1283_21# _076_ 0.00101f
C5943 output22/a_27_47# net43 1.91e-19
C5944 trim_mask\[4\] _279_/a_396_47# 6.28e-19
C5945 VPWR _336_/a_1217_47# 5.34e-19
C5946 _053_ _284_/a_68_297# 0.171f
C5947 VPWR _127_ 0.264f
C5948 mask\[6\] _018_ 3.93e-20
C5949 _000_ _041_ 0.2f
C5950 VPWR _329_/a_1270_413# 8.28e-19
C5951 _117_ _057_ 7.58e-20
C5952 net8 _334_/a_639_47# 7.53e-19
C5953 _319_/a_1108_47# _049_ 0.00215f
C5954 VPWR result[7] 0.646f
C5955 _321_/a_27_47# mask\[1\] 3.14e-21
C5956 _036_ net17 0.00164f
C5957 _074_ _146_/a_68_297# 4.36e-21
C5958 _050_ _337_/a_1108_47# 3.29e-20
C5959 output23/a_27_47# clknet_2_0__leaf_clk 0.00967f
C5960 _313_/a_27_47# net29 0.00312f
C5961 _237_/a_76_199# _241_/a_297_47# 7.48e-20
C5962 _195_/a_76_199# clkbuf_2_3__f_clk/a_110_47# 1.49e-19
C5963 _167_/a_161_47# _050_ 1.97e-20
C5964 _051_ _166_/a_161_47# 0.0551f
C5965 _323_/a_27_47# mask\[5\] 9.28e-19
C5966 _012_ _315_/a_651_413# 1.08e-20
C5967 calibrate _315_/a_805_47# 3.62e-20
C5968 _200_/a_80_21# clknet_2_3__leaf_clk 0.00128f
C5969 _331_/a_193_47# _330_/a_193_47# 0.00469f
C5970 _322_/a_448_47# _320_/a_1283_21# 2.48e-20
C5971 VPWR _168_/a_27_413# 0.235f
C5972 _326_/a_543_47# mask\[6\] 1.16e-21
C5973 _212_/a_113_297# net14 0.0087f
C5974 fanout44/a_27_47# _337_/a_761_289# 4.89e-20
C5975 _324_/a_27_47# _324_/a_193_47# 0.906f
C5976 state\[0\] _316_/a_543_47# 1.56e-19
C5977 _246_/a_373_47# net52 0.00141f
C5978 _308_/a_193_47# net23 4.14e-19
C5979 _308_/a_1283_21# net43 0.294f
C5980 VPWR net22 0.751f
C5981 _308_/a_1108_47# _005_ 1.51e-19
C5982 net10 net9 2.17e-19
C5983 _328_/a_1108_47# _025_ 7.13e-20
C5984 trim_mask\[2\] _025_ 1.26e-19
C5985 VPWR _126_ 0.852f
C5986 net45 _315_/a_805_47# 0.00316f
C5987 _002_ _203_/a_59_75# 5.1e-20
C5988 _189_/a_27_47# wire42/a_75_212# 4.96e-20
C5989 net2 _065_ 1.15f
C5990 net2 _135_ 0.0394f
C5991 _305_/a_1283_21# _065_ 6.43e-20
C5992 _339_/a_1032_413# cal_count\[2\] 3.38e-21
C5993 mask\[4\] net19 0.0812f
C5994 _110_ _330_/a_1270_413# 1.46e-19
C5995 _327_/a_27_47# _256_/a_109_297# 3.33e-19
C5996 _327_/a_193_47# _256_/a_27_297# 2.86e-20
C5997 _327_/a_543_47# net18 0.00215f
C5998 net43 _320_/a_639_47# 5.05e-20
C5999 _097_ _317_/a_193_47# 4.42e-21
C6000 _323_/a_1270_413# mask\[4\] 2.86e-20
C6001 _321_/a_1283_21# mask\[3\] 5.87e-20
C6002 _305_/a_27_47# _305_/a_1217_47# 2.56e-19
C6003 _305_/a_761_289# _305_/a_639_47# 3.16e-19
C6004 calibrate _232_/a_32_297# 2.97e-19
C6005 _281_/a_253_47# _090_ 0.00432f
C6006 _110_ _267_/a_59_75# 0.17f
C6007 _309_/a_193_47# _309_/a_1108_47# 0.119f
C6008 _309_/a_27_47# _309_/a_448_47# 0.0931f
C6009 VPWR _313_/a_1108_47# 0.31f
C6010 comp net34 0.108f
C6011 _312_/a_27_47# _084_ 0.0128f
C6012 net5 comp 6.19e-20
C6013 _146_/a_68_297# _146_/a_150_297# 0.00477f
C6014 _256_/a_27_297# _058_ 0.0068f
C6015 _241_/a_388_297# _241_/a_297_47# 0.0023f
C6016 _305_/a_761_289# clknet_2_1__leaf_clk 3.05e-20
C6017 VPWR _172_/a_68_297# 0.156f
C6018 _259_/a_27_297# _259_/a_109_297# 0.171f
C6019 _081_ _017_ 8.78e-21
C6020 _149_/a_68_297# _311_/a_1108_47# 4.14e-20
C6021 _309_/a_1283_21# _040_ 3.64e-19
C6022 _030_ net49 4.69e-20
C6023 _182_/a_27_47# _047_ 4.27e-20
C6024 _113_ _112_ 0.11f
C6025 clkbuf_0_clk/a_110_47# _062_ 0.00163f
C6026 cal_count\[3\] _062_ 0.0484f
C6027 cal_itt\[1\] _304_/a_805_47# 8.64e-20
C6028 VPWR _284_/a_68_297# 0.165f
C6029 _050_ _331_/a_543_47# 0.00129f
C6030 clkbuf_2_1__f_clk/a_110_47# _319_/a_193_47# 0.0204f
C6031 _155_/a_68_297# _045_ 0.106f
C6032 comp _299_/a_298_297# 2.03e-19
C6033 _325_/a_193_47# _101_ 5.62e-19
C6034 _324_/a_1108_47# _152_/a_68_297# 4.78e-20
C6035 _036_ _339_/a_193_47# 0.0549f
C6036 net42 _262_/a_27_47# 0.0928f
C6037 mask\[7\] _085_ 2e-19
C6038 _128_ _339_/a_1032_413# 0.0126f
C6039 _119_ _330_/a_448_47# 4.88e-19
C6040 net52 rebuffer5/a_161_47# 0.306f
C6041 _313_/a_1108_47# _009_ 4.04e-20
C6042 _072_ _202_/a_297_47# 0.00672f
C6043 _232_/a_32_297# _065_ 0.00109f
C6044 _053_ _230_/a_59_75# 0.0834f
C6045 VPWR output5/a_27_47# 0.283f
C6046 _125_ _122_ 8.39e-20
C6047 _058_ _302_/a_109_47# 6.13e-20
C6048 net46 clknet_2_3__leaf_clk 0.375f
C6049 _303_/a_761_289# _303_/a_639_47# 3.16e-19
C6050 _303_/a_27_47# _303_/a_1217_47# 2.56e-19
C6051 _047_ net37 0.454f
C6052 _102_ _216_/a_113_297# 3.99e-20
C6053 _089_ _226_/a_27_47# 2.73e-19
C6054 _020_ net19 0.0017f
C6055 net15 _316_/a_27_47# 2.99e-20
C6056 clkbuf_0_clk/a_110_47# _195_/a_76_199# 0.011f
C6057 _104_ calibrate 0.145f
C6058 _292_/a_78_199# _292_/a_493_297# 3.15e-19
C6059 _337_/a_27_47# _244_/a_27_297# 4.58e-20
C6060 output40/a_27_47# net40 0.246f
C6061 _295_/a_113_47# _131_ 0.00951f
C6062 _097_ net30 4.53e-21
C6063 _053_ _098_ 4.65e-21
C6064 _110_ net37 5.19e-20
C6065 _071_ clknet_2_3__leaf_clk 7.99e-20
C6066 _123_ _065_ 0.0142f
C6067 _337_/a_1462_47# _075_ 6.2e-19
C6068 _125_ _299_/a_27_413# 1.04e-19
C6069 _101_ _076_ 0.036f
C6070 _185_/a_68_297# _051_ 1.82e-20
C6071 VPWR _316_/a_761_289# 0.213f
C6072 net28 _158_/a_68_297# 0.0184f
C6073 _041_ _077_ 5.12e-20
C6074 net12 _228_/a_79_21# 0.00707f
C6075 _259_/a_109_297# trim_mask\[1\] 1.38e-20
C6076 _093_ _096_ 0.119f
C6077 _324_/a_761_289# _324_/a_805_47# 3.69e-19
C6078 _324_/a_193_47# _324_/a_1217_47# 2.36e-20
C6079 _324_/a_543_47# _324_/a_639_47# 0.0138f
C6080 _306_/a_27_47# _073_ 2.64e-20
C6081 calibrate net55 0.404f
C6082 net13 mask\[4\] 0.0131f
C6083 net13 _322_/a_639_47# 0.00121f
C6084 _300_/a_129_47# net16 4.35e-20
C6085 _104_ net45 2.79e-21
C6086 state\[2\] _048_ 0.0104f
C6087 _103_ _227_/a_209_311# 0.046f
C6088 _104_ rebuffer3/a_75_212# 2.43e-21
C6089 _316_/a_1283_21# net41 0.0673f
C6090 _322_/a_448_47# _040_ 2.36e-19
C6091 _232_/a_32_297# _243_/a_109_297# 8.58e-19
C6092 _053_ clknet_0_clk 0.0952f
C6093 _329_/a_27_47# _259_/a_27_297# 7.3e-21
C6094 cal_itt\[2\] trim_mask\[0\] 1.07e-20
C6095 VPWR _079_ 0.122f
C6096 _309_/a_651_413# net43 0.0149f
C6097 _309_/a_1283_21# net23 0.00142f
C6098 net45 net55 1.01e-19
C6099 VPWR trimb[3] 0.553f
C6100 net13 _220_/a_199_47# 2.21e-20
C6101 _325_/a_543_47# net21 0.00162f
C6102 net14 _310_/a_761_289# 0.0115f
C6103 _258_/a_27_297# _327_/a_27_47# 2.01e-21
C6104 _116_ net46 3.1e-19
C6105 _117_ _027_ 1.84e-20
C6106 _327_/a_543_47# trim_mask\[0\] 5.05e-19
C6107 _327_/a_27_47# _024_ 0.213f
C6108 _053_ _304_/a_651_413# 0.00352f
C6109 _238_/a_75_212# clknet_2_0__leaf_clk 0.00103f
C6110 mask\[7\] _314_/a_543_47# 0.00299f
C6111 _305_/a_1108_47# _002_ 0.0343f
C6112 _283_/a_75_212# _034_ 0.109f
C6113 comp _133_ 5.22e-20
C6114 _250_/a_27_297# _250_/a_109_47# 0.00393f
C6115 net9 _300_/a_285_47# 8.04e-19
C6116 net42 wire42/a_75_212# 0.147f
C6117 _152_/a_150_297# _044_ 4.96e-19
C6118 _232_/a_32_297# _232_/a_304_297# 0.00167f
C6119 trim_val\[3\] trim_mask\[4\] 3.15e-20
C6120 _051_ _088_ 2.97e-19
C6121 _320_/a_27_47# _076_ 2.2e-21
C6122 _190_/a_465_47# _190_/a_655_47# 0.0905f
C6123 en_co_clk net19 0.00479f
C6124 _321_/a_193_47# _247_/a_109_297# 1.21e-19
C6125 _248_/a_109_297# mask\[4\] 0.0105f
C6126 _322_/a_193_47# mask\[4\] 0.0011f
C6127 trim_mask\[0\] net35 0.012f
C6128 _095_ _092_ 0.533f
C6129 _322_/a_543_47# _322_/a_651_413# 0.0572f
C6130 _322_/a_761_289# _322_/a_1270_413# 2.6e-19
C6131 _322_/a_193_47# _322_/a_639_47# 2.28e-19
C6132 _104_ _105_ 8.7e-20
C6133 _065_ net55 7.5e-20
C6134 _250_/a_373_47# clknet_2_1__leaf_clk 2.72e-19
C6135 _251_/a_109_297# clknet_2_1__leaf_clk 1.3e-19
C6136 _320_/a_651_413# mask\[2\] 4.21e-20
C6137 _320_/a_1283_21# _017_ 3.61e-20
C6138 cal net14 0.0197f
C6139 net49 net33 1.57e-20
C6140 trim_val\[2\] _176_/a_27_47# 0.0044f
C6141 _078_ _315_/a_193_47# 1.25e-19
C6142 net22 _315_/a_543_47# 8.02e-19
C6143 trim_val\[1\] _112_ 0.00578f
C6144 trim_mask\[1\] net49 0.17f
C6145 _042_ clknet_2_1__leaf_clk 0.665f
C6146 output21/a_27_47# ctlp[7] 0.373f
C6147 _253_/a_299_297# _310_/a_1108_47# 6.39e-20
C6148 _290_/a_207_413# net33 0.00314f
C6149 _327_/a_448_47# _136_ 5.57e-19
C6150 trim_mask\[1\] _336_/a_543_47# 5.37e-21
C6151 _200_/a_209_47# _063_ 0.00187f
C6152 _105_ net55 0.112f
C6153 _329_/a_27_47# trim_mask\[1\] 8.3e-22
C6154 _336_/a_761_289# _336_/a_543_47# 0.21f
C6155 _336_/a_193_47# _336_/a_1283_21# 0.0424f
C6156 _336_/a_27_47# _336_/a_1108_47# 0.102f
C6157 _303_/a_651_413# mask\[4\] 4.61e-20
C6158 cal_itt\[0\] _338_/a_193_47# 6.21e-19
C6159 _040_ _246_/a_109_297# 7.16e-19
C6160 _050_ _260_/a_256_47# 0.00128f
C6161 _319_/a_543_47# _319_/a_1108_47# 7.99e-20
C6162 _319_/a_193_47# _319_/a_651_413# 0.0346f
C6163 VPWR _230_/a_59_75# 0.205f
C6164 _290_/a_27_413# _290_/a_207_413# 0.185f
C6165 result[4] _253_/a_384_47# 1.3e-20
C6166 mask\[3\] _101_ 0.341f
C6167 net16 _269_/a_299_297# 0.00983f
C6168 _237_/a_505_21# _048_ 0.0416f
C6169 trim_mask\[0\] _332_/a_761_289# 0.0255f
C6170 _119_ _027_ 6.44e-20
C6171 _293_/a_299_297# _293_/a_384_47# 1.48e-19
C6172 _211_/a_109_297# net30 5.38e-19
C6173 net43 mask\[4\] 9.74e-20
C6174 net43 _322_/a_639_47# 1.83e-20
C6175 _169_/a_109_53# net4 0.0193f
C6176 _074_ _078_ 0.166f
C6177 _303_/a_1108_47# _000_ 5.47e-21
C6178 _067_ _065_ 0.0259f
C6179 VPWR _299_/a_382_47# 3.78e-19
C6180 _065_ _070_ 0.657f
C6181 _243_/a_109_47# _096_ 0.00145f
C6182 _243_/a_109_297# net55 0.0477f
C6183 _090_ _075_ 6.42e-21
C6184 VPWR _098_ 0.184f
C6185 _322_/a_1283_21# _008_ 4.31e-20
C6186 _324_/a_1108_47# mask\[5\] 0.00427f
C6187 _317_/a_651_413# _316_/a_543_47# 3.6e-21
C6188 _292_/a_215_47# cal_count\[1\] 0.05f
C6189 _051_ _108_ 1.4e-20
C6190 _110_ _332_/a_651_413# 2.02e-20
C6191 _015_ _185_/a_68_297# 0.00565f
C6192 _188_/a_27_47# _187_/a_212_413# 0.00133f
C6193 clk cal 2.95e-20
C6194 mask\[0\] net45 0.203f
C6195 _328_/a_27_47# net46 0.301f
C6196 _110_ _053_ 4.68e-19
C6197 _267_/a_59_75# clknet_2_2__leaf_clk 0.0181f
C6198 VPWR clknet_0_clk 3.19f
C6199 _104_ _336_/a_1283_21# 0.0587f
C6200 ctln[1] _317_/a_27_47# 1.75e-20
C6201 _237_/a_505_21# _120_ 0.00182f
C6202 net13 _222_/a_199_47# 3.31e-21
C6203 _322_/a_1283_21# mask\[5\] 5.3e-21
C6204 _019_ _040_ 8.42e-20
C6205 _232_/a_304_297# net55 4.17e-20
C6206 _329_/a_193_47# _104_ 5.06e-20
C6207 _330_/a_805_47# net19 3.89e-19
C6208 trim_mask\[2\] _334_/a_1283_21# 4.78e-20
C6209 VPWR _304_/a_651_413# 0.143f
C6210 _050_ _107_ 0.0466f
C6211 _049_ _003_ 1.6e-19
C6212 _325_/a_27_47# net13 0.00283f
C6213 _104_ _239_/a_27_297# 1.47e-22
C6214 net13 en_co_clk 0.0537f
C6215 _089_ _052_ 0.00686f
C6216 _026_ fanout46/a_27_47# 4.89e-21
C6217 _053_ net47 0.0146f
C6218 mask\[0\] _065_ 6.95e-19
C6219 _266_/a_68_297# net46 2.34e-20
C6220 net23 _246_/a_109_297# 7.55e-20
C6221 _200_/a_303_47# net19 0.00109f
C6222 _304_/a_543_47# _286_/a_76_199# 3.01e-20
C6223 _251_/a_109_47# mask\[6\] 0.00286f
C6224 clknet_2_0__leaf_clk output30/a_27_47# 0.0847f
C6225 _250_/a_109_297# _021_ 0.0018f
C6226 _288_/a_59_75# _297_/a_47_47# 0.00179f
C6227 _308_/a_761_289# mask\[1\] 5.96e-19
C6228 _321_/a_193_47# _018_ 0.223f
C6229 _328_/a_448_47# _058_ 0.00115f
C6230 _309_/a_1108_47# mask\[2\] 6.47e-20
C6231 _239_/a_277_297# net42 2.29e-19
C6232 _022_ clknet_2_1__leaf_clk 0.144f
C6233 _341_/a_193_47# net46 0.0241f
C6234 _088_ _242_/a_79_21# 1.81e-20
C6235 _194_/a_113_297# _067_ 0.103f
C6236 mask\[0\] _319_/a_27_47# 0.23f
C6237 _272_/a_299_297# _114_ 2.49e-19
C6238 _309_/a_27_47# _212_/a_113_297# 1.24e-20
C6239 _040_ _208_/a_218_47# 3.98e-20
C6240 net24 clkbuf_2_1__f_clk/a_110_47# 0.00181f
C6241 net12 _053_ 0.00965f
C6242 _321_/a_27_47# net26 4.33e-20
C6243 _320_/a_651_413# mask\[1\] 0.0278f
C6244 clkbuf_2_2__f_clk/a_110_47# net30 5.18e-19
C6245 _200_/a_303_47# _107_ 8.43e-20
C6246 _336_/a_1283_21# _336_/a_1462_47# 0.0074f
C6247 _336_/a_1108_47# _336_/a_1217_47# 0.00742f
C6248 _079_ _315_/a_543_47# 8.18e-20
C6249 _336_/a_761_289# _106_ 6.44e-20
C6250 _040_ _017_ 0.0831f
C6251 net44 _311_/a_543_47# 0.156f
C6252 _107_ _228_/a_297_47# 7.76e-19
C6253 net13 _050_ 0.00894f
C6254 _334_/a_1108_47# _175_/a_68_297# 2.85e-20
C6255 _093_ _316_/a_761_289# 8.41e-20
C6256 _267_/a_59_75# trim_val\[0\] 3.87e-19
C6257 _117_ _032_ 0.278f
C6258 _327_/a_1283_21# _341_/a_1283_21# 1.03e-20
C6259 _235_/a_297_47# _337_/a_543_47# 1.22e-20
C6260 _329_/a_543_47# _329_/a_651_413# 0.0572f
C6261 _329_/a_761_289# _329_/a_1270_413# 2.6e-19
C6262 _329_/a_193_47# _329_/a_639_47# 2.28e-19
C6263 VPWR _321_/a_651_413# 0.143f
C6264 mask\[1\] _140_/a_68_297# 0.132f
C6265 _035_ _286_/a_76_199# 1.97e-19
C6266 output29/a_27_47# result[7] 0.159f
C6267 _073_ cal_itt\[3\] 0.0366f
C6268 _188_/a_27_47# net2 0.00103f
C6269 _167_/a_161_47# net15 1.04e-19
C6270 clknet_2_1__leaf_clk _313_/a_1283_21# 0.0609f
C6271 net43 _222_/a_199_47# 2.03e-19
C6272 _253_/a_81_21# net29 8.48e-19
C6273 _284_/a_150_297# _065_ 0.00156f
C6274 VPWR _337_/a_651_413# 0.143f
C6275 VPWR _047_ 0.374f
C6276 _286_/a_218_374# net18 7.07e-19
C6277 _281_/a_103_199# _281_/a_253_297# 0.0148f
C6278 trim[4] _136_ 7.1e-20
C6279 _300_/a_285_47# _122_ 9.84e-21
C6280 clknet_2_0__leaf_clk _316_/a_1108_47# 2.11e-21
C6281 _014_ _316_/a_1283_21# 3.34e-20
C6282 net45 _316_/a_543_47# 0.156f
C6283 fanout43/a_27_47# _101_ 0.00344f
C6284 net34 _132_ 0.0169f
C6285 _074_ _004_ 0.136f
C6286 _325_/a_27_47# net43 0.308f
C6287 VPWR _110_ 3.18f
C6288 net5 _132_ 0.00278f
C6289 state\[2\] _169_/a_373_53# 1.35e-19
C6290 net43 en_co_clk 1.22e-20
C6291 state\[2\] net54 0.00408f
C6292 _101_ _311_/a_448_47# 2.57e-21
C6293 _058_ _333_/a_543_47# 0.00144f
C6294 _328_/a_1217_47# net46 0.00112f
C6295 net27 _101_ 1.61e-19
C6296 _337_/a_27_47# _192_/a_174_21# 1.43e-21
C6297 _008_ _083_ 0.129f
C6298 _058_ _265_/a_384_47# 1.18e-19
C6299 _182_/a_27_47# trim_val\[0\] 0.0344f
C6300 _064_ _033_ 0.00276f
C6301 fanout45/a_27_47# _317_/a_193_47# 1.34e-19
C6302 _329_/a_1108_47# net9 0.0115f
C6303 _301_/a_47_47# _332_/a_651_413# 5.55e-20
C6304 _012_ sample 3.98e-19
C6305 VPWR _245_/a_27_297# 0.213f
C6306 _327_/a_1270_413# clknet_2_2__leaf_clk 2.27e-20
C6307 VPWR _143_/a_150_297# 0.00128f
C6308 VPWR net47 2.15f
C6309 _262_/a_27_47# _098_ 1.07e-20
C6310 net28 _085_ 0.127f
C6311 _032_ _119_ 2.87e-21
C6312 _226_/a_27_47# _092_ 0.0669f
C6313 _299_/a_298_297# _132_ 8.29e-19
C6314 _341_/a_1283_21# _108_ 1.43e-20
C6315 net52 net51 0.229f
C6316 _325_/a_1217_47# net13 1.36e-19
C6317 _326_/a_193_47# _253_/a_299_297# 3.25e-19
C6318 _326_/a_761_289# _253_/a_81_21# 1.8e-19
C6319 _047_ _161_/a_68_297# 0.11f
C6320 VPWR _340_/a_1140_413# 0.00306f
C6321 _121_ net45 2.82e-20
C6322 _275_/a_299_297# trim_val\[3\] 0.00937f
C6323 _275_/a_81_21# trim_mask\[3\] 0.062f
C6324 _083_ mask\[5\] 0.00101f
C6325 _341_/a_27_47# _053_ 0.017f
C6326 _333_/a_27_47# _332_/a_543_47# 2.44e-21
C6327 _333_/a_27_47# _108_ 0.00562f
C6328 net23 _017_ 1.83e-20
C6329 trim_val\[3\] _178_/a_68_297# 0.191f
C6330 trim_val\[0\] net37 0.0153f
C6331 _158_/a_68_297# _085_ 1.59e-19
C6332 _323_/a_651_413# _068_ 1.1e-21
C6333 result[1] result[2] 0.0367f
C6334 _265_/a_81_21# _332_/a_761_289# 3.19e-19
C6335 _265_/a_299_297# _332_/a_193_47# 4.56e-20
C6336 _337_/a_1108_47# _049_ 0.0107f
C6337 clknet_0_clk _262_/a_27_47# 0.00311f
C6338 output23/a_27_47# _004_ 9.22e-20
C6339 _125_ _297_/a_285_47# 1.08e-20
C6340 _337_/a_543_47# net30 1.27e-19
C6341 net43 _050_ 1.75e-20
C6342 _335_/a_543_47# trim_mask\[4\] 4.33e-20
C6343 _270_/a_59_75# net49 3.31e-19
C6344 trim_mask\[0\] _227_/a_296_53# 4.03e-19
C6345 _341_/a_1462_47# net46 0.00225f
C6346 VPWR net12 1.57f
C6347 _121_ _065_ 0.273f
C6348 _306_/a_27_47# _101_ 0.01f
C6349 mask\[0\] _319_/a_1217_47# 8.79e-19
C6350 _309_/a_1108_47# mask\[1\] 1.15e-19
C6351 _333_/a_1270_413# net46 2.06e-19
C6352 output36/a_27_47# net33 0.0323f
C6353 net54 _237_/a_505_21# 1.53e-19
C6354 _307_/a_761_289# _039_ 0.00152f
C6355 _327_/a_27_47# _257_/a_27_297# 0.00109f
C6356 VPWR _331_/a_1108_47# 0.31f
C6357 _322_/a_27_47# mask\[3\] 0.307f
C6358 mask\[3\] _248_/a_27_297# 0.0669f
C6359 mask\[6\] _313_/a_1108_47# 2.19e-20
C6360 net12 net53 0.0178f
C6361 VPWR _159_/a_27_47# 0.243f
C6362 _307_/a_193_47# fanout43/a_27_47# 1.71e-21
C6363 _062_ _190_/a_215_47# 7.64e-19
C6364 _199_/a_193_297# _001_ 0.0158f
C6365 net27 _312_/a_448_47# 5.98e-20
C6366 _053_ clknet_2_2__leaf_clk 0.00227f
C6367 output37/a_27_47# _125_ 0.0117f
C6368 _311_/a_1108_47# net19 5.66e-19
C6369 cal_itt\[0\] _303_/a_761_289# 1.93e-19
C6370 _329_/a_1283_21# _026_ 1.29e-20
C6371 _233_/a_27_297# net14 0.00997f
C6372 _094_ _337_/a_639_47# 0.00511f
C6373 net13 _169_/a_301_53# 2.46e-19
C6374 _035_ cal_count\[0\] 2.29e-19
C6375 _059_ _089_ 0.0142f
C6376 net28 _314_/a_543_47# 0.0102f
C6377 result[6] _314_/a_193_47# 0.00342f
C6378 _309_/a_761_289# _310_/a_27_47# 1.76e-19
C6379 _309_/a_193_47# _310_/a_193_47# 8.2e-21
C6380 _093_ clknet_0_clk 3.8e-20
C6381 VPWR net44 3.87f
C6382 result[3] _216_/a_199_47# 5.04e-20
C6383 _043_ _150_/a_27_47# 0.194f
C6384 _087_ net41 1.99e-19
C6385 _281_/a_253_297# _120_ 6.75e-19
C6386 _281_/a_337_297# en_co_clk 0.00424f
C6387 _327_/a_1108_47# _109_ 2.67e-20
C6388 wire42/a_75_212# _098_ 0.191f
C6389 _133_ _132_ 0.00744f
C6390 _103_ _100_ 3.7e-20
C6391 net12 _306_/a_1270_413# 3.74e-20
C6392 _257_/a_27_297# _335_/a_27_47# 2.3e-20
C6393 net12 _009_ 8.32e-19
C6394 _326_/a_639_47# net14 0.00129f
C6395 _325_/a_1217_47# net43 2.95e-19
C6396 net43 net25 0.261f
C6397 _119_ _171_/a_27_47# 2.72e-19
C6398 _313_/a_193_47# _313_/a_543_47# 0.22f
C6399 _313_/a_27_47# _313_/a_1283_21# 0.0436f
C6400 net44 net53 0.123f
C6401 cal_itt\[2\] _190_/a_27_47# 0.0929f
C6402 clk _318_/a_193_47# 0.546f
C6403 _111_ clknet_2_3__leaf_clk 2.64e-20
C6404 clknet_0_clk wire42/a_75_212# 8.82e-22
C6405 net12 _318_/a_27_47# 8.01e-19
C6406 _000_ _076_ 1.78e-20
C6407 VPWR _301_/a_47_47# 0.341f
C6408 _208_/a_76_199# rebuffer5/a_161_47# 0.00349f
C6409 _023_ net26 0.0652f
C6410 _187_/a_27_413# trim_mask\[0\] 5.9e-21
C6411 _331_/a_193_47# _054_ 1.63e-22
C6412 net8 _272_/a_299_297# 6.57e-19
C6413 _331_/a_543_47# _049_ 1.15e-19
C6414 ctlp[6] net20 0.0904f
C6415 VPWR _338_/a_562_413# 0.00414f
C6416 VPWR _263_/a_79_21# 0.252f
C6417 _306_/a_1270_413# net44 2.98e-19
C6418 VPWR _341_/a_27_47# 0.456f
C6419 _304_/a_27_47# _123_ 1.94e-19
C6420 net44 _009_ 0.0049f
C6421 _326_/a_1108_47# _102_ 0.00202f
C6422 _326_/a_448_47# mask\[7\] 8.14e-20
C6423 _326_/a_1283_21# _023_ 4.1e-20
C6424 trim_mask\[0\] _268_/a_75_212# 6.85e-19
C6425 ctlp[5] net19 0.00847f
C6426 VPWR _274_/a_75_212# 0.281f
C6427 _214_/a_113_297# net15 1.13e-20
C6428 _333_/a_1217_47# _108_ 2.9e-19
C6429 _255_/a_27_47# _106_ 5.59e-19
C6430 net4 _318_/a_193_47# 1.57e-19
C6431 _294_/a_68_297# _288_/a_59_75# 1.56e-20
C6432 _041_ _286_/a_76_199# 0.0591f
C6433 net37 _131_ 0.00604f
C6434 _286_/a_76_199# _338_/a_1182_261# 7.41e-21
C6435 _067_ _278_/a_27_47# 6.89e-19
C6436 trim_val\[0\] _332_/a_651_413# 4.58e-20
C6437 _330_/a_27_47# _330_/a_193_47# 0.614f
C6438 net43 _314_/a_651_413# 0.0139f
C6439 clk _317_/a_639_47# 5.58e-19
C6440 net47 _300_/a_47_47# 1.31e-20
C6441 _315_/a_1283_21# net14 1.52e-19
C6442 clknet_2_3__leaf_clk rebuffer3/a_75_212# 1.9e-19
C6443 _110_ _029_ 1.78e-19
C6444 trim[1] _112_ 4.99e-21
C6445 _340_/a_476_47# net2 2.46e-19
C6446 _320_/a_193_47# net15 1.55e-19
C6447 _123_ _298_/a_292_297# 0.00285f
C6448 _319_/a_193_47# clknet_0_clk 0.00163f
C6449 cal_itt\[1\] _092_ 0.00235f
C6450 net3 en_co_clk 0.0269f
C6451 VPWR _320_/a_543_47# 0.197f
C6452 _052_ _092_ 3.03e-19
C6453 _097_ _316_/a_27_47# 0.00526f
C6454 VPWR clknet_2_2__leaf_clk 4.34f
C6455 net8 output9/a_27_47# 3.66e-19
C6456 mask\[1\] _246_/a_109_47# 7.12e-19
C6457 VPWR _260_/a_584_47# 4.8e-20
C6458 net43 _310_/a_543_47# 0.156f
C6459 _086_ net14 0.0147f
C6460 _336_/a_27_47# net18 7.34e-22
C6461 _198_/a_27_47# _072_ 8.68e-20
C6462 _232_/a_32_297# _337_/a_27_47# 5.83e-20
C6463 mask\[0\] _282_/a_68_297# 3.54e-19
C6464 _065_ clknet_2_3__leaf_clk 0.305f
C6465 VPWR _328_/a_805_47# 2.71e-19
C6466 _324_/a_193_47# net27 2.33e-19
C6467 _324_/a_543_47# _311_/a_1283_21# 0.00122f
C6468 _135_ clknet_2_3__leaf_clk 0.194f
C6469 _125_ _339_/a_1602_47# 1.71e-20
C6470 _323_/a_543_47# net26 8.13e-19
C6471 _015_ _317_/a_1283_21# 9.37e-19
C6472 _167_/a_161_47# state\[1\] 0.284f
C6473 _325_/a_27_47# _325_/a_543_47# 0.115f
C6474 _325_/a_193_47# _325_/a_761_289# 0.186f
C6475 cal_count\[1\] net37 6.29e-19
C6476 _305_/a_193_47# _198_/a_27_47# 6.08e-20
C6477 VPWR net11 0.572f
C6478 _064_ clkbuf_2_3__f_clk/a_110_47# 0.0533f
C6479 VPWR _307_/a_1283_21# 0.389f
C6480 VPWR _323_/a_805_47# 3.81e-19
C6481 fanout46/a_27_47# _280_/a_75_212# 0.0197f
C6482 _226_/a_27_47# _226_/a_197_47# 0.00167f
C6483 clknet_0_clk _202_/a_79_21# 2.29e-19
C6484 trim_val\[3\] _334_/a_27_47# 9.05e-23
C6485 _068_ _190_/a_655_47# 0.0412f
C6486 _313_/a_448_47# _313_/a_639_47# 4.61e-19
C6487 _050_ net3 0.148f
C6488 net9 _122_ 0.0809f
C6489 _080_ _212_/a_199_47# 0.00151f
C6490 mask\[7\] _074_ 0.156f
C6491 trimb[1] trimb[4] 0.0486f
C6492 _043_ _042_ 0.019f
C6493 net12 _318_/a_1217_47# 9.9e-20
C6494 _015_ _192_/a_174_21# 1.97e-19
C6495 _304_/a_27_47# _067_ 1.01e-19
C6496 net45 _245_/a_109_297# 0.0535f
C6497 net43 _039_ 0.0278f
C6498 _321_/a_761_289# _042_ 0.00526f
C6499 VPWR _209_/a_27_47# 0.396f
C6500 _189_/a_27_47# trim_mask\[0\] 3.41e-19
C6501 _005_ fanout43/a_27_47# 4.32e-19
C6502 cal_itt\[0\] _199_/a_193_297# 3.23e-19
C6503 trim_mask\[4\] _170_/a_81_21# 1.48e-20
C6504 _260_/a_93_21# _054_ 0.00149f
C6505 _260_/a_256_47# _049_ 0.00435f
C6506 _321_/a_448_47# clknet_2_1__leaf_clk 1.61e-19
C6507 VPWR _341_/a_1217_47# 3.07e-20
C6508 net47 _285_/a_113_47# 3.32e-19
C6509 trim[2] _055_ 1.84e-20
C6510 net34 net32 0.459f
C6511 VPWR _333_/a_651_413# 0.144f
C6512 _340_/a_476_47# _123_ 0.0324f
C6513 _041_ _072_ 5.23e-20
C6514 _189_/a_218_47# _051_ 0.00187f
C6515 clknet_0_clk _206_/a_27_93# 0.0422f
C6516 _041_ cal_count\[0\] 0.419f
C6517 VPWR trim_val\[0\] 0.354f
C6518 cal_count\[0\] _338_/a_1182_261# 0.00246f
C6519 _270_/a_59_75# _270_/a_145_75# 0.00658f
C6520 _008_ _311_/a_27_47# 0.279f
C6521 _330_/a_543_47# _330_/a_639_47# 0.0138f
C6522 _330_/a_193_47# _330_/a_1217_47# 2.36e-20
C6523 _330_/a_761_289# _330_/a_805_47# 3.69e-19
C6524 _077_ _076_ 0.0132f
C6525 _301_/a_47_47# _300_/a_47_47# 0.0163f
C6526 _194_/a_113_297# clknet_2_3__leaf_clk 0.0227f
C6527 _337_/a_193_47# _096_ 6.48e-19
C6528 _337_/a_27_47# net55 2.11e-19
C6529 net19 _049_ 1.21e-20
C6530 VPWR _308_/a_639_47# 7.36e-19
C6531 en_co_clk _062_ 0.114f
C6532 _237_/a_218_374# net15 1.97e-19
C6533 clknet_2_1__leaf_clk net14 0.0168f
C6534 state\[2\] _318_/a_543_47# 7.62e-19
C6535 _064_ _302_/a_109_297# 0.00114f
C6536 _341_/a_27_47# _300_/a_47_47# 1.01e-20
C6537 _125_ cal_count\[2\] 2.52e-20
C6538 fanout44/a_27_47# en_co_clk 1.91e-21
C6539 _305_/a_193_47# _041_ 7.19e-21
C6540 _264_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 4.03e-20
C6541 _307_/a_27_47# net30 1.97e-19
C6542 _262_/a_109_297# _063_ 8.95e-19
C6543 VPWR _237_/a_218_47# 4.61e-20
C6544 VPWR _309_/a_193_47# 0.291f
C6545 net45 _331_/a_448_47# 2.56e-19
C6546 _081_ net45 6.44e-20
C6547 net13 _235_/a_79_21# 0.0118f
C6548 net13 net15 0.00271f
C6549 _074_ _312_/a_27_47# 7.4e-19
C6550 VPWR _339_/a_956_413# 0.00405f
C6551 _143_/a_68_297# clknet_2_1__leaf_clk 4.36e-21
C6552 _328_/a_761_289# _030_ 7.31e-20
C6553 mask\[7\] _146_/a_150_297# 1.25e-20
C6554 _102_ _146_/a_68_297# 1.65e-19
C6555 trim_mask\[0\] _336_/a_27_47# 8.59e-20
C6556 _058_ _048_ 2.11e-19
C6557 VPWR ctln[7] 0.391f
C6558 _000_ _068_ 0.101f
C6559 en_co_clk _195_/a_76_199# 0.0344f
C6560 _107_ _049_ 0.0962f
C6561 _051_ _232_/a_32_297# 1.22e-21
C6562 output39/a_27_47# trimb[3] 0.34f
C6563 _161_/a_68_297# trim_val\[0\] 0.215f
C6564 VPWR _279_/a_204_297# 0.237f
C6565 net50 net46 0.0769f
C6566 _127_ _129_ 1.48e-19
C6567 _335_/a_27_47# _330_/a_193_47# 0.00461f
C6568 _259_/a_109_297# _119_ 1.16e-20
C6569 _051_ _336_/a_193_47# 0.00327f
C6570 net7 output6/a_27_47# 1.39e-19
C6571 output34/a_27_47# _334_/a_193_47# 2.12e-19
C6572 _211_/a_109_297# sample 3.96e-19
C6573 _004_ output30/a_27_47# 0.0445f
C6574 _050_ _062_ 0.504f
C6575 _293_/a_384_47# _125_ 0.0015f
C6576 _019_ _141_/a_27_47# 4.93e-20
C6577 VPWR _324_/a_1283_21# 0.371f
C6578 net31 output35/a_27_47# 0.00667f
C6579 _110_ _336_/a_1108_47# 0.0126f
C6580 _064_ cal_count\[3\] 0.297f
C6581 output14/a_27_47# result[6] 6.17e-19
C6582 ctlp[0] output28/a_27_47# 0.0347f
C6583 _050_ fanout44/a_27_47# 1.33e-21
C6584 calibrate _263_/a_382_297# 8.7e-21
C6585 _282_/a_68_297# _121_ 0.106f
C6586 _302_/a_109_47# _066_ 3.82e-20
C6587 _329_/a_761_289# _110_ 7.05e-19
C6588 _128_ _125_ 8.35e-19
C6589 VPWR net6 0.495f
C6590 _262_/a_27_47# clknet_2_2__leaf_clk 7.63e-20
C6591 state\[0\] _164_/a_161_47# 0.234f
C6592 _313_/a_639_47# _010_ 5e-19
C6593 _322_/a_193_47# net15 1.58e-21
C6594 _060_ _048_ 0.392f
C6595 _324_/a_1283_21# net53 2.43e-21
C6596 _321_/a_761_289# _022_ 7.48e-20
C6597 net8 _179_/a_27_47# 0.00169f
C6598 _323_/a_1108_47# _150_/a_27_47# 2.94e-19
C6599 _304_/a_1217_47# _067_ 1.37e-19
C6600 net45 _016_ 0.0528f
C6601 VPWR _322_/a_543_47# 0.197f
C6602 VPWR _248_/a_373_47# 3.11e-19
C6603 mask\[3\] _077_ 6.46e-21
C6604 _304_/a_193_47# _284_/a_68_297# 7.13e-21
C6605 VPWR _257_/a_373_47# 5.17e-20
C6606 _083_ _311_/a_761_289# 1.99e-20
C6607 _303_/a_761_289# net26 0.00133f
C6608 _059_ _092_ 0.289f
C6609 _308_/a_27_47# _074_ 0.0183f
C6610 mask\[0\] _337_/a_27_47# 7.17e-20
C6611 _029_ clknet_2_2__leaf_clk 0.0802f
C6612 net31 _125_ 0.00536f
C6613 _126_ _129_ 0.0109f
C6614 _113_ _333_/a_27_47# 0.0141f
C6615 _338_/a_193_47# _123_ 0.00678f
C6616 net13 _049_ 0.127f
C6617 ctln[7] _318_/a_27_47# 2.13e-19
C6618 net13 _318_/a_761_289# 0.00583f
C6619 _316_/a_193_47# _316_/a_1270_413# 1.46e-19
C6620 _316_/a_27_47# _316_/a_639_47# 3.82e-19
C6621 _316_/a_543_47# _316_/a_448_47# 0.0498f
C6622 _316_/a_761_289# _316_/a_651_413# 0.0977f
C6623 _316_/a_1283_21# _316_/a_1108_47# 0.234f
C6624 _248_/a_373_47# net53 0.00406f
C6625 VPWR _303_/a_639_47# 4.33e-19
C6626 net43 net15 0.0355f
C6627 _200_/a_303_47# _062_ 3.3e-19
C6628 net50 _335_/a_651_413# 0.0012f
C6629 trim_val\[3\] _335_/a_639_47# 2.33e-20
C6630 _104_ _051_ 0.00947f
C6631 net44 _319_/a_193_47# 4.35e-20
C6632 _210_/a_113_297# net14 0.00505f
C6633 _308_/a_193_47# clknet_2_0__leaf_clk 0.00336f
C6634 VPWR _131_ 0.563f
C6635 cal_count\[0\] _338_/a_1296_47# 9.23e-20
C6636 _340_/a_1602_47# net16 0.00324f
C6637 trim_mask\[0\] net42 3.74e-20
C6638 _330_/a_1108_47# net46 0.231f
C6639 _330_/a_448_47# _027_ 0.17f
C6640 _301_/a_377_297# _135_ 0.00605f
C6641 output32/a_27_47# net34 0.0191f
C6642 calibrate _028_ 1.24e-19
C6643 _341_/a_193_47# _065_ 0.0116f
C6644 trim[1] _188_/a_27_47# 8.91e-21
C6645 _341_/a_193_47# _135_ 0.00145f
C6646 _341_/a_1283_21# net2 0.00641f
C6647 _106_ _261_/a_113_47# 7.22e-21
C6648 _051_ net55 0.121f
C6649 _250_/a_109_297# _101_ 0.0119f
C6650 _306_/a_1108_47# _092_ 1.92e-19
C6651 _053_ _231_/a_161_47# 8.17e-19
C6652 net1 net3 8.1e-20
C6653 _320_/a_448_47# clknet_2_0__leaf_clk 0.00139f
C6654 _320_/a_1283_21# net45 4.09e-19
C6655 _107_ _262_/a_193_297# 0.00229f
C6656 VPWR _044_ 0.512f
C6657 VPWR _309_/a_1462_47# 3.65e-19
C6658 net45 _028_ 0.0288f
C6659 net34 clkc 0.00407f
C6660 net5 clkc 0.0669f
C6661 _328_/a_27_47# _112_ 2.47e-21
C6662 _328_/a_761_289# trim_mask\[1\] 0.0188f
C6663 _200_/a_209_47# cal_itt\[2\] 3.56e-19
C6664 _200_/a_80_21# cal_itt\[1\] 0.0396f
C6665 _200_/a_209_297# cal_itt\[0\] 0.066f
C6666 clknet_2_1__leaf_clk net52 0.743f
C6667 net51 _208_/a_76_199# 0.00203f
C6668 net12 _239_/a_277_297# 0.00306f
C6669 net9 _340_/a_381_47# 0.003f
C6670 output23/a_27_47# _308_/a_27_47# 0.0112f
C6671 _319_/a_27_47# _016_ 0.156f
C6672 _284_/a_68_297# net18 0.00837f
C6673 _319_/a_1283_21# _101_ 8.24e-20
C6674 _327_/a_1283_21# _267_/a_59_75# 0.0141f
C6675 _307_/a_448_47# _074_ 0.00471f
C6676 _241_/a_388_297# net30 3.79e-19
C6677 net4 _336_/a_448_47# 2.01e-20
C6678 _334_/a_27_47# _334_/a_1108_47# 0.102f
C6679 _334_/a_193_47# _334_/a_1283_21# 0.0424f
C6680 _334_/a_761_289# _334_/a_543_47# 0.21f
C6681 _329_/a_27_47# _328_/a_193_47# 9.64e-20
C6682 _314_/a_27_47# _314_/a_448_47# 0.0931f
C6683 _314_/a_193_47# _314_/a_1108_47# 0.125f
C6684 fanout46/a_27_47# _107_ 1.45e-20
C6685 net27 _156_/a_27_47# 3.71e-20
C6686 _228_/a_79_21# _088_ 0.0908f
C6687 _122_ _299_/a_27_413# 1.63e-20
C6688 net44 _202_/a_79_21# 0.00333f
C6689 _339_/a_1032_413# cal_count\[0\] 0.0796f
C6690 net12 _206_/a_27_93# 1.95e-19
C6691 _320_/a_1283_21# _065_ 0.00212f
C6692 _327_/a_27_47# _327_/a_193_47# 0.863f
C6693 _053_ _001_ 5.28e-19
C6694 net12 mask\[6\] 0.00824f
C6695 _053_ _166_/a_161_47# 0.0314f
C6696 VPWR cal_count\[1\] 1.03f
C6697 net25 _082_ 0.415f
C6698 _239_/a_694_21# _087_ 0.0132f
C6699 _307_/a_1108_47# net45 0.237f
C6700 _169_/a_215_311# _185_/a_68_297# 3.85e-19
C6701 result[0] net45 3.23e-19
C6702 net43 _049_ 0.006f
C6703 trim_mask\[0\] _168_/a_27_413# 1.5e-20
C6704 _302_/a_27_297# _284_/a_68_297# 5.22e-19
C6705 mask\[6\] _159_/a_27_47# 2.6e-19
C6706 _251_/a_373_47# _046_ 2.01e-19
C6707 _094_ _099_ 5.11e-20
C6708 _327_/a_27_47# _058_ 0.033f
C6709 _042_ net21 4.64e-20
C6710 _259_/a_373_47# clknet_2_2__leaf_clk 3.54e-21
C6711 _258_/a_27_297# net9 6.46e-19
C6712 net9 _024_ 2.6e-20
C6713 net9 _147_/a_27_47# 6.92e-19
C6714 net44 _206_/a_27_93# 2.28e-19
C6715 _056_ _175_/a_68_297# 0.105f
C6716 _218_/a_113_297# net26 0.0486f
C6717 _064_ trim_mask\[2\] 0.525f
C6718 output15/a_27_47# net52 1.33e-21
C6719 _325_/a_761_289# net27 3.28e-20
C6720 _267_/a_59_75# _108_ 9.5e-19
C6721 _168_/a_207_413# _051_ 0.21f
C6722 mask\[6\] net44 2.19e-21
C6723 _269_/a_81_21# _333_/a_448_47# 8.84e-19
C6724 trim_val\[1\] _333_/a_27_47# 0.008f
C6725 net15 _281_/a_337_297# 9.27e-19
C6726 _316_/a_543_47# _013_ 9.07e-19
C6727 net16 _041_ 0.0115f
C6728 _323_/a_1108_47# _042_ 0.0531f
C6729 _192_/a_476_47# _095_ 2.62e-21
C6730 _192_/a_27_47# _092_ 0.0198f
C6731 _309_/a_543_47# _074_ 0.00391f
C6732 _090_ _096_ 0.372f
C6733 _335_/a_27_47# _335_/a_193_47# 0.906f
C6734 _326_/a_805_47# net43 0.00316f
C6735 _032_ _057_ 3.05e-20
C6736 _007_ _310_/a_1108_47# 9.3e-21
C6737 output26/a_27_47# _310_/a_27_47# 0.0131f
C6738 _106_ _119_ 0.00412f
C6739 clk _033_ 2.05e-20
C6740 VPWR _231_/a_161_47# 0.582f
C6741 _263_/a_79_21# _206_/a_27_93# 4.86e-19
C6742 _015_ net55 0.00176f
C6743 trimb[1] net33 6.99e-19
C6744 _337_/a_27_47# _121_ 0.0509f
C6745 _021_ _101_ 1.28e-19
C6746 output10/a_27_47# net50 0.00167f
C6747 _309_/a_761_289# net45 1.46e-19
C6748 _182_/a_27_47# _108_ 0.00233f
C6749 VPWR trim_mask\[3\] 0.53f
C6750 _304_/a_193_47# clknet_0_clk 5.02e-20
C6751 _334_/a_651_413# net46 0.0122f
C6752 VPWR _208_/a_505_21# 0.166f
C6753 net28 _074_ 0.0147f
C6754 mask\[3\] _310_/a_1108_47# 0.00101f
C6755 net25 _310_/a_448_47# 4.37e-20
C6756 _082_ _310_/a_543_47# 9.92e-20
C6757 net24 _245_/a_27_297# 0.00126f
C6758 _053_ _181_/a_68_297# 5.41e-22
C6759 _290_/a_27_413# trimb[1] 0.00504f
C6760 _315_/a_193_47# _099_ 7.61e-21
C6761 _315_/a_761_289# _095_ 1.86e-20
C6762 _300_/a_285_47# cal_count\[2\] 1.85e-20
C6763 net2 _295_/a_113_47# 1.11e-19
C6764 net55 _242_/a_79_21# 0.048f
C6765 _327_/a_1108_47# net46 0.252f
C6766 net9 _338_/a_1032_413# 0.00191f
C6767 _336_/a_27_47# trim_mask\[4\] 0.229f
C6768 _336_/a_1108_47# clknet_2_2__leaf_clk 0.00144f
C6769 cal_itt\[1\] _195_/a_439_47# 9.57e-19
C6770 net13 state\[1\] 0.144f
C6771 cal_itt\[1\] _071_ 6.15e-19
C6772 result[1] _308_/a_1108_47# 3.76e-19
C6773 _329_/a_761_289# clknet_2_2__leaf_clk 4.82e-20
C6774 VPWR mask\[2\] 0.609f
C6775 _102_ _078_ 0.00123f
C6776 net34 _130_ 0.0128f
C6777 _304_/a_543_47# _304_/a_1108_47# 7.99e-20
C6778 _304_/a_193_47# _304_/a_651_413# 0.0346f
C6779 ctlp[1] _046_ 0.00205f
C6780 net5 _130_ 2.21e-19
C6781 _339_/a_652_21# _123_ 0.0317f
C6782 _048_ _227_/a_109_93# 0.0208f
C6783 _040_ net45 0.0264f
C6784 _149_/a_150_297# _043_ 4.96e-19
C6785 _190_/a_655_47# cal_itt\[3\] 3.11e-19
C6786 net4 _033_ 0.0333f
C6787 _334_/a_1108_47# _334_/a_1217_47# 0.00742f
C6788 _334_/a_1283_21# _334_/a_1462_47# 0.0074f
C6789 _340_/a_27_47# _304_/a_27_47# 0.00162f
C6790 VPWR _001_ 1.83f
C6791 net37 _108_ 1.02e-19
C6792 VPWR _166_/a_161_47# 0.629f
C6793 _065_ _205_/a_27_47# 0.246f
C6794 mask\[2\] net53 0.0021f
C6795 _327_/a_761_289# _327_/a_805_47# 3.69e-19
C6796 _327_/a_543_47# _327_/a_639_47# 0.0138f
C6797 _327_/a_193_47# _327_/a_1217_47# 2.36e-20
C6798 _235_/a_297_47# _048_ 0.0341f
C6799 _336_/a_651_413# net19 0.00269f
C6800 _254_/a_109_297# _107_ 6.64e-19
C6801 _335_/a_1108_47# net46 0.268f
C6802 _322_/a_1108_47# _074_ 6.87e-19
C6803 calibrate _095_ 0.00101f
C6804 net3 net15 0.0611f
C6805 _235_/a_79_21# net3 0.0348f
C6806 _293_/a_299_297# cal_count\[0\] 0.0903f
C6807 state\[0\] _185_/a_150_297# 0.00186f
C6808 net54 _060_ 0.214f
C6809 _306_/a_193_47# _076_ 0.0151f
C6810 _299_/a_298_297# _130_ 0.0553f
C6811 _299_/a_382_47# _129_ 5.63e-19
C6812 _040_ _065_ 8.69e-19
C6813 _304_/a_27_47# clknet_2_3__leaf_clk 0.469f
C6814 _333_/a_193_47# _173_/a_27_47# 1.92e-19
C6815 output26/a_27_47# output27/a_27_47# 0.00269f
C6816 _006_ _078_ 3.87e-19
C6817 clkbuf_2_1__f_clk/a_110_47# _283_/a_75_212# 2.04e-21
C6818 _309_/a_27_47# clknet_2_1__leaf_clk 0.264f
C6819 _327_/a_1217_47# _058_ 1.84e-19
C6820 net46 rebuffer2/a_75_212# 2.15e-19
C6821 net45 _095_ 0.0222f
C6822 _014_ _099_ 0.0885f
C6823 clknet_2_0__leaf_clk _092_ 0.144f
C6824 result[3] _074_ 6.03e-19
C6825 VPWR _330_/a_1283_21# 0.384f
C6826 _103_ clk 0.00537f
C6827 _332_/a_1283_21# net46 0.282f
C6828 _292_/a_215_47# net2 0.0383f
C6829 _328_/a_651_413# net9 0.00125f
C6830 _304_/a_1108_47# _035_ 3.54e-20
C6831 _033_ _063_ 1.18e-21
C6832 _137_/a_68_297# _039_ 0.106f
C6833 _336_/a_651_413# _107_ 5.99e-19
C6834 clknet_2_1__leaf_clk _155_/a_150_297# 0.00148f
C6835 _337_/a_193_47# clknet_0_clk 0.0128f
C6836 net48 _333_/a_193_47# 4.16e-21
C6837 _304_/a_651_413# net18 9.07e-20
C6838 _324_/a_193_47# _250_/a_109_297# 4.14e-19
C6839 _109_ net33 9.17e-21
C6840 _298_/a_215_47# _133_ 0.0104f
C6841 net24 net44 2.51e-21
C6842 trim_mask\[1\] _109_ 1.61e-20
C6843 _310_/a_193_47# _310_/a_1270_413# 1.46e-19
C6844 _310_/a_27_47# _310_/a_639_47# 0.00188f
C6845 _310_/a_543_47# _310_/a_448_47# 0.0498f
C6846 _310_/a_761_289# _310_/a_651_413# 0.0977f
C6847 _310_/a_1283_21# _310_/a_1108_47# 0.234f
C6848 _314_/a_193_47# _224_/a_113_297# 1.97e-19
C6849 mask\[4\] _150_/a_27_47# 0.049f
C6850 cal_itt\[0\] _053_ 0.037f
C6851 VPWR _325_/a_1108_47# 0.309f
C6852 _322_/a_1283_21# _065_ 0.00339f
C6853 _065_ _095_ 0.178f
C6854 _053_ _088_ 0.00465f
C6855 net21 _313_/a_1283_21# 0.00744f
C6856 _046_ _313_/a_448_47# 1.64e-19
C6857 _335_/a_543_47# _335_/a_639_47# 0.0138f
C6858 _335_/a_193_47# _335_/a_1217_47# 2.36e-20
C6859 _335_/a_761_289# _335_/a_805_47# 3.69e-19
C6860 net23 net45 0.0169f
C6861 _324_/a_543_47# clknet_2_1__leaf_clk 8.78e-19
C6862 net16 _333_/a_543_47# 0.0106f
C6863 output11/a_27_47# ctln[5] 0.16f
C6864 result[4] _310_/a_1108_47# 2.85e-19
C6865 net16 _265_/a_384_47# 8.6e-20
C6866 _311_/a_27_47# _311_/a_761_289# 0.0701f
C6867 _325_/a_1108_47# net53 2.71e-20
C6868 _048_ _054_ 1.46e-19
C6869 VPWR _181_/a_68_297# 0.16f
C6870 net35 _332_/a_1270_413# 8.41e-20
C6871 _058_ _332_/a_805_47# 4.09e-19
C6872 _304_/a_651_413# _302_/a_27_297# 9.19e-21
C6873 _048_ net30 0.468f
C6874 output23/a_27_47# result[3] 0.00101f
C6875 net9 _134_ 8.17e-20
C6876 _050_ _227_/a_209_311# 0.00104f
C6877 _189_/a_408_47# _092_ 0.00778f
C6878 net3 _049_ 0.0661f
C6879 clknet_2_0__leaf_clk _246_/a_109_297# 1.16e-20
C6880 _315_/a_1462_47# _099_ 5.67e-20
C6881 _130_ _133_ 3.75e-19
C6882 net9 _341_/a_1270_413# 9.87e-20
C6883 _336_/a_1217_47# trim_mask\[4\] 9.77e-19
C6884 output21/a_27_47# clknet_2_1__leaf_clk 7.72e-20
C6885 _330_/a_27_47# net30 6.12e-20
C6886 _304_/a_193_47# net47 0.0345f
C6887 _243_/a_27_297# _099_ 9.67e-21
C6888 _243_/a_109_297# _095_ 8.87e-21
C6889 _164_/a_161_47# calibrate 0.0444f
C6890 net43 _305_/a_805_47# 0.0019f
C6891 _256_/a_27_297# _256_/a_109_47# 0.00393f
C6892 _026_ _328_/a_448_47# 2.79e-19
C6893 net43 _250_/a_27_297# 4.17e-21
C6894 clk _316_/a_1270_413# 2.55e-20
C6895 _336_/a_448_47# _279_/a_396_47# 6.19e-19
C6896 VPWR _314_/a_193_47# 0.59f
C6897 net16 _339_/a_1032_413# 0.00115f
C6898 _308_/a_543_47# net22 5.67e-19
C6899 _308_/a_193_47# _078_ 0.00934f
C6900 VPWR mask\[1\] 2.43f
C6901 _332_/a_651_413# _108_ 0.00129f
C6902 _321_/a_543_47# _321_/a_1108_47# 7.99e-20
C6903 _321_/a_193_47# _321_/a_651_413# 0.0346f
C6904 _340_/a_193_47# _340_/a_652_21# 0.0849f
C6905 _340_/a_27_47# _340_/a_476_47# 0.211f
C6906 _332_/a_193_47# _332_/a_639_47# 2.28e-19
C6907 _332_/a_761_289# _332_/a_1270_413# 2.6e-19
C6908 _332_/a_543_47# _332_/a_651_413# 0.0572f
C6909 _136_ _298_/a_78_199# 0.00209f
C6910 VPWR _185_/a_68_297# 0.176f
C6911 net25 net29 7.99e-20
C6912 _053_ _108_ 0.00353f
C6913 _032_ _027_ 5.79e-20
C6914 _164_/a_161_47# net45 6.11e-19
C6915 _186_/a_109_297# _060_ 0.00175f
C6916 _292_/a_215_47# _123_ 0.025f
C6917 trim_mask\[0\] _098_ 0.00401f
C6918 _120_ net30 1.38e-19
C6919 _168_/a_27_413# trim_mask\[4\] 0.0309f
C6920 net43 _319_/a_543_47# 0.153f
C6921 net23 _319_/a_27_47# 6.85e-20
C6922 _041_ net40 5.18e-22
C6923 _110_ net18 0.0157f
C6924 _337_/a_543_47# _337_/a_1108_47# 7.99e-20
C6925 _337_/a_193_47# _337_/a_651_413# 0.0346f
C6926 output31/a_27_47# trim_val\[1\] 0.00829f
C6927 trim[0] _269_/a_81_21# 1.8e-19
C6928 net2 _199_/a_193_297# 3.07e-19
C6929 _333_/a_448_47# net32 6.05e-20
C6930 _297_/a_129_47# net40 0.00189f
C6931 _340_/a_1032_413# _133_ 0.0121f
C6932 _340_/a_476_47# clknet_2_3__leaf_clk 6.56e-19
C6933 _074_ _084_ 0.0777f
C6934 trim_mask\[0\] clknet_0_clk 0.00637f
C6935 _042_ _045_ 1.83e-21
C6936 _175_/a_68_297# _172_/a_68_297# 0.0129f
C6937 _326_/a_193_47# _007_ 1.42e-19
C6938 _333_/a_193_47# _172_/a_68_297# 3.32e-19
C6939 _308_/a_27_47# output30/a_27_47# 3.05e-21
C6940 _042_ _249_/a_109_297# 0.0425f
C6941 mask\[0\] _140_/a_68_297# 0.00105f
C6942 _338_/a_1032_413# _122_ 0.0012f
C6943 _076_ net30 0.0106f
C6944 _276_/a_59_75# _110_ 0.134f
C6945 VPWR _195_/a_218_374# 1.7e-19
C6946 _097_ _237_/a_218_374# 9.3e-19
C6947 clone1/a_27_47# _092_ 1.19e-19
C6948 VPWR cal_itt\[0\] 2.46f
C6949 net47 net18 0.283f
C6950 state\[2\] clone7/a_27_47# 9.29e-19
C6951 _324_/a_193_47# _021_ 0.234f
C6952 _239_/a_694_21# _099_ 1.37e-20
C6953 net42 _190_/a_27_47# 1.25e-19
C6954 VPWR _334_/a_448_47# 0.0857f
C6955 _326_/a_193_47# mask\[3\] 2.68e-20
C6956 _326_/a_761_289# net25 1.58e-19
C6957 VPWR _088_ 0.704f
C6958 _314_/a_651_413# net29 9.55e-19
C6959 VPWR _327_/a_1283_21# 0.411f
C6960 _307_/a_639_47# net22 9.4e-19
C6961 _307_/a_1270_413# mask\[0\] 4.86e-21
C6962 net47 _129_ 1.66e-19
C6963 _046_ _010_ 9.53e-19
C6964 _335_/a_448_47# _032_ 0.16f
C6965 _313_/a_193_47# _155_/a_68_297# 5.89e-21
C6966 _167_/a_161_47# fanout45/a_27_47# 1.28e-19
C6967 net1 output41/a_27_47# 0.189f
C6968 _299_/a_27_413# _297_/a_285_47# 4.23e-20
C6969 _062_ _049_ 0.0151f
C6970 _311_/a_1108_47# _311_/a_1270_413# 0.00645f
C6971 _311_/a_761_289# _311_/a_1217_47# 4.2e-19
C6972 _311_/a_543_47# _311_/a_805_47# 0.00171f
C6973 fanout44/a_27_47# _049_ 0.0028f
C6974 net50 rebuffer3/a_75_212# 0.109f
C6975 _042_ mask\[4\] 0.0476f
C6976 output10/a_27_47# _335_/a_1108_47# 2.48e-20
C6977 net47 _302_/a_27_297# 4.88e-20
C6978 _304_/a_805_47# _136_ 1.62e-19
C6979 trim_mask\[2\] net34 2.69e-19
C6980 _310_/a_543_47# net29 4.49e-22
C6981 net4 clkbuf_2_3__f_clk/a_110_47# 0.0209f
C6982 VPWR _335_/a_1283_21# 0.362f
C6983 _071_ _306_/a_1108_47# 1.73e-20
C6984 _253_/a_81_21# net14 0.00317f
C6985 clknet_2_0__leaf_clk _017_ 0.123f
C6986 _319_/a_639_47# _092_ 1.66e-20
C6987 trim[4] _332_/a_1108_47# 5.6e-19
C6988 calibrate _226_/a_27_47# 8.89e-21
C6989 _307_/a_27_47# sample 0.00361f
C6990 _304_/a_1462_47# net47 0.00288f
C6991 _326_/a_761_289# _314_/a_651_413# 1.09e-20
C6992 _076_ _072_ 0.00276f
C6993 _341_/a_27_47# _304_/a_193_47# 3.33e-21
C6994 _341_/a_193_47# _304_/a_27_47# 5.81e-21
C6995 _051_ clknet_2_3__leaf_clk 4.57e-19
C6996 _256_/a_109_297# _024_ 0.00732f
C6997 net54 _235_/a_297_47# 0.00733f
C6998 _340_/a_1182_261# net47 0.119f
C6999 net9 cal_count\[2\] 1.69e-20
C7000 _037_ _304_/a_761_289# 1.29e-19
C7001 _033_ _279_/a_396_47# 0.00101f
C7002 VPWR _314_/a_1462_47# 0.00178f
C7003 _012_ net3 2.04e-20
C7004 _043_ net4 1.61e-20
C7005 _065_ _208_/a_218_374# 0.00203f
C7006 VPWR _108_ 1.68f
C7007 VPWR _332_/a_543_47# 0.207f
C7008 _340_/a_476_47# _340_/a_586_47# 0.00807f
C7009 _340_/a_1032_413# _340_/a_956_413# 0.00212f
C7010 _340_/a_27_47# _340_/a_1224_47# 1.63e-19
C7011 _340_/a_652_21# _340_/a_796_47# 0.00196f
C7012 net2 _208_/a_439_47# 0.00537f
C7013 VPWR _244_/a_27_297# 0.404f
C7014 _293_/a_299_297# net16 0.00195f
C7015 net26 _310_/a_193_47# 8.49e-20
C7016 _327_/a_27_47# net30 9.27e-21
C7017 trim_mask\[0\] _047_ 2.97e-19
C7018 _305_/a_193_47# _076_ 6.5e-19
C7019 clkbuf_2_0__f_clk/a_110_47# en_co_clk 0.0217f
C7020 _308_/a_193_47# _004_ 1.44e-20
C7021 _291_/a_35_297# net33 0.00618f
C7022 VPWR _288_/a_145_75# 4.87e-19
C7023 _090_ _098_ 1.75e-19
C7024 _309_/a_1108_47# mask\[0\] 3.55e-19
C7025 _309_/a_1283_21# _078_ 0.0767f
C7026 _074_ _085_ 0.0914f
C7027 _259_/a_109_47# net50 9.28e-19
C7028 _064_ _275_/a_384_47# 8.95e-20
C7029 _104_ _275_/a_81_21# 6.99e-22
C7030 net3 state\[1\] 0.00998f
C7031 _259_/a_373_47# trim_mask\[3\] 0.00366f
C7032 _110_ trim_mask\[0\] 0.0683f
C7033 _326_/a_193_47# _310_/a_1283_21# 3.39e-19
C7034 _326_/a_761_289# _310_/a_543_47# 0.00116f
C7035 _326_/a_27_47# _310_/a_1108_47# 4.22e-22
C7036 _309_/a_193_47# net24 0.551f
C7037 _063_ clkbuf_2_3__f_clk/a_110_47# 0.0504f
C7038 _337_/a_193_47# net44 0.0282f
C7039 _303_/a_1462_47# _069_ 7.35e-20
C7040 _338_/a_193_47# clknet_2_3__leaf_clk 0.352f
C7041 _137_/a_68_297# _049_ 1.37e-19
C7042 VPWR _310_/a_1270_413# 5.57e-19
C7043 _037_ _298_/a_215_47# 0.00228f
C7044 clknet_2_1__leaf_clk _208_/a_76_199# 0.00533f
C7045 net43 _313_/a_193_47# 0.0345f
C7046 _133_ _297_/a_377_297# 0.00272f
C7047 _134_ _122_ 0.084f
C7048 net34 _175_/a_150_297# 2.58e-19
C7049 _113_ _267_/a_59_75# 6.11e-20
C7050 _333_/a_1283_21# _055_ 0.0274f
C7051 clknet_0_clk _090_ 9.53e-21
C7052 _042_ _020_ 0.0462f
C7053 _035_ _338_/a_1602_47# 6.62e-21
C7054 VPWR output19/a_27_47# 0.298f
C7055 _270_/a_59_75# _109_ 1.23e-19
C7056 _321_/a_1283_21# _101_ 0.0616f
C7057 _306_/a_543_47# net51 1.5e-19
C7058 _338_/a_562_413# net18 5.82e-19
C7059 _341_/a_27_47# net18 0.017f
C7060 _128_ net9 0.00665f
C7061 clkbuf_2_2__f_clk/a_110_47# net19 0.0269f
C7062 clkbuf_0_clk/a_110_47# clk 0.315f
C7063 clk cal_count\[3\] 1.09e-20
C7064 VPWR _031_ 0.426f
C7065 _134_ _299_/a_27_413# 4.24e-20
C7066 _301_/a_47_47# _129_ 6.02e-20
C7067 output34/a_27_47# _176_/a_27_47# 0.00787f
C7068 _337_/a_1283_21# _101_ 4.33e-21
C7069 _050_ clkbuf_2_0__f_clk/a_110_47# 0.0678f
C7070 net13 _313_/a_1462_47# 3.89e-20
C7071 net15 _247_/a_27_297# 0.00809f
C7072 _107_ _240_/a_109_297# 2.8e-19
C7073 _053_ _170_/a_299_297# 0.00863f
C7074 _339_/a_1032_413# net40 2.31e-19
C7075 clk _331_/a_27_47# 0.0236f
C7076 _169_/a_215_311# _318_/a_651_413# 8.32e-20
C7077 _110_ _191_/a_27_297# 4.33e-20
C7078 _198_/a_27_47# _198_/a_181_47# 0.00401f
C7079 _199_/a_109_297# _069_ 0.0097f
C7080 _314_/a_27_47# _086_ 0.00916f
C7081 _311_/a_543_47# net26 0.0301f
C7082 _271_/a_75_212# _058_ 0.00186f
C7083 _303_/a_193_47# fanout47/a_27_47# 2.48e-19
C7084 _306_/a_27_47# _306_/a_193_47# 0.906f
C7085 _074_ _314_/a_543_47# 0.00163f
C7086 clkbuf_0_clk/a_110_47# net4 0.0159f
C7087 net12 trim_mask\[0\] 5.52e-21
C7088 net4 cal_count\[3\] 0.0122f
C7089 _329_/a_761_289# trim_mask\[3\] 8.85e-19
C7090 _329_/a_193_47# net50 3.78e-20
C7091 _341_/a_27_47# _302_/a_27_297# 4.17e-19
C7092 clkbuf_2_2__f_clk/a_110_47# _107_ 0.00242f
C7093 trimb[2] trimb[3] 0.0408f
C7094 cal_itt\[2\] _262_/a_109_297# 7.66e-20
C7095 _326_/a_193_47# net27 3.19e-20
C7096 _287_/a_75_212# _339_/a_193_47# 4.91e-21
C7097 _331_/a_193_47# _331_/a_543_47# 0.223f
C7098 _331_/a_27_47# _331_/a_1283_21# 0.0435f
C7099 _339_/a_1602_47# _122_ 9.53e-20
C7100 _329_/a_27_47# _057_ 1.44e-20
C7101 _185_/a_68_297# _093_ 7.18e-20
C7102 VPWR _311_/a_805_47# 1.18e-19
C7103 _001_ _202_/a_79_21# 3.4e-20
C7104 _199_/a_193_297# _070_ 1.01e-19
C7105 clknet_2_2__leaf_clk net18 0.123f
C7106 _325_/a_27_47# _042_ 1.4e-19
C7107 net4 _331_/a_27_47# 1.01e-19
C7108 net47 _338_/a_652_21# 0.174f
C7109 _258_/a_27_297# _024_ 8.17e-20
C7110 _323_/a_543_47# clknet_2_3__leaf_clk 2.78e-20
C7111 _282_/a_68_297# _095_ 4.78e-19
C7112 _340_/a_1296_47# net47 0.00232f
C7113 _064_ en_co_clk 3.22e-20
C7114 _068_ net30 0.00285f
C7115 state\[0\] _317_/a_1108_47# 1.75e-19
C7116 _325_/a_1283_21# clknet_2_1__leaf_clk 5.54e-20
C7117 _253_/a_81_21# net52 1.82e-19
C7118 _311_/a_805_47# net53 2.96e-19
C7119 net47 _297_/a_47_47# 1.21e-19
C7120 trim_mask\[4\] _098_ 1.66e-20
C7121 _340_/a_1032_413# _037_ 1.39e-19
C7122 trim[0] net32 0.00352f
C7123 ctlp[7] _313_/a_1108_47# 1.83e-19
C7124 net43 result[2] 5.53e-20
C7125 _327_/a_1108_47# _111_ 0.00162f
C7126 _276_/a_59_75# clknet_2_2__leaf_clk 8.39e-22
C7127 _008_ _078_ 0.165f
C7128 VPWR output14/a_27_47# 0.432f
C7129 en_co_clk _100_ 8.95e-19
C7130 mask\[7\] _102_ 0.206f
C7131 clkbuf_0_clk/a_110_47# _063_ 0.013f
C7132 _110_ _328_/a_1283_21# 5.34e-21
C7133 cal_count\[3\] _063_ 0.168f
C7134 mask\[6\] mask\[2\] 1.18e-20
C7135 _337_/a_1462_47# net44 0.00312f
C7136 _302_/a_27_297# clknet_2_2__leaf_clk 2.3e-20
C7137 clknet_0_clk trim_mask\[4\] 0.0177f
C7138 _291_/a_285_297# _127_ 0.0557f
C7139 net2 net37 0.61f
C7140 _341_/a_1283_21# clknet_2_3__leaf_clk 0.0722f
C7141 calibrate _052_ 0.233f
C7142 _037_ cal_count\[3\] 4.07e-20
C7143 _336_/a_1283_21# _330_/a_1108_47# 8.54e-21
C7144 calibrate input1/a_75_212# 0.00115f
C7145 _336_/a_1108_47# _330_/a_1283_21# 1.45e-19
C7146 state\[0\] _192_/a_27_47# 1.55e-21
C7147 _030_ net46 0.0539f
C7148 net43 _313_/a_1462_47# 0.00196f
C7149 _329_/a_193_47# _330_/a_1108_47# 1.79e-21
C7150 fanout46/a_27_47# _335_/a_761_289# 0.00111f
C7151 _078_ mask\[5\] 0.281f
C7152 _276_/a_59_75# net11 9.67e-20
C7153 clkbuf_2_2__f_clk/a_110_47# _279_/a_27_47# 8.19e-20
C7154 VPWR _306_/a_1283_21# 0.377f
C7155 trim_mask\[0\] _301_/a_47_47# 3.95e-20
C7156 _051_ _266_/a_68_297# 4.76e-20
C7157 _340_/a_193_47# _339_/a_193_47# 4.41e-21
C7158 net15 net29 0.0176f
C7159 net45 _052_ 1.21e-19
C7160 clknet_2_1__leaf_clk _314_/a_27_47# 0.395f
C7161 _307_/a_193_47# _138_/a_27_47# 0.00105f
C7162 cal_itt\[0\] _285_/a_113_47# 6.84e-20
C7163 output22/a_27_47# net14 1.67e-19
C7164 _122_ cal_count\[2\] 0.224f
C7165 _068_ _072_ 0.015f
C7166 _288_/a_59_75# _132_ 9.11e-19
C7167 VPWR _170_/a_299_297# 0.238f
C7168 _029_ _108_ 0.104f
C7169 _029_ _332_/a_543_47# 5.32e-19
C7170 _050_ _100_ 8.69e-21
C7171 _195_/a_535_374# _065_ 1.25e-20
C7172 _146_/a_68_297# _310_/a_27_47# 4.56e-21
C7173 _316_/a_1283_21# _092_ 4.55e-19
C7174 _291_/a_285_297# _126_ 0.00108f
C7175 cal_itt\[1\] _065_ 0.00318f
C7176 _162_/a_27_47# _333_/a_1108_47# 0.00116f
C7177 ctlp[0] net29 4.27e-19
C7178 _323_/a_1283_21# net47 0.294f
C7179 _312_/a_761_289# net20 0.0042f
C7180 ctln[6] _331_/a_1270_413# 1.07e-21
C7181 _299_/a_27_413# cal_count\[2\] 0.0242f
C7182 _305_/a_193_47# _068_ 2.12e-20
C7183 _019_ _078_ 5.23e-20
C7184 _136_ _301_/a_285_47# 0.0495f
C7185 _141_/a_27_47# net45 0.0379f
C7186 _259_/a_27_297# net46 0.00358f
C7187 _259_/a_109_297# _027_ 0.00475f
C7188 _306_/a_761_289# _306_/a_805_47# 3.69e-19
C7189 _306_/a_193_47# _306_/a_1217_47# 2.36e-20
C7190 _306_/a_543_47# _306_/a_639_47# 0.0138f
C7191 _293_/a_299_297# net40 0.0103f
C7192 _071_ _305_/a_1108_47# 2.83e-19
C7193 VPWR _227_/a_368_53# 1.14e-19
C7194 _341_/a_543_47# _136_ 0.0067f
C7195 _235_/a_382_297# _235_/a_297_47# 8.13e-19
C7196 cal_itt\[1\] _105_ 4.25e-19
C7197 _035_ _339_/a_381_47# 9.09e-21
C7198 clkbuf_2_3__f_clk/a_110_47# _279_/a_396_47# 6.1e-19
C7199 net12 _090_ 0.0052f
C7200 _110_ _265_/a_81_21# 0.00533f
C7201 _331_/a_448_47# _331_/a_639_47# 4.61e-19
C7202 net7 _317_/a_27_47# 1.44e-20
C7203 net15 _317_/a_761_289# 0.0136f
C7204 _331_/a_543_47# _260_/a_93_21# 7.88e-19
C7205 VPWR net26 2.42f
C7206 _325_/a_1108_47# mask\[6\] 0.0417f
C7207 _325_/a_27_47# _022_ 0.396f
C7208 _317_/a_27_47# _317_/a_193_47# 0.9f
C7209 _326_/a_27_47# _326_/a_193_47# 0.889f
C7210 _097_ net3 5.88e-20
C7211 trim_mask\[0\] clknet_2_2__leaf_clk 0.0931f
C7212 trim_val\[1\] net37 8.1e-20
C7213 _306_/a_761_289# _049_ 4.88e-20
C7214 _169_/a_215_311# _232_/a_32_297# 1.86e-20
C7215 net25 _042_ 9.06e-19
C7216 _104_ _228_/a_79_21# 0.0025f
C7217 net47 _338_/a_1056_47# 0.00264f
C7218 _041_ _338_/a_1602_47# 2.1e-19
C7219 _338_/a_652_21# _338_/a_562_413# 9.35e-20
C7220 _338_/a_1182_261# _338_/a_1602_47# 0.144f
C7221 _338_/a_476_47# _338_/a_381_47# 0.0356f
C7222 VPWR _317_/a_1283_21# 0.353f
C7223 VPWR _326_/a_1283_21# 0.43f
C7224 _328_/a_27_47# _328_/a_543_47# 0.111f
C7225 _328_/a_193_47# _328_/a_761_289# 0.171f
C7226 _306_/a_27_47# net30 6.46e-21
C7227 _198_/a_27_47# net19 0.00225f
C7228 cal _315_/a_639_47# 3.17e-19
C7229 trim_mask\[2\] net4 9.27e-20
C7230 state\[0\] clknet_2_0__leaf_clk 2.17e-20
C7231 _128_ _122_ 0.0325f
C7232 _074_ _310_/a_805_47# 7.09e-19
C7233 output29/a_27_47# _314_/a_193_47# 0.00864f
C7234 net26 net53 0.132f
C7235 _331_/a_193_47# net19 0.00104f
C7236 _087_ _089_ 0.162f
C7237 _321_/a_27_47# _040_ 1.17e-21
C7238 net13 _337_/a_543_47# 0.014f
C7239 _228_/a_79_21# net55 3.8e-20
C7240 _051_ _028_ 0.156f
C7241 _110_ trim_mask\[4\] 0.0431f
C7242 _293_/a_81_21# _299_/a_298_297# 2.3e-21
C7243 cal_itt\[0\] _197_/a_113_297# 0.114f
C7244 _283_/a_75_212# clknet_0_clk 0.00409f
C7245 _040_ _337_/a_27_47# 4.82e-21
C7246 net31 _055_ 0.131f
C7247 VPWR _286_/a_535_374# 1e-19
C7248 clknet_0_clk _190_/a_27_47# 0.0106f
C7249 trim[0] output32/a_27_47# 1.44e-19
C7250 net33 net46 0.0155f
C7251 output31/a_27_47# trim[1] 0.00179f
C7252 _325_/a_543_47# _313_/a_193_47# 3.45e-20
C7253 _325_/a_193_47# _313_/a_543_47# 2.85e-21
C7254 _325_/a_761_289# _313_/a_761_289# 3.75e-20
C7255 VPWR _192_/a_174_21# 0.31f
C7256 trim_mask\[1\] net46 0.046f
C7257 net44 _312_/a_543_47# 0.155f
C7258 _312_/a_27_47# _312_/a_193_47# 0.897f
C7259 _078_ _017_ 1.16e-19
C7260 _061_ output35/a_27_47# 7.29e-19
C7261 _336_/a_761_289# net46 0.159f
C7262 _125_ cal_count\[0\] 0.504f
C7263 _227_/a_209_311# _049_ 0.0102f
C7264 net24 mask\[2\] 0.725f
C7265 _320_/a_27_47# _101_ 7.48e-21
C7266 _303_/a_761_289# clknet_2_3__leaf_clk 0.0429f
C7267 _053_ net2 8.1e-20
C7268 _329_/a_27_47# _027_ 2.54e-19
C7269 _320_/a_193_47# _041_ 0.00174f
C7270 cal_itt\[0\] _194_/a_199_47# 2.4e-19
C7271 _212_/a_113_297# net22 4.11e-19
C7272 _149_/a_150_297# mask\[4\] 5.78e-19
C7273 net47 _339_/a_476_47# 0.206f
C7274 cal_itt\[2\] _202_/a_382_297# 2.25e-19
C7275 _305_/a_543_47# net51 0.00137f
C7276 _257_/a_373_47# net18 1.51e-19
C7277 _257_/a_27_297# _256_/a_109_297# 8.48e-20
C7278 _075_ _206_/a_206_47# 0.00673f
C7279 _322_/a_27_47# _321_/a_1283_21# 1.92e-19
C7280 _321_/a_1283_21# _248_/a_27_297# 0.0186f
C7281 net48 _334_/a_27_47# 0.00996f
C7282 trim_val\[2\] _334_/a_761_289# 0.00131f
C7283 _323_/a_27_47# _323_/a_543_47# 0.115f
C7284 _323_/a_193_47# _323_/a_761_289# 0.181f
C7285 _002_ rebuffer4/a_27_47# 1.05e-19
C7286 VPWR _187_/a_212_413# 0.209f
C7287 _327_/a_27_47# _066_ 1.59e-20
C7288 _140_/a_68_297# _245_/a_109_297# 5.91e-20
C7289 _306_/a_193_47# cal_itt\[3\] 4.34e-19
C7290 _306_/a_27_47# _072_ 2.88e-19
C7291 _263_/a_79_21# _090_ 0.022f
C7292 _337_/a_27_47# _095_ 0.00525f
C7293 net50 _278_/a_27_47# 1.62e-19
C7294 _189_/a_218_47# _053_ 1.22e-19
C7295 _328_/a_27_47# _333_/a_27_47# 1.45e-19
C7296 trim_mask\[2\] _273_/a_145_75# 0.00278f
C7297 _319_/a_193_47# _244_/a_27_297# 3.22e-20
C7298 VPWR _318_/a_651_413# 0.136f
C7299 _315_/a_193_47# net41 2.66e-21
C7300 _041_ net19 0.013f
C7301 trim_mask\[0\] trim_val\[0\] 0.551f
C7302 _308_/a_27_47# _006_ 1.37e-20
C7303 _308_/a_761_289# _081_ 9.1e-22
C7304 _042_ _310_/a_543_47# 5.03e-21
C7305 _239_/a_27_297# _052_ 2.78e-19
C7306 _169_/a_215_311# net55 1.35e-20
C7307 _169_/a_109_53# _096_ 8.02e-19
C7308 _306_/a_27_47# _305_/a_193_47# 1.34e-19
C7309 _306_/a_193_47# _305_/a_27_47# 1.92e-19
C7310 net43 _321_/a_543_47# 0.188f
C7311 net12 trim_mask\[4\] 0.0958f
C7312 _129_ _131_ 0.00886f
C7313 clknet_2_1__leaf_clk _310_/a_651_413# 0.0278f
C7314 net12 output13/a_27_47# 0.00349f
C7315 _293_/a_81_21# _133_ 1.84e-20
C7316 _059_ calibrate 0.0092f
C7317 net43 _337_/a_543_47# 3.35e-20
C7318 _341_/a_805_47# _038_ 7.31e-19
C7319 cal_count\[3\] _279_/a_396_47# 9.29e-19
C7320 _331_/a_639_47# _028_ 0.00129f
C7321 _331_/a_805_47# clknet_2_2__leaf_clk 8.94e-20
C7322 _331_/a_1108_47# trim_mask\[4\] 0.0036f
C7323 _260_/a_93_21# _260_/a_256_47# 0.0114f
C7324 _317_/a_543_47# _317_/a_639_47# 0.0138f
C7325 _317_/a_193_47# _317_/a_1217_47# 2.36e-20
C7326 _317_/a_761_289# _317_/a_805_47# 3.69e-19
C7327 net9 _334_/a_543_47# 4.91e-19
C7328 _074_ net41 2.02e-19
C7329 _328_/a_1283_21# clknet_2_2__leaf_clk 0.0763f
C7330 _012_ output41/a_27_47# 9.78e-19
C7331 _341_/a_1108_47# _301_/a_47_47# 4.46e-20
C7332 _258_/a_373_47# trim_mask\[4\] 1.19e-19
C7333 _112_ rebuffer2/a_75_212# 1.37e-19
C7334 _326_/a_761_289# _326_/a_805_47# 3.69e-19
C7335 _326_/a_193_47# _326_/a_1217_47# 2.36e-20
C7336 _326_/a_543_47# _326_/a_639_47# 0.0138f
C7337 _337_/a_761_289# _034_ 3.46e-19
C7338 _327_/a_193_47# net9 9.64e-20
C7339 trim_mask\[1\] _332_/a_448_47# 1.91e-20
C7340 net49 _332_/a_1108_47# 2.02e-19
C7341 _136_ _109_ 0.00114f
C7342 trim_val\[2\] rebuffer1/a_75_212# 0.00255f
C7343 _341_/a_761_289# _341_/a_543_47# 0.21f
C7344 _341_/a_193_47# _341_/a_1283_21# 0.0424f
C7345 _341_/a_27_47# _341_/a_1108_47# 0.102f
C7346 _081_ _140_/a_68_297# 0.0504f
C7347 _059_ net45 1.18e-20
C7348 VPWR _113_ 0.355f
C7349 _336_/a_1108_47# _108_ 2.38e-19
C7350 _320_/a_1270_413# net44 1.7e-19
C7351 net47 _303_/a_543_47# 0.155f
C7352 _301_/a_47_47# _265_/a_81_21# 1.43e-20
C7353 _303_/a_27_47# _338_/a_27_47# 1.71e-19
C7354 _256_/a_27_297# _118_ 2.6e-19
C7355 _256_/a_109_297# trim_val\[4\] 9.23e-20
C7356 trim_mask\[0\] _279_/a_204_297# 0.0551f
C7357 _014_ net41 0.00917f
C7358 _309_/a_651_413# net14 0.00184f
C7359 state\[2\] _260_/a_250_297# 0.00858f
C7360 _094_ _192_/a_505_280# 5.63e-20
C7361 _273_/a_145_75# _115_ 5.76e-19
C7362 net16 rebuffer1/a_75_212# 0.0176f
C7363 _053_ _123_ 0.181f
C7364 _318_/a_27_47# _318_/a_651_413# 9.73e-19
C7365 _318_/a_761_289# _318_/a_1108_47# 0.0512f
C7366 _318_/a_193_47# _318_/a_448_47# 0.0594f
C7367 _340_/a_381_47# cal_count\[2\] 1.81e-20
C7368 _071_ _069_ 4.41e-20
C7369 net9 _058_ 0.0376f
C7370 clknet_2_1__leaf_clk _247_/a_109_297# 0.00436f
C7371 net27 _251_/a_27_297# 2.01e-19
C7372 cal_count\[1\] _129_ 0.0153f
C7373 _059_ _065_ 0.00213f
C7374 VPWR net2 2.05f
C7375 _312_/a_543_47# _312_/a_639_47# 0.0138f
C7376 _312_/a_193_47# _312_/a_1217_47# 2.36e-20
C7377 _312_/a_761_289# _312_/a_805_47# 3.69e-19
C7378 net43 _253_/a_299_297# 6.99e-20
C7379 _309_/a_1108_47# _245_/a_109_297# 6.06e-22
C7380 _312_/a_1108_47# net19 6.62e-19
C7381 _286_/a_505_21# _124_ 1.38e-20
C7382 calibrate _170_/a_384_47# 7.93e-19
C7383 VPWR _305_/a_1283_21# 0.349f
C7384 _329_/a_805_47# net46 0.00316f
C7385 _308_/a_27_47# _308_/a_193_47# 0.864f
C7386 _323_/a_448_47# net19 0.00137f
C7387 ctln[2] _057_ 0.0674f
C7388 _258_/a_27_297# _257_/a_27_297# 8.59e-20
C7389 _041_ _339_/a_381_47# 0.0194f
C7390 _025_ _256_/a_27_297# 2.61e-20
C7391 net47 _339_/a_1224_47# 4.9e-19
C7392 net34 en_co_clk 1.13e-19
C7393 _107_ _260_/a_93_21# 0.00214f
C7394 _192_/a_174_21# _192_/a_548_47# 0.00101f
C7395 net9 _332_/a_27_47# 4.94e-19
C7396 _307_/a_27_47# _307_/a_761_289# 0.0626f
C7397 net5 en_co_clk 6.94e-19
C7398 net13 _041_ 0.0129f
C7399 net24 mask\[1\] 0.00304f
C7400 VPWR _189_/a_218_47# 0.00252f
C7401 _304_/a_193_47# _001_ 0.236f
C7402 _333_/a_193_47# clknet_2_2__leaf_clk 8.94e-19
C7403 clkbuf_2_0__f_clk/a_110_47# net15 0.0194f
C7404 VPWR _315_/a_805_47# 4.89e-19
C7405 net35 net32 2.58e-19
C7406 _306_/a_1462_47# cal_itt\[3\] 6.42e-19
C7407 _104_ _053_ 0.802f
C7408 _329_/a_761_289# _031_ 1.76e-19
C7409 _328_/a_1108_47# _333_/a_448_47# 6.86e-21
C7410 net43 _198_/a_27_47# 7.84e-20
C7411 _265_/a_81_21# clknet_2_2__leaf_clk 0.00101f
C7412 _026_ _327_/a_27_47# 2.01e-20
C7413 _051_ _095_ 6.97e-20
C7414 _303_/a_1283_21# net4 0.00105f
C7415 _324_/a_193_47# _101_ 5.02e-20
C7416 _078_ _310_/a_27_47# 0.00749f
C7417 _036_ _340_/a_476_47# 6.1e-19
C7418 _053_ net55 0.0461f
C7419 _326_/a_543_47# _086_ 0.00197f
C7420 _326_/a_193_47# _011_ 0.00135f
C7421 clkbuf_2_2__f_clk/a_110_47# _330_/a_761_289# 0.00656f
C7422 output24/a_27_47# _310_/a_193_47# 5.71e-21
C7423 _303_/a_543_47# net44 5.09e-19
C7424 _306_/a_1108_47# _305_/a_651_413# 1.35e-19
C7425 _231_/a_161_47# net18 1.49e-19
C7426 _243_/a_27_297# net41 2.57e-19
C7427 _136_ _092_ 0.222f
C7428 _326_/a_448_47# _074_ 0.00612f
C7429 net30 cal_itt\[3\] 0.176f
C7430 _320_/a_27_47# _320_/a_1217_47# 2.56e-19
C7431 _320_/a_761_289# _320_/a_639_47# 3.16e-19
C7432 _119_ _279_/a_490_47# 3.7e-19
C7433 _309_/a_543_47# _006_ 5.1e-19
C7434 _323_/a_193_47# _303_/a_193_47# 7.45e-21
C7435 _323_/a_27_47# _303_/a_761_289# 1.76e-20
C7436 _323_/a_761_289# _303_/a_27_47# 9.42e-21
C7437 _309_/a_1108_47# _081_ 0.00126f
C7438 _033_ _335_/a_543_47# 1.35e-19
C7439 trim_mask\[3\] net18 0.692f
C7440 mask\[7\] _158_/a_150_297# 9.44e-19
C7441 _076_ _003_ 0.149f
C7442 net12 _249_/a_27_297# 0.00691f
C7443 _248_/a_27_297# _101_ 0.176f
C7444 _322_/a_27_47# _101_ 0.0181f
C7445 _339_/a_27_47# _339_/a_193_47# 0.549f
C7446 clknet_2_2__leaf_clk trim_mask\[4\] 0.559f
C7447 trim_mask\[4\] _260_/a_584_47# 1.83e-20
C7448 _322_/a_193_47# _041_ 1.44e-20
C7449 _306_/a_543_47# clknet_2_1__leaf_clk 1.07e-19
C7450 VPWR _232_/a_32_297# 0.367f
C7451 _317_/a_761_289# state\[1\] 2.01e-19
C7452 _317_/a_651_413# clknet_2_0__leaf_clk 0.0267f
C7453 _317_/a_1108_47# net45 0.245f
C7454 _317_/a_448_47# _014_ 0.16f
C7455 _305_/a_27_47# net30 4.23e-20
C7456 VPWR trim_val\[1\] 0.815f
C7457 net44 _283_/a_75_212# 3.92e-21
C7458 _321_/a_193_47# mask\[2\] 0.00833f
C7459 _262_/a_205_47# net30 1.49e-19
C7460 _315_/a_27_47# _315_/a_761_289# 0.0701f
C7461 _093_ _192_/a_174_21# 8.93e-19
C7462 calibrate _192_/a_27_47# 2.36e-20
C7463 _341_/a_1283_21# _341_/a_1462_47# 0.0074f
C7464 _341_/a_1108_47# _341_/a_1217_47# 0.00742f
C7465 VPWR _336_/a_193_47# 0.591f
C7466 _053_ _067_ 0.0272f
C7467 _110_ _275_/a_299_297# 0.0517f
C7468 _276_/a_145_75# trim_val\[3\] 1.39e-20
C7469 _276_/a_59_75# trim_mask\[3\] 2e-20
C7470 _116_ _275_/a_81_21# 0.115f
C7471 _001_ net18 0.00937f
C7472 _053_ _070_ 1.58e-19
C7473 _110_ _178_/a_68_297# 0.0586f
C7474 _024_ trim_val\[4\] 1.29e-20
C7475 VPWR _123_ 3.25f
C7476 _323_/a_193_47# _152_/a_68_297# 1.58e-20
C7477 _333_/a_193_47# _333_/a_651_413# 0.0346f
C7478 _333_/a_543_47# _333_/a_1108_47# 7.99e-20
C7479 clkbuf_2_0__f_clk/a_110_47# _049_ 0.0271f
C7480 _005_ _101_ 2.24e-20
C7481 net44 _249_/a_27_297# 2.04e-19
C7482 _270_/a_59_75# net46 1.89e-20
C7483 net43 _041_ 5.66e-19
C7484 trim_val\[0\] _333_/a_193_47# 1.49e-20
C7485 output14/a_27_47# output29/a_27_47# 0.00355f
C7486 clknet_2_1__leaf_clk _018_ 0.0945f
C7487 _297_/a_47_47# _131_ 3.37e-19
C7488 net28 _312_/a_193_47# 1.5e-20
C7489 _078_ _311_/a_761_289# 1.33e-20
C7490 net8 trim[3] 2.86e-19
C7491 _219_/a_109_297# _101_ 9.22e-19
C7492 _251_/a_109_297# net15 0.00109f
C7493 _074_ _315_/a_193_47# 0.0166f
C7494 _265_/a_81_21# trim_val\[0\] 0.189f
C7495 calibrate _315_/a_27_47# 0.00333f
C7496 cal_itt\[3\] _072_ 0.352f
C7497 net16 _125_ 0.0151f
C7498 _326_/a_27_47# _251_/a_27_297# 5.41e-21
C7499 _042_ net15 0.00595f
C7500 _327_/a_27_47# net40 8.8e-20
C7501 _324_/a_639_47# net44 0.00198f
C7502 output36/a_27_47# net36 0.218f
C7503 _324_/a_543_47# _312_/a_1283_21# 0.00141f
C7504 _063_ _190_/a_215_47# 0.131f
C7505 _334_/a_193_47# net34 2.5e-19
C7506 _324_/a_27_47# net19 3.72e-19
C7507 VPWR _251_/a_373_47# 3.06e-19
C7508 _048_ _337_/a_1108_47# 2.81e-21
C7509 net12 _218_/a_199_47# 1.39e-19
C7510 _308_/a_761_289# _308_/a_805_47# 3.69e-19
C7511 _308_/a_193_47# _308_/a_1217_47# 2.36e-20
C7512 _308_/a_543_47# _308_/a_639_47# 0.0138f
C7513 trim_mask\[2\] _257_/a_109_47# 4.58e-19
C7514 output21/a_27_47# net21 0.201f
C7515 net3 _337_/a_543_47# 1.35e-21
C7516 net15 _319_/a_448_47# 0.00961f
C7517 net4 mask\[4\] 1.18e-20
C7518 _060_ clone7/a_27_47# 0.078f
C7519 _192_/a_27_47# _065_ 0.131f
C7520 _014_ _315_/a_193_47# 0.00248f
C7521 clknet_2_0__leaf_clk _315_/a_761_289# 0.00145f
C7522 _089_ _099_ 9.94e-20
C7523 _087_ _092_ 0.0261f
C7524 _307_/a_543_47# _307_/a_805_47# 0.00171f
C7525 _307_/a_761_289# _307_/a_1217_47# 4.2e-19
C7526 _307_/a_1108_47# _307_/a_1270_413# 0.00645f
C7527 net45 _315_/a_27_47# 0.298f
C7528 _326_/a_543_47# clknet_2_1__leaf_clk 6.62e-19
C7529 _305_/a_27_47# _072_ 0.0117f
C7530 _305_/a_193_47# cal_itt\[3\] 6.76e-21
C7531 VPWR _104_ 1.95f
C7532 _249_/a_373_47# _101_ 5.79e-19
C7533 _235_/a_79_21# _100_ 3.23e-20
C7534 result[0] _307_/a_1270_413# 7.73e-21
C7535 VPWR _319_/a_1270_413# 7.67e-19
C7536 _322_/a_1270_413# net44 1.67e-20
C7537 _300_/a_47_47# net2 0.398f
C7538 _318_/a_1270_413# net45 1.7e-19
C7539 net27 _313_/a_543_47# 2.25e-20
C7540 _309_/a_27_47# _308_/a_1283_21# 6.42e-21
C7541 _309_/a_193_47# _308_/a_543_47# 8.5e-21
C7542 _113_ _029_ 5.19e-19
C7543 _159_/a_27_47# _220_/a_113_297# 1.62e-21
C7544 _276_/a_59_75# _330_/a_1283_21# 7.73e-20
C7545 _015_ _095_ 1.44e-20
C7546 _128_ _338_/a_1032_413# 2.37e-20
C7547 VPWR net55 1.78f
C7548 _325_/a_193_47# _321_/a_1108_47# 3.1e-20
C7549 _305_/a_27_47# _305_/a_193_47# 0.578f
C7550 VPWR _223_/a_109_297# 0.00643f
C7551 trim[1] _182_/a_27_47# 0.00212f
C7552 output32/a_27_47# net35 0.00348f
C7553 _078_ _310_/a_1217_47# 3.02e-19
C7554 _237_/a_76_199# _237_/a_218_374# 0.00557f
C7555 _314_/a_1108_47# _010_ 1.93e-21
C7556 cal_count\[1\] _297_/a_47_47# 5.21e-20
C7557 _061_ _300_/a_285_47# 2.76e-20
C7558 trim_mask\[0\] _231_/a_161_47# 0.0047f
C7559 _337_/a_448_47# en_co_clk 5.36e-19
C7560 calibrate clknet_2_0__leaf_clk 0.0216f
C7561 _074_ _014_ 1.05e-21
C7562 _303_/a_1108_47# net19 0.00455f
C7563 fanout45/a_27_47# net3 0.0249f
C7564 _238_/a_75_212# net41 1.43e-19
C7565 trim_mask\[3\] trim_mask\[0\] 3.32e-21
C7566 cal _316_/a_761_289# 2.1e-20
C7567 net1 _316_/a_193_47# 6.22e-20
C7568 _322_/a_1217_47# _101_ 2.21e-19
C7569 net2 _029_ 1.01e-24
C7570 _339_/a_193_47# _339_/a_586_47# 0.00127f
C7571 _270_/a_59_75# _332_/a_448_47# 4.39e-20
C7572 _263_/a_297_47# _092_ 0.0243f
C7573 _341_/a_761_289# _092_ 1.29e-21
C7574 trim[1] net37 0.0301f
C7575 clknet_2_0__leaf_clk net45 0.854f
C7576 net43 _307_/a_27_47# 4.95e-19
C7577 _005_ _307_/a_193_47# 4.58e-20
C7578 comp output5/a_27_47# 0.00409f
C7579 VPWR _067_ 0.829f
C7580 cal_itt\[1\] _304_/a_27_47# 1.28e-19
C7581 output13/a_27_47# ctln[7] 0.362f
C7582 cal_itt\[0\] _304_/a_193_47# 2.67e-20
C7583 VPWR _070_ 0.673f
C7584 VPWR _114_ 0.274f
C7585 _315_/a_1108_47# _315_/a_1270_413# 0.00645f
C7586 _315_/a_761_289# _315_/a_1217_47# 4.2e-19
C7587 _315_/a_543_47# _315_/a_805_47# 0.00171f
C7588 _337_/a_1108_47# _076_ 0.00105f
C7589 trim_mask\[4\] _279_/a_204_297# 5.72e-20
C7590 VPWR _336_/a_1462_47# 8.89e-19
C7591 VPWR ctlp[1] 0.348f
C7592 output23/a_27_47# _074_ 0.00436f
C7593 _190_/a_465_47# net19 0.00242f
C7594 _053_ _284_/a_150_297# 3.68e-19
C7595 _134_ cal_count\[2\] 0.0359f
C7596 VPWR _329_/a_639_47# 2.96e-19
C7597 net8 _334_/a_805_47# 4.44e-19
C7598 _313_/a_193_47# _221_/a_109_297# 6.1e-21
C7599 _321_/a_193_47# mask\[1\] 4.19e-21
C7600 _140_/a_68_297# _040_ 0.106f
C7601 _319_/a_1283_21# net30 1.19e-19
C7602 _303_/a_27_47# _303_/a_193_47# 0.584f
C7603 _038_ _193_/a_109_297# 0.00313f
C7604 _100_ _049_ 0.0119f
C7605 mask\[5\] _312_/a_27_47# 1.04e-19
C7606 clknet_2_0__leaf_clk _065_ 0.113f
C7607 mask\[6\] net26 1.39e-19
C7608 _313_/a_193_47# net29 0.0017f
C7609 net31 output37/a_27_47# 0.0146f
C7610 _323_/a_193_47# mask\[5\] 6.07e-19
C7611 _022_ net15 0.00821f
C7612 _048_ _229_/a_27_297# 0.00561f
C7613 cal_itt\[2\] clkbuf_2_3__f_clk/a_110_47# 0.00843f
C7614 _322_/a_651_413# _320_/a_1283_21# 2.66e-20
C7615 VPWR _168_/a_207_413# 0.166f
C7616 _326_/a_1283_21# mask\[6\] 2.47e-19
C7617 _300_/a_47_47# _123_ 7.17e-20
C7618 fanout44/a_27_47# _337_/a_543_47# 0.00143f
C7619 _212_/a_199_47# net14 3.92e-19
C7620 _257_/a_373_47# trim_mask\[4\] 1.57e-19
C7621 _051_ _226_/a_27_47# 0.0397f
C7622 clk en_co_clk 0.00988f
C7623 _324_/a_27_47# _324_/a_761_289# 0.0701f
C7624 _308_/a_448_47# _005_ 0.168f
C7625 _308_/a_1108_47# net43 0.264f
C7626 state\[0\] _316_/a_1283_21# 0.062f
C7627 _308_/a_761_289# net23 2.72e-19
C7628 VPWR mask\[0\] 1.44f
C7629 _015_ _164_/a_161_47# 0.0142f
C7630 _328_/a_448_47# _025_ 0.158f
C7631 net12 rebuffer5/a_161_47# 0.00721f
C7632 VPWR output24/a_27_47# 0.438f
C7633 net45 _315_/a_1217_47# 6.03e-19
C7634 _319_/a_27_47# clknet_2_0__leaf_clk 0.854f
C7635 _305_/a_1217_47# _072_ 5.94e-21
C7636 _189_/a_218_47# wire42/a_75_212# 8.25e-21
C7637 cal_itt\[0\] net18 4.6e-19
C7638 _339_/a_1602_47# cal_count\[2\] 8.14e-20
C7639 _327_/a_1283_21# net18 2.81e-19
C7640 net43 _320_/a_805_47# 7.98e-21
C7641 output35/a_27_47# net40 0.0147f
C7642 _323_/a_639_47# mask\[4\] 4.1e-19
C7643 _321_/a_1108_47# mask\[3\] 1.86e-21
C7644 _321_/a_448_47# net25 8.78e-21
C7645 net4 en_co_clk 0.125f
C7646 _093_ _232_/a_32_297# 0.37f
C7647 _305_/a_761_289# _305_/a_805_47# 3.69e-19
C7648 _305_/a_193_47# _305_/a_1217_47# 2.36e-20
C7649 _305_/a_543_47# _305_/a_639_47# 0.0138f
C7650 _110_ _267_/a_145_75# 5.4e-19
C7651 VPWR _313_/a_448_47# 0.0836f
C7652 _309_/a_193_47# _309_/a_448_47# 0.0594f
C7653 _309_/a_761_289# _309_/a_1108_47# 0.0512f
C7654 _309_/a_27_47# _309_/a_651_413# 9.73e-19
C7655 _312_/a_193_47# _084_ 2.63e-19
C7656 _110_ _334_/a_27_47# 0.00314f
C7657 net23 _140_/a_68_297# 0.17f
C7658 net44 rebuffer5/a_161_47# 6.17e-19
C7659 net31 _134_ 4.59e-22
C7660 _178_/a_68_297# clknet_2_2__leaf_clk 3.17e-20
C7661 _144_/a_27_47# net37 1.83e-21
C7662 _256_/a_109_297# _058_ 0.00327f
C7663 _322_/a_27_47# _248_/a_27_297# 2.75e-19
C7664 trim_mask\[0\] _181_/a_68_297# 0.0193f
C7665 trim_val\[3\] trim_mask\[2\] 3.18e-19
C7666 _305_/a_543_47# clknet_2_1__leaf_clk 6.69e-20
C7667 _104_ _262_/a_27_47# 8.47e-20
C7668 clk _050_ 0.0344f
C7669 input1/a_75_212# _013_ 2.53e-20
C7670 _335_/a_1283_21# net18 0.00776f
C7671 net25 net14 0.00744f
C7672 _259_/a_27_297# _259_/a_109_47# 0.00393f
C7673 VPWR _172_/a_150_297# 0.00191f
C7674 calibrate clone1/a_27_47# 0.0484f
C7675 net31 _333_/a_1283_21# 0.0177f
C7676 trim_mask\[1\] rebuffer3/a_75_212# 8.85e-19
C7677 _125_ net40 0.227f
C7678 _030_ _112_ 0.0213f
C7679 _262_/a_27_47# net55 0.133f
C7680 cal_itt\[1\] _304_/a_1217_47# 1.09e-19
C7681 VPWR _284_/a_150_297# 0.00135f
C7682 clkbuf_2_1__f_clk/a_110_47# clknet_2_1__leaf_clk 1.63f
C7683 _064_ fanout46/a_27_47# 0.00164f
C7684 clkbuf_2_1__f_clk/a_110_47# _319_/a_761_289# 0.00668f
C7685 _155_/a_150_297# _045_ 4.96e-19
C7686 _198_/a_27_47# _062_ 6.55e-20
C7687 _325_/a_27_47# net52 0.00612f
C7688 _325_/a_761_289# _101_ 1.37e-19
C7689 net42 _262_/a_109_297# 0.0131f
C7690 _128_ _339_/a_1602_47# 0.00794f
C7691 _036_ _339_/a_652_21# 2.56e-19
C7692 en_co_clk _063_ 0.0175f
C7693 _108_ net18 0.192f
C7694 _315_/a_1283_21# _096_ 8.71e-21
C7695 _050_ net4 0.773f
C7696 _294_/a_68_297# _131_ 0.0477f
C7697 _166_/a_161_47# _090_ 1.39e-20
C7698 _053_ _230_/a_145_75# 4.01e-19
C7699 _285_/a_113_47# _123_ 0.0096f
C7700 _058_ _302_/a_373_47# 3.46e-20
C7701 _037_ en_co_clk 3.09e-20
C7702 _303_/a_761_289# _303_/a_805_47# 3.69e-19
C7703 _303_/a_543_47# _303_/a_639_47# 0.0138f
C7704 _303_/a_193_47# _303_/a_1217_47# 2.36e-20
C7705 _135_ net33 2.17e-20
C7706 _103_ _170_/a_81_21# 3.65e-19
C7707 _087_ _226_/a_197_47# 3.03e-20
C7708 net15 _316_/a_193_47# 2.68e-19
C7709 net2 _202_/a_79_21# 0.0392f
C7710 cal_itt\[2\] clkbuf_0_clk/a_110_47# 0.0416f
C7711 _317_/a_27_47# _316_/a_27_47# 5.3e-21
C7712 net54 _337_/a_1108_47# 1.55e-20
C7713 _060_ _337_/a_1283_21# 3.9e-20
C7714 _292_/a_78_199# _292_/a_215_47# 0.0907f
C7715 _337_/a_193_47# _244_/a_27_297# 2.43e-20
C7716 _235_/a_297_47# clone7/a_27_47# 8.79e-20
C7717 _305_/a_1283_21# _202_/a_79_21# 0.0114f
C7718 _314_/a_651_413# net14 0.00311f
C7719 _101_ _077_ 0.00277f
C7720 _019_ _320_/a_1108_47# 5.18e-20
C7721 net24 net26 6.35e-21
C7722 _288_/a_59_75# _130_ 8.84e-22
C7723 VPWR _316_/a_543_47# 0.209f
C7724 net28 _158_/a_150_297# 3.76e-19
C7725 _326_/a_651_413# _078_ 9.07e-20
C7726 net34 output40/a_27_47# 0.0147f
C7727 _324_/a_543_47# _324_/a_805_47# 0.00171f
C7728 _324_/a_761_289# _324_/a_1217_47# 4.2e-19
C7729 _324_/a_1108_47# _324_/a_1270_413# 0.00645f
C7730 _093_ net55 0.0155f
C7731 _306_/a_27_47# _003_ 0.169f
C7732 net13 _322_/a_805_47# 5.18e-19
C7733 _306_/a_193_47# _073_ 0.00579f
C7734 _048_ net19 0.0218f
C7735 _300_/a_285_47# net16 2.73e-19
C7736 _302_/a_27_297# _108_ 6.25e-19
C7737 _103_ _227_/a_296_53# 1.66e-19
C7738 _316_/a_1108_47# net41 0.0403f
C7739 _238_/a_75_212# _074_ 1.47e-21
C7740 _158_/a_68_297# _158_/a_150_297# 0.00477f
C7741 output21/a_27_47# _045_ 0.0124f
C7742 clknet_0_clk net51 1.07e-20
C7743 _329_/a_193_47# _259_/a_27_297# 3.28e-19
C7744 _257_/a_27_297# trim_val\[4\] 0.00148f
C7745 cal_itt\[0\] trim_mask\[0\] 7.46e-19
C7746 _330_/a_27_47# net19 0.0187f
C7747 state\[1\] _100_ 0.0265f
C7748 _335_/a_27_47# _280_/a_75_212# 2.42e-20
C7749 _309_/a_1270_413# net43 1.7e-19
C7750 trim_mask\[0\] _088_ 0.0317f
C7751 _325_/a_1283_21# net21 0.0015f
C7752 net14 _310_/a_543_47# 0.00416f
C7753 _309_/a_1108_47# net23 0.00161f
C7754 _258_/a_109_297# _327_/a_27_47# 6.37e-21
C7755 _258_/a_27_297# _327_/a_193_47# 7.13e-19
C7756 _117_ net46 5.03e-19
C7757 _327_/a_1283_21# trim_mask\[0\] 0.129f
C7758 _327_/a_193_47# _024_ 0.303f
C7759 _324_/a_543_47# mask\[4\] 1.92e-20
C7760 net9 cal_count\[0\] 0.045f
C7761 _294_/a_68_297# cal_count\[1\] 4.41e-21
C7762 VPWR net8 0.557f
C7763 mask\[7\] _314_/a_1283_21# 0.00165f
C7764 _238_/a_75_212# _014_ 0.00786f
C7765 net55 wire42/a_75_212# 0.00638f
C7766 _305_/a_448_47# _002_ 0.183f
C7767 _053_ _340_/a_27_47# 0.00282f
C7768 VPWR _121_ 0.395f
C7769 _250_/a_27_297# _250_/a_373_47# 0.0134f
C7770 fanout44/a_27_47# _041_ 4.69e-21
C7771 _136_ net46 0.0557f
C7772 VPWR _010_ 0.372f
C7773 _048_ _107_ 0.176f
C7774 _250_/a_27_297# _042_ 5.22e-20
C7775 trim_mask\[3\] trim_mask\[4\] 0.352f
C7776 _051_ _052_ 0.0393f
C7777 _320_/a_27_47# _077_ 3.13e-20
C7778 _128_ cal_count\[2\] 0.00309f
C7779 _258_/a_27_297# _058_ 7.2e-19
C7780 _024_ _058_ 0.047f
C7781 _322_/a_27_47# _322_/a_1217_47# 2.56e-19
C7782 _322_/a_761_289# _322_/a_639_47# 3.16e-19
C7783 _248_/a_109_47# mask\[4\] 0.00184f
C7784 _322_/a_761_289# mask\[4\] 2.91e-20
C7785 _099_ _092_ 0.341f
C7786 _126_ _132_ 9.98e-21
C7787 _320_/a_1108_47# _017_ 1.49e-19
C7788 _320_/a_1270_413# mask\[2\] 1.03e-21
C7789 net1 net14 0.0299f
C7790 trim_mask\[1\] _112_ 0.216f
C7791 _272_/a_299_297# trim_mask\[1\] 1.52e-20
C7792 _259_/a_373_47# _104_ 0.00178f
C7793 _053_ clknet_2_3__leaf_clk 1.13f
C7794 trim_mask\[1\] _336_/a_1283_21# 3.51e-19
C7795 VPWR trim[1] 0.488f
C7796 _069_ _065_ 0.131f
C7797 _200_/a_303_47# _063_ 0.00116f
C7798 _336_/a_193_47# _336_/a_1108_47# 0.125f
C7799 _336_/a_27_47# _336_/a_448_47# 0.0897f
C7800 _322_/a_1283_21# _218_/a_113_297# 1.4e-19
C7801 _285_/a_113_47# _067_ 1.96e-20
C7802 _040_ _246_/a_109_47# 0.00443f
C7803 _050_ _260_/a_346_47# 8.98e-19
C7804 _319_/a_543_47# _319_/a_448_47# 0.0498f
C7805 _319_/a_27_47# _319_/a_639_47# 3.82e-19
C7806 _319_/a_193_47# _319_/a_1270_413# 1.46e-19
C7807 _319_/a_761_289# _319_/a_651_413# 0.0977f
C7808 _319_/a_1283_21# _319_/a_1108_47# 0.234f
C7809 net14 _039_ 0.00319f
C7810 VPWR _230_/a_145_75# 1.91e-19
C7811 net25 net52 3.65e-19
C7812 output26/a_27_47# _023_ 0.00178f
C7813 net16 _269_/a_384_47# 4.9e-19
C7814 _237_/a_218_374# _048_ 7.33e-19
C7815 _209_/a_27_47# rebuffer5/a_161_47# 0.0197f
C7816 _117_ _335_/a_651_413# 1.39e-19
C7817 _119_ net46 0.0655f
C7818 trim_mask\[0\] _332_/a_543_47# 0.00719f
C7819 trim_mask\[0\] _108_ 0.295f
C7820 _274_/a_75_212# _334_/a_27_47# 6.05e-21
C7821 _237_/a_76_199# net3 9.98e-19
C7822 _286_/a_76_199# _122_ 0.0652f
C7823 calibrate _078_ 2.42e-20
C7824 _303_/a_448_47# _000_ 0.16f
C7825 _185_/a_68_297# _090_ 1.5e-21
C7826 _243_/a_109_47# net55 8.55e-19
C7827 _059_ _337_/a_27_47# 2.77e-19
C7828 net13 _048_ 0.00631f
C7829 _322_/a_1108_47# _008_ 0.00155f
C7830 net15 _316_/a_1462_47# 2.71e-19
C7831 _324_/a_448_47# mask\[5\] 7.84e-20
C7832 _324_/a_543_47# _020_ 7.24e-20
C7833 _097_ clkbuf_2_0__f_clk/a_110_47# 2.21e-19
C7834 _239_/a_27_297# clone1/a_27_47# 7.83e-20
C7835 _292_/a_215_47# _036_ 0.00228f
C7836 clknet_2_2__leaf_clk _330_/a_639_47# 0.00497f
C7837 trim_mask\[4\] _330_/a_1283_21# 4.53e-19
C7838 _015_ _185_/a_150_297# 5.02e-19
C7839 clk net1 2.9e-20
C7840 trim[1] _161_/a_68_297# 2.18e-19
C7841 _078_ net45 0.412f
C7842 _107_ _076_ 2.89e-19
C7843 _328_/a_193_47# net46 0.0269f
C7844 _267_/a_145_75# clknet_2_2__leaf_clk 3.94e-19
C7845 _136_ _332_/a_448_47# 0.00156f
C7846 ctln[1] net7 0.0117f
C7847 _104_ _336_/a_1108_47# 0.0578f
C7848 _334_/a_27_47# clknet_2_2__leaf_clk 0.254f
C7849 _320_/a_193_47# mask\[3\] 9.22e-21
C7850 mask\[7\] output27/a_27_47# 1.11e-19
C7851 _074_ output30/a_27_47# 0.0204f
C7852 trim_mask\[2\] _334_/a_1108_47# 8.01e-19
C7853 VPWR _304_/a_1270_413# 7.67e-19
C7854 _187_/a_27_413# clkc 3.36e-19
C7855 result[7] clknet_2_1__leaf_clk 0.00252f
C7856 _325_/a_193_47# net13 0.00405f
C7857 _328_/a_1283_21# _327_/a_1283_21# 1.65e-19
C7858 VPWR _340_/a_27_47# 0.437f
C7859 net30 _073_ 0.348f
C7860 _090_ _088_ 1.46e-20
C7861 _078_ _065_ 0.274f
C7862 _282_/a_68_297# clknet_2_0__leaf_clk 0.0127f
C7863 net23 _246_/a_109_47# 3.31e-21
C7864 _197_/a_113_297# _067_ 0.0492f
C7865 _251_/a_373_47# mask\[6\] 0.00286f
C7866 _250_/a_109_47# _021_ 6.05e-20
C7867 _181_/a_68_297# trim_mask\[4\] 0.135f
C7868 _101_ _310_/a_1108_47# 1.33e-21
C7869 _308_/a_543_47# mask\[1\] 1.21e-19
C7870 _321_/a_761_289# _018_ 1.1e-20
C7871 _269_/a_81_21# _172_/a_68_297# 0.00128f
C7872 _328_/a_651_413# _058_ 5.41e-19
C7873 VPWR _144_/a_27_47# 0.242f
C7874 _239_/a_474_297# net42 3.84e-19
C7875 net13 _076_ 1.04e-20
C7876 VPWR clknet_2_3__leaf_clk 3.33f
C7877 _341_/a_761_289# net46 0.162f
C7878 _194_/a_199_47# _067_ 0.00191f
C7879 _052_ _242_/a_79_21# 0.154f
C7880 _246_/a_27_297# _246_/a_109_297# 0.171f
C7881 mask\[0\] _319_/a_193_47# 0.0252f
C7882 _078_ _319_/a_27_47# 1.06e-21
C7883 net55 _206_/a_27_93# 1.27e-19
C7884 _202_/a_79_21# _070_ 0.0951f
C7885 _309_/a_193_47# _212_/a_113_297# 2.38e-20
C7886 _040_ _208_/a_439_47# 2.37e-20
C7887 net12 net51 0.0437f
C7888 VPWR _153_/a_27_47# 0.293f
C7889 _321_/a_193_47# net26 1.99e-19
C7890 _320_/a_1270_413# mask\[1\] 4.37e-19
C7891 _307_/a_27_47# _137_/a_68_297# 3.94e-21
C7892 _336_/a_27_47# _033_ 0.168f
C7893 _321_/a_448_47# net15 0.00623f
C7894 _336_/a_543_47# _106_ 7.17e-19
C7895 clknet_2_3__leaf_clk net53 1.23e-20
C7896 _335_/a_27_47# net19 0.00104f
C7897 _255_/a_27_47# _105_ 1.18e-19
C7898 net44 _311_/a_1283_21# 0.284f
C7899 _328_/a_1283_21# _108_ 5.16e-21
C7900 _327_/a_27_47# _107_ 0.00192f
C7901 ctlp[1] output29/a_27_47# 1.47e-19
C7902 output15/a_27_47# result[7] 4.15e-20
C7903 calibrate _316_/a_1283_21# 5.86e-20
C7904 _093_ _316_/a_543_47# 5.04e-20
C7905 _189_/a_27_47# _103_ 1.28e-19
C7906 _329_/a_27_47# _329_/a_1217_47# 2.56e-19
C7907 _329_/a_761_289# _329_/a_639_47# 3.16e-19
C7908 VPWR _321_/a_1270_413# 7.5e-19
C7909 mask\[1\] _140_/a_150_297# 2.2e-19
C7910 _035_ _286_/a_505_21# 2.02e-20
C7911 cal_count\[0\] _122_ 0.0604f
C7912 _073_ _072_ 0.00309f
C7913 _003_ cal_itt\[3\] 2.56e-19
C7914 _218_/a_113_297# _083_ 0.0912f
C7915 _329_/a_1108_47# net16 6.01e-21
C7916 clknet_2_1__leaf_clk _313_/a_1108_47# 0.0614f
C7917 VPWR _337_/a_1270_413# 7.85e-19
C7918 _236_/a_109_297# _092_ 0.00351f
C7919 _059_ _337_/a_1217_47# 1.23e-19
C7920 _281_/a_103_199# _281_/a_337_297# 0.0101f
C7921 net15 net14 6.76e-20
C7922 _058_ _134_ 4.45e-19
C7923 clknet_2_0__leaf_clk _316_/a_448_47# 9.35e-19
C7924 _014_ _316_/a_1108_47# 0.00182f
C7925 net45 _316_/a_1283_21# 0.275f
C7926 net44 net51 0.158f
C7927 calibrate _004_ 2.09e-19
C7928 VPWR _116_ 0.299f
C7929 _059_ _051_ 0.0305f
C7930 _325_/a_193_47# net43 0.0382f
C7931 _048_ _118_ 3.3e-20
C7932 state\[2\] _060_ 1.84e-19
C7933 net43 _120_ 5.67e-20
C7934 cal_count\[0\] _299_/a_27_413# 4.7e-20
C7935 net9 _066_ 2.45e-20
C7936 _328_/a_1462_47# net46 0.00426f
C7937 _101_ _311_/a_651_413# 2.69e-21
C7938 _337_/a_27_47# _192_/a_27_47# 3.85e-20
C7939 ctlp[0] net14 0.0159f
C7940 fanout47/a_27_47# _065_ 1e-19
C7941 _034_ en_co_clk 5.03e-19
C7942 _329_/a_448_47# net9 0.00125f
C7943 _309_/a_27_47# net25 2.54e-19
C7944 _004_ net45 0.00493f
C7945 trim_mask\[4\] _088_ 1.03e-19
C7946 _134_ _332_/a_27_47# 2.04e-20
C7947 VPWR _245_/a_109_297# 0.194f
C7948 _173_/a_27_47# net32 0.129f
C7949 net9 net16 0.00341f
C7950 net43 _076_ 0.00837f
C7951 output16/a_27_47# net16 0.174f
C7952 _325_/a_1462_47# net13 4.27e-19
C7953 net13 mask\[3\] 0.109f
C7954 _326_/a_543_47# _253_/a_81_21# 0.00344f
C7955 _333_/a_27_47# rebuffer2/a_75_212# 4.72e-20
C7956 _175_/a_68_297# _108_ 0.0279f
C7957 _047_ _161_/a_150_297# 4.96e-19
C7958 _187_/a_212_413# _129_ 7.67e-22
C7959 VPWR _340_/a_586_47# 2.04e-19
C7960 net54 _107_ 9.96e-19
C7961 _275_/a_384_47# trim_val\[3\] 3.91e-19
C7962 _333_/a_193_47# _108_ 0.00776f
C7963 _275_/a_81_21# net50 0.00491f
C7964 _275_/a_299_297# trim_mask\[3\] 0.059f
C7965 mask\[5\] _084_ 0.143f
C7966 _068_ net19 0.276f
C7967 _341_/a_193_47# _053_ 0.0171f
C7968 _091_ net30 1.3e-19
C7969 VPWR net20 0.582f
C7970 trim_val\[3\] _178_/a_150_297# 1.12e-19
C7971 trim_mask\[3\] _178_/a_68_297# 0.103f
C7972 trim[2] trim_val\[2\] 0.00257f
C7973 _041_ rebuffer6/a_27_47# 0.0359f
C7974 output17/a_27_47# net17 0.174f
C7975 clk net15 0.0472f
C7976 _265_/a_81_21# _332_/a_543_47# 0.00114f
C7977 _265_/a_81_21# _108_ 0.00934f
C7978 _337_/a_448_47# _049_ 0.009f
C7979 net34 _176_/a_27_47# 0.0156f
C7980 _210_/a_113_297# net22 0.00758f
C7981 clknet_0_clk _262_/a_109_297# 0.00374f
C7982 _188_/a_27_47# net33 0.00552f
C7983 _304_/a_193_47# net2 1.14e-20
C7984 _335_/a_1283_21# trim_mask\[4\] 7.62e-19
C7985 _270_/a_145_75# net49 2.9e-19
C7986 _270_/a_59_75# _112_ 0.171f
C7987 net20 net53 3.24e-20
C7988 trim_mask\[0\] _227_/a_368_53# 0.00514f
C7989 trim[2] net16 4.03e-19
C7990 _306_/a_193_47# _101_ 0.00382f
C7991 _246_/a_27_297# _017_ 0.117f
C7992 _246_/a_373_47# mask\[2\] 0.00122f
C7993 net3 _281_/a_103_199# 1.3e-20
C7994 mask\[0\] _319_/a_1462_47# 0.00198f
C7995 _050_ _034_ 2.82e-20
C7996 _138_/a_27_47# net30 9.28e-20
C7997 _333_/a_639_47# net46 0.00328f
C7998 _307_/a_543_47# _039_ 6.6e-19
C7999 VPWR _331_/a_448_47# 0.0844f
C8000 net4 net15 0.384f
C8001 _327_/a_193_47# _257_/a_27_297# 2.21e-20
C8002 VPWR _081_ 0.676f
C8003 _322_/a_193_47# mask\[3\] 0.625f
C8004 mask\[3\] _248_/a_109_297# 0.0051f
C8005 _325_/a_1283_21# mask\[4\] 3.75e-20
C8006 trim_mask\[4\] _108_ 0.183f
C8007 net20 _009_ 0.0217f
C8008 ctln[5] net11 0.0102f
C8009 VPWR _328_/a_27_47# 0.411f
C8010 _062_ _190_/a_465_47# 0.00215f
C8011 _053_ _028_ 2.45e-19
C8012 net27 _312_/a_651_413# 2.35e-19
C8013 _290_/a_207_413# output36/a_27_47# 2.71e-21
C8014 cal_itt\[0\] _303_/a_543_47# 1.64e-19
C8015 _071_ _303_/a_27_47# 1.33e-19
C8016 net2 _298_/a_493_297# 2.43e-20
C8017 _233_/a_109_297# net14 0.00183f
C8018 net27 net19 0.0249f
C8019 _329_/a_1108_47# _026_ 3.46e-19
C8020 _300_/a_47_47# clknet_2_3__leaf_clk 0.0435f
C8021 _094_ _337_/a_805_47# 0.00271f
C8022 net13 _169_/a_373_53# 6.93e-19
C8023 net13 net54 0.0449f
C8024 _337_/a_27_47# clknet_2_0__leaf_clk 0.404f
C8025 net28 _314_/a_1283_21# 2.21e-19
C8026 result[6] _314_/a_761_289# 4.99e-19
C8027 net43 _007_ 7.35e-19
C8028 _309_/a_543_47# _310_/a_27_47# 1.16e-20
C8029 _309_/a_27_47# _310_/a_543_47# 1.17e-20
C8030 _319_/a_193_47# _121_ 3.72e-20
C8031 output25/a_27_47# _082_ 3.65e-19
C8032 _262_/a_27_47# clknet_2_3__leaf_clk 1.87e-19
C8033 _257_/a_27_297# _058_ 3.18e-19
C8034 _281_/a_337_297# _120_ 8.29e-19
C8035 _281_/a_253_47# en_co_clk 0.0136f
C8036 _089_ net41 4.47e-19
C8037 net12 _306_/a_639_47# 0.00108f
C8038 _257_/a_27_297# _335_/a_193_47# 3.18e-22
C8039 clknet_2_0__leaf_clk _013_ 0.0347f
C8040 _326_/a_805_47# net14 6.71e-19
C8041 _189_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.01f
C8042 _168_/a_27_413# _033_ 2.41e-20
C8043 VPWR _323_/a_27_47# 0.484f
C8044 _325_/a_1462_47# net43 0.00196f
C8045 net43 mask\[3\] 0.0301f
C8046 net2 net18 0.0112f
C8047 _103_ net42 0.127f
C8048 VPWR _266_/a_68_297# 0.174f
C8049 _313_/a_27_47# _313_/a_1108_47# 0.102f
C8050 _313_/a_193_47# _313_/a_1283_21# 0.0423f
C8051 _313_/a_761_289# _313_/a_543_47# 0.21f
C8052 clk _049_ 0.483f
C8053 _051_ _203_/a_59_75# 7.77e-20
C8054 cal_itt\[2\] _190_/a_215_47# 0.12f
C8055 cal_itt\[0\] _190_/a_27_47# 2.61e-20
C8056 clk _318_/a_761_289# 0.0185f
C8057 _268_/a_75_212# cal_count\[3\] 2.44e-19
C8058 net15 net52 0.228f
C8059 net2 _129_ 0.0365f
C8060 net12 _318_/a_193_47# 8.6e-19
C8061 _051_ _192_/a_27_47# 3.56e-21
C8062 _323_/a_27_47# net53 0.00178f
C8063 _308_/a_1270_413# _039_ 1.6e-20
C8064 _026_ net9 0.0184f
C8065 _321_/a_27_47# _146_/a_68_297# 8.23e-19
C8066 VPWR _301_/a_377_297# 0.00924f
C8067 VPWR _016_ 0.714f
C8068 _048_ net3 1.05f
C8069 output8/a_27_47# trim_val\[2\] 1.29e-20
C8070 net8 _272_/a_384_47# 3.26e-19
C8071 VPWR _263_/a_382_297# 0.00532f
C8072 VPWR _338_/a_956_413# 0.0046f
C8073 _306_/a_639_47# net44 9.54e-19
C8074 VPWR _341_/a_193_47# 0.262f
C8075 net51 _209_/a_27_47# 0.00296f
C8076 _304_/a_193_47# _123_ 0.00196f
C8077 _326_/a_448_47# _102_ 3.52e-20
C8078 _326_/a_1108_47# _023_ 1.26e-19
C8079 _333_/a_1462_47# _108_ 3.59e-19
C8080 net4 _049_ 2.26e-19
C8081 _327_/a_27_47# _118_ 1.7e-20
C8082 _024_ net30 1.38e-20
C8083 output32/a_27_47# _173_/a_27_47# 5.36e-21
C8084 _050_ _281_/a_253_47# 8.07e-19
C8085 _041_ _286_/a_505_21# 0.0215f
C8086 _286_/a_505_21# _338_/a_1182_261# 6.11e-20
C8087 output8/a_27_47# net16 2.4e-20
C8088 _330_/a_27_47# _330_/a_761_289# 0.0535f
C8089 _304_/a_639_47# _065_ 1.91e-19
C8090 clk _317_/a_805_47# 2.74e-19
C8091 net43 _314_/a_1270_413# 3.18e-19
C8092 _227_/a_209_311# _260_/a_93_21# 4.03e-19
C8093 _100_ _240_/a_109_297# 6.37e-19
C8094 _315_/a_1108_47# net14 0.00637f
C8095 _340_/a_193_47# _065_ 1.53e-20
C8096 trim_val\[2\] _055_ 5.25e-19
C8097 net24 mask\[0\] 3.77e-20
C8098 _064_ clkbuf_2_2__f_clk/a_110_47# 2.53e-20
C8099 _340_/a_1182_261# net2 3.27e-20
C8100 output24/a_27_47# net24 0.221f
C8101 clknet_2_1__leaf_clk clknet_0_clk 0.00737f
C8102 _058_ trim_val\[4\] 0.0193f
C8103 _079_ _210_/a_113_297# 0.0909f
C8104 _319_/a_761_289# clknet_0_clk 0.00127f
C8105 net13 net27 0.074f
C8106 result[3] _310_/a_27_47# 0.00348f
C8107 net3 _120_ 2.04e-19
C8108 net27 _155_/a_68_297# 3.65e-20
C8109 _103_ _168_/a_27_413# 3.34e-21
C8110 net47 _132_ 4.97e-20
C8111 _136_ _111_ 0.0028f
C8112 VPWR _320_/a_1283_21# 0.366f
C8113 _097_ _316_/a_193_47# 0.00178f
C8114 net16 _055_ 8.2e-22
C8115 VPWR _028_ 0.442f
C8116 state\[2\] _227_/a_109_93# 8.42e-20
C8117 _327_/a_27_47# _025_ 5.29e-19
C8118 net43 _310_/a_1283_21# 0.337f
C8119 net27 output28/a_27_47# 1.41e-19
C8120 mask\[1\] _246_/a_373_47# 1.91e-20
C8121 _336_/a_193_47# net18 8.89e-21
C8122 mask\[6\] _010_ 3.7e-19
C8123 trim_mask\[0\] _113_ 3.43e-19
C8124 _232_/a_32_297# _337_/a_193_47# 3.63e-22
C8125 mask\[0\] _282_/a_150_297# 6.75e-20
C8126 _303_/a_651_413# _068_ 2.26e-19
C8127 VPWR _328_/a_1217_47# 1.2e-20
C8128 net52 _049_ 2.01e-19
C8129 _063_ _049_ 9.1e-20
C8130 _078_ _313_/a_639_47# 1.01e-19
C8131 _012_ net14 0.0159f
C8132 _324_/a_1283_21# _311_/a_1283_21# 3.86e-20
C8133 net16 _122_ 0.0236f
C8134 _101_ net30 4.32e-20
C8135 ctlp[6] _312_/a_27_47# 6.16e-19
C8136 _123_ net18 0.00946f
C8137 _320_/a_1283_21# net53 4.06e-21
C8138 _337_/a_639_47# net45 3.56e-20
C8139 net31 _058_ 5.96e-20
C8140 net43 result[4] 7.88e-19
C8141 net43 _068_ 1.05e-19
C8142 _015_ _317_/a_1108_47# 5.52e-19
C8143 _325_/a_27_47# _325_/a_1283_21# 0.0436f
C8144 _325_/a_193_47# _325_/a_543_47# 0.23f
C8145 net9 net40 0.0692f
C8146 _105_ _261_/a_113_47# 0.0096f
C8147 _051_ clknet_2_0__leaf_clk 3.44e-19
C8148 _110_ _269_/a_81_21# 0.00291f
C8149 _053_ _279_/a_314_297# 1.27e-20
C8150 _123_ _129_ 8.37e-20
C8151 _147_/a_27_47# cal_count\[0\] 2.04e-19
C8152 net4 _124_ 0.00181f
C8153 net16 _299_/a_27_413# 0.00306f
C8154 VPWR _307_/a_1108_47# 0.298f
C8155 _090_ _192_/a_174_21# 4.94e-20
C8156 net38 net33 0.126f
C8157 VPWR _323_/a_1217_47# 1.75e-19
C8158 trim_mask\[0\] net2 1.07e-20
C8159 _239_/a_474_297# _098_ 0.126f
C8160 _226_/a_27_47# _226_/a_303_47# 0.00119f
C8161 _042_ _035_ 2.32e-20
C8162 VPWR result[0] 0.335f
C8163 _136_ rebuffer3/a_75_212# 0.0027f
C8164 _313_/a_1108_47# _313_/a_1217_47# 0.00742f
C8165 _313_/a_1283_21# _313_/a_1462_47# 0.0074f
C8166 clkbuf_2_2__f_clk/a_110_47# _264_/a_27_297# 5.39e-21
C8167 _048_ _062_ 0.118f
C8168 _102_ _074_ 0.415f
C8169 net12 _318_/a_1462_47# 3.18e-19
C8170 _015_ _192_/a_27_47# 3.58e-20
C8171 _304_/a_193_47# _067_ 2.16e-19
C8172 _321_/a_543_47# _042_ 0.0026f
C8173 _218_/a_113_297# _311_/a_27_47# 3e-20
C8174 _104_ net18 0.0279f
C8175 _189_/a_218_47# trim_mask\[0\] 8.43e-21
C8176 _064_ _256_/a_27_297# 0.0912f
C8177 _277_/a_75_212# fanout46/a_27_47# 3e-19
C8178 net42 clkbuf_2_3__f_clk/a_110_47# 0.00341f
C8179 net43 fanout43/a_27_47# 0.35f
C8180 state\[0\] _099_ 3.09e-20
C8181 comp _131_ 0.00527f
C8182 _260_/a_346_47# _049_ 0.00256f
C8183 _321_/a_651_413# clknet_2_1__leaf_clk 0.0045f
C8184 VPWR _341_/a_1462_47# 6.25e-20
C8185 _136_ _065_ 0.0334f
C8186 net43 net27 0.021f
C8187 VPWR _333_/a_1270_413# 7.19e-19
C8188 fanout46/a_27_47# net4 0.208f
C8189 _136_ _135_ 0.189f
C8190 _340_/a_1182_261# _123_ 0.0391f
C8191 _275_/a_299_297# _335_/a_1283_21# 7.21e-20
C8192 _189_/a_408_47# _051_ 5.25e-20
C8193 clknet_0_clk _206_/a_206_47# 4.75e-19
C8194 cal_count\[0\] _338_/a_1032_413# 0.00966f
C8195 _008_ _311_/a_193_47# 0.301f
C8196 _330_/a_1108_47# _330_/a_1270_413# 0.00645f
C8197 _330_/a_761_289# _330_/a_1217_47# 4.2e-19
C8198 _330_/a_543_47# _330_/a_805_47# 0.00171f
C8199 clk state\[1\] 0.00418f
C8200 _074_ _006_ 0.274f
C8201 VPWR _308_/a_805_47# 4.2e-19
C8202 _194_/a_199_47# clknet_2_3__leaf_clk 5.14e-19
C8203 _337_/a_193_47# net55 1.84e-19
C8204 cal_count\[0\] _297_/a_285_47# 2.37e-20
C8205 en_co_clk _075_ 0.17f
C8206 state\[2\] _054_ 1.37e-20
C8207 _341_/a_193_47# _300_/a_47_47# 2.39e-19
C8208 _104_ _302_/a_27_297# 4.46e-22
C8209 state\[2\] _318_/a_1283_21# 0.0638f
C8210 state\[2\] net30 9.58e-20
C8211 calibrate _087_ 0.0116f
C8212 _307_/a_193_47# net30 1.28e-19
C8213 _262_/a_193_297# _063_ 0.0324f
C8214 net2 _297_/a_47_47# 0.00997f
C8215 VPWR _237_/a_439_47# 1.95e-19
C8216 VPWR _309_/a_761_289# 0.204f
C8217 net45 _331_/a_651_413# 0.0135f
C8218 VPWR _205_/a_27_47# 0.475f
C8219 _074_ _312_/a_193_47# 2.25e-19
C8220 clknet_2_1__leaf_clk _245_/a_27_297# 0.00291f
C8221 _097_ _316_/a_1462_47# 1.03e-19
C8222 trim_mask\[0\] trim_val\[1\] 8.27e-22
C8223 _067_ net18 0.0225f
C8224 VPWR _339_/a_1140_413# 0.00296f
C8225 net47 clknet_2_1__leaf_clk 6.21e-20
C8226 _328_/a_543_47# _030_ 2.04e-20
C8227 _328_/a_1283_21# _113_ 0.0215f
C8228 net4 state\[1\] 0.483f
C8229 en_co_clk _195_/a_505_21# 0.0307f
C8230 _161_/a_150_297# trim_val\[0\] 7.82e-19
C8231 cal_itt\[2\] en_co_clk 0.253f
C8232 _205_/a_27_47# net53 3.34e-19
C8233 VPWR _040_ 0.344f
C8234 _212_/a_113_297# mask\[1\] 0.0552f
C8235 net43 _306_/a_27_47# 1.21e-19
C8236 VPWR _279_/a_314_297# 0.0647f
C8237 output5/a_27_47# clkc 0.11f
C8238 _015_ clknet_2_0__leaf_clk 0.0843f
C8239 _325_/a_448_47# _325_/a_639_47# 4.61e-19
C8240 VPWR _292_/a_78_199# 0.278f
C8241 _051_ _336_/a_761_289# 1.05e-20
C8242 _057_ net46 1.95e-19
C8243 _050_ _075_ 0.059f
C8244 VPWR _324_/a_1108_47# 0.303f
C8245 _329_/a_543_47# _110_ 9.34e-19
C8246 _302_/a_373_47# _066_ 6.81e-19
C8247 _282_/a_150_297# _121_ 4.96e-19
C8248 mask\[4\] _311_/a_639_47# 0.00428f
C8249 _302_/a_27_297# _067_ 0.00366f
C8250 _051_ clone1/a_27_47# 5.88e-20
C8251 net12 clknet_2_1__leaf_clk 1.46f
C8252 net19 cal_itt\[3\] 4.96e-20
C8253 _313_/a_805_47# _010_ 2.14e-19
C8254 _120_ _137_/a_68_297# 2.11e-20
C8255 _033_ clknet_0_clk 0.00723f
C8256 _324_/a_1108_47# net53 1.86e-21
C8257 _321_/a_543_47# _022_ 8.25e-19
C8258 net54 net3 0.195f
C8259 _321_/a_27_47# _078_ 6.69e-19
C8260 _304_/a_1462_47# _067_ 4.31e-19
C8261 VPWR _322_/a_1283_21# 0.404f
C8262 _304_/a_761_289# _284_/a_68_297# 1.96e-20
C8263 VPWR _095_ 0.967f
C8264 net42 cal_count\[3\] 9.22e-20
C8265 _104_ trim_mask\[0\] 0.348f
C8266 _303_/a_543_47# net26 3.75e-20
C8267 _083_ _311_/a_543_47# 5.28e-20
C8268 clknet_2_1__leaf_clk _159_/a_27_47# 8.29e-20
C8269 _305_/a_639_47# net44 7.55e-19
C8270 _308_/a_193_47# _074_ 0.028f
C8271 mask\[0\] _337_/a_193_47# 5.23e-20
C8272 _113_ _333_/a_193_47# 6.65e-20
C8273 _030_ _333_/a_27_47# 0.381f
C8274 _092_ net41 5.14e-20
C8275 ctln[7] _318_/a_193_47# 3.63e-20
C8276 net13 _318_/a_543_47# 0.0122f
C8277 _316_/a_193_47# _316_/a_639_47# 2.28e-19
C8278 _316_/a_761_289# _316_/a_1270_413# 2.6e-19
C8279 _316_/a_543_47# _316_/a_651_413# 0.0572f
C8280 _322_/a_1283_21# net53 3.23e-20
C8281 trim_mask\[0\] net55 0.0775f
C8282 VPWR _303_/a_805_47# 2.3e-19
C8283 clknet_2_1__leaf_clk net44 0.0466f
C8284 net50 _335_/a_1270_413# 1.41e-19
C8285 trim_val\[3\] _335_/a_805_47# 2.13e-20
C8286 _049_ _279_/a_396_47# 1.43e-19
C8287 net44 _319_/a_761_289# 5.86e-20
C8288 _210_/a_199_47# net14 1.81e-19
C8289 _308_/a_761_289# clknet_2_0__leaf_clk 6.24e-20
C8290 _308_/a_27_47# net45 2.93e-20
C8291 _326_/a_27_47# net43 0.304f
C8292 _330_/a_651_413# _027_ 8.49e-19
C8293 _330_/a_448_47# net46 2.46e-19
C8294 _122_ net40 5.85e-20
C8295 _301_/a_129_47# _135_ 0.00236f
C8296 _341_/a_761_289# _065_ 4.41e-19
C8297 VPWR net23 0.72f
C8298 _244_/a_27_297# rebuffer5/a_161_47# 8.58e-19
C8299 net15 _034_ 1.23e-19
C8300 _341_/a_761_289# _135_ 1.11e-20
C8301 _341_/a_1108_47# net2 2.97e-19
C8302 _103_ _098_ 0.0872f
C8303 _251_/a_27_297# _101_ 0.118f
C8304 _250_/a_109_47# _101_ 0.00328f
C8305 _320_/a_1108_47# net45 1.03e-19
C8306 _107_ _262_/a_205_47# 1.29e-19
C8307 _042_ _041_ 4.99e-19
C8308 _299_/a_27_413# net40 0.00526f
C8309 _061_ _134_ 0.0033f
C8310 trim_mask\[2\] _056_ 6.23e-19
C8311 _047_ net32 0.147f
C8312 _249_/a_27_297# net26 8.35e-19
C8313 _232_/a_32_297# _090_ 0.164f
C8314 mask\[6\] net20 1.84e-19
C8315 _328_/a_543_47# trim_mask\[1\] 0.03f
C8316 _097_ net14 1.49e-20
C8317 trim_mask\[0\] _067_ 0.0937f
C8318 net51 _208_/a_505_21# 0.144f
C8319 net12 _239_/a_474_297# 0.0104f
C8320 _200_/a_209_297# cal_itt\[1\] 0.0437f
C8321 _073_ _003_ 0.00241f
C8322 output23/a_27_47# _308_/a_193_47# 2.18e-19
C8323 _319_/a_193_47# _016_ 0.289f
C8324 net9 _340_/a_562_413# 6.51e-19
C8325 _319_/a_1108_47# _101_ 7.56e-20
C8326 _319_/a_543_47# net52 6.98e-19
C8327 _284_/a_150_297# net18 4.94e-19
C8328 _328_/a_27_47# _336_/a_1108_47# 3.63e-20
C8329 _103_ clknet_0_clk 0.00673f
C8330 trim_mask\[2\] _336_/a_27_47# 2.46e-19
C8331 _110_ net32 4.19e-20
C8332 _327_/a_1108_47# _267_/a_59_75# 3.19e-19
C8333 _007_ _082_ 0.113f
C8334 _140_/a_68_297# clknet_2_0__leaf_clk 5.04e-20
C8335 _307_/a_651_413# _074_ 0.00467f
C8336 _241_/a_297_47# net30 7.26e-20
C8337 net4 _336_/a_651_413# 0.00382f
C8338 _334_/a_27_47# _334_/a_448_47# 0.0856f
C8339 _334_/a_193_47# _334_/a_1108_47# 0.125f
C8340 _314_/a_27_47# _314_/a_651_413# 9.73e-19
C8341 _314_/a_761_289# _314_/a_1108_47# 0.0512f
C8342 _314_/a_193_47# _314_/a_448_47# 0.0642f
C8343 _326_/a_651_413# net28 7.39e-20
C8344 _122_ _299_/a_215_297# 1.87e-19
C8345 _228_/a_79_21# _052_ 0.0101f
C8346 _228_/a_382_297# _088_ 0.0156f
C8347 net44 _202_/a_382_297# 2.86e-19
C8348 _339_/a_1602_47# cal_count\[0\] 0.0475f
C8349 fanout43/a_27_47# _080_ 8.51e-19
C8350 net12 _206_/a_206_47# 1.84e-20
C8351 _320_/a_1108_47# _065_ 6.09e-19
C8352 _327_/a_27_47# _327_/a_761_289# 0.0701f
C8353 VPWR _036_ 0.975f
C8354 mask\[3\] _082_ 0.0846f
C8355 _307_/a_448_47# net45 2.47e-19
C8356 _239_/a_694_21# _089_ 1.88e-19
C8357 net2 _339_/a_476_47# 1.28e-19
C8358 _308_/a_27_47# _319_/a_27_47# 1.75e-19
C8359 trim[3] _334_/a_651_413# 5.61e-20
C8360 _169_/a_109_53# _185_/a_68_297# 0.00167f
C8361 _168_/a_27_413# _331_/a_27_47# 6.84e-19
C8362 _110_ _033_ 0.00853f
C8363 VPWR _164_/a_161_47# 0.613f
C8364 _299_/a_27_413# _299_/a_215_297# 0.141f
C8365 _005_ net30 5.05e-20
C8366 _094_ _092_ 0.105f
C8367 _327_/a_193_47# _058_ 0.042f
C8368 _320_/a_193_47# _319_/a_1283_21# 8.37e-21
C8369 _034_ _049_ 0.0137f
C8370 _237_/a_76_199# clkbuf_2_0__f_clk/a_110_47# 8.03e-19
C8371 _258_/a_109_297# net9 7.53e-20
C8372 clone1/a_27_47# _242_/a_79_21# 7.45e-19
C8373 net44 _206_/a_206_47# 1.57e-19
C8374 _056_ _175_/a_150_297# 4.96e-19
C8375 _218_/a_199_47# net26 1.86e-19
C8376 _333_/a_27_47# net33 2.82e-20
C8377 _325_/a_543_47# net27 1.05e-19
C8378 _115_ _056_ 4.69e-21
C8379 _267_/a_145_75# _108_ 1.73e-19
C8380 trim_val\[1\] _175_/a_68_297# 5.65e-19
C8381 trim_mask\[1\] _333_/a_27_47# 0.0168f
C8382 trim_val\[1\] _333_/a_193_47# 6.71e-19
C8383 net15 _281_/a_253_47# 0.00261f
C8384 _334_/a_1283_21# rebuffer1/a_75_212# 6.81e-19
C8385 _269_/a_81_21# trim_val\[0\] 2.93e-19
C8386 _068_ _062_ 0.0311f
C8387 VPWR _083_ 0.172f
C8388 _192_/a_505_280# _092_ 5.22e-19
C8389 _192_/a_548_47# _095_ 1.35e-20
C8390 _323_/a_448_47# _042_ 0.0161f
C8391 _159_/a_27_47# _313_/a_27_47# 3.54e-20
C8392 _090_ net55 0.339f
C8393 _335_/a_27_47# _335_/a_761_289# 0.0701f
C8394 _308_/a_1217_47# net45 6.07e-20
C8395 net30 trim_val\[4\] 6.05e-20
C8396 _326_/a_1217_47# net43 6.03e-19
C8397 _027_ net46 0.283f
C8398 result[2] net14 6.6e-20
C8399 _007_ _310_/a_448_47# 0.158f
C8400 _097_ net4 0.00243f
C8401 output26/a_27_47# _310_/a_193_47# 2.68e-19
C8402 _284_/a_68_297# cal_count\[3\] 2.16e-19
C8403 _294_/a_68_297# net2 0.177f
C8404 _083_ net53 0.0625f
C8405 _211_/a_109_297# net14 9.08e-19
C8406 _337_/a_193_47# _121_ 7.28e-19
C8407 _230_/a_59_75# clkbuf_2_3__f_clk/a_110_47# 0.0067f
C8408 output28/a_27_47# _011_ 0.00175f
C8409 _309_/a_543_47# net45 1.49e-19
C8410 _255_/a_27_47# _051_ 6.49e-19
C8411 _182_/a_27_47# _332_/a_1283_21# 0.0125f
C8412 _058_ _332_/a_27_47# 0.00986f
C8413 VPWR net50 0.429f
C8414 net43 cal_itt\[3\] 1.33e-20
C8415 output10/a_27_47# _057_ 4.11e-19
C8416 _110_ _103_ 4.07e-20
C8417 _334_/a_1270_413# net46 2.06e-19
C8418 _082_ _310_/a_1283_21# 3.18e-19
C8419 VPWR _208_/a_218_374# 0.00215f
C8420 _195_/a_76_199# _068_ 0.0783f
C8421 VPWR _207_/a_109_297# 0.00439f
C8422 _290_/a_207_413# trimb[1] 7.14e-19
C8423 net55 _242_/a_382_297# 0.00129f
C8424 net9 _338_/a_1602_47# 0.00333f
C8425 _327_/a_448_47# net46 8.97e-19
C8426 input2/a_27_47# net37 4.62e-20
C8427 _336_/a_193_47# trim_mask\[4\] 0.0256f
C8428 trim_mask\[2\] net48 0.139f
C8429 result[1] _308_/a_448_47# 6.45e-20
C8430 _329_/a_543_47# clknet_2_2__leaf_clk 2.28e-19
C8431 _304_/a_1283_21# _304_/a_1108_47# 0.234f
C8432 _304_/a_761_289# _304_/a_651_413# 0.0977f
C8433 _304_/a_543_47# _304_/a_448_47# 0.0498f
C8434 _304_/a_27_47# _304_/a_639_47# 0.00188f
C8435 _304_/a_193_47# _304_/a_1270_413# 1.46e-19
C8436 _023_ _078_ 3.55e-19
C8437 _162_/a_27_47# net34 2.42e-20
C8438 _339_/a_476_47# _123_ 0.0325f
C8439 _048_ _227_/a_209_311# 0.0748f
C8440 net43 _305_/a_27_47# 0.921f
C8441 output32/a_27_47# _047_ 0.0241f
C8442 _334_/a_27_47# _031_ 0.167f
C8443 _076_ rebuffer6/a_27_47# 0.212f
C8444 net37 rebuffer2/a_75_212# 1.32e-20
C8445 _026_ _258_/a_27_297# 0.11f
C8446 _132_ _131_ 0.119f
C8447 output20/a_27_47# _156_/a_27_47# 5.42e-20
C8448 _327_/a_543_47# _327_/a_805_47# 0.00171f
C8449 _327_/a_761_289# _327_/a_1217_47# 4.2e-19
C8450 _327_/a_1108_47# _327_/a_1270_413# 0.00645f
C8451 mask\[1\] net51 5.71e-20
C8452 clknet_0_clk clkbuf_2_3__f_clk/a_110_47# 0.327f
C8453 _335_/a_448_47# net46 0.0054f
C8454 _281_/a_253_47# _049_ 8.9e-20
C8455 _093_ _095_ 1.33e-19
C8456 calibrate _099_ 4.75e-19
C8457 VPWR _226_/a_27_47# 0.422f
C8458 _188_/a_27_47# _136_ 3.66e-21
C8459 _308_/a_1108_47# _319_/a_448_47# 4.21e-21
C8460 _235_/a_382_297# net3 2.21e-19
C8461 _293_/a_384_47# cal_count\[0\] 0.00958f
C8462 net3 _317_/a_27_47# 1.33e-19
C8463 _306_/a_761_289# _076_ 3.26e-20
C8464 _038_ _284_/a_68_297# 0.00282f
C8465 _304_/a_193_47# clknet_2_3__leaf_clk 0.161f
C8466 _128_ cal_count\[0\] 0.0184f
C8467 mask\[3\] _247_/a_27_297# 0.197f
C8468 _327_/a_1462_47# _058_ 2.66e-19
C8469 _309_/a_193_47# clknet_2_1__leaf_clk 0.00269f
C8470 _078_ _046_ 0.357f
C8471 net45 _099_ 0.0026f
C8472 _014_ _092_ 0.00462f
C8473 net24 _081_ 0.277f
C8474 _104_ trim_mask\[4\] 0.297f
C8475 VPWR _330_/a_1108_47# 0.318f
C8476 _332_/a_1108_47# net46 0.286f
C8477 _328_/a_1270_413# net9 1.5e-19
C8478 net43 _011_ 6.44e-19
C8479 net12 _103_ 8.81e-21
C8480 VPWR _217_/a_109_297# 0.00478f
C8481 _137_/a_150_297# _039_ 4.96e-19
C8482 net13 _319_/a_1283_21# 5.1e-19
C8483 _112_ _333_/a_639_47# 6.26e-19
C8484 net49 _333_/a_805_47# 6.71e-19
C8485 _021_ _312_/a_651_413# 6.03e-21
C8486 _340_/a_562_413# _122_ 7.19e-20
C8487 _337_/a_761_289# clknet_0_clk 2.53e-20
C8488 net48 _333_/a_761_289# 6.02e-21
C8489 trim_val\[2\] _333_/a_1283_21# 1.8e-20
C8490 _115_ net48 0.0183f
C8491 trim_mask\[4\] net55 6.4e-20
C8492 net31 cal_count\[0\] 6.25e-20
C8493 _134_ net16 0.335f
C8494 cal_count\[1\] _132_ 1.61e-19
C8495 _310_/a_193_47# _310_/a_639_47# 2.28e-19
C8496 _310_/a_761_289# _310_/a_1270_413# 2.6e-19
C8497 _310_/a_543_47# _310_/a_651_413# 0.0572f
C8498 _324_/a_27_47# _042_ 7.87e-20
C8499 _008_ _074_ 0.0504f
C8500 cal_itt\[1\] _053_ 0.00161f
C8501 _306_/a_27_47# fanout44/a_27_47# 3.47e-21
C8502 _307_/a_1283_21# _210_/a_113_297# 3.48e-20
C8503 _059_ _228_/a_79_21# 2.24e-19
C8504 _327_/a_639_47# _108_ 3.69e-19
C8505 VPWR _216_/a_113_297# 0.264f
C8506 VPWR _325_/a_448_47# 0.0857f
C8507 _065_ _099_ 3.14e-19
C8508 _322_/a_1108_47# _065_ 3.11e-20
C8509 _050_ _170_/a_81_21# 0.0186f
C8510 _053_ _052_ 0.0087f
C8511 _046_ _313_/a_651_413# 4.33e-19
C8512 net21 _313_/a_1108_47# 0.00661f
C8513 _335_/a_1108_47# _335_/a_1270_413# 0.00645f
C8514 _335_/a_761_289# _335_/a_1217_47# 4.2e-19
C8515 _335_/a_543_47# _335_/a_805_47# 0.00171f
C8516 output22/a_27_47# net22 0.171f
C8517 _324_/a_1283_21# clknet_2_1__leaf_clk 9.42e-19
C8518 _340_/a_27_47# _129_ 1.16e-20
C8519 result[4] _310_/a_448_47# 6.75e-19
C8520 _000_ _072_ 6.77e-22
C8521 _305_/a_448_47# _092_ 4.12e-20
C8522 _311_/a_193_47# _311_/a_761_289# 0.181f
C8523 _311_/a_27_47# _311_/a_543_47# 0.111f
C8524 _024_ net40 5.23e-20
C8525 clkbuf_0_clk/a_110_47# _230_/a_59_75# 8.11e-20
C8526 _230_/a_59_75# cal_count\[3\] 3.92e-20
C8527 net31 _061_ 1.31e-19
C8528 VPWR _181_/a_150_297# 0.00144f
C8529 _074_ mask\[5\] 5.12e-19
C8530 clknet_2_3__leaf_clk net18 0.0822f
C8531 _058_ _332_/a_1217_47# 9.77e-20
C8532 _304_/a_27_47# _136_ 0.00313f
C8533 trim_mask\[2\] _172_/a_68_297# 1.33e-19
C8534 _067_ trim_mask\[4\] 6.2e-21
C8535 _144_/a_27_47# _129_ 0.00317f
C8536 trim[1] trim_mask\[0\] 6.55e-19
C8537 _336_/a_1462_47# trim_mask\[4\] 0.00226f
C8538 _033_ clknet_2_2__leaf_clk 0.759f
C8539 clknet_2_3__leaf_clk _129_ 3e-21
C8540 net15 _314_/a_27_47# 1.97e-21
C8541 cal_count\[3\] _098_ 1.22e-20
C8542 result[1] _005_ 0.077f
C8543 _304_/a_761_289# net47 0.166f
C8544 _096_ _241_/a_105_352# 1.46e-19
C8545 _164_/a_161_47# _093_ 0.0694f
C8546 net43 _305_/a_1217_47# 6.59e-20
C8547 _256_/a_27_297# _256_/a_373_47# 0.0134f
C8548 _110_ clkbuf_2_3__f_clk/a_110_47# 1.11e-20
C8549 net16 _339_/a_1602_47# 0.00389f
C8550 _336_/a_651_413# _279_/a_396_47# 6.53e-20
C8551 _187_/a_27_413# en_co_clk 0.0927f
C8552 VPWR _314_/a_761_289# 0.212f
C8553 _308_/a_761_289# _078_ 3.77e-19
C8554 _308_/a_1283_21# net22 8.92e-21
C8555 _321_/a_1283_21# _321_/a_1108_47# 0.234f
C8556 _321_/a_761_289# _321_/a_651_413# 0.0977f
C8557 _321_/a_543_47# _321_/a_448_47# 0.0498f
C8558 _321_/a_27_47# _321_/a_639_47# 3.82e-19
C8559 _321_/a_193_47# _321_/a_1270_413# 1.46e-19
C8560 _332_/a_761_289# _332_/a_639_47# 3.16e-19
C8561 _332_/a_27_47# _332_/a_1217_47# 2.56e-19
C8562 _340_/a_27_47# _340_/a_1182_261# 0.0608f
C8563 _340_/a_193_47# _340_/a_476_47# 0.215f
C8564 _228_/a_382_297# _170_/a_299_297# 3.58e-19
C8565 _136_ _298_/a_292_297# 6.7e-20
C8566 clk clkbuf_2_2__f_clk/a_110_47# 0.00318f
C8567 clkbuf_0_clk/a_110_47# clknet_0_clk 1.74f
C8568 clknet_0_clk cal_count\[3\] 1.76e-20
C8569 VPWR _185_/a_150_297# 0.00214f
C8570 _302_/a_27_297# clknet_2_3__leaf_clk 0.0472f
C8571 ctlp[0] _314_/a_27_47# 0.00196f
C8572 _032_ net46 0.0299f
C8573 clkbuf_2_0__f_clk/a_110_47# _281_/a_103_199# 0.0142f
C8574 _019_ _074_ 7.53e-20
C8575 trim[4] net46 5.7e-19
C8576 net43 _319_/a_1283_21# 0.313f
C8577 _244_/a_27_297# net51 0.049f
C8578 net23 _319_/a_193_47# 8.7e-20
C8579 _168_/a_207_413# trim_mask\[4\] 0.0619f
C8580 input3/a_75_212# clknet_2_0__leaf_clk 1.56e-19
C8581 output31/a_27_47# net33 0.0052f
C8582 _116_ net18 0.0016f
C8583 _337_/a_1283_21# _337_/a_1108_47# 0.234f
C8584 _337_/a_761_289# _337_/a_651_413# 0.0977f
C8585 _337_/a_543_47# _337_/a_448_47# 0.0498f
C8586 _337_/a_27_47# _337_/a_639_47# 3.82e-19
C8587 _337_/a_193_47# _337_/a_1270_413# 1.46e-19
C8588 clknet_0_clk _331_/a_27_47# 0.0133f
C8589 output31/a_27_47# trim_mask\[1\] 0.00105f
C8590 trim[0] _269_/a_299_297# 1.79e-19
C8591 net25 _018_ 0.00104f
C8592 result[4] result[5] 0.049f
C8593 _340_/a_1602_47# _133_ 0.00808f
C8594 _297_/a_285_47# net40 0.00447f
C8595 net9 _339_/a_381_47# 0.00292f
C8596 trim_val\[0\] net32 1.68e-19
C8597 net4 clkbuf_2_2__f_clk/a_110_47# 0.214f
C8598 _270_/a_59_75# _333_/a_27_47# 0.00308f
C8599 _308_/a_193_47# output30/a_27_47# 1.86e-20
C8600 _287_/a_75_212# _338_/a_193_47# 0.00801f
C8601 _078_ _140_/a_68_297# 0.00199f
C8602 _101_ _003_ 5.74e-19
C8603 _276_/a_145_75# _110_ 0.00165f
C8604 VPWR output26/a_27_47# 0.322f
C8605 _276_/a_59_75# _116_ 0.185f
C8606 VPWR _195_/a_535_374# 8.98e-19
C8607 _301_/a_47_47# clkc 7.43e-20
C8608 _097_ _237_/a_535_374# 1.33e-19
C8609 VPWR cal_itt\[1\] 0.95f
C8610 net47 _043_ 0.0686f
C8611 _324_/a_761_289# _021_ 1.27e-19
C8612 _239_/a_694_21# _092_ 0.0334f
C8613 VPWR _334_/a_651_413# 0.155f
C8614 net37 trimb[4] 0.00207f
C8615 VPWR _052_ 0.357f
C8616 VPWR input1/a_75_212# 0.259f
C8617 _314_/a_1270_413# net29 1.14e-19
C8618 _307_/a_805_47# net22 7.15e-19
C8619 VPWR _327_/a_1108_47# 0.309f
C8620 _307_/a_1270_413# _078_ 1.06e-19
C8621 output37/a_27_47# net40 2.1e-20
C8622 output16/a_27_47# net39 0.01f
C8623 input1/a_75_212# valid 1.27e-19
C8624 _075_ _049_ 0.178f
C8625 net16 cal_count\[2\] 0.0127f
C8626 net27 result[5] 0.00579f
C8627 clkbuf_2_0__f_clk/a_110_47# _048_ 0.012f
C8628 trim_mask\[0\] clknet_2_3__leaf_clk 0.324f
C8629 ctln[4] _335_/a_27_47# 3.44e-19
C8630 _304_/a_651_413# _038_ 2.17e-20
C8631 _304_/a_1217_47# _136_ 1.02e-19
C8632 VPWR _141_/a_27_47# 0.258f
C8633 _310_/a_1283_21# net29 1.08e-21
C8634 VPWR _335_/a_1108_47# 0.305f
C8635 net2 rebuffer5/a_161_47# 5.89e-19
C8636 _319_/a_805_47# _092_ 2.63e-21
C8637 trimb[0] output37/a_27_47# 0.00178f
C8638 output36/a_27_47# trimb[1] 6.66e-20
C8639 VPWR input2/a_27_47# 0.407f
C8640 VPWR _311_/a_27_47# 0.423f
C8641 _305_/a_543_47# en_co_clk 4.11e-21
C8642 net4 _035_ 3.57e-20
C8643 _341_/a_193_47# _304_/a_193_47# 1.89e-21
C8644 _341_/a_27_47# _304_/a_761_289# 9.3e-20
C8645 _328_/a_27_47# net18 2.45e-21
C8646 _110_ cal_count\[3\] 4.11e-20
C8647 _060_ _235_/a_297_47# 1.12e-19
C8648 _340_/a_1032_413# net47 0.217f
C8649 VPWR rebuffer2/a_75_212# 0.28f
C8650 _037_ _304_/a_543_47# 2.7e-19
C8651 _189_/a_27_47# en_co_clk 4.84e-21
C8652 _311_/a_27_47# net53 0.0225f
C8653 _065_ _208_/a_535_374# 0.00104f
C8654 output31/a_27_47# output33/a_27_47# 0.0523f
C8655 VPWR _332_/a_1283_21# 0.37f
C8656 _340_/a_652_21# _340_/a_1056_47# 3.94e-19
C8657 _340_/a_476_47# _340_/a_796_47# 0.00184f
C8658 _340_/a_1032_413# _340_/a_1140_413# 0.00523f
C8659 _340_/a_381_47# _340_/a_562_413# 8.75e-19
C8660 _043_ net44 1.13e-20
C8661 _293_/a_384_47# net16 2.61e-19
C8662 _059_ _053_ 4.32e-20
C8663 _134_ net40 1.8e-19
C8664 clkbuf_2_0__f_clk/a_110_47# _120_ 0.0439f
C8665 _291_/a_117_297# net33 0.00159f
C8666 mask\[0\] _283_/a_75_212# 4.16e-20
C8667 _309_/a_1108_47# _078_ 0.0499f
C8668 _128_ net16 0.0758f
C8669 clk fanout45/a_27_47# 0.00263f
C8670 state\[0\] net41 0.272f
C8671 _323_/a_27_47# net18 6.31e-21
C8672 _326_/a_193_47# _310_/a_1108_47# 4.77e-21
C8673 _326_/a_761_289# _310_/a_1283_21# 1.09e-20
C8674 _326_/a_543_47# _310_/a_543_47# 1.3e-20
C8675 clkbuf_0_clk/a_110_47# net47 3.95e-19
C8676 _337_/a_761_289# net44 0.167f
C8677 _309_/a_761_289# net24 0.0191f
C8678 net47 cal_count\[3\] 9.79e-21
C8679 _338_/a_652_21# clknet_2_3__leaf_clk 0.0268f
C8680 _062_ cal_itt\[3\] 2.91e-19
C8681 _291_/a_35_297# _290_/a_207_413# 0.0019f
C8682 net13 clone7/a_27_47# 0.00466f
C8683 VPWR _310_/a_639_47# 7.41e-19
C8684 clknet_2_1__leaf_clk _208_/a_505_21# 0.00601f
C8685 net43 _313_/a_761_289# 0.162f
C8686 _058_ net30 0.00133f
C8687 _333_/a_1108_47# _055_ 0.00518f
C8688 _106_ _092_ 2.91e-20
C8689 _035_ _063_ 8.42e-20
C8690 clknet_2_1__leaf_clk mask\[2\] 0.387f
C8691 _304_/a_27_47# _339_/a_27_47# 2.67e-20
C8692 _035_ _338_/a_381_47# 0.144f
C8693 _293_/a_81_21# _126_ 8.39e-19
C8694 net27 net29 0.284f
C8695 net31 net16 4.4e-20
C8696 net24 _040_ 1.22e-19
C8697 _242_/a_297_47# _098_ 0.0523f
C8698 _161_/a_68_297# _332_/a_1283_21# 0.00113f
C8699 _189_/a_27_47# _050_ 0.216f
C8700 _321_/a_1108_47# _101_ 0.0581f
C8701 trim[1] _265_/a_81_21# 4.51e-20
C8702 output32/a_27_47# trim_val\[0\] 0.00905f
C8703 _338_/a_956_413# net18 7.18e-19
C8704 fanout45/a_27_47# net4 0.213f
C8705 _341_/a_193_47# net18 0.00307f
C8706 _134_ _299_/a_215_297# 0.082f
C8707 _306_/a_27_47# rebuffer6/a_27_47# 2.16e-21
C8708 _195_/a_76_199# cal_itt\[3\] 4.72e-20
C8709 _337_/a_1108_47# _101_ 1.38e-19
C8710 _337_/a_543_47# net52 3.49e-21
C8711 _337_/a_27_47# _263_/a_297_47# 1.6e-20
C8712 _064_ _048_ 7.4e-21
C8713 net15 _247_/a_109_297# 0.00362f
C8714 _313_/a_1108_47# _045_ 7.2e-20
C8715 _053_ _170_/a_384_47# 1.26e-19
C8716 _291_/a_35_297# _289_/a_68_297# 3.32e-19
C8717 _339_/a_1602_47# net40 1.88e-20
C8718 clk _331_/a_193_47# 0.0195f
C8719 _199_/a_193_297# _069_ 0.0012f
C8720 _258_/a_27_297# _280_/a_75_212# 0.02f
C8721 _314_/a_193_47# _086_ 8.56e-20
C8722 net12 _331_/a_27_47# 1.36e-19
C8723 _311_/a_1283_21# net26 0.11f
C8724 net28 _313_/a_639_47# 0.00432f
C8725 _339_/a_1032_413# net34 4.15e-21
C8726 _064_ _330_/a_27_47# 5.22e-21
C8727 net50 _336_/a_1108_47# 1.67e-20
C8728 _306_/a_27_47# _306_/a_761_289# 0.0701f
C8729 net9 _025_ 9.33e-19
C8730 _048_ _100_ 0.21f
C8731 ctln[4] _335_/a_1217_47# 6.4e-20
C8732 _329_/a_543_47# trim_mask\[3\] 0.00103f
C8733 net47 _038_ 4.05e-20
C8734 _341_/a_193_47# _302_/a_27_297# 4.26e-20
C8735 _341_/a_27_47# _302_/a_109_297# 5.29e-20
C8736 cal_itt\[2\] _262_/a_193_297# 2.71e-19
C8737 _326_/a_761_289# net27 4.37e-19
C8738 _326_/a_27_47# result[5] 0.00691f
C8739 _329_/a_193_47# _057_ 3.06e-19
C8740 _331_/a_27_47# _331_/a_1108_47# 0.102f
C8741 _331_/a_193_47# _331_/a_1283_21# 0.0424f
C8742 _331_/a_761_289# _331_/a_543_47# 0.21f
C8743 VPWR _311_/a_1217_47# 4.26e-20
C8744 _083_ mask\[6\] 6.36e-20
C8745 net4 _198_/a_27_47# 0.0121f
C8746 clkbuf_0_clk/a_110_47# net44 0.00349f
C8747 _051_ _119_ 4.4e-20
C8748 _218_/a_113_297# _078_ 0.0791f
C8749 _321_/a_1283_21# _320_/a_193_47# 1.97e-19
C8750 _321_/a_1108_47# _320_/a_27_47# 3.64e-21
C8751 _143_/a_68_297# _041_ 0.109f
C8752 _325_/a_193_47# _042_ 2.83e-19
C8753 _001_ _202_/a_382_297# 1.78e-20
C8754 net4 _331_/a_193_47# 1.66e-19
C8755 net47 _338_/a_476_47# 0.254f
C8756 _258_/a_27_297# _258_/a_109_297# 0.171f
C8757 _328_/a_27_47# trim_mask\[0\] 1.21e-20
C8758 _258_/a_109_297# _024_ 6.81e-20
C8759 _050_ _336_/a_27_47# 2.14e-19
C8760 _323_/a_1283_21# clknet_2_3__leaf_clk 7.04e-22
C8761 input1/a_75_212# _315_/a_543_47# 2.16e-20
C8762 _311_/a_1217_47# net53 5.17e-20
C8763 _325_/a_1108_47# clknet_2_1__leaf_clk 5.88e-20
C8764 _074_ _310_/a_27_47# 0.0175f
C8765 VPWR _059_ 0.816f
C8766 _340_/a_1602_47# _037_ 5.93e-20
C8767 net23 net24 3.22e-19
C8768 _051_ _331_/a_651_413# 2.87e-19
C8769 _327_/a_448_47# _111_ 9.03e-20
C8770 _257_/a_27_297# net40 5.9e-22
C8771 mask\[7\] _023_ 4.85e-19
C8772 en_co_clk _096_ 0.0308f
C8773 _301_/a_47_47# cal_count\[3\] 3.02e-19
C8774 _048_ _264_/a_27_297# 0.00146f
C8775 _110_ _328_/a_1108_47# 3.3e-20
C8776 _110_ trim_mask\[2\] 0.515f
C8777 output9/a_27_47# _057_ 0.0557f
C8778 _051_ _087_ 0.316f
C8779 _097_ _281_/a_253_47# 2.12e-19
C8780 net42 en_co_clk 2.04e-20
C8781 _302_/a_109_297# clknet_2_2__leaf_clk 5.41e-20
C8782 trim_mask\[0\] _266_/a_68_297# 9.75e-19
C8783 _341_/a_27_47# cal_count\[3\] 0.0348f
C8784 _338_/a_1056_47# clknet_2_3__leaf_clk 2.82e-19
C8785 _291_/a_285_47# _127_ 3.98e-19
C8786 _341_/a_1108_47# clknet_2_3__leaf_clk 0.0465f
C8787 _336_/a_1108_47# _330_/a_1108_47# 6.38e-21
C8788 state\[0\] _192_/a_505_280# 3.6e-21
C8789 _198_/a_27_47# _063_ 0.0778f
C8790 trim_mask\[1\] _267_/a_59_75# 2.13e-21
C8791 _065_ rebuffer4/a_27_47# 0.0332f
C8792 cal_count\[2\] net40 0.00976f
C8793 state\[2\] _167_/a_161_47# 7.2e-19
C8794 fanout46/a_27_47# _335_/a_543_47# 1.78e-19
C8795 clkbuf_2_2__f_clk/a_110_47# _279_/a_396_47# 0.00226f
C8796 VPWR _306_/a_1108_47# 0.306f
C8797 _265_/a_81_21# clknet_2_3__leaf_clk 3.16e-21
C8798 _226_/a_27_47# _206_/a_27_93# 6.99e-19
C8799 _283_/a_75_212# _121_ 0.188f
C8800 _340_/a_27_47# _339_/a_476_47# 1.06e-20
C8801 _340_/a_476_47# _339_/a_27_47# 8.3e-21
C8802 _091_ _107_ 0.00135f
C8803 clknet_2_1__leaf_clk _314_/a_193_47# 0.0242f
C8804 _307_/a_27_47# net14 0.0096f
C8805 mask\[1\] clknet_2_1__leaf_clk 0.00928f
C8806 _041_ net4 0.0577f
C8807 _326_/a_27_47# net29 1.88e-19
C8808 VPWR trimb[4] 0.577f
C8809 mask\[7\] _046_ 0.0168f
C8810 trim[3] net33 0.00119f
C8811 VPWR _170_/a_384_47# 5.39e-20
C8812 _337_/a_1283_21# _107_ 2.03e-19
C8813 _029_ _332_/a_1283_21# 1.04e-20
C8814 _050_ _096_ 0.0653f
C8815 net15 _018_ 0.00157f
C8816 _182_/a_27_47# net33 0.00559f
C8817 output27/a_27_47# _074_ 2.17e-20
C8818 _146_/a_68_297# _310_/a_193_47# 2.8e-20
C8819 net43 _073_ 1.23e-19
C8820 _339_/a_1032_413# _133_ 7.58e-21
C8821 clk _260_/a_93_21# 2.46e-19
C8822 _323_/a_1108_47# net47 0.24f
C8823 net42 _050_ 0.00488f
C8824 trim_mask\[4\] clknet_2_3__leaf_clk 1.03e-21
C8825 _312_/a_543_47# net20 0.00959f
C8826 _299_/a_215_297# cal_count\[2\] 0.0799f
C8827 _259_/a_109_297# net46 0.00236f
C8828 trim_mask\[3\] _033_ 4.38e-20
C8829 _306_/a_543_47# _306_/a_805_47# 0.00171f
C8830 _306_/a_761_289# _306_/a_1217_47# 4.2e-19
C8831 _306_/a_1108_47# _306_/a_1270_413# 0.00645f
C8832 net12 net21 2.37e-20
C8833 _007_ _042_ 0.00131f
C8834 trim_val\[4\] net40 1.61e-20
C8835 _110_ _115_ 0.00253f
C8836 _341_/a_27_47# _038_ 0.218f
C8837 _341_/a_1283_21# _136_ 0.00872f
C8838 clkbuf_2_3__f_clk/a_110_47# _279_/a_204_297# 2.91e-21
C8839 _128_ net40 2.4e-21
C8840 _110_ _265_/a_299_297# 0.00182f
C8841 _331_/a_1108_47# _331_/a_1217_47# 0.00742f
C8842 _331_/a_1283_21# _331_/a_1462_47# 0.0074f
C8843 _331_/a_27_47# clknet_2_2__leaf_clk 0.274f
C8844 net7 _317_/a_193_47# 1.8e-20
C8845 net15 _317_/a_543_47# 0.00815f
C8846 _325_/a_193_47# _022_ 0.329f
C8847 _317_/a_27_47# _317_/a_761_289# 0.0701f
C8848 _325_/a_448_47# mask\[6\] 0.0248f
C8849 net33 net37 0.841f
C8850 _041_ net52 0.00218f
C8851 _326_/a_27_47# _326_/a_761_289# 0.0701f
C8852 _041_ _063_ 1.61e-20
C8853 _159_/a_27_47# net21 0.111f
C8854 _306_/a_543_47# _049_ 3.01e-20
C8855 _169_/a_109_53# _232_/a_32_297# 1.51e-20
C8856 mask\[3\] _042_ 0.768f
C8857 _308_/a_1108_47# net14 4.01e-19
C8858 _338_/a_652_21# _338_/a_956_413# 3.11e-19
C8859 _338_/a_1032_413# _338_/a_1602_47# 0.111f
C8860 _338_/a_476_47# _338_/a_562_413# 0.00972f
C8861 net47 _338_/a_1224_47# 0.00173f
C8862 VPWR _317_/a_1108_47# 0.277f
C8863 net4 _260_/a_93_21# 7.28e-20
C8864 _328_/a_27_47# _328_/a_1283_21# 0.0435f
C8865 _328_/a_193_47# _328_/a_543_47# 0.207f
C8866 _064_ _327_/a_27_47# 4.55e-19
C8867 VPWR _326_/a_1108_47# 0.328f
C8868 _258_/a_373_47# trim_mask\[2\] 0.00175f
C8869 net10 ctln[4] 0.0067f
C8870 _306_/a_193_47# net30 2.7e-20
C8871 net13 _321_/a_1283_21# 0.0043f
C8872 _037_ _041_ 1.72e-20
C8873 cal _315_/a_805_47# 4.66e-20
C8874 _290_/a_27_413# net37 3.35e-19
C8875 state\[0\] _014_ 1.06e-20
C8876 net31 net40 2.27e-19
C8877 net13 _337_/a_1283_21# 2.47e-19
C8878 net12 _242_/a_297_47# 4.52e-19
C8879 _214_/a_113_297# _101_ 0.00483f
C8880 net2 comp 0.0198f
C8881 _170_/a_81_21# _049_ 0.105f
C8882 cal_itt\[1\] _197_/a_113_297# 0.00924f
C8883 cal_itt\[0\] _197_/a_199_47# 0.0109f
C8884 VPWR _203_/a_59_75# 0.222f
C8885 _040_ _337_/a_193_47# 4.4e-20
C8886 VPWR _286_/a_218_47# 9.7e-20
C8887 clknet_0_clk _190_/a_215_47# 2.56e-19
C8888 _325_/a_761_289# _313_/a_543_47# 4.07e-20
C8889 _325_/a_543_47# _313_/a_761_289# 3.29e-20
C8890 VPWR _192_/a_27_47# 0.329f
C8891 _064_ _335_/a_27_47# 4.61e-20
C8892 _038_ clknet_2_2__leaf_clk 1.8e-20
C8893 net49 net46 0.0204f
C8894 _272_/a_81_21# net46 0.00853f
C8895 net44 _312_/a_1283_21# 0.287f
C8896 _312_/a_27_47# _312_/a_761_289# 0.0701f
C8897 _033_ _330_/a_1283_21# 1.15e-20
C8898 _336_/a_543_47# net46 0.152f
C8899 _168_/a_27_413# _050_ 0.236f
C8900 _227_/a_109_93# _054_ 7.34e-20
C8901 _227_/a_296_53# _049_ 1.28e-19
C8902 _320_/a_193_47# _101_ 3.1e-20
C8903 _087_ _242_/a_79_21# 5.14e-20
C8904 _323_/a_1108_47# net44 5.49e-20
C8905 _329_/a_193_47# _027_ 0.00194f
C8906 _329_/a_27_47# net46 0.308f
C8907 _303_/a_543_47# clknet_2_3__leaf_clk 0.0335f
C8908 net2 net51 0.0602f
C8909 net31 trimb[0] 0.00722f
C8910 _227_/a_109_93# net30 0.00138f
C8911 _298_/a_215_47# _131_ 0.00144f
C8912 output33/a_27_47# trim[3] 6.66e-20
C8913 trim[2] output34/a_27_47# 0.00212f
C8914 net47 _339_/a_1182_261# 0.116f
C8915 cal_itt\[2\] _202_/a_297_47# 0.0563f
C8916 _321_/a_1108_47# _248_/a_27_297# 7.15e-19
C8917 _114_ _334_/a_27_47# 8.99e-20
C8918 net48 _334_/a_193_47# 6.36e-19
C8919 trim_val\[2\] _334_/a_543_47# 0.00627f
C8920 _323_/a_27_47# _323_/a_1283_21# 0.0436f
C8921 _323_/a_193_47# _323_/a_543_47# 0.217f
C8922 _200_/a_80_21# _106_ 1.09e-20
C8923 _024_ _107_ 6.14e-21
C8924 _305_/a_27_47# rebuffer6/a_27_47# 6.02e-20
C8925 _307_/a_1217_47# net14 2.97e-20
C8926 VPWR _315_/a_27_47# 0.537f
C8927 _263_/a_382_297# _090_ 0.00164f
C8928 _306_/a_193_47# _072_ 3.02e-19
C8929 _306_/a_761_289# cal_itt\[3\] 3.97e-19
C8930 _337_/a_27_47# _099_ 8.76e-22
C8931 _337_/a_193_47# _095_ 0.00207f
C8932 _284_/a_68_297# en_co_clk 0.0135f
C8933 _189_/a_408_47# _053_ 1.94e-19
C8934 net14 output6/a_27_47# 0.0251f
C8935 _328_/a_27_47# _333_/a_193_47# 2.74e-21
C8936 trim_mask\[2\] _274_/a_75_212# 0.036f
C8937 result[5] _011_ 5.91e-19
C8938 net3 clone7/a_27_47# 1.92e-20
C8939 VPWR _318_/a_1270_413# 6.47e-19
C8940 _315_/a_27_47# valid 0.0101f
C8941 _308_/a_193_47# _006_ 4.59e-21
C8942 _308_/a_543_47# _081_ 7.83e-20
C8943 _042_ _310_/a_1283_21# 2.13e-19
C8944 en_co_clk output5/a_27_47# 2.25e-19
C8945 _239_/a_277_297# _052_ 2.72e-19
C8946 _292_/a_78_199# _340_/a_1182_261# 0.00813f
C8947 _190_/a_27_47# clknet_2_3__leaf_clk 3.8e-20
C8948 _179_/a_27_47# _057_ 0.206f
C8949 _169_/a_109_53# net55 1.7e-20
C8950 state\[0\] _243_/a_27_297# 0.0209f
C8951 net54 _100_ 0.0442f
C8952 _058_ _066_ 0.00225f
C8953 _306_/a_193_47# _305_/a_193_47# 3.79e-20
C8954 _306_/a_761_289# _305_/a_27_47# 1.38e-19
C8955 net43 _321_/a_1283_21# 0.291f
C8956 VPWR _225_/a_109_297# 0.00508f
C8957 output33/a_27_47# net37 6.98e-21
C8958 _130_ _131_ 0.203f
C8959 _181_/a_68_297# _033_ 3.76e-22
C8960 clknet_2_1__leaf_clk _310_/a_1270_413# 6.5e-19
C8961 _320_/a_27_47# _320_/a_193_47# 0.85f
C8962 _071_ _002_ 3.17e-21
C8963 _059_ _093_ 9.99e-21
C8964 _341_/a_1217_47# _038_ 1.94e-20
C8965 output14/a_27_47# _086_ 0.00109f
C8966 _331_/a_448_47# trim_mask\[4\] 1.05e-19
C8967 _331_/a_805_47# _028_ 6.71e-19
C8968 _331_/a_1217_47# clknet_2_2__leaf_clk 2.72e-20
C8969 _237_/a_76_199# net4 5.62e-20
C8970 _058_ net16 0.0446f
C8971 _260_/a_93_21# _260_/a_346_47# 0.0119f
C8972 _317_/a_1108_47# _317_/a_1270_413# 0.00645f
C8973 _317_/a_761_289# _317_/a_1217_47# 4.2e-19
C8974 _317_/a_543_47# _317_/a_805_47# 0.00171f
C8975 _328_/a_27_47# trim_mask\[4\] 9.71e-19
C8976 trim_mask\[2\] clknet_2_2__leaf_clk 0.59f
C8977 _328_/a_1108_47# clknet_2_2__leaf_clk 0.0568f
C8978 calibrate net41 0.0278f
C8979 _326_/a_543_47# _326_/a_805_47# 0.00171f
C8980 _326_/a_761_289# _326_/a_1217_47# 4.2e-19
C8981 _326_/a_1108_47# _326_/a_1270_413# 0.00645f
C8982 _325_/a_639_47# _078_ 1.55e-19
C8983 net17 _339_/a_193_47# 1.07e-20
C8984 _337_/a_543_47# _034_ 0.00142f
C8985 VPWR clknet_2_0__leaf_clk 7.25f
C8986 net43 _138_/a_27_47# 0.0341f
C8987 _328_/a_448_47# _328_/a_639_47# 4.61e-19
C8988 _341_/a_193_47# _341_/a_1108_47# 0.119f
C8989 _341_/a_27_47# _341_/a_448_47# 0.0866f
C8990 _081_ _140_/a_150_297# 0.00117f
C8991 VPWR _030_ 0.405f
C8992 clk output6/a_27_47# 0.00421f
C8993 _320_/a_639_47# net44 1.79e-19
C8994 net47 _303_/a_1283_21# 0.344f
C8995 _303_/a_193_47# _338_/a_27_47# 0.00228f
C8996 _303_/a_27_47# _338_/a_193_47# 7.98e-21
C8997 _091_ _118_ 1.49e-21
C8998 _256_/a_109_297# _118_ 5.6e-20
C8999 trim_mask\[0\] _279_/a_314_297# 0.0472f
C9000 _024_ _279_/a_27_47# 1.08e-20
C9001 net45 net41 0.413f
C9002 clknet_2_0__leaf_clk valid 0.00553f
C9003 _010_ _222_/a_113_297# 0.00151f
C9004 _257_/a_27_297# _280_/a_75_212# 1.85e-19
C9005 _274_/a_75_212# _115_ 0.187f
C9006 net16 _332_/a_27_47# 0.0122f
C9007 _318_/a_193_47# _318_/a_651_413# 0.0276f
C9008 _318_/a_543_47# _318_/a_1108_47# 7.99e-20
C9009 net30 _054_ 0.0194f
C9010 _340_/a_562_413# cal_count\[2\] 6.34e-21
C9011 _053_ clone1/a_27_47# 0.0101f
C9012 _266_/a_68_297# trim_mask\[4\] 1.75e-20
C9013 clknet_2_1__leaf_clk _247_/a_109_47# 3.7e-19
C9014 cal_count\[1\] _130_ 0.00126f
C9015 _064_ _335_/a_1217_47# 3.56e-20
C9016 _104_ _335_/a_639_47# 7.42e-20
C9017 net27 _042_ 9.12e-20
C9018 _011_ net29 0.00552f
C9019 _312_/a_1108_47# _312_/a_1270_413# 0.00645f
C9020 _312_/a_761_289# _312_/a_1217_47# 4.2e-19
C9021 _312_/a_543_47# _312_/a_805_47# 0.00171f
C9022 input4/a_27_47# ctln[0] 3.49e-19
C9023 net4 output6/a_27_47# 0.0302f
C9024 _106_ net46 9.94e-21
C9025 _286_/a_76_199# cal_count\[0\] 0.319f
C9026 _286_/a_218_374# _124_ 2.88e-19
C9027 VPWR _305_/a_1108_47# 0.28f
C9028 _306_/a_448_47# net45 4.42e-22
C9029 _329_/a_1217_47# net46 6.97e-19
C9030 calibrate _171_/a_27_47# 1.26e-19
C9031 _078_ _314_/a_1108_47# 7.59e-21
C9032 _308_/a_27_47# _308_/a_761_289# 0.0701f
C9033 _323_/a_651_413# net19 0.00193f
C9034 _258_/a_109_297# _257_/a_27_297# 1.18e-19
C9035 net47 _339_/a_1296_47# 8.83e-19
C9036 VPWR _146_/a_68_297# 0.159f
C9037 clkbuf_2_1__f_clk/a_110_47# net15 0.11f
C9038 _107_ _260_/a_250_297# 0.0013f
C9039 net13 _101_ 0.0171f
C9040 _307_/a_27_47# _307_/a_543_47# 0.114f
C9041 _307_/a_193_47# _307_/a_761_289# 0.18f
C9042 _192_/a_505_280# _192_/a_476_47# 9.37e-20
C9043 _192_/a_174_21# _192_/a_639_47# 2.58e-19
C9044 net9 _332_/a_193_47# 2.35e-19
C9045 _323_/a_448_47# _323_/a_639_47# 4.61e-19
C9046 VPWR _259_/a_27_297# 0.277f
C9047 VPWR _189_/a_408_47# 0.00334f
C9048 _333_/a_761_289# clknet_2_2__leaf_clk 1.54e-20
C9049 _115_ clknet_2_2__leaf_clk 8.04e-20
C9050 _304_/a_761_289# _001_ 6.85e-20
C9051 VPWR _315_/a_1217_47# 2.13e-19
C9052 _293_/a_81_21# net47 1.83e-20
C9053 _329_/a_543_47# _031_ 1.22e-19
C9054 _318_/a_27_47# clknet_2_0__leaf_clk 0.248f
C9055 net26 _086_ 6.86e-21
C9056 _230_/a_59_75# en_co_clk 0.0101f
C9057 _051_ _099_ 0.012f
C9058 _306_/a_448_47# _065_ 2.9e-20
C9059 _303_/a_1108_47# net4 1.61e-19
C9060 _078_ _310_/a_193_47# 0.00812f
C9061 _186_/a_109_297# _100_ 0.00279f
C9062 state\[2\] _107_ 0.0225f
C9063 _036_ _340_/a_1182_261# 7.23e-19
C9064 _023_ net28 2.04e-20
C9065 clkbuf_2_2__f_clk/a_110_47# _330_/a_543_47# 0.00978f
C9066 _093_ _317_/a_1108_47# 8.22e-22
C9067 _326_/a_651_413# _074_ 0.0022f
C9068 net30 _072_ 0.00455f
C9069 _320_/a_761_289# _320_/a_805_47# 3.69e-19
C9070 _320_/a_193_47# _320_/a_1217_47# 2.36e-20
C9071 _320_/a_543_47# _320_/a_639_47# 0.0138f
C9072 _309_/a_448_47# _081_ 2.48e-21
C9073 _309_/a_1283_21# _006_ 4.1e-20
C9074 _001_ _298_/a_215_47# 2.78e-21
C9075 net32 _108_ 2.14e-19
C9076 _323_/a_193_47# _303_/a_761_289# 4e-21
C9077 _323_/a_27_47# _303_/a_543_47# 1.23e-20
C9078 _323_/a_543_47# _303_/a_27_47# 1.92e-20
C9079 _323_/a_761_289# _303_/a_193_47# 1.8e-21
C9080 _026_ _058_ 4.85e-19
C9081 _053_ _069_ 0.00188f
C9082 net50 net18 1.09f
C9083 net12 _249_/a_109_297# 0.00238f
C9084 _339_/a_27_47# _339_/a_652_21# 0.181f
C9085 _248_/a_109_297# _101_ 0.0373f
C9086 _322_/a_193_47# _101_ 0.0138f
C9087 _028_ trim_mask\[4\] 0.0918f
C9088 net13 _320_/a_27_47# 0.00721f
C9089 _322_/a_761_289# _041_ 5.07e-21
C9090 _187_/a_212_413# _132_ 8.94e-20
C9091 _237_/a_439_47# _090_ 0.00553f
C9092 net47 mask\[4\] 0.243f
C9093 _094_ net45 1.73e-20
C9094 VPWR _232_/a_114_297# 0.0058f
C9095 _317_/a_543_47# state\[1\] 1.69e-19
C9096 _317_/a_1270_413# clknet_2_0__leaf_clk 6.2e-19
C9097 _317_/a_448_47# net45 2.47e-19
C9098 net4 _190_/a_465_47# 1.89e-21
C9099 VPWR net33 1.02f
C9100 _308_/a_1283_21# _307_/a_1283_21# 5.14e-19
C9101 _305_/a_193_47# net30 1.22e-19
C9102 clknet_0_clk en_co_clk 0.0377f
C9103 VPWR trim_mask\[1\] 1.98f
C9104 _321_/a_761_289# mask\[2\] 2.7e-19
C9105 _315_/a_193_47# _315_/a_761_289# 0.181f
C9106 _315_/a_27_47# _315_/a_543_47# 0.115f
C9107 _093_ _192_/a_27_47# 1.76e-20
C9108 VPWR _336_/a_761_289# 0.211f
C9109 _189_/a_27_47# _049_ 4.05e-19
C9110 _033_ _108_ 6.2e-21
C9111 _116_ _275_/a_299_297# 5.83e-20
C9112 _110_ _275_/a_384_47# 7.91e-21
C9113 _276_/a_59_75# net50 4.67e-19
C9114 _117_ _275_/a_81_21# 0.014f
C9115 ctlp[7] net20 4.56e-19
C9116 VPWR _290_/a_27_413# 0.219f
C9117 _303_/a_1108_47# _063_ 1.29e-21
C9118 net51 _070_ 1.36e-20
C9119 clkbuf_2_1__f_clk/a_110_47# _049_ 0.00147f
C9120 net28 _046_ 0.389f
C9121 _303_/a_1108_47# _338_/a_381_47# 5.79e-20
C9122 output8/a_27_47# _334_/a_1283_21# 9.9e-19
C9123 net8 _334_/a_27_47# 0.013f
C9124 _024_ _118_ 1.14e-20
C9125 _110_ _178_/a_150_297# 0.00108f
C9126 _116_ _178_/a_68_297# 3.67e-20
C9127 net22 _039_ 0.412f
C9128 _333_/a_193_47# _333_/a_1270_413# 1.46e-19
C9129 _333_/a_543_47# _333_/a_448_47# 0.0498f
C9130 _333_/a_761_289# _333_/a_651_413# 0.0977f
C9131 _333_/a_1283_21# _333_/a_1108_47# 0.234f
C9132 VPWR clone1/a_27_47# 0.26f
C9133 _062_ _073_ 5.27e-20
C9134 net44 _045_ 2.82e-20
C9135 _094_ _065_ 0.191f
C9136 _103_ _088_ 0.121f
C9137 net16 _332_/a_1217_47# 1.59e-19
C9138 net43 _101_ 0.139f
C9139 state\[2\] net13 0.127f
C9140 net44 _249_/a_109_297# 2.66e-20
C9141 _046_ _158_/a_68_297# 0.106f
C9142 net12 mask\[4\] 0.105f
C9143 _050_ _098_ 0.201f
C9144 _078_ _311_/a_543_47# 4.13e-20
C9145 _074_ _315_/a_761_289# 0.00545f
C9146 _093_ _315_/a_27_47# 8.32e-20
C9147 _265_/a_299_297# trim_val\[0\] 0.00926f
C9148 calibrate _315_/a_193_47# 0.26f
C9149 _326_/a_193_47# _251_/a_27_297# 5.49e-20
C9150 _327_/a_193_47# net40 2.47e-20
C9151 _324_/a_805_47# net44 0.00374f
C9152 _161_/a_68_297# net33 0.00612f
C9153 _324_/a_1283_21# _312_/a_1283_21# 9.77e-20
C9154 _324_/a_543_47# _312_/a_1108_47# 4.48e-20
C9155 _334_/a_761_289# net34 5.32e-21
C9156 _063_ _190_/a_465_47# 0.0185f
C9157 _324_/a_193_47# net19 5.02e-19
C9158 _059_ _206_/a_27_93# 0.00252f
C9159 _330_/a_1108_47# net18 1.78e-36
C9160 clknet_2_1__leaf_clk net26 0.105f
C9161 _308_/a_543_47# _308_/a_805_47# 0.00171f
C9162 _308_/a_761_289# _308_/a_1217_47# 4.2e-19
C9163 _308_/a_1108_47# _308_/a_1270_413# 0.00645f
C9164 net12 _220_/a_199_47# 2.76e-19
C9165 _050_ clknet_0_clk 0.783f
C9166 _258_/a_27_297# _025_ 0.00121f
C9167 net3 _337_/a_1283_21# 6.01e-19
C9168 _025_ _024_ 6.82e-20
C9169 net15 _319_/a_651_413# 0.00187f
C9170 _094_ _319_/a_27_47# 3.12e-21
C9171 clknet_2_0__leaf_clk _315_/a_543_47# 0.00107f
C9172 _014_ _315_/a_761_289# 1.89e-20
C9173 net45 _315_/a_193_47# 0.0259f
C9174 _192_/a_505_280# _065_ 0.00195f
C9175 _090_ _095_ 0.132f
C9176 _089_ _092_ 1.2e-20
C9177 _326_/a_1283_21# clknet_2_1__leaf_clk 4.23e-20
C9178 _305_/a_193_47# _072_ 0.134f
C9179 mask\[0\] net51 6.26e-20
C9180 _231_/a_161_47# cal_count\[3\] 0.0022f
C9181 net15 _096_ 0.00182f
C9182 _235_/a_79_21# _096_ 0.00268f
C9183 net47 _020_ 0.00472f
C9184 _058_ net40 0.00678f
C9185 _300_/a_377_297# net2 0.00683f
C9186 _322_/a_639_47# net44 0.00274f
C9187 net44 mask\[4\] 0.42f
C9188 VPWR _319_/a_639_47# 2.37e-19
C9189 _318_/a_639_47# net45 9.54e-19
C9190 net27 _313_/a_1283_21# 1.17e-20
C9191 _309_/a_193_47# _308_/a_1283_21# 5.28e-20
C9192 _309_/a_27_47# _308_/a_1108_47# 4.8e-19
C9193 _074_ calibrate 0.299f
C9194 _030_ _029_ 3.04e-21
C9195 _015_ _099_ 3.09e-20
C9196 net43 _320_/a_27_47# 2.28e-20
C9197 _128_ _338_/a_1602_47# 3.23e-20
C9198 _325_/a_448_47# _321_/a_193_47# 6.78e-20
C9199 _305_/a_27_47# _305_/a_761_289# 0.0535f
C9200 _078_ _310_/a_1462_47# 2.33e-19
C9201 _237_/a_76_199# _237_/a_535_374# 6.64e-19
C9202 net2 _132_ 0.00922f
C9203 _242_/a_79_21# _099_ 5.38e-19
C9204 _255_/a_27_47# _053_ 0.00554f
C9205 _093_ clknet_2_0__leaf_clk 0.0107f
C9206 calibrate _014_ 0.00963f
C9207 VPWR _069_ 0.288f
C9208 _074_ net45 0.0117f
C9209 _337_/a_651_413# en_co_clk 1.93e-19
C9210 _303_/a_448_47# net19 0.0028f
C9211 VPWR output33/a_27_47# 0.384f
C9212 ctlp[3] net16 2.35e-19
C9213 _291_/a_285_47# net47 1.21e-20
C9214 clkbuf_0_clk/a_110_47# _001_ 6.44e-21
C9215 _001_ cal_count\[3\] 3.63e-20
C9216 _332_/a_27_47# net40 0.0196f
C9217 net50 trim_mask\[0\] 0.00851f
C9218 cal _316_/a_543_47# 5.95e-20
C9219 net12 _020_ 5.58e-20
C9220 _339_/a_27_47# _339_/a_1056_47# 0.00248f
C9221 net13 _320_/a_1217_47# 1.84e-20
C9222 net34 rebuffer1/a_75_212# 4.93e-19
C9223 _126_ output40/a_27_47# 0.0463f
C9224 _341_/a_543_47# _092_ 4.93e-21
C9225 _014_ net45 0.346f
C9226 net43 _307_/a_193_47# 2.76e-19
C9227 _078_ _224_/a_113_297# 0.05f
C9228 cal_itt\[1\] _304_/a_193_47# 3.34e-19
C9229 result[7] net15 1.8e-20
C9230 _122_ _332_/a_193_47# 8.3e-20
C9231 clk _048_ 0.137f
C9232 _337_/a_448_47# _076_ 3.97e-20
C9233 trim_mask\[4\] _279_/a_314_297# 1.27e-19
C9234 _074_ _065_ 0.0585f
C9235 _190_/a_655_47# net19 0.00661f
C9236 _038_ _231_/a_161_47# 1.62e-19
C9237 VPWR _329_/a_805_47# 1.87e-19
C9238 net8 _334_/a_1217_47# 5.59e-19
C9239 _319_/a_651_413# _049_ 2.26e-19
C9240 net47 en_co_clk 1.35e-19
C9241 clk _330_/a_27_47# 0.00365f
C9242 _140_/a_150_297# _040_ 4.96e-19
C9243 _319_/a_1108_47# net30 1.04e-20
C9244 _303_/a_27_47# _303_/a_761_289# 0.0535f
C9245 _091_ _062_ 0.00153f
C9246 _312_/a_639_47# _045_ 1.15e-19
C9247 _096_ _049_ 0.0741f
C9248 net44 _020_ 0.0153f
C9249 mask\[5\] _312_/a_193_47# 1.47e-20
C9250 ctlp[0] result[7] 0.144f
C9251 output23/a_27_47# net45 6.32e-21
C9252 net42 _049_ 0.0459f
C9253 _164_/a_161_47# _090_ 0.00462f
C9254 _048_ net4 0.00405f
C9255 cal_itt\[0\] clkbuf_2_3__f_clk/a_110_47# 0.00811f
C9256 _337_/a_1283_21# _062_ 4.43e-19
C9257 net15 net22 4.98e-20
C9258 VPWR _168_/a_297_47# 1.7e-19
C9259 _326_/a_1108_47# mask\[6\] 6.58e-20
C9260 _326_/a_27_47# _022_ 6.41e-22
C9261 calibrate _243_/a_27_297# 0.0313f
C9262 _324_/a_27_47# _324_/a_543_47# 0.115f
C9263 _324_/a_193_47# _324_/a_761_289# 0.186f
C9264 net13 _248_/a_27_297# 0.0128f
C9265 net13 _322_/a_27_47# 0.0193f
C9266 net4 _330_/a_27_47# 2.28e-19
C9267 state\[0\] _316_/a_1108_47# 0.00316f
C9268 VPWR _078_ 4.55f
C9269 _308_/a_448_47# net43 5.45e-19
C9270 _308_/a_543_47# net23 6.34e-19
C9271 _308_/a_651_413# _005_ 1.23e-20
C9272 net10 ctln[3] 3.57e-21
C9273 net12 en_co_clk 0.013f
C9274 net45 _315_/a_1462_47# 0.00342f
C9275 _319_/a_193_47# clknet_2_0__leaf_clk 0.606f
C9276 _123_ _132_ 9.06e-21
C9277 cal_itt\[1\] net18 2.96e-20
C9278 trim_mask\[1\] _029_ 5.78e-21
C9279 _338_/a_476_47# _001_ 2.17e-20
C9280 _107_ trim_val\[4\] 9.3e-19
C9281 _181_/a_68_297# cal_count\[3\] 1.25e-21
C9282 _078_ net53 0.229f
C9283 _325_/a_27_47# _159_/a_27_47# 4.34e-20
C9284 net9 _286_/a_505_21# 2.47e-19
C9285 _327_/a_1108_47# net18 5.62e-19
C9286 _253_/a_81_21# _314_/a_193_47# 2.75e-22
C9287 _323_/a_805_47# mask\[4\] 2.83e-19
C9288 _321_/a_448_47# mask\[3\] 1.66e-20
C9289 _305_/a_543_47# _305_/a_805_47# 0.00171f
C9290 _305_/a_761_289# _305_/a_1217_47# 4.2e-19
C9291 _305_/a_1108_47# _305_/a_1270_413# 0.00645f
C9292 VPWR _255_/a_27_47# 0.00295f
C9293 net36 net38 0.0522f
C9294 _048_ _063_ 0.268f
C9295 VPWR _313_/a_651_413# 0.143f
C9296 _007_ net14 7.62e-19
C9297 output35/a_27_47# net34 0.018f
C9298 _309_/a_543_47# _309_/a_1108_47# 7.99e-20
C9299 _309_/a_193_47# _309_/a_651_413# 0.0276f
C9300 net5 output35/a_27_47# 0.00159f
C9301 _312_/a_761_289# _084_ 2.17e-20
C9302 net44 en_co_clk 0.165f
C9303 _110_ _334_/a_193_47# 0.00154f
C9304 _000_ net19 0.0338f
C9305 net2 clknet_2_1__leaf_clk 0.0109f
C9306 _136_ _267_/a_59_75# 7.02e-19
C9307 _248_/a_27_297# _248_/a_109_297# 0.171f
C9308 _176_/a_27_47# _056_ 0.208f
C9309 trim_mask\[0\] _181_/a_150_297# 9.24e-19
C9310 _322_/a_27_47# _322_/a_193_47# 0.737f
C9311 _322_/a_193_47# _248_/a_27_297# 3.05e-19
C9312 _322_/a_27_47# _248_/a_109_297# 2.38e-19
C9313 trim_mask\[3\] trim_mask\[2\] 0.0993f
C9314 _104_ _262_/a_109_297# 4.63e-19
C9315 _065_ _243_/a_27_297# 1.46e-19
C9316 _257_/a_27_297# _257_/a_109_297# 0.171f
C9317 _168_/a_27_413# _049_ 1.45e-19
C9318 _335_/a_1108_47# net18 0.00662f
C9319 clkbuf_2_3__f_clk/a_110_47# _108_ 1.24e-19
C9320 mask\[3\] net14 2.84e-21
C9321 net12 _050_ 0.0242f
C9322 _269_/a_81_21# trim_val\[1\] 0.184f
C9323 VPWR _270_/a_59_75# 0.25f
C9324 _259_/a_27_297# _259_/a_373_47# 0.0134f
C9325 net31 _333_/a_1108_47# 0.00298f
C9326 _239_/a_694_21# calibrate 9.72e-20
C9327 net35 _162_/a_27_47# 6.06e-22
C9328 net22 _049_ 2.83e-19
C9329 cal_itt\[1\] _304_/a_1462_47# 4.99e-19
C9330 _262_/a_109_297# net55 0.0133f
C9331 _140_/a_68_297# _246_/a_27_297# 7.2e-21
C9332 _050_ _331_/a_1108_47# 7.7e-19
C9333 clkbuf_2_1__f_clk/a_110_47# _319_/a_543_47# 0.0132f
C9334 _081_ _212_/a_113_297# 1.76e-20
C9335 _125_ net34 0.0132f
C9336 input2/a_27_47# _129_ 3.05e-19
C9337 _325_/a_543_47# _101_ 2.6e-19
C9338 _325_/a_193_47# net52 5.69e-20
C9339 _305_/a_1108_47# _197_/a_113_297# 8.6e-23
C9340 _301_/a_47_47# en_co_clk 0.00143f
C9341 net42 _262_/a_193_297# 0.0041f
C9342 _036_ _339_/a_476_47# 9.17e-19
C9343 cal_count\[1\] _339_/a_1182_261# 0.00358f
C9344 mask\[3\] _143_/a_68_297# 3.51e-21
C9345 _315_/a_1108_47# _096_ 4.88e-19
C9346 clkbuf_2_0__f_clk/a_110_47# _319_/a_1283_21# 0.00124f
C9347 en_co_clk _263_/a_79_21# 3.16e-19
C9348 net43 _248_/a_27_297# 8.88e-19
C9349 _341_/a_27_47# en_co_clk 2.39e-19
C9350 _279_/a_27_47# trim_val\[4\] 0.085f
C9351 _303_/a_543_47# _303_/a_805_47# 0.00171f
C9352 _303_/a_761_289# _303_/a_1217_47# 4.2e-19
C9353 _303_/a_1108_47# _303_/a_1270_413# 0.00645f
C9354 _291_/a_35_297# trimb[1] 6.6e-19
C9355 net28 result[6] 0.0457f
C9356 _243_/a_27_297# _243_/a_109_297# 0.171f
C9357 _050_ net44 4.63e-19
C9358 _087_ _226_/a_303_47# 9.6e-20
C9359 _090_ _226_/a_27_47# 8.61e-20
C9360 net2 _202_/a_382_297# 7.04e-20
C9361 _317_/a_193_47# _316_/a_27_47# 6.94e-21
C9362 _317_/a_27_47# _316_/a_193_47# 1.35e-20
C9363 VPWR fanout47/a_27_47# 0.339f
C9364 cal_itt\[0\] clkbuf_0_clk/a_110_47# 0.0265f
C9365 net54 _337_/a_448_47# 5.27e-21
C9366 _060_ _337_/a_1108_47# 3.21e-21
C9367 clknet_2_0__leaf_clk _206_/a_27_93# 5.13e-20
C9368 cal_itt\[0\] cal_count\[3\] 8.11e-20
C9369 _305_/a_1108_47# _202_/a_79_21# 6.84e-19
C9370 net16 cal_count\[0\] 0.081f
C9371 net52 _076_ 0.0165f
C9372 VPWR _316_/a_1283_21# 0.375f
C9373 net12 _228_/a_297_47# 8.49e-19
C9374 _136_ net37 2.66e-20
C9375 _306_/a_193_47# _003_ 0.221f
C9376 _327_/a_639_47# clknet_2_3__leaf_clk 3.69e-20
C9377 _302_/a_109_297# _108_ 9.02e-19
C9378 _005_ net43 9e-19
C9379 _103_ _227_/a_368_53# 2.7e-19
C9380 _237_/a_76_199# _281_/a_253_47# 9.7e-19
C9381 _046_ _085_ 0.0687f
C9382 _322_/a_1283_21# _249_/a_27_297# 1.05e-20
C9383 _316_/a_448_47# net41 0.0212f
C9384 _238_/a_75_212# calibrate 0.0273f
C9385 _329_/a_193_47# _259_/a_109_297# 3.97e-19
C9386 state\[2\] net3 6.86e-20
C9387 cal_itt\[1\] trim_mask\[0\] 7.2e-20
C9388 _212_/a_113_297# _016_ 5.52e-20
C9389 _330_/a_193_47# net19 0.0203f
C9390 _058_ _280_/a_75_212# 1.64e-19
C9391 VPWR output7/a_27_47# 0.292f
C9392 VPWR _004_ 0.353f
C9393 _002_ _065_ 0.0293f
C9394 _050_ _263_/a_79_21# 5.24e-20
C9395 state\[1\] _096_ 2.16e-19
C9396 _335_/a_193_47# _280_/a_75_212# 5.89e-20
C9397 _309_/a_639_47# net43 0.00156f
C9398 trim_mask\[0\] _052_ 1.94e-25
C9399 _325_/a_1108_47# net21 0.00558f
C9400 _325_/a_651_413# _046_ 4.66e-20
C9401 _094_ _282_/a_68_297# 0.0449f
C9402 _061_ net16 2.82e-19
C9403 _327_/a_761_289# _024_ 0.00253f
C9404 _327_/a_1108_47# trim_mask\[0\] 0.00583f
C9405 clk _335_/a_27_47# 1.35e-21
C9406 _087_ _228_/a_79_21# 0.0111f
C9407 _053_ _304_/a_639_47# 8.12e-19
C9408 _101_ _062_ 3.72e-20
C9409 _238_/a_75_212# net45 0.0324f
C9410 mask\[7\] _314_/a_1108_47# 8.56e-19
C9411 fanout44/a_27_47# _101_ 8.89e-19
C9412 output11/a_27_47# output12/a_27_47# 4.72e-21
C9413 _053_ _340_/a_193_47# 1.6e-19
C9414 result[4] net14 8.01e-20
C9415 _320_/a_193_47# _077_ 0.00176f
C9416 net50 trim_mask\[4\] 0.0786f
C9417 _277_/a_75_212# _335_/a_27_47# 2.48e-20
C9418 _320_/a_761_289# _076_ 3.49e-21
C9419 _258_/a_109_297# _058_ 2.93e-19
C9420 _248_/a_373_47# mask\[4\] 5.55e-19
C9421 _322_/a_761_289# _322_/a_805_47# 3.69e-19
C9422 _322_/a_193_47# _322_/a_1217_47# 2.36e-20
C9423 _322_/a_543_47# _322_/a_639_47# 0.0138f
C9424 cal_itt\[0\] _038_ 6.38e-20
C9425 _257_/a_27_297# _025_ 0.116f
C9426 _320_/a_448_47# _017_ 0.158f
C9427 cal_count\[3\] _108_ 0.00102f
C9428 net22 _315_/a_1108_47# 8.95e-21
C9429 net4 _335_/a_27_47# 2.87e-19
C9430 net49 _112_ 5.7e-19
C9431 net48 _269_/a_299_297# 1.06e-19
C9432 _272_/a_299_297# net49 9.52e-20
C9433 _272_/a_81_21# _272_/a_299_297# 0.0821f
C9434 mask\[5\] _152_/a_68_297# 0.231f
C9435 trim_mask\[1\] _336_/a_1108_47# 2.78e-19
C9436 _125_ _133_ 4.17e-21
C9437 cal_itt\[2\] _041_ 5.23e-20
C9438 VPWR _287_/a_75_212# 0.209f
C9439 _336_/a_193_47# _336_/a_448_47# 0.0642f
C9440 _336_/a_761_289# _336_/a_1108_47# 0.0512f
C9441 _336_/a_27_47# _336_/a_651_413# 9.73e-19
C9442 cal_itt\[0\] _338_/a_476_47# 3.8e-19
C9443 _050_ clknet_2_2__leaf_clk 0.00221f
C9444 _040_ _246_/a_373_47# 0.00356f
C9445 _050_ _260_/a_584_47# 1.85e-20
C9446 _319_/a_193_47# _319_/a_639_47# 2.28e-19
C9447 _319_/a_761_289# _319_/a_1270_413# 2.6e-19
C9448 _319_/a_543_47# _319_/a_651_413# 0.0572f
C9449 _308_/a_448_47# _080_ 7.37e-19
C9450 trim_mask\[0\] rebuffer2/a_75_212# 2.87e-20
C9451 _290_/a_207_413# _290_/a_297_47# 0.00476f
C9452 mask\[3\] net52 0.261f
C9453 _082_ _101_ 8.79e-21
C9454 _237_/a_535_374# _048_ 3.1e-19
C9455 trim_mask\[0\] _332_/a_1283_21# 0.107f
C9456 fanout43/a_27_47# net14 0.00189f
C9457 _329_/a_27_47# _329_/a_193_47# 0.906f
C9458 _273_/a_59_75# _334_/a_543_47# 2.63e-20
C9459 _237_/a_505_21# net3 0.0158f
C9460 _286_/a_505_21# _122_ 0.039f
C9461 trim_val\[4\] _118_ 0.385f
C9462 _093_ _078_ 4.53e-21
C9463 _012_ net22 9.79e-21
C9464 net54 net4 1.14e-19
C9465 net27 net14 0.00986f
C9466 _293_/a_81_21# cal_count\[1\] 0.00317f
C9467 _243_/a_373_47# net55 0.00122f
C9468 _059_ _337_/a_193_47# 3.64e-19
C9469 clk _068_ 2.05e-20
C9470 _324_/a_1283_21# _020_ 8.91e-19
C9471 _006_ _310_/a_27_47# 1.34e-21
C9472 trim_val\[0\] en_co_clk 7.78e-20
C9473 clknet_2_2__leaf_clk _330_/a_805_47# 0.00252f
C9474 trim_mask\[4\] _330_/a_1108_47# 1.95e-22
C9475 _048_ _279_/a_396_47# 0.00276f
C9476 net15 clknet_0_clk 0.0846f
C9477 _235_/a_79_21# clknet_0_clk 8.61e-20
C9478 net30 sample 0.017f
C9479 state\[2\] _062_ 2.69e-21
C9480 _254_/a_109_297# net42 5.63e-19
C9481 _328_/a_761_289# net46 0.169f
C9482 net30 net40 0.0489f
C9483 _106_ _105_ 0.14f
C9484 net24 clknet_2_0__leaf_clk 1.23e-19
C9485 _038_ _108_ 1.47e-19
C9486 _270_/a_59_75# _029_ 7.15e-20
C9487 _197_/a_113_297# _069_ 0.1f
C9488 _104_ _336_/a_448_47# 2.61e-19
C9489 ctln[1] _317_/a_761_289# 2.4e-20
C9490 _013_ net41 0.107f
C9491 _074_ _313_/a_639_47# 1.35e-20
C9492 _334_/a_193_47# clknet_2_2__leaf_clk 0.00461f
C9493 _053_ _136_ 0.0545f
C9494 input2/a_27_47# _297_/a_47_47# 1.11e-19
C9495 _025_ trim_val\[4\] 1.11e-20
C9496 net4 _068_ 0.00707f
C9497 VPWR _304_/a_639_47# 3.32e-19
C9498 _205_/a_27_47# rebuffer5/a_161_47# 1.96e-19
C9499 _187_/a_212_413# clkc 7.77e-19
C9500 _328_/a_1108_47# _327_/a_1283_21# 2.15e-22
C9501 _325_/a_761_289# net13 0.00324f
C9502 VPWR _340_/a_193_47# 0.311f
C9503 net30 _003_ 0.0681f
C9504 _090_ _052_ 1.32e-19
C9505 _282_/a_150_297# clknet_2_0__leaf_clk 8.17e-21
C9506 output15/a_27_47# _223_/a_109_297# 5.98e-20
C9507 _197_/a_199_47# _067_ 6.92e-19
C9508 _129_ trimb[4] 0.00203f
C9509 _197_/a_199_47# _070_ 3.51e-21
C9510 _250_/a_373_47# _021_ 0.00133f
C9511 _040_ rebuffer5/a_161_47# 1.1e-20
C9512 trim_val\[1\] net32 0.00288f
C9513 net52 _310_/a_1283_21# 3.73e-19
C9514 _308_/a_1283_21# mask\[1\] 0.00118f
C9515 _098_ _049_ 0.0909f
C9516 _269_/a_299_297# _172_/a_68_297# 0.00615f
C9517 _321_/a_543_47# _018_ 2.86e-19
C9518 _328_/a_1270_413# _058_ 3.74e-20
C9519 _289_/a_68_297# _289_/a_150_297# 0.00477f
C9520 _322_/a_448_47# _019_ 0.159f
C9521 net9 _042_ 3.59e-19
C9522 VPWR _261_/a_113_47# 1.32e-19
C9523 net24 _146_/a_68_297# 0.00108f
C9524 net13 _077_ 2.18e-20
C9525 trim_mask\[2\] _335_/a_1283_21# 2.02e-20
C9526 _053_ _119_ 0.00168f
C9527 _008_ mask\[5\] 1.37e-19
C9528 _341_/a_543_47# net46 0.153f
C9529 _052_ _242_/a_382_297# 0.00147f
C9530 _246_/a_27_297# _246_/a_109_47# 0.00393f
C9531 clknet_2_1__leaf_clk mask\[0\] 1.88e-19
C9532 mask\[0\] _319_/a_761_289# 0.0221f
C9533 _078_ _319_/a_193_47# 1.47e-21
C9534 _020_ _044_ 1.01e-19
C9535 _043_ net26 9.81e-19
C9536 _202_/a_382_297# _070_ 0.0149f
C9537 output24/a_27_47# clknet_2_1__leaf_clk 2.58e-19
C9538 _068_ _063_ 0.647f
C9539 cal_count\[0\] net40 0.0315f
C9540 clknet_0_clk _049_ 0.0925f
C9541 _320_/a_639_47# mask\[1\] 7.19e-21
C9542 _058_ net19 2.29e-20
C9543 _307_/a_193_47# _137_/a_68_297# 1.18e-19
C9544 _336_/a_193_47# _033_ 0.259f
C9545 _321_/a_651_413# net15 1.36e-20
C9546 cal_itt\[0\] _341_/a_448_47# 7.48e-21
C9547 output15/a_27_47# ctlp[1] 0.166f
C9548 _335_/a_193_47# net19 2.89e-20
C9549 net44 _311_/a_1108_47# 0.235f
C9550 _005_ _080_ 0.156f
C9551 _322_/a_1283_21# rebuffer5/a_161_47# 1.06e-20
C9552 trim_mask\[2\] _108_ 0.167f
C9553 trim_val\[2\] net16 0.111f
C9554 _327_/a_193_47# _107_ 5.4e-21
C9555 _048_ _034_ 2.06e-21
C9556 _093_ _316_/a_1283_21# 9.52e-20
C9557 _094_ _337_/a_27_47# 0.222f
C9558 _329_/a_761_289# _329_/a_805_47# 3.69e-19
C9559 _329_/a_193_47# _329_/a_1217_47# 2.36e-20
C9560 _329_/a_543_47# _329_/a_639_47# 0.0138f
C9561 VPWR _321_/a_639_47# 2.07e-19
C9562 _115_ _334_/a_448_47# 5.13e-19
C9563 _323_/a_27_47# _311_/a_1283_21# 9.27e-19
C9564 _003_ _072_ 6.33e-20
C9565 _218_/a_199_47# _083_ 0.003f
C9566 clknet_2_1__leaf_clk _313_/a_448_47# 0.0149f
C9567 _053_ _087_ 3.09e-20
C9568 mask\[7\] _224_/a_113_297# 0.0502f
C9569 _306_/a_27_47# clk 1.37e-20
C9570 VPWR _337_/a_639_47# 2.44e-19
C9571 _247_/a_27_297# _101_ 0.132f
C9572 _286_/a_218_47# net18 3.63e-19
C9573 _327_/a_1108_47# _265_/a_81_21# 4.92e-20
C9574 _281_/a_103_199# _281_/a_253_47# 0.0606f
C9575 _061_ net40 0.0224f
C9576 _317_/a_27_47# net14 8.86e-19
C9577 en_co_clk _131_ 0.00178f
C9578 _014_ _316_/a_448_47# 0.00439f
C9579 net45 _316_/a_1108_47# 0.236f
C9580 fanout43/a_27_47# net52 6.06e-19
C9581 _097_ _096_ 0.0117f
C9582 _326_/a_27_47# net14 0.00737f
C9583 _058_ _107_ 4.44e-19
C9584 _325_/a_761_289# net43 0.164f
C9585 VPWR _117_ 0.231f
C9586 _309_/a_27_47# _007_ 1.26e-19
C9587 _305_/a_761_289# _073_ 2.27e-20
C9588 _322_/a_639_47# mask\[2\] 4.73e-19
C9589 _058_ _333_/a_1108_47# 3.95e-19
C9590 net27 net52 3.96e-19
C9591 net2 clkc 3.18e-19
C9592 _051_ net41 0.116f
C9593 VPWR _136_ 0.642f
C9594 net15 _245_/a_27_297# 6.52e-19
C9595 _104_ _033_ 0.0252f
C9596 output29/a_27_47# _078_ 1.41e-19
C9597 _309_/a_193_47# net25 3.78e-20
C9598 _309_/a_27_47# mask\[3\] 1.75e-19
C9599 _329_/a_651_413# net9 0.00203f
C9600 trim_mask\[4\] _052_ 0.144f
C9601 _253_/a_81_21# net26 0.0495f
C9602 _134_ _332_/a_193_47# 4.73e-20
C9603 VPWR _245_/a_109_47# 6.05e-19
C9604 trim_mask\[2\] _031_ 0.12f
C9605 _333_/a_193_47# rebuffer2/a_75_212# 3.4e-20
C9606 VPWR _340_/a_796_47# 3.86e-19
C9607 _175_/a_150_297# _108_ 5.09e-19
C9608 _060_ _107_ 0.00674f
C9609 _333_/a_193_47# _332_/a_1283_21# 5.72e-21
C9610 _333_/a_761_289# _108_ 0.00569f
C9611 _275_/a_384_47# trim_mask\[3\] 0.0101f
C9612 _275_/a_299_297# net50 0.0493f
C9613 _115_ _108_ 0.00253f
C9614 VPWR mask\[7\] 0.736f
C9615 _101_ rebuffer6/a_27_47# 3.72e-21
C9616 net50 _178_/a_68_297# 8.75e-19
C9617 _275_/a_81_21# _057_ 1.13e-19
C9618 _034_ _076_ 1.79e-20
C9619 _265_/a_299_297# _332_/a_543_47# 9.16e-20
C9620 _265_/a_299_297# _108_ 0.0687f
C9621 mask\[6\] _078_ 0.307f
C9622 _337_/a_651_413# _049_ 0.00244f
C9623 clk _317_/a_27_47# 0.00834f
C9624 clknet_0_clk _262_/a_193_297# 7.06e-19
C9625 _210_/a_199_47# net22 1.55e-19
C9626 _210_/a_113_297# mask\[0\] 0.0502f
C9627 net23 _212_/a_113_297# 0.00889f
C9628 _335_/a_1108_47# trim_mask\[4\] 4.24e-19
C9629 VPWR _119_ 0.494f
C9630 _270_/a_145_75# _112_ 6.69e-19
C9631 _051_ _171_/a_27_47# 0.0094f
C9632 output32/a_27_47# trim_val\[1\] 1.5e-19
C9633 net9 ctln[3] 0.0104f
C9634 _048_ _281_/a_253_47# 0.00302f
C9635 _321_/a_27_47# _074_ 2.72e-20
C9636 VPWR ctln[6] 0.364f
C9637 _306_/a_27_47# net52 2.88e-20
C9638 _306_/a_761_289# _101_ 1.05e-20
C9639 _246_/a_109_297# _017_ 0.00387f
C9640 _306_/a_543_47# _041_ 1.18e-21
C9641 _200_/a_80_21# _092_ 0.0621f
C9642 _333_/a_805_47# net46 0.00322f
C9643 _100_ clone7/a_27_47# 0.0701f
C9644 _307_/a_1283_21# _039_ 0.0346f
C9645 VPWR _331_/a_651_413# 0.144f
C9646 _325_/a_1108_47# mask\[4\] 7.84e-19
C9647 _332_/a_639_47# clknet_2_2__leaf_clk 5.75e-19
C9648 _109_ net46 3.12e-20
C9649 mask\[3\] _248_/a_109_47# 4.58e-19
C9650 _322_/a_761_289# mask\[3\] 0.0505f
C9651 net4 _317_/a_27_47# 0.0101f
C9652 _321_/a_193_47# clknet_2_0__leaf_clk 9.79e-21
C9653 _320_/a_1283_21# net51 2e-20
C9654 VPWR _328_/a_193_47# 0.269f
C9655 net27 _312_/a_1270_413# 8.03e-20
C9656 _062_ _190_/a_655_47# 0.0401f
C9657 net2 _298_/a_215_47# 0.00118f
C9658 net31 output34/a_27_47# 1.78e-19
C9659 cal_itt\[0\] _303_/a_1283_21# 0.102f
C9660 _233_/a_109_47# net14 9.7e-20
C9661 _074_ _013_ 1.14e-20
C9662 _104_ _103_ 0.0652f
C9663 net15 net44 2.1e-21
C9664 _094_ _337_/a_1217_47# 3.29e-19
C9665 _329_/a_448_47# _026_ 0.16f
C9666 _300_/a_377_297# clknet_2_3__leaf_clk 2.43e-21
C9667 VPWR _087_ 0.506f
C9668 net13 _060_ 0.202f
C9669 _337_/a_193_47# clknet_2_0__leaf_clk 0.11f
C9670 _115_ _031_ 0.00257f
C9671 _059_ _090_ 0.0303f
C9672 net28 _314_/a_1108_47# 1.46e-19
C9673 result[6] _314_/a_543_47# 8.65e-19
C9674 _051_ _094_ 9.78e-22
C9675 _309_/a_27_47# _310_/a_1283_21# 1.17e-19
C9676 clknet_2_1__leaf_clk _010_ 0.0338f
C9677 VPWR _312_/a_27_47# 0.43f
C9678 _257_/a_109_297# _058_ 2.86e-19
C9679 _281_/a_253_47# _120_ 3.38e-19
C9680 _103_ net55 0.0766f
C9681 _062_ trim_val\[4\] 8.95e-19
C9682 net12 _306_/a_805_47# 4.47e-19
C9683 _257_/a_109_297# _335_/a_193_47# 5.17e-22
C9684 _014_ _013_ 0.0694f
C9685 _314_/a_1108_47# _158_/a_68_297# 7.54e-20
C9686 VPWR _323_/a_193_47# 0.274f
C9687 VPWR _266_/a_150_297# 0.00152f
C9688 _231_/a_161_47# en_co_clk 0.00148f
C9689 _195_/a_76_199# _190_/a_655_47# 6.49e-20
C9690 _313_/a_27_47# _313_/a_448_47# 0.0867f
C9691 _313_/a_193_47# _313_/a_1108_47# 0.125f
C9692 _015_ net41 0.00932f
C9693 _336_/a_27_47# clkbuf_2_2__f_clk/a_110_47# 0.0189f
C9694 _312_/a_27_47# net53 1.2e-19
C9695 clk _318_/a_543_47# 0.0298f
C9696 cal_itt\[2\] _190_/a_465_47# 0.012f
C9697 cal_itt\[1\] _190_/a_27_47# 7.64e-19
C9698 cal_itt\[0\] _190_/a_215_47# 1.53e-19
C9699 net12 _049_ 0.214f
C9700 net12 _318_/a_761_289# 9.81e-19
C9701 net2 _130_ 0.137f
C9702 _323_/a_193_47# net53 0.00126f
C9703 _321_/a_193_47# _146_/a_68_297# 4.27e-20
C9704 _326_/a_27_47# net52 3.61e-19
C9705 _259_/a_27_297# net18 0.00703f
C9706 VPWR _301_/a_129_47# 1.83e-19
C9707 _331_/a_543_47# _054_ 1.12e-20
C9708 _169_/a_215_311# _099_ 1.08e-21
C9709 _325_/a_27_47# mask\[2\] 1.68e-19
C9710 _260_/a_93_21# _170_/a_81_21# 4.36e-19
C9711 VPWR _338_/a_1140_413# 0.00336f
C9712 VPWR _263_/a_297_47# 0.00535f
C9713 _306_/a_805_47# net44 0.00316f
C9714 VPWR _341_/a_761_289# 0.213f
C9715 en net3 0.0045f
C9716 _312_/a_27_47# _009_ 0.345f
C9717 _326_/a_448_47# _023_ 0.16f
C9718 _326_/a_1270_413# mask\[7\] 1.46e-19
C9719 _326_/a_651_413# _102_ 1.19e-19
C9720 _340_/a_193_47# _285_/a_113_47# 5.7e-21
C9721 _001_ en_co_clk 6.44e-20
C9722 _136_ _300_/a_47_47# 0.0118f
C9723 net4 _318_/a_543_47# 1.8e-20
C9724 _309_/a_27_47# fanout43/a_27_47# 1.41e-19
C9725 _041_ _286_/a_218_374# 9.13e-19
C9726 output15/a_27_47# _010_ 0.0629f
C9727 _286_/a_505_21# _338_/a_1032_413# 0.00227f
C9728 net47 _124_ 0.0145f
C9729 _330_/a_193_47# _330_/a_761_289# 0.176f
C9730 _330_/a_27_47# _330_/a_543_47# 0.106f
C9731 _208_/a_76_199# _076_ 0.342f
C9732 _066_ net40 4.32e-20
C9733 net43 _314_/a_639_47# 9.54e-19
C9734 _304_/a_805_47# _065_ 3.02e-20
C9735 net44 _049_ 0.0558f
C9736 clk _317_/a_1217_47# 5.25e-20
C9737 VPWR _308_/a_27_47# 0.509f
C9738 net46 _092_ 9.46e-20
C9739 _068_ _201_/a_113_47# 1.96e-19
C9740 _110_ fanout46/a_27_47# 0.00447f
C9741 net24 _078_ 0.506f
C9742 _320_/a_543_47# net15 6.38e-19
C9743 _340_/a_1032_413# net2 1.06e-19
C9744 _123_ _298_/a_215_47# 0.0215f
C9745 _254_/a_109_297# _098_ 0.002f
C9746 _058_ _118_ 0.00858f
C9747 _079_ _210_/a_199_47# 0.0016f
C9748 net21 net26 2.96e-20
C9749 net16 net40 0.129f
C9750 _319_/a_543_47# clknet_0_clk 8.27e-19
C9751 _071_ _092_ 0.0264f
C9752 _249_/a_27_297# _311_/a_27_47# 0.0111f
C9753 clk cal_itt\[3\] 0.0472f
C9754 VPWR _320_/a_1108_47# 0.294f
C9755 _136_ _029_ 0.0046f
C9756 _097_ _316_/a_761_289# 1.11e-19
C9757 _238_/a_75_212# _316_/a_448_47# 5.77e-19
C9758 _227_/a_109_93# net19 5.86e-21
C9759 trim_mask\[1\] net18 0.204f
C9760 VPWR _339_/a_27_47# 0.404f
C9761 state\[2\] _227_/a_209_311# 4.33e-19
C9762 _327_/a_193_47# _025_ 8.86e-20
C9763 _325_/a_1270_413# _019_ 8.1e-21
C9764 net43 _310_/a_1108_47# 0.257f
C9765 _011_ net14 0.00251f
C9766 net51 _205_/a_27_47# 9.02e-20
C9767 net4 _317_/a_1217_47# 5.18e-19
C9768 net33 _129_ 2.66e-19
C9769 VPWR _328_/a_1462_47# 1.46e-19
C9770 clkbuf_0_clk/a_110_47# net2 3.61e-20
C9771 net2 cal_count\[3\] 0.29f
C9772 output20/a_27_47# _312_/a_651_413# 2.85e-19
C9773 ctlp[6] _312_/a_193_47# 1.31e-19
C9774 _324_/a_543_47# net27 2e-19
C9775 _324_/a_1108_47# _311_/a_1283_21# 1.27e-20
C9776 _263_/a_79_21# _049_ 9.78e-19
C9777 _305_/a_1283_21# clkbuf_0_clk/a_110_47# 0.00428f
C9778 _305_/a_27_47# clk 0.00415f
C9779 _166_/a_161_47# _050_ 0.327f
C9780 _337_/a_805_47# net45 5.61e-21
C9781 _323_/a_1108_47# net26 7.59e-19
C9782 trimb[0] net16 1.1e-19
C9783 _325_/a_761_289# _325_/a_543_47# 0.21f
C9784 _325_/a_193_47# _325_/a_1283_21# 0.0424f
C9785 _325_/a_27_47# _325_/a_1108_47# 0.102f
C9786 _040_ net51 0.00283f
C9787 _110_ _269_/a_299_297# 4.72e-19
C9788 net4 cal_itt\[3\] 7.46e-21
C9789 _025_ _058_ 0.00193f
C9790 _104_ clkbuf_2_3__f_clk/a_110_47# 1.77e-19
C9791 net16 _299_/a_215_297# 0.0116f
C9792 VPWR _307_/a_448_47# 0.0834f
C9793 VPWR _323_/a_1462_47# 1.98e-19
C9794 _302_/a_27_297# trim_mask\[1\] 1.57e-21
C9795 _090_ _192_/a_27_47# 5.02e-20
C9796 _107_ _227_/a_109_93# 0.00575f
C9797 output21/a_27_47# net27 6.42e-21
C9798 _313_/a_27_47# _010_ 0.168f
C9799 _305_/a_27_47# net4 3.13e-22
C9800 _048_ _075_ 0.0203f
C9801 _023_ _074_ 0.175f
C9802 _290_/a_207_413# net38 4.06e-21
C9803 net55 clkbuf_2_3__f_clk/a_110_47# 1.03e-19
C9804 _321_/a_1283_21# _042_ 0.0066f
C9805 _064_ _091_ 0.003f
C9806 _259_/a_27_297# trim_mask\[0\] 4.06e-21
C9807 _064_ _256_/a_109_297# 0.0118f
C9808 _278_/a_109_297# _278_/a_27_47# 5.37e-19
C9809 _321_/a_1270_413# clknet_2_1__leaf_clk 6.85e-20
C9810 trim[3] _057_ 3.31e-19
C9811 trim[2] net34 0.0157f
C9812 VPWR _333_/a_639_47# 8.68e-19
C9813 VPWR _303_/a_27_47# 0.49f
C9814 _340_/a_1032_413# _123_ 0.0867f
C9815 _063_ cal_itt\[3\] 0.0056f
C9816 trim[1] net32 0.16f
C9817 trim_val\[3\] _335_/a_27_47# 0.0124f
C9818 net28 _224_/a_113_297# 0.0628f
C9819 cal_count\[0\] _338_/a_1602_47# 0.0857f
C9820 _008_ _311_/a_761_289# 6.55e-19
C9821 cal_itt\[2\] _048_ 2.04e-20
C9822 calibrate _331_/a_1270_413# 2.39e-20
C9823 _338_/a_27_47# _065_ 1.44e-20
C9824 _069_ net18 1.21e-20
C9825 _337_/a_543_47# _096_ 4.24e-19
C9826 _067_ clkbuf_2_3__f_clk/a_110_47# 0.00377f
C9827 _337_/a_761_289# net55 0.00343f
C9828 VPWR _308_/a_1217_47# 5.6e-20
C9829 _074_ _046_ 5.07e-20
C9830 net2 _338_/a_476_47# 2.54e-20
C9831 _303_/a_27_47# net53 1.37e-21
C9832 net30 net19 0.00891f
C9833 state\[2\] _318_/a_1108_47# 0.00311f
C9834 _305_/a_27_47# net52 5.39e-21
C9835 _341_/a_193_47# _300_/a_377_297# 1.22e-20
C9836 _051_ _243_/a_27_297# 2.4e-20
C9837 _305_/a_27_47# _063_ 4.88e-21
C9838 _307_/a_1283_21# _049_ 1.66e-19
C9839 calibrate _089_ 0.0219f
C9840 _307_/a_761_289# net30 4.59e-21
C9841 _123_ cal_count\[3\] 1.48e-19
C9842 VPWR _309_/a_543_47# 0.195f
C9843 net45 _331_/a_1270_413# 3.47e-19
C9844 net13 _235_/a_297_47# 0.00116f
C9845 trim_mask\[0\] net33 0.0121f
C9846 _074_ _312_/a_761_289# 1.75e-20
C9847 trim_mask\[0\] trim_mask\[1\] 0.0496f
C9848 _238_/a_75_212# _013_ 0.109f
C9849 VPWR _339_/a_586_47# 5.47e-20
C9850 _211_/a_109_297# _079_ 1.66e-20
C9851 _328_/a_1108_47# _113_ 0.00303f
C9852 _328_/a_1283_21# _030_ 6.43e-19
C9853 trim_mask\[2\] _113_ 2.11e-19
C9854 _075_ _076_ 0.0525f
C9855 trim_mask\[0\] _336_/a_761_289# 1.49e-20
C9856 clknet_2_0__leaf_clk _090_ 0.00154f
C9857 en_co_clk _195_/a_218_374# 0.0029f
C9858 _107_ _054_ 0.00434f
C9859 fanout45/a_27_47# _096_ 5.43e-19
C9860 clknet_2_1__leaf_clk net20 0.0971f
C9861 cal_itt\[0\] en_co_clk 0.426f
C9862 _212_/a_199_47# mask\[1\] 0.00963f
C9863 _107_ net30 0.239f
C9864 VPWR _279_/a_206_47# 0.00298f
C9865 net43 _306_/a_193_47# 5.95e-20
C9866 trim_mask\[0\] clone1/a_27_47# 9.29e-20
C9867 VPWR net28 2.08f
C9868 en_co_clk _088_ 9.79e-21
C9869 output40/a_27_47# _131_ 3.38e-21
C9870 _325_/a_1283_21# _325_/a_1462_47# 0.0074f
C9871 _325_/a_1108_47# _325_/a_1217_47# 0.00742f
C9872 VPWR _292_/a_292_297# 0.00902f
C9873 net12 _250_/a_27_297# 0.0117f
C9874 _051_ _336_/a_543_47# 4.44e-21
C9875 net9 _133_ 1.33e-19
C9876 VPWR _324_/a_448_47# 0.0859f
C9877 _104_ cal_count\[3\] 1.88e-20
C9878 VPWR _158_/a_68_297# 0.178f
C9879 _302_/a_109_297# _067_ 0.00139f
C9880 _136_ _194_/a_199_47# 1.49e-19
C9881 _329_/a_1283_21# _110_ 2.51e-19
C9882 mask\[4\] _311_/a_805_47# 0.00207f
C9883 VPWR ctln[0] 0.194f
C9884 net19 _072_ 7.43e-19
C9885 _313_/a_1217_47# _010_ 4.2e-20
C9886 _239_/a_694_21# _051_ 0.116f
C9887 _104_ _331_/a_27_47# 1.07e-19
C9888 cal_count\[3\] net55 6.92e-20
C9889 _324_/a_448_47# net53 7.43e-19
C9890 ctln[2] _179_/a_27_47# 0.00504f
C9891 output8/a_27_47# net34 8.93e-19
C9892 _060_ net3 0.0282f
C9893 _147_/a_27_47# _042_ 0.222f
C9894 _321_/a_193_47# _078_ 3.45e-20
C9895 _304_/a_543_47# _284_/a_68_297# 4.89e-19
C9896 VPWR _322_/a_1108_47# 0.31f
C9897 VPWR _099_ 0.234f
C9898 _081_ clknet_2_1__leaf_clk 1e-19
C9899 _064_ _258_/a_27_297# 0.0867f
C9900 _083_ _311_/a_1283_21# 7.61e-22
C9901 _064_ _024_ 1.83e-19
C9902 _305_/a_805_47# net44 4.25e-19
C9903 _250_/a_27_297# net44 9.27e-20
C9904 _314_/a_1108_47# _085_ 1.44e-20
C9905 net33 _297_/a_47_47# 0.0046f
C9906 _308_/a_761_289# _074_ 0.00835f
C9907 _305_/a_193_47# net19 1.43e-20
C9908 fanout46/a_27_47# clknet_2_2__leaf_clk 0.105f
C9909 net28 _009_ 8.18e-21
C9910 _113_ _333_/a_761_289# 7.33e-21
C9911 _030_ _333_/a_193_47# 0.329f
C9912 _338_/a_476_47# _123_ 9.46e-22
C9913 _316_/a_761_289# _316_/a_639_47# 3.16e-19
C9914 _316_/a_27_47# _316_/a_1217_47# 2.56e-19
C9915 ctln[7] _318_/a_761_289# 8.2e-20
C9916 net13 _318_/a_1283_21# 0.00214f
C9917 net13 net30 0.0102f
C9918 _322_/a_1108_47# net53 9.34e-20
C9919 _050_ _088_ 0.121f
C9920 VPWR _303_/a_1217_47# 1.15e-19
C9921 _030_ _265_/a_81_21# 2.45e-19
C9922 VPWR result[3] 0.268f
C9923 _275_/a_81_21# _032_ 6.04e-19
C9924 net50 _335_/a_639_47# 3.14e-19
C9925 en_co_clk _108_ 7.36e-21
C9926 net44 _319_/a_543_47# 2.16e-20
C9927 mask\[7\] output29/a_27_47# 1.67e-19
C9928 _308_/a_543_47# clknet_2_0__leaf_clk 7.75e-19
C9929 _308_/a_193_47# net45 9.57e-19
C9930 _326_/a_193_47# net43 0.0348f
C9931 net30 _279_/a_27_47# 7.15e-20
C9932 net34 _055_ 0.161f
C9933 _330_/a_1270_413# _027_ 3.05e-19
C9934 _330_/a_651_413# net46 0.0122f
C9935 _301_/a_285_47# _135_ 0.0675f
C9936 clkbuf_0_clk/a_110_47# _067_ 0.00733f
C9937 en_co_clk _244_/a_27_297# 3.94e-20
C9938 _336_/a_1108_47# _119_ 3.82e-20
C9939 _323_/a_27_47# clknet_2_1__leaf_clk 0.243f
C9940 clkbuf_0_clk/a_110_47# _070_ 0.00201f
C9941 _067_ cal_count\[3\] 0.0363f
C9942 _341_/a_543_47# _065_ 0.00413f
C9943 output32/a_27_47# trim[1] 0.343f
C9944 _000_ rebuffer6/a_27_47# 2.8e-20
C9945 _015_ _243_/a_27_297# 0.113f
C9946 _251_/a_109_297# _101_ 0.0603f
C9947 _074_ _140_/a_68_297# 1.04e-20
C9948 _042_ _101_ 0.0277f
C9949 _107_ _262_/a_465_47# 3.06e-19
C9950 _299_/a_215_297# net40 0.00375f
C9951 _249_/a_109_297# net26 6.35e-20
C9952 _232_/a_114_297# _090_ 0.0179f
C9953 trim_mask\[2\] trim_val\[1\] 1.73e-20
C9954 _328_/a_1283_21# trim_mask\[1\] 0.0871f
C9955 mask\[7\] mask\[6\] 0.224f
C9956 _200_/a_303_47# cal_itt\[0\] 3.38e-19
C9957 _200_/a_80_21# _071_ 0.0776f
C9958 clknet_2_1__leaf_clk _016_ 0.0775f
C9959 net9 _340_/a_956_413# 3.42e-19
C9960 VPWR _246_/a_27_297# 0.217f
C9961 _319_/a_761_289# _016_ 3.37e-19
C9962 _328_/a_193_47# _336_/a_1108_47# 2.05e-20
C9963 trim_mask\[2\] _336_/a_193_47# 6.73e-20
C9964 _024_ _264_/a_27_297# 2.56e-20
C9965 _190_/a_27_47# _203_/a_59_75# 0.0134f
C9966 _334_/a_27_47# _334_/a_651_413# 9.73e-19
C9967 _334_/a_761_289# _334_/a_1108_47# 0.0512f
C9968 _334_/a_193_47# _334_/a_448_47# 0.0642f
C9969 _314_/a_193_47# _314_/a_651_413# 0.0346f
C9970 _314_/a_543_47# _314_/a_1108_47# 7.99e-20
C9971 _296_/a_113_47# cal_count\[2\] 2.23e-20
C9972 _228_/a_297_47# _088_ 0.0482f
C9973 _228_/a_382_297# _052_ 0.00165f
C9974 _339_/a_381_47# cal_count\[0\] 0.0167f
C9975 _327_/a_193_47# _327_/a_761_289# 0.186f
C9976 _327_/a_27_47# _327_/a_543_47# 0.115f
C9977 _307_/a_651_413# net45 0.0122f
C9978 trim[3] _334_/a_1270_413# 1.63e-20
C9979 _168_/a_207_413# _331_/a_27_47# 1.17e-19
C9980 _051_ _106_ 5.03e-19
C9981 net2 _339_/a_1182_261# 3.73e-21
C9982 _308_/a_27_47# _319_/a_193_47# 1.77e-21
C9983 _308_/a_193_47# _319_/a_27_47# 8.25e-20
C9984 _111_ _109_ 9.95e-19
C9985 _306_/a_27_47# _208_/a_76_199# 1.43e-20
C9986 _060_ _062_ 0.0644f
C9987 _299_/a_27_413# _299_/a_298_297# 0.00498f
C9988 _304_/a_27_47# _298_/a_78_199# 6.77e-20
C9989 _038_ _067_ 3.04e-20
C9990 mask\[4\] net26 0.718f
C9991 net43 net30 0.156f
C9992 net36 net37 0.00645f
C9993 _327_/a_761_289# _058_ 0.0126f
C9994 _259_/a_27_297# trim_mask\[4\] 0.0667f
C9995 output36/a_27_47# net38 0.0398f
C9996 _320_/a_193_47# _319_/a_1108_47# 9.6e-21
C9997 _237_/a_505_21# clkbuf_2_0__f_clk/a_110_47# 0.00244f
C9998 clone1/a_27_47# _242_/a_382_297# 2.88e-19
C9999 _304_/a_448_47# _122_ 0.0014f
C10000 net33 _175_/a_68_297# 0.0158f
C10001 en output41/a_27_47# 0.00805f
C10002 _104_ trim_mask\[2\] 0.553f
C10003 _333_/a_193_47# net33 1.54e-19
C10004 _325_/a_1283_21# net27 6.09e-20
C10005 trim_mask\[1\] _175_/a_68_297# 1.33e-19
C10006 mask\[6\] _312_/a_27_47# 5.53e-20
C10007 trim_mask\[1\] _333_/a_193_47# 0.00414f
C10008 net49 _333_/a_27_47# 0.0136f
C10009 trim_val\[1\] _333_/a_761_289# 9.6e-19
C10010 _273_/a_59_75# trim_val\[2\] 6.49e-19
C10011 _298_/a_78_199# _298_/a_292_297# 0.013f
C10012 _334_/a_1108_47# rebuffer1/a_75_212# 3.8e-20
C10013 _316_/a_1108_47# _013_ 4.03e-21
C10014 _329_/a_1283_21# _274_/a_75_212# 0.0112f
C10015 net42 _260_/a_93_21# 5.04e-19
C10016 VPWR _084_ 0.346f
C10017 _323_/a_651_413# _042_ 0.0262f
C10018 _192_/a_639_47# _095_ 1.24e-19
C10019 _054_ _118_ 8.99e-21
C10020 trim_mask\[0\] _255_/a_27_47# 0.0762f
C10021 _159_/a_27_47# _313_/a_193_47# 6.61e-20
C10022 _335_/a_193_47# _335_/a_761_289# 0.186f
C10023 _335_/a_27_47# _335_/a_543_47# 0.113f
C10024 _308_/a_1462_47# net45 5.4e-19
C10025 _326_/a_1462_47# net43 0.00288f
C10026 net30 _118_ 0.222f
C10027 _273_/a_59_75# net16 3.67e-19
C10028 clkbuf_2_2__f_clk/a_110_47# clknet_0_clk 0.326f
C10029 _122_ _133_ 0.11f
C10030 _084_ net53 6.92e-21
C10031 mask\[1\] _039_ 1.8e-20
C10032 state\[2\] _100_ 0.00152f
C10033 net31 _296_/a_113_47# 1.37e-19
C10034 _048_ _170_/a_81_21# 2.47e-19
C10035 _283_/a_75_212# clknet_2_0__leaf_clk 0.0101f
C10036 _022_ _101_ 0.0144f
C10037 VPWR _236_/a_109_297# 0.0042f
C10038 _303_/a_193_47# _065_ 1.73e-20
C10039 net10 trim_val\[3\] 5.28e-22
C10040 _309_/a_1283_21# net45 1.36e-20
C10041 _058_ _332_/a_193_47# 0.00777f
C10042 net43 _072_ 0.0964f
C10043 trim_mask\[0\] _270_/a_59_75# 2.23e-19
C10044 _334_/a_639_47# net46 0.00418f
C10045 net15 mask\[2\] 0.291f
C10046 trim_mask\[1\] trim_mask\[4\] 0.0742f
C10047 net25 _310_/a_1270_413# 2.35e-19
C10048 clknet_2_3__leaf_clk clkc 1.48e-19
C10049 VPWR _057_ 1.86f
C10050 VPWR _208_/a_535_374# 7.28e-19
C10051 _315_/a_1283_21# _095_ 8.55e-19
C10052 net55 _242_/a_297_47# 2.28e-19
C10053 _327_/a_651_413# net46 0.0133f
C10054 net27 _314_/a_27_47# 0.00152f
C10055 _020_ net26 3.23e-19
C10056 _299_/a_27_413# _133_ 3.3e-19
C10057 _336_/a_448_47# _028_ 4.1e-20
C10058 _336_/a_761_289# trim_mask\[4\] 0.0221f
C10059 cal_itt\[2\] _068_ 0.0725f
C10060 trim_mask\[2\] _114_ 0.154f
C10061 _287_/a_75_212# net18 2.08e-19
C10062 net9 _037_ 0.11f
C10063 _329_/a_1283_21# clknet_2_2__leaf_clk 0.0163f
C10064 _304_/a_543_47# _304_/a_651_413# 0.0572f
C10065 _304_/a_761_289# _304_/a_1270_413# 2.6e-19
C10066 _304_/a_193_47# _304_/a_639_47# 2.28e-19
C10067 clkbuf_2_0__f_clk/a_110_47# _241_/a_297_47# 1.08e-19
C10068 _339_/a_1182_261# _123_ 0.0138f
C10069 _009_ _084_ 0.189f
C10070 _048_ _227_/a_296_53# 1.17e-19
C10071 net43 _305_/a_193_47# 0.639f
C10072 _334_/a_193_47# _031_ 0.222f
C10073 _329_/a_639_47# trim_mask\[2\] 1.57e-19
C10074 trim_mask\[4\] clone1/a_27_47# 9.23e-21
C10075 _026_ _258_/a_109_297# 0.00169f
C10076 _332_/a_1108_47# net37 4.63e-20
C10077 _066_ net19 8.99e-21
C10078 _332_/a_27_47# _332_/a_193_47# 0.685f
C10079 input1/a_75_212# cal 0.196f
C10080 _336_/a_639_47# net19 7.16e-19
C10081 _335_/a_651_413# net46 0.0168f
C10082 _322_/a_651_413# _074_ 0.00182f
C10083 _093_ _099_ 0.0555f
C10084 calibrate _092_ 0.0617f
C10085 VPWR _226_/a_109_47# 1.4e-19
C10086 _305_/a_1108_47# _190_/a_27_47# 4.06e-20
C10087 _235_/a_297_47# net3 0.0409f
C10088 net3 _317_/a_193_47# 8.87e-20
C10089 _306_/a_543_47# _076_ 0.00105f
C10090 output33/a_27_47# _175_/a_68_297# 0.001f
C10091 _304_/a_761_289# clknet_2_3__leaf_clk 0.00101f
C10092 mask\[3\] _247_/a_109_297# 0.0583f
C10093 _293_/a_81_21# net2 5.27e-19
C10094 _309_/a_761_289# clknet_2_1__leaf_clk 9.01e-21
C10095 _218_/a_113_297# _074_ 1.16e-20
C10096 net45 _092_ 0.00188f
C10097 _294_/a_68_297# net33 0.00445f
C10098 net4 clone7/a_27_47# 2.18e-20
C10099 VPWR _330_/a_448_47# 0.0851f
C10100 _332_/a_448_47# net46 0.0165f
C10101 _237_/a_76_199# _096_ 0.318f
C10102 _306_/a_1283_21# _050_ 5.67e-21
C10103 _333_/a_1462_47# net33 7.82e-19
C10104 _325_/a_27_47# net26 9.87e-21
C10105 _336_/a_639_47# _107_ 2.69e-19
C10106 VPWR _085_ 0.278f
C10107 _340_/a_956_413# _122_ 3.06e-19
C10108 net13 _319_/a_1108_47# 3.56e-36
C10109 net49 _333_/a_1217_47# 1.84e-19
C10110 _337_/a_543_47# clknet_0_clk 1.84e-19
C10111 _115_ _114_ 0.142f
C10112 clknet_2_1__leaf_clk _040_ 0.00956f
C10113 _112_ _109_ 0.00155f
C10114 _310_/a_761_289# _310_/a_639_47# 3.16e-19
C10115 _310_/a_27_47# _310_/a_1217_47# 2.56e-19
C10116 _324_/a_193_47# _042_ 8.79e-20
C10117 _340_/a_193_47# net18 1.81e-20
C10118 _314_/a_543_47# _224_/a_113_297# 9.8e-19
C10119 clknet_2_3__leaf_clk _298_/a_215_47# 1.91e-20
C10120 _110_ clkbuf_2_2__f_clk/a_110_47# 0.0083f
C10121 _307_/a_27_47# net22 0.175f
C10122 clkbuf_2_3__f_clk/a_110_47# clknet_2_3__leaf_clk 1.62f
C10123 VPWR _325_/a_651_413# 0.144f
C10124 _050_ _170_/a_299_297# 0.00539f
C10125 _327_/a_805_47# _108_ 1.45e-19
C10126 VPWR _216_/a_199_47# 1.28e-19
C10127 _065_ _092_ 0.0108f
C10128 output35/a_27_47# net35 0.265f
C10129 net21 _313_/a_448_47# 5.49e-20
C10130 _046_ _313_/a_1270_413# 7.93e-21
C10131 _324_/a_1108_47# clknet_2_1__leaf_clk 0.00114f
C10132 _340_/a_193_47# _129_ 0.00163f
C10133 _228_/a_79_21# net41 9.74e-20
C10134 output22/a_27_47# output24/a_27_47# 9.71e-21
C10135 clk _073_ 0.00414f
C10136 input2/a_27_47# comp 0.233f
C10137 _311_/a_193_47# _311_/a_543_47# 0.217f
C10138 _311_/a_27_47# _311_/a_1283_21# 0.0436f
C10139 _105_ _092_ 2.75e-20
C10140 _042_ _248_/a_27_297# 5.2e-19
C10141 _322_/a_27_47# _042_ 4.43e-19
C10142 en_co_clk _192_/a_174_21# 0.0229f
C10143 _304_/a_193_47# _136_ 0.00208f
C10144 _064_ _257_/a_27_297# 0.109f
C10145 cal_itt\[2\] _306_/a_27_47# 2.48e-21
C10146 _322_/a_1283_21# clknet_2_1__leaf_clk 5.83e-20
C10147 trim[4] net37 0.00207f
C10148 _033_ _028_ 7.86e-20
C10149 _141_/a_27_47# net51 3.52e-20
C10150 _227_/a_109_93# _062_ 6.61e-21
C10151 result[1] net43 1.33e-19
C10152 mask\[1\] net15 0.00484f
C10153 _304_/a_543_47# net47 0.153f
C10154 _326_/a_27_47# _314_/a_27_47# 0.002f
C10155 net43 _305_/a_1462_47# 0.00288f
C10156 net43 _251_/a_27_297# 1.31e-19
C10157 net43 _250_/a_109_47# 1.33e-20
C10158 VPWR _314_/a_543_47# 0.209f
C10159 _187_/a_212_413# en_co_clk 0.195f
C10160 _308_/a_1283_21# mask\[0\] 0.0103f
C10161 _308_/a_543_47# _078_ 0.00147f
C10162 _332_/a_639_47# _108_ 0.00129f
C10163 _321_/a_543_47# _321_/a_651_413# 0.0572f
C10164 _321_/a_761_289# _321_/a_1270_413# 2.6e-19
C10165 _321_/a_193_47# _321_/a_639_47# 2.28e-19
C10166 _340_/a_27_47# _340_/a_1032_413# 0.178f
C10167 _340_/a_193_47# _340_/a_1182_261# 0.0728f
C10168 _340_/a_652_21# _340_/a_476_47# 0.26f
C10169 _332_/a_543_47# _332_/a_639_47# 0.0138f
C10170 _332_/a_193_47# _332_/a_1217_47# 2.36e-20
C10171 _332_/a_761_289# _332_/a_805_47# 3.69e-19
C10172 _308_/a_27_47# net24 8.97e-21
C10173 _136_ _298_/a_493_297# 1.66e-20
C10174 _302_/a_109_297# clknet_2_3__leaf_clk 7.57e-20
C10175 VPWR rebuffer4/a_27_47# 0.261f
C10176 output14/a_27_47# _314_/a_651_413# 1.74e-19
C10177 ctlp[0] _314_/a_193_47# 0.00268f
C10178 net23 clknet_2_1__leaf_clk 0.00695f
C10179 _168_/a_297_47# trim_mask\[4\] 3.87e-19
C10180 net43 _319_/a_1108_47# 0.219f
C10181 _198_/a_27_47# clknet_0_clk 1.31e-19
C10182 ctln[1] clk 0.00132f
C10183 _199_/a_109_297# _065_ 0.00221f
C10184 _117_ net18 8.86e-19
C10185 _169_/a_215_311# net41 3.77e-20
C10186 _050_ _192_/a_174_21# 0.00179f
C10187 _337_/a_543_47# _337_/a_651_413# 0.0572f
C10188 _337_/a_761_289# _337_/a_1270_413# 2.6e-19
C10189 _337_/a_193_47# _337_/a_639_47# 2.28e-19
C10190 clknet_0_clk _331_/a_193_47# 0.00248f
C10191 _162_/a_27_47# _047_ 0.191f
C10192 mask\[3\] _018_ 0.163f
C10193 _288_/a_59_75# _125_ 0.122f
C10194 _126_ _339_/a_1032_413# 1.28e-21
C10195 _319_/a_1283_21# _034_ 1.22e-20
C10196 _340_/a_27_47# cal_count\[3\] 1.3e-20
C10197 _316_/a_1283_21# _090_ 9.09e-20
C10198 VPWR net36 0.383f
C10199 net39 net16 0.0166f
C10200 net9 _339_/a_562_413# 4.34e-19
C10201 output10/a_27_47# net46 1.46e-20
C10202 _340_/a_1032_413# clknet_2_3__leaf_clk 9.51e-21
C10203 _136_ net18 0.0321f
C10204 trim_mask\[3\] fanout46/a_27_47# 0.0016f
C10205 VPWR _027_ 0.706f
C10206 _110_ _162_/a_27_47# 9.22e-20
C10207 net47 _035_ 0.144f
C10208 net28 mask\[6\] 0.365f
C10209 _287_/a_75_212# _338_/a_652_21# 7.07e-19
C10210 _078_ _140_/a_150_297# 1.95e-19
C10211 _063_ _073_ 1.41e-19
C10212 net25 net26 0.00158f
C10213 _015_ _316_/a_1108_47# 3.41e-20
C10214 _270_/a_59_75# _265_/a_81_21# 0.00111f
C10215 _276_/a_59_75# _117_ 0.114f
C10216 VPWR _195_/a_218_47# 8.79e-20
C10217 _037_ _122_ 0.00898f
C10218 _097_ _237_/a_218_47# 2.88e-19
C10219 _301_/a_377_297# clkc 7.52e-20
C10220 _064_ trim_val\[4\] 0.0378f
C10221 _303_/a_1283_21# _067_ 2.4e-21
C10222 _324_/a_448_47# mask\[6\] 2.48e-21
C10223 _303_/a_1283_21# _070_ 2.2e-20
C10224 ctln[1] net4 0.0343f
C10225 _324_/a_543_47# _021_ 5.07e-19
C10226 _321_/a_1283_21# _143_/a_68_297# 0.00127f
C10227 _239_/a_474_297# _095_ 2.97e-20
C10228 _239_/a_27_297# _092_ 0.0722f
C10229 VPWR _334_/a_1270_413# 7.7e-19
C10230 mask\[6\] _158_/a_68_297# 6.03e-19
C10231 _326_/a_1283_21# net25 2.65e-21
C10232 net8 trim_mask\[2\] 0.0279f
C10233 net14 _138_/a_27_47# 0.113f
C10234 clkbuf_0_clk/a_110_47# clknet_2_3__leaf_clk 5.7e-20
C10235 clknet_2_0__leaf_clk rebuffer5/a_161_47# 0.005f
C10236 cal_count\[3\] clknet_2_3__leaf_clk 0.519f
C10237 _307_/a_1217_47# net22 1.27e-19
C10238 VPWR _327_/a_448_47# 0.0851f
C10239 _189_/a_27_47# _048_ 0.0893f
C10240 _185_/a_68_297# _049_ 3.65e-19
C10241 _302_/a_27_297# _136_ 0.0986f
C10242 _037_ _299_/a_27_413# 5.48e-21
C10243 output37/a_27_47# net34 0.0167f
C10244 _307_/a_27_47# _079_ 2.27e-19
C10245 _062_ _054_ 1.53e-22
C10246 _119_ net18 1.51e-19
C10247 _062_ net30 0.148f
C10248 _311_/a_448_47# _311_/a_639_47# 4.61e-19
C10249 fanout44/a_27_47# net30 1.5e-19
C10250 ctln[4] _335_/a_193_47# 3.05e-19
C10251 _041_ clknet_0_clk 2.41e-20
C10252 output19/a_27_47# ctlp[5] 0.168f
C10253 VPWR _335_/a_448_47# 0.1f
C10254 net2 en_co_clk 0.09f
C10255 fanout46/a_27_47# _330_/a_1283_21# 0.00774f
C10256 trim[4] _332_/a_651_413# 1.32e-19
C10257 VPWR _311_/a_193_47# 0.287f
C10258 _304_/a_1283_21# _063_ 0.00322f
C10259 _000_ _042_ 1.3e-20
C10260 _276_/a_59_75# _119_ 6.99e-22
C10261 _341_/a_193_47# _304_/a_761_289# 1.36e-20
C10262 _341_/a_27_47# _304_/a_543_47# 8.14e-19
C10263 _018_ _310_/a_1283_21# 3.75e-19
C10264 _256_/a_373_47# _024_ 1.97e-19
C10265 _340_/a_1602_47# net47 0.00218f
C10266 _037_ _304_/a_1283_21# 1.58e-20
C10267 _293_/a_299_297# _127_ 2.03e-20
C10268 _091_ net4 0.0128f
C10269 _195_/a_76_199# net30 8.82e-21
C10270 _083_ clknet_2_1__leaf_clk 0.0112f
C10271 _065_ _208_/a_218_47# 0.00117f
C10272 _264_/a_27_297# trim_val\[4\] 3.83e-19
C10273 _311_/a_193_47# net53 0.0181f
C10274 _266_/a_68_297# clkbuf_2_3__f_clk/a_110_47# 9.54e-19
C10275 VPWR _332_/a_1108_47# 0.292f
C10276 clkbuf_2_1__f_clk/a_110_47# _120_ 4.98e-20
C10277 _340_/a_652_21# _340_/a_1224_47# 1.57e-19
C10278 _088_ _049_ 0.0514f
C10279 _260_/a_93_21# _098_ 2.07e-21
C10280 net8 _115_ 2.98e-19
C10281 _038_ clknet_2_3__leaf_clk 0.0816f
C10282 _017_ _065_ 6.2e-21
C10283 net26 _310_/a_543_47# 2.08e-19
C10284 _149_/a_68_297# net19 0.013f
C10285 _281_/a_103_199# _096_ 2.67e-20
C10286 _291_/a_285_297# net33 0.00361f
C10287 _309_/a_448_47# _078_ 3.69e-19
C10288 _215_/a_109_297# net14 0.00101f
C10289 _323_/a_27_47# _043_ 3.7e-19
C10290 _323_/a_193_47# net18 6.64e-20
C10291 _053_ net41 8.1e-20
C10292 _134_ net34 1.5e-20
C10293 _309_/a_543_47# net24 0.0302f
C10294 _337_/a_543_47# net44 0.153f
C10295 net5 _134_ 0.00203f
C10296 clkbuf_2_2__f_clk/a_110_47# clknet_2_2__leaf_clk 1.71f
C10297 _338_/a_476_47# clknet_2_3__leaf_clk 0.0467f
C10298 _062_ _072_ 5.18e-20
C10299 VPWR _310_/a_805_47# 4.15e-19
C10300 _336_/a_27_47# _330_/a_27_47# 4.35e-20
C10301 _233_/a_27_297# input1/a_75_212# 3.78e-19
C10302 _181_/a_68_297# fanout46/a_27_47# 0.00121f
C10303 net30 _137_/a_68_297# 0.00208f
C10304 net47 _198_/a_27_47# 1.02e-19
C10305 net43 _313_/a_543_47# 0.159f
C10306 _133_ _297_/a_285_47# 0.0439f
C10307 trim_mask\[0\] _136_ 0.00162f
C10308 comp trimb[4] 0.0482f
C10309 net34 _333_/a_1283_21# 0.00138f
C10310 _078_ _249_/a_27_297# 9.33e-19
C10311 _333_/a_448_47# _055_ 8.27e-22
C10312 _035_ _338_/a_562_413# 3.7e-19
C10313 _293_/a_299_297# _126_ 0.0549f
C10314 _232_/a_32_297# en_co_clk 0.00613f
C10315 _091_ _063_ 0.0171f
C10316 _161_/a_68_297# _332_/a_1108_47# 5.3e-19
C10317 _189_/a_218_47# _050_ 0.0867f
C10318 _306_/a_1108_47# net51 1.37e-21
C10319 _321_/a_448_47# _101_ 0.0198f
C10320 trim[1] _265_/a_299_297# 7.76e-20
C10321 _338_/a_1140_413# net18 3.91e-19
C10322 clkbuf_2_2__f_clk/a_110_47# net11 2.35e-20
C10323 _134_ _299_/a_298_297# 4.26e-21
C10324 result[1] _080_ 8.38e-19
C10325 _306_/a_193_47# rebuffer6/a_27_47# 3.16e-21
C10326 _108_ _049_ 2.47e-20
C10327 cal_itt\[2\] cal_itt\[3\] 0.00647f
C10328 output12/a_27_47# net12 0.24f
C10329 _337_/a_193_47# _263_/a_297_47# 1.46e-20
C10330 cal_itt\[0\] _124_ 7.19e-19
C10331 net15 _247_/a_109_47# 9.36e-19
C10332 _123_ en_co_clk 5.23e-20
C10333 _304_/a_1108_47# net19 1.83e-21
C10334 VPWR output17/a_27_47# 0.301f
C10335 _244_/a_27_297# _049_ 7.59e-19
C10336 clk _331_/a_761_289# 0.00262f
C10337 _053_ _171_/a_27_47# 0.0358f
C10338 _307_/a_639_47# _004_ 2.31e-19
C10339 trim_mask\[0\] _119_ 0.0387f
C10340 _314_/a_27_47# _011_ 0.167f
C10341 _314_/a_761_289# _086_ 1.62e-19
C10342 net12 _331_/a_193_47# 1.35e-19
C10343 _311_/a_1108_47# net26 0.0587f
C10344 net28 _313_/a_805_47# 0.0021f
C10345 _322_/a_1270_413# _078_ 1.91e-19
C10346 _064_ _330_/a_193_47# 2.68e-21
C10347 _306_/a_27_47# _306_/a_543_47# 0.115f
C10348 _306_/a_193_47# _306_/a_761_289# 0.186f
C10349 cal_itt\[2\] _305_/a_27_47# 0.00131f
C10350 clk rstn 0.0354f
C10351 _048_ _096_ 0.0551f
C10352 ctlp[7] _078_ 5.41e-19
C10353 cal_itt\[2\] _262_/a_205_47# 3.12e-20
C10354 VPWR _032_ 0.398f
C10355 _326_/a_543_47# net27 5.3e-20
C10356 _326_/a_193_47# result[5] 7.03e-19
C10357 _331_/a_27_47# _331_/a_448_47# 0.0902f
C10358 _331_/a_193_47# _331_/a_1108_47# 0.125f
C10359 VPWR trim[4] 0.585f
C10360 net42 _048_ 0.454f
C10361 _217_/a_109_297# clknet_2_1__leaf_clk 8.92e-19
C10362 VPWR _311_/a_1462_47# 7.21e-20
C10363 net4 _198_/a_109_47# 1.92e-19
C10364 _050_ _232_/a_32_297# 6.01e-21
C10365 _111_ net46 0.00637f
C10366 mask\[6\] _084_ 0.0364f
C10367 _325_/a_1108_47# _250_/a_27_297# 8.86e-20
C10368 _143_/a_68_297# _101_ 1.1e-20
C10369 _321_/a_1108_47# _320_/a_193_47# 4.8e-21
C10370 _256_/a_27_297# clknet_2_2__leaf_clk 0.0116f
C10371 _078_ _220_/a_113_297# 0.0637f
C10372 net13 _003_ 1.12e-20
C10373 _143_/a_150_297# _041_ 4.96e-19
C10374 net47 _041_ 0.611f
C10375 net47 _338_/a_1182_261# 0.143f
C10376 _338_/a_27_47# _338_/a_193_47# 0.55f
C10377 _258_/a_27_297# _258_/a_109_47# 0.00393f
C10378 _050_ _336_/a_193_47# 9.32e-20
C10379 cal _315_/a_27_47# 0.00255f
C10380 _266_/a_68_297# cal_count\[3\] 8.9e-19
C10381 _325_/a_448_47# clknet_2_1__leaf_clk 0.00239f
C10382 _253_/a_384_47# net52 8.16e-20
C10383 _074_ _310_/a_193_47# 0.015f
C10384 _339_/a_27_47# _129_ 4.2e-20
C10385 _185_/a_68_297# state\[1\] 2.14e-19
C10386 trim_mask\[0\] _087_ 3.44e-21
C10387 net47 _297_/a_129_47# 2.49e-20
C10388 mask\[3\] clkbuf_2_1__f_clk/a_110_47# 8.09e-21
C10389 trim[0] trim[2] 0.0391f
C10390 rstn net4 0.00313f
C10391 _340_/a_381_47# _037_ 0.149f
C10392 VPWR net41 0.501f
C10393 en_co_clk net55 0.0459f
C10394 _102_ _023_ 2.21e-19
C10395 _134_ _133_ 0.00631f
C10396 trim_val\[3\] net9 4.6e-19
C10397 _301_/a_377_297# cal_count\[3\] 6.02e-20
C10398 _051_ _089_ 0.00231f
C10399 _341_/a_193_47# cal_count\[3\] 0.547f
C10400 net12 _041_ 0.00956f
C10401 trim[4] _161_/a_68_297# 0.00111f
C10402 output14/a_27_47# ctlp[0] 0.338f
C10403 _338_/a_1224_47# clknet_2_3__leaf_clk 1.82e-19
C10404 input2/a_27_47# _132_ 0.00127f
C10405 _341_/a_448_47# clknet_2_3__leaf_clk 0.016f
C10406 net41 valid 0.0214f
C10407 net46 rebuffer3/a_75_212# 8.12e-20
C10408 state\[0\] _192_/a_476_47# 3.57e-20
C10409 _320_/a_27_47# _143_/a_68_297# 8.61e-19
C10410 clkbuf_2_2__f_clk/a_110_47# _279_/a_204_297# 6.65e-21
C10411 VPWR _306_/a_448_47# 0.0849f
C10412 trim_mask\[1\] _334_/a_27_47# 1.41e-20
C10413 trim_val\[1\] _334_/a_193_47# 5.84e-22
C10414 _026_ _025_ 0.00206f
C10415 net34 cal_count\[2\] 7.97e-20
C10416 _340_/a_193_47# _339_/a_476_47# 5.41e-19
C10417 _340_/a_1182_261# _339_/a_27_47# 2.07e-19
C10418 _340_/a_476_47# _339_/a_193_47# 3.29e-21
C10419 _168_/a_27_413# _048_ 3.58e-20
C10420 _104_ _050_ 0.0258f
C10421 _307_/a_193_47# net14 0.0105f
C10422 clknet_2_1__leaf_clk _314_/a_761_289# 4.07e-20
C10423 cal clknet_2_0__leaf_clk 0.00552f
C10424 output29/a_27_47# _085_ 9.81e-20
C10425 en_co_clk _067_ 0.0436f
C10426 _326_/a_193_47# net29 1.03e-19
C10427 en_co_clk _070_ 4.53e-21
C10428 _065_ net46 0.00145f
C10429 _227_/a_109_93# _227_/a_209_311# 0.168f
C10430 net21 net20 0.00154f
C10431 fanout46/a_27_47# _108_ 1.48e-20
C10432 _135_ net46 6e-20
C10433 _041_ net44 0.0236f
C10434 _029_ _332_/a_1108_47# 5.34e-21
C10435 output34/a_27_47# trim_val\[2\] 0.0717f
C10436 VPWR _171_/a_27_47# 0.344f
C10437 _050_ net55 0.128f
C10438 _146_/a_150_297# _310_/a_193_47# 1.9e-20
C10439 net43 _003_ 0.00181f
C10440 fanout44/a_27_47# _319_/a_1108_47# 7.24e-20
C10441 _071_ _065_ 6.44e-20
C10442 _339_/a_1602_47# _133_ 6.44e-21
C10443 _323_/a_448_47# net47 2.46e-19
C10444 _318_/a_27_47# net41 1.75e-20
C10445 _312_/a_1283_21# net20 9.79e-19
C10446 _299_/a_298_297# cal_count\[2\] 3.59e-19
C10447 _259_/a_373_47# _027_ 1.97e-19
C10448 net50 _033_ 2.07e-20
C10449 _162_/a_27_47# trim_val\[0\] 6.71e-21
C10450 mask\[6\] _085_ 0.104f
C10451 cal_itt\[2\] _305_/a_1217_47# 1.19e-20
C10452 net15 net26 0.0071f
C10453 _078_ _222_/a_113_297# 0.05f
C10454 _118_ net40 0.129f
C10455 _341_/a_193_47# _038_ 0.207f
C10456 _341_/a_1108_47# _136_ 0.00705f
C10457 clkbuf_2_3__f_clk/a_110_47# _279_/a_314_297# 2.66e-21
C10458 _331_/a_27_47# _028_ 0.458f
C10459 _331_/a_193_47# clknet_2_2__leaf_clk 0.00247f
C10460 net7 _317_/a_761_289# 4.61e-20
C10461 state\[0\] calibrate 0.00673f
C10462 _280_/a_75_212# net19 1.78e-22
C10463 _326_/a_1283_21# net15 9.71e-21
C10464 _101_ net52 0.874f
C10465 _317_/a_193_47# _317_/a_761_289# 0.181f
C10466 _317_/a_27_47# _317_/a_543_47# 0.115f
C10467 _325_/a_761_289# _022_ 7.67e-19
C10468 output26/a_27_47# clknet_2_1__leaf_clk 0.0227f
C10469 _326_/a_27_47# _326_/a_543_47# 0.115f
C10470 _326_/a_193_47# _326_/a_761_289# 0.186f
C10471 state\[2\] clk 0.0574f
C10472 net49 net37 1.62e-19
C10473 VPWR _094_ 0.382f
C10474 net22 _120_ 0.00171f
C10475 output12/a_27_47# net11 0.00102f
C10476 _104_ _228_/a_297_47# 0.03f
C10477 _269_/a_299_297# _108_ 9.71e-20
C10478 net47 _338_/a_1296_47# 0.0028f
C10479 _136_ _265_/a_81_21# 8.24e-20
C10480 _338_/a_193_47# _338_/a_586_47# 0.00127f
C10481 VPWR _317_/a_448_47# 0.0794f
C10482 _078_ rebuffer5/a_161_47# 5.39e-19
C10483 _328_/a_27_47# trim_mask\[2\] 3.93e-19
C10484 VPWR _326_/a_448_47# 0.0859f
C10485 _328_/a_761_289# _328_/a_543_47# 0.21f
C10486 _328_/a_193_47# _328_/a_1283_21# 0.0424f
C10487 _328_/a_27_47# _328_/a_1108_47# 0.102f
C10488 _328_/a_1462_47# trim_mask\[0\] 8.3e-20
C10489 net13 _321_/a_1108_47# 0.00106f
C10490 _290_/a_207_413# net37 0.0104f
C10491 state\[0\] net45 0.00525f
C10492 clknet_2_0__leaf_clk net51 0.0639f
C10493 _066_ _062_ 0.0114f
C10494 _087_ _090_ 0.0952f
C10495 state\[2\] _331_/a_1283_21# 6.97e-19
C10496 net13 _337_/a_1108_47# 0.00163f
C10497 _214_/a_199_47# _101_ 3.77e-19
C10498 _170_/a_299_297# _049_ 0.0588f
C10499 VPWR _203_/a_145_75# 1.48e-19
C10500 net13 _167_/a_161_47# 1.79e-19
C10501 net31 net34 0.966f
C10502 trim[0] _055_ 0.0624f
C10503 VPWR _286_/a_439_47# 6.47e-20
C10504 net31 net5 0.0416f
C10505 _064_ _058_ 0.12f
C10506 state\[2\] net4 0.325f
C10507 _325_/a_543_47# _313_/a_543_47# 0.00153f
C10508 VPWR _192_/a_505_280# 0.234f
C10509 _064_ _335_/a_193_47# 5e-19
C10510 fanout43/a_27_47# clkbuf_2_1__f_clk/a_110_47# 1.43e-20
C10511 _272_/a_299_297# net46 0.00102f
C10512 _112_ net46 0.00936f
C10513 net44 _312_/a_1108_47# 0.247f
C10514 _312_/a_193_47# _312_/a_761_289# 0.186f
C10515 _312_/a_27_47# _312_/a_543_47# 0.115f
C10516 clknet_2_1__leaf_clk _141_/a_27_47# 4.73e-19
C10517 _168_/a_207_413# _050_ 0.0617f
C10518 _033_ _330_/a_1108_47# 5.66e-20
C10519 _336_/a_1108_47# _027_ 1.01e-21
C10520 _336_/a_1283_21# net46 0.319f
C10521 state\[0\] _065_ 2.46e-21
C10522 _320_/a_27_47# net52 0.00489f
C10523 _227_/a_368_53# _049_ 2.88e-19
C10524 _227_/a_209_311# _054_ 5.12e-20
C10525 clknet_2_1__leaf_clk _311_/a_27_47# 0.266f
C10526 _323_/a_448_47# net44 0.00175f
C10527 _329_/a_193_47# net46 0.0283f
C10528 _303_/a_1283_21# clknet_2_3__leaf_clk 0.0739f
C10529 _227_/a_209_311# net30 1.72e-20
C10530 _133_ cal_count\[2\] 0.308f
C10531 _212_/a_113_297# _078_ 0.0661f
C10532 _050_ mask\[0\] 9.79e-21
C10533 net47 _339_/a_1032_413# 0.216f
C10534 _321_/a_1108_47# _248_/a_109_297# 2.52e-19
C10535 _114_ _334_/a_193_47# 5.54e-20
C10536 _323_/a_761_289# _323_/a_543_47# 0.21f
C10537 _323_/a_193_47# _323_/a_1283_21# 0.0424f
C10538 _323_/a_27_47# _323_/a_1108_47# 0.102f
C10539 trim_val\[2\] _334_/a_1283_21# 0.0646f
C10540 _336_/a_448_47# _052_ 1.24e-20
C10541 VPWR _315_/a_193_47# 0.452f
C10542 _306_/a_761_289# _072_ 1.19e-19
C10543 _306_/a_543_47# cal_itt\[3\] 3.33e-19
C10544 _263_/a_297_47# _090_ 1.29e-19
C10545 _107_ _229_/a_27_297# 7.58e-19
C10546 _284_/a_150_297# en_co_clk 8.78e-19
C10547 _337_/a_193_47# _099_ 7.41e-21
C10548 _337_/a_27_47# _092_ 0.00189f
C10549 net3 _316_/a_27_47# 1.24e-19
C10550 VPWR _318_/a_639_47# 0.001f
C10551 net16 _334_/a_1283_21# 0.00492f
C10552 _315_/a_193_47# valid 0.00582f
C10553 _119_ trim_mask\[4\] 0.00837f
C10554 _042_ _310_/a_1108_47# 1.99e-19
C10555 _292_/a_78_199# _340_/a_1032_413# 6.61e-19
C10556 _239_/a_474_297# _052_ 1.88e-19
C10557 state\[0\] _243_/a_109_297# 1.27e-19
C10558 net54 _096_ 0.376f
C10559 _060_ _100_ 0.312f
C10560 _306_/a_543_47# _305_/a_27_47# 0.00347f
C10561 net43 _321_/a_1108_47# 0.252f
C10562 output9/a_27_47# net46 1.71e-19
C10563 comp net33 3.24e-19
C10564 clknet_2_1__leaf_clk _310_/a_639_47# 9.94e-19
C10565 _058_ _264_/a_27_297# 0.0014f
C10566 net2 output40/a_27_47# 0.0013f
C10567 output12/a_27_47# ctln[7] 4.45e-20
C10568 ctln[6] output13/a_27_47# 1.71e-19
C10569 _192_/a_174_21# _049_ 0.00495f
C10570 _320_/a_27_47# _320_/a_761_289# 0.0701f
C10571 _293_/a_81_21# _144_/a_27_47# 0.0184f
C10572 _336_/a_1108_47# _335_/a_448_47# 3.67e-21
C10573 VPWR _074_ 3.7f
C10574 _341_/a_1462_47# _038_ 3.39e-20
C10575 _331_/a_1217_47# _028_ 1.84e-19
C10576 _331_/a_1462_47# clknet_2_2__leaf_clk 3.64e-20
C10577 clknet_2_2__leaf_clk _260_/a_93_21# 1.05e-20
C10578 _260_/a_93_21# _260_/a_584_47# 0.00278f
C10579 _128_ _133_ 5.69e-19
C10580 _041_ _209_/a_27_47# 3.39e-20
C10581 net9 _334_/a_1108_47# 2.52e-20
C10582 _093_ net41 1.4e-19
C10583 _328_/a_448_47# clknet_2_2__leaf_clk 0.0164f
C10584 _074_ valid 0.0171f
C10585 _337_/a_1283_21# _034_ 7.08e-20
C10586 _074_ net53 0.0143f
C10587 _005_ net14 8.37e-20
C10588 _112_ _332_/a_448_47# 1.93e-19
C10589 VPWR _014_ 1f
C10590 net48 rebuffer1/a_75_212# 0.109f
C10591 _341_/a_193_47# _341_/a_448_47# 0.0564f
C10592 _341_/a_761_289# _341_/a_1108_47# 0.0512f
C10593 _341_/a_27_47# _341_/a_651_413# 9.73e-19
C10594 _328_/a_1283_21# _328_/a_1462_47# 0.0074f
C10595 _328_/a_1108_47# _328_/a_1217_47# 0.00742f
C10596 net12 _324_/a_27_47# 5.32e-19
C10597 _006_ _140_/a_68_297# 4.01e-20
C10598 output24/a_27_47# net25 2.02e-20
C10599 _336_/a_651_413# _108_ 3.38e-20
C10600 _320_/a_805_47# net44 0.0019f
C10601 _341_/a_1270_413# _037_ 8.1e-21
C10602 net47 _303_/a_1108_47# 0.251f
C10603 _010_ _222_/a_199_47# 1.01e-19
C10604 net31 _133_ 1.06e-20
C10605 _309_/a_639_47# net14 0.00144f
C10606 _308_/a_1283_21# _016_ 1.83e-20
C10607 trim_mask\[3\] clkbuf_2_2__f_clk/a_110_47# 1.5e-20
C10608 net16 _332_/a_193_47# 0.0169f
C10609 _318_/a_193_47# _318_/a_1270_413# 1.46e-19
C10610 _318_/a_27_47# _318_/a_639_47# 0.00188f
C10611 _318_/a_543_47# _318_/a_448_47# 0.0498f
C10612 _318_/a_761_289# _318_/a_651_413# 0.0977f
C10613 _318_/a_1283_21# _318_/a_1108_47# 0.234f
C10614 _340_/a_956_413# cal_count\[2\] 1.2e-20
C10615 _074_ _009_ 0.0558f
C10616 mask\[4\] clknet_2_3__leaf_clk 1.27e-19
C10617 clknet_2_1__leaf_clk _247_/a_373_47# 1.25e-19
C10618 _121_ en_co_clk 0.00168f
C10619 _325_/a_27_47# _010_ 5.33e-19
C10620 _104_ _335_/a_805_47# 1.17e-20
C10621 _233_/a_27_297# _315_/a_27_47# 1.81e-19
C10622 VPWR output23/a_27_47# 0.252f
C10623 _309_/a_27_47# _101_ 5.47e-20
C10624 _324_/a_27_47# net44 0.316f
C10625 _286_/a_505_21# cal_count\[0\] 0.258f
C10626 VPWR _305_/a_448_47# 0.0851f
C10627 _329_/a_1462_47# net46 0.00339f
C10628 _308_/a_27_47# _308_/a_543_47# 0.115f
C10629 _308_/a_193_47# _308_/a_761_289# 0.186f
C10630 _048_ _098_ 0.24f
C10631 _323_/a_1270_413# net19 1.39e-19
C10632 trim_mask\[0\] _099_ 8.74e-21
C10633 VPWR _146_/a_150_297# 0.00131f
C10634 _107_ _260_/a_256_47# 2.35e-19
C10635 _192_/a_505_280# _192_/a_548_47# 8.61e-19
C10636 _019_ _321_/a_27_47# 7.83e-21
C10637 _307_/a_27_47# _307_/a_1283_21# 0.0435f
C10638 _307_/a_193_47# _307_/a_543_47# 0.227f
C10639 net9 _332_/a_761_289# 8.16e-20
C10640 _323_/a_1283_21# _323_/a_1462_47# 0.0074f
C10641 _323_/a_1108_47# _323_/a_1217_47# 0.00742f
C10642 result[2] mask\[1\] 0.00154f
C10643 VPWR _259_/a_109_297# 0.197f
C10644 _333_/a_543_47# clknet_2_2__leaf_clk 4.83e-20
C10645 _304_/a_543_47# _001_ 0.0119f
C10646 VPWR _315_/a_1462_47# 4.59e-19
C10647 _293_/a_299_297# net47 2.46e-20
C10648 _329_/a_1283_21# _031_ 0.00166f
C10649 _318_/a_193_47# clknet_2_0__leaf_clk 0.00447f
C10650 output22/a_27_47# result[0] 0.158f
C10651 _048_ clknet_0_clk 0.0719f
C10652 net20 _045_ 0.014f
C10653 _230_/a_145_75# en_co_clk 1.15e-19
C10654 _051_ _092_ 0.0918f
C10655 VPWR _243_/a_27_297# 0.176f
C10656 _078_ _310_/a_761_289# 1.96e-19
C10657 _107_ net19 0.0393f
C10658 cal_count\[1\] _340_/a_1602_47# 0.00724f
C10659 _050_ _121_ 4.53e-21
C10660 clknet_0_clk _330_/a_27_47# 5.66e-19
C10661 clkbuf_2_2__f_clk/a_110_47# _330_/a_1283_21# 0.0109f
C10662 _303_/a_1108_47# net44 1.56e-20
C10663 _235_/a_79_21# _232_/a_32_297# 3.62e-19
C10664 _320_/a_543_47# _320_/a_805_47# 0.00171f
C10665 _320_/a_761_289# _320_/a_1217_47# 4.2e-19
C10666 _320_/a_1108_47# _320_/a_1270_413# 0.00645f
C10667 _309_/a_651_413# _081_ 8.91e-20
C10668 _309_/a_1108_47# _006_ 1.26e-19
C10669 _336_/a_1108_47# _032_ 3.86e-21
C10670 _323_/a_193_47# _303_/a_543_47# 3.24e-19
C10671 _323_/a_543_47# _303_/a_193_47# 2.56e-20
C10672 _323_/a_1283_21# _303_/a_27_47# 2.93e-20
C10673 _323_/a_761_289# _303_/a_761_289# 7e-20
C10674 trim_mask\[3\] _256_/a_27_297# 3.89e-20
C10675 _020_ clknet_2_3__leaf_clk 0.00112f
C10676 net12 _249_/a_109_47# 8.77e-19
C10677 _248_/a_109_47# _101_ 0.00145f
C10678 _322_/a_761_289# _101_ 0.00355f
C10679 _322_/a_27_47# net52 1.87e-19
C10680 _057_ net18 0.026f
C10681 _339_/a_193_47# _339_/a_652_21# 0.078f
C10682 _339_/a_27_47# _339_/a_476_47# 0.198f
C10683 net13 _320_/a_193_47# 0.00871f
C10684 VPWR _232_/a_220_297# 0.00569f
C10685 _062_ net40 0.122f
C10686 _251_/a_27_297# net29 5.81e-21
C10687 _317_/a_1283_21# state\[1\] 0.0668f
C10688 _317_/a_651_413# net45 0.0122f
C10689 net4 _190_/a_655_47# 0.00167f
C10690 _308_/a_1283_21# _307_/a_1108_47# 1.05e-20
C10691 _305_/a_761_289# net30 1.72e-20
C10692 net27 result[7] 8.81e-19
C10693 _035_ _001_ 1.09e-19
C10694 VPWR net49 0.357f
C10695 clknet_0_clk _120_ 8.5e-19
C10696 VPWR _272_/a_81_21# 0.239f
C10697 _315_/a_193_47# _315_/a_543_47# 0.229f
C10698 _315_/a_27_47# _315_/a_1283_21# 0.0435f
C10699 _321_/a_543_47# mask\[2\] 6.01e-19
C10700 mask\[4\] net20 1.68e-22
C10701 VPWR _336_/a_543_47# 0.209f
C10702 _117_ _275_/a_299_297# 2.22e-19
C10703 _276_/a_145_75# net50 1.8e-20
C10704 VPWR _290_/a_207_413# 0.166f
C10705 VPWR _329_/a_27_47# 0.518f
C10706 output8/a_27_47# _334_/a_1108_47# 0.00177f
C10707 net8 _334_/a_193_47# 0.0163f
C10708 _117_ _178_/a_68_297# 7.35e-20
C10709 _053_ _106_ 0.00112f
C10710 mask\[0\] _039_ 0.0319f
C10711 net4 trim_val\[4\] 0.0023f
C10712 _333_/a_193_47# _333_/a_639_47# 2.28e-19
C10713 _333_/a_761_289# _333_/a_1270_413# 2.6e-19
C10714 _333_/a_543_47# _333_/a_651_413# 0.0572f
C10715 _062_ _003_ 1.18e-20
C10716 fanout43/a_27_47# net22 4.37e-22
C10717 _103_ _052_ 9.12e-20
C10718 net16 _332_/a_1462_47# 2.04e-19
C10719 VPWR _239_/a_694_21# 0.194f
C10720 fanout44/a_27_47# _003_ 1.15e-19
C10721 _249_/a_27_297# _312_/a_27_47# 3.88e-21
C10722 _127_ _125_ 0.0731f
C10723 _037_ cal_count\[2\] 2.99e-19
C10724 clkbuf_2_0__f_clk/a_110_47# net30 0.0321f
C10725 _109_ _333_/a_27_47# 1.75e-20
C10726 _046_ _158_/a_150_297# 4.96e-19
C10727 _250_/a_27_297# net26 2.73e-20
C10728 ctln[2] trim[3] 2.75e-19
C10729 _251_/a_373_47# net15 5.93e-19
C10730 _323_/a_193_47# _249_/a_27_297# 1.81e-20
C10731 calibrate _315_/a_761_289# 0.0238f
C10732 _093_ _315_/a_193_47# 1.05e-19
C10733 _265_/a_384_47# trim_val\[0\] 3.13e-19
C10734 _074_ _315_/a_543_47# 0.016f
C10735 _326_/a_193_47# _251_/a_109_297# 1.92e-20
C10736 _309_/a_1217_47# _101_ 9.27e-21
C10737 _324_/a_1217_47# net44 8.4e-19
C10738 _161_/a_150_297# net33 3.83e-19
C10739 _063_ _190_/a_655_47# 0.0339f
C10740 _334_/a_543_47# net34 3.03e-21
C10741 VPWR _002_ 0.414f
C10742 _324_/a_761_289# net19 2.59e-19
C10743 en_co_clk clknet_2_3__leaf_clk 0.0129f
C10744 net3 _337_/a_1108_47# 6.9e-20
C10745 VPWR _289_/a_68_297# 0.176f
C10746 _232_/a_32_297# _049_ 0.0563f
C10747 _225_/a_109_297# _086_ 0.00114f
C10748 _192_/a_476_47# _065_ 7.4e-21
C10749 clknet_2_0__leaf_clk _315_/a_1283_21# 0.00635f
C10750 _014_ _315_/a_543_47# 4.82e-21
C10751 _090_ _099_ 0.07f
C10752 _307_/a_448_47# _307_/a_639_47# 4.61e-19
C10753 net45 _315_/a_761_289# 0.166f
C10754 _326_/a_1108_47# clknet_2_1__leaf_clk 0.00135f
C10755 _110_ _048_ 0.017f
C10756 _305_/a_761_289# _072_ 0.0264f
C10757 _305_/a_543_47# cal_itt\[3\] 6.56e-19
C10758 net13 _107_ 5.96e-20
C10759 _078_ net51 0.00111f
C10760 _167_/a_161_47# net3 0.0394f
C10761 _321_/a_193_47# _085_ 3.94e-21
C10762 net15 net55 1.07e-20
C10763 _235_/a_79_21# net55 0.0138f
C10764 _063_ trim_val\[4\] 6.93e-21
C10765 _322_/a_805_47# net44 0.0043f
C10766 VPWR _319_/a_805_47# 1.2e-19
C10767 _300_/a_129_47# net2 0.00236f
C10768 _107_ _279_/a_27_47# 0.0022f
C10769 _111_ rebuffer3/a_75_212# 1.05e-21
C10770 _318_/a_805_47# net45 0.00316f
C10771 _309_/a_27_47# _308_/a_448_47# 5.28e-21
C10772 _309_/a_543_47# _308_/a_543_47# 5.29e-20
C10773 _309_/a_193_47# _308_/a_1108_47# 7.29e-21
C10774 en net14 0.0186f
C10775 _074_ _093_ 3.37e-19
C10776 _126_ _125_ 0.272f
C10777 _110_ _330_/a_27_47# 0.00698f
C10778 net50 cal_count\[3\] 0.0229f
C10779 _189_/a_27_47# cal_itt\[3\] 2.17e-19
C10780 _015_ _092_ 4.53e-21
C10781 net43 _320_/a_193_47# 0.00113f
C10782 cal_count\[1\] _041_ 0.0426f
C10783 _058_ net34 7.39e-20
C10784 _020_ net20 2.56e-22
C10785 _323_/a_27_47# mask\[4\] 0.00766f
C10786 _305_/a_27_47# _305_/a_543_47# 0.106f
C10787 _305_/a_193_47# _305_/a_761_289# 0.172f
C10788 _237_/a_76_199# _237_/a_218_47# 0.00783f
C10789 VPWR _238_/a_75_212# 0.24f
C10790 _242_/a_79_21# _092_ 3.06e-20
C10791 _093_ _014_ 0.0073f
C10792 calibrate net45 0.158f
C10793 _303_/a_651_413# net19 0.00477f
C10794 _337_/a_1270_413# en_co_clk 7.91e-20
C10795 _332_/a_193_47# net40 0.0137f
C10796 trim_val\[3\] _258_/a_27_297# 1.39e-19
C10797 net1 _316_/a_543_47# 1.71e-20
C10798 _024_ _193_/a_109_297# 1.86e-19
C10799 _339_/a_476_47# _339_/a_586_47# 0.00807f
C10800 _339_/a_1032_413# _339_/a_956_413# 0.00212f
C10801 _339_/a_27_47# _339_/a_1224_47# 1.63e-19
C10802 _339_/a_652_21# _339_/a_796_47# 0.00196f
C10803 net43 net19 4.36e-20
C10804 net13 _320_/a_1462_47# 5.11e-19
C10805 net34 _332_/a_27_47# 2.82e-21
C10806 _309_/a_1283_21# _140_/a_68_297# 0.00109f
C10807 _341_/a_1283_21# _092_ 1.81e-21
C10808 _030_ _269_/a_81_21# 0.00419f
C10809 ctlp[1] net15 0.037f
C10810 net43 _307_/a_761_289# 3.38e-19
C10811 _078_ _224_/a_199_47# 7.62e-19
C10812 output35/a_27_47# output5/a_27_47# 3.56e-20
C10813 _320_/a_639_47# _040_ 0.00474f
C10814 input2/a_27_47# clkc 5.42e-19
C10815 cal_itt\[1\] _304_/a_761_289# 1.88e-19
C10816 _315_/a_448_47# _315_/a_639_47# 4.61e-19
C10817 output22/a_27_47# net23 3.74e-20
C10818 _337_/a_651_413# _076_ 1.38e-19
C10819 calibrate _065_ 3.98e-20
C10820 trim_mask\[4\] _279_/a_206_47# 0.00114f
C10821 _104_ _049_ 0.307f
C10822 net12 _048_ 0.489f
C10823 VPWR _106_ 0.516f
C10824 clk en 0.0348f
C10825 _064_ net30 0.184f
C10826 _292_/a_78_199# _339_/a_1182_261# 0.0121f
C10827 VPWR _329_/a_1217_47# 6.3e-20
C10828 net8 _334_/a_1462_47# 4.63e-19
C10829 _319_/a_1270_413# _049_ 3.27e-20
C10830 clk _330_/a_193_47# 0.00144f
C10831 _288_/a_59_75# _122_ 5.33e-20
C10832 _319_/a_448_47# net30 5.56e-19
C10833 _303_/a_193_47# _303_/a_761_289# 0.176f
C10834 _303_/a_27_47# _303_/a_543_47# 0.111f
C10835 _312_/a_805_47# _045_ 5.01e-20
C10836 net55 _049_ 0.0429f
C10837 net45 _065_ 6.92e-19
C10838 _065_ rebuffer3/a_75_212# 9.5e-22
C10839 clknet_2_1__leaf_clk _225_/a_109_297# 4.44e-19
C10840 _094_ _206_/a_27_93# 3.47e-19
C10841 net19 _118_ 3.87e-20
C10842 _313_/a_543_47# net29 1.85e-22
C10843 _124_ _123_ 0.0129f
C10844 _323_/a_27_47# _020_ 0.288f
C10845 _323_/a_543_47# mask\[5\] 4.63e-19
C10846 cal_itt\[1\] clkbuf_2_3__f_clk/a_110_47# 0.0102f
C10847 net54 _098_ 1.04e-19
C10848 _337_/a_1108_47# _062_ 9.67e-20
C10849 _320_/a_1283_21# mask\[4\] 7.02e-20
C10850 _101_ _208_/a_76_199# 0.00106f
C10851 net15 mask\[0\] 0.124f
C10852 _337_/a_1283_21# _075_ 0.0308f
C10853 _321_/a_27_47# _310_/a_27_47# 5.48e-21
C10854 _041_ _208_/a_505_21# 3.19e-20
C10855 net33 _132_ 0.00629f
C10856 _051_ _226_/a_197_47# 2.74e-19
C10857 _027_ net18 1.1e-19
C10858 _324_/a_27_47# _324_/a_1283_21# 0.0436f
C10859 _324_/a_193_47# _324_/a_543_47# 0.23f
C10860 _048_ net44 2e-20
C10861 _093_ _243_/a_27_297# 0.0328f
C10862 calibrate _243_/a_109_297# 0.0473f
C10863 net13 _248_/a_109_297# 0.00833f
C10864 net13 _322_/a_193_47# 0.0153f
C10865 state\[0\] _316_/a_448_47# 1.44e-20
C10866 net4 _330_/a_193_47# 2.27e-19
C10867 _308_/a_651_413# net43 0.0122f
C10868 _308_/a_1283_21# net23 0.0612f
C10869 clkbuf_2_2__f_clk/a_110_47# _108_ 7.12e-19
C10870 cal_itt\[0\] _035_ 0.0171f
C10871 _041_ mask\[2\] 0.284f
C10872 _316_/a_27_47# output41/a_27_47# 1.6e-21
C10873 _091_ _195_/a_505_21# 0.00583f
C10874 clknet_2_1__leaf_clk clknet_2_0__leaf_clk 0.028f
C10875 _319_/a_761_289# clknet_2_0__leaf_clk 0.0526f
C10876 _319_/a_27_47# net45 3.7e-19
C10877 net54 clknet_0_clk 4.49e-20
C10878 VPWR ctlp[2] 0.274f
C10879 _041_ _001_ 8.1e-20
C10880 _338_/a_1182_261# _001_ 5.8e-20
C10881 output6/a_27_47# net6 0.211f
C10882 _107_ _118_ 0.0151f
C10883 _325_/a_193_47# _159_/a_27_47# 2.65e-20
C10884 _309_/a_27_47# _005_ 9.51e-20
C10885 _110_ _330_/a_1217_47# 4.53e-19
C10886 _276_/a_59_75# _027_ 1.64e-21
C10887 _327_/a_448_47# net18 0.0021f
C10888 net43 _320_/a_1462_47# 1.48e-19
C10889 _264_/a_27_297# net30 0.0977f
C10890 _253_/a_81_21# _314_/a_761_289# 1.88e-22
C10891 _323_/a_1217_47# mask\[4\] 5.2e-19
C10892 net12 _076_ 0.619f
C10893 net43 net13 0.126f
C10894 VPWR _313_/a_1270_413# 7.57e-19
C10895 _309_/a_1283_21# _309_/a_1108_47# 0.234f
C10896 _309_/a_761_289# _309_/a_651_413# 0.0977f
C10897 _309_/a_543_47# _309_/a_448_47# 0.0498f
C10898 _309_/a_27_47# _309_/a_639_47# 0.00188f
C10899 _309_/a_193_47# _309_/a_1270_413# 1.46e-19
C10900 _048_ _263_/a_79_21# 0.154f
C10901 _152_/a_68_297# _152_/a_150_297# 0.00477f
C10902 _319_/a_27_47# _065_ 2.03e-19
C10903 _312_/a_543_47# _084_ 1.05e-19
C10904 _320_/a_27_47# _208_/a_76_199# 3.03e-21
C10905 VPWR output30/a_27_47# 0.403f
C10906 _110_ _334_/a_761_289# 6.43e-21
C10907 _136_ _267_/a_145_75# 1.14e-19
C10908 VPWR _278_/a_109_297# 0.00384f
C10909 _256_/a_373_47# _058_ 2.63e-19
C10910 _322_/a_27_47# _322_/a_761_289# 0.0532f
C10911 _248_/a_27_297# _248_/a_109_47# 0.00393f
C10912 _322_/a_193_47# _248_/a_109_297# 3.84e-19
C10913 _322_/a_761_289# _248_/a_27_297# 0.00173f
C10914 net50 trim_mask\[2\] 0.00675f
C10915 _110_ _327_/a_27_47# 1.76e-20
C10916 _241_/a_105_352# _095_ 0.211f
C10917 clknet_0_clk _068_ 0.0251f
C10918 _305_/a_1108_47# clknet_2_1__leaf_clk 9.63e-21
C10919 net42 cal_itt\[3\] 2.24e-19
C10920 _232_/a_32_297# state\[1\] 8.56e-19
C10921 _257_/a_27_297# _257_/a_109_47# 0.00393f
C10922 _168_/a_207_413# _049_ 0.00139f
C10923 _210_/a_113_297# _315_/a_27_47# 3.34e-20
C10924 _269_/a_299_297# trim_val\[1\] 0.0585f
C10925 _269_/a_81_21# trim_mask\[1\] 0.118f
C10926 VPWR _270_/a_145_75# 0.00207f
C10927 _146_/a_68_297# clknet_2_1__leaf_clk 0.0653f
C10928 _043_ _311_/a_27_47# 8.03e-22
C10929 _239_/a_27_297# calibrate 0.113f
C10930 mask\[0\] _049_ 0.0782f
C10931 _262_/a_193_297# net55 0.00126f
C10932 net9 _268_/a_75_212# 0.00327f
C10933 net44 _076_ 0.148f
C10934 _104_ fanout46/a_27_47# 0.0101f
C10935 clkbuf_2_1__f_clk/a_110_47# _319_/a_1283_21# 0.00615f
C10936 input2/a_27_47# _130_ 0.0114f
C10937 _301_/a_377_297# en_co_clk 5.5e-20
C10938 _325_/a_1283_21# _101_ 0.00102f
C10939 _325_/a_761_289# net52 1.3e-20
C10940 mask\[3\] _245_/a_27_297# 1.03e-19
C10941 cal_count\[1\] _339_/a_1032_413# 0.0161f
C10942 _036_ _339_/a_1182_261# 9.37e-20
C10943 _276_/a_59_75# _335_/a_448_47# 4.67e-19
C10944 _110_ _335_/a_27_47# 0.0268f
C10945 _256_/a_27_297# _108_ 1.48e-19
C10946 VPWR output36/a_27_47# 0.497f
C10947 clkbuf_2_0__f_clk/a_110_47# _319_/a_1108_47# 1.63e-20
C10948 en_co_clk _263_/a_382_297# 1.73e-19
C10949 _341_/a_193_47# en_co_clk 5.4e-20
C10950 mask\[6\] _074_ 0.491f
C10951 _279_/a_27_47# _118_ 0.0492f
C10952 _279_/a_396_47# trim_val\[4\] 0.00958f
C10953 _048_ clknet_2_2__leaf_clk 2.04e-20
C10954 _291_/a_117_297# trimb[1] 2.67e-19
C10955 _243_/a_27_297# _243_/a_109_47# 0.00393f
C10956 _162_/a_27_47# _108_ 0.00185f
C10957 net2 _202_/a_297_47# 0.0404f
C10958 cal_itt\[1\] clkbuf_0_clk/a_110_47# 0.0143f
C10959 _317_/a_193_47# _316_/a_193_47# 9.38e-21
C10960 _317_/a_27_47# _316_/a_761_289# 0.00112f
C10961 _292_/a_493_297# _292_/a_215_47# 3.25e-19
C10962 cal_itt\[1\] cal_count\[3\] 7.38e-21
C10963 _305_/a_1283_21# _202_/a_297_47# 3e-19
C10964 clknet_2_2__leaf_clk _330_/a_27_47# 0.514f
C10965 _110_ rebuffer1/a_75_212# 9.81e-20
C10966 mask\[4\] _205_/a_27_47# 1.07e-21
C10967 net52 _077_ 5.79e-19
C10968 VPWR _316_/a_1108_47# 0.314f
C10969 _321_/a_448_47# _310_/a_1108_47# 2e-21
C10970 _210_/a_113_297# clknet_2_0__leaf_clk 0.0654f
C10971 cal_itt\[0\] _198_/a_27_47# 0.0715f
C10972 _324_/a_448_47# _324_/a_639_47# 4.61e-19
C10973 _106_ _262_/a_27_47# 0.0964f
C10974 _306_/a_761_289# _003_ 2.33e-20
C10975 _306_/a_543_47# _073_ 9.17e-19
C10976 state\[0\] _013_ 7.07e-20
C10977 net12 mask\[3\] 0.011f
C10978 _238_/a_75_212# _093_ 0.0377f
C10979 _257_/a_109_47# trim_val\[4\] 4.68e-19
C10980 _330_/a_27_47# net11 1.44e-20
C10981 _330_/a_761_289# net19 0.00452f
C10982 _338_/a_1296_47# _001_ 1.29e-19
C10983 _041_ mask\[1\] 0.0171f
C10984 ctlp[7] net28 0.00152f
C10985 _051_ net46 1.84e-21
C10986 state\[1\] net55 0.0176f
C10987 _335_/a_761_289# _280_/a_75_212# 1.36e-21
C10988 _309_/a_805_47# net43 0.00378f
C10989 net14 _310_/a_1108_47# 4.01e-19
C10990 net15 _121_ 0.0264f
C10991 _094_ _282_/a_150_297# 7.8e-19
C10992 _258_/a_27_297# _327_/a_543_47# 1.14e-20
C10993 _327_/a_448_47# trim_mask\[0\] 7.47e-20
C10994 _327_/a_543_47# _024_ 0.00409f
C10995 VPWR ctln[2] 0.182f
C10996 _089_ _228_/a_79_21# 0.111f
C10997 net15 _010_ 0.00749f
C10998 _053_ _304_/a_805_47# 6.41e-19
C10999 _053_ _340_/a_652_21# 2.67e-20
C11000 _251_/a_27_297# _251_/a_109_297# 0.171f
C11001 mask\[3\] net44 0.295f
C11002 _320_/a_761_289# _077_ 4.25e-20
C11003 _277_/a_75_212# _335_/a_193_47# 0.00452f
C11004 _030_ net32 3.33e-21
C11005 _306_/a_27_47# clknet_0_clk 1.07e-20
C11006 result[7] _011_ 0.00565f
C11007 _322_/a_543_47# _322_/a_805_47# 0.00171f
C11008 _322_/a_761_289# _322_/a_1217_47# 4.2e-19
C11009 _322_/a_1108_47# _322_/a_1270_413# 0.00645f
C11010 _322_/a_1283_21# mask\[4\] 0.0114f
C11011 VPWR _298_/a_78_199# 0.298f
C11012 _058_ net4 4.91e-20
C11013 _257_/a_109_297# _025_ 0.00186f
C11014 _114_ _176_/a_27_47# 1.25e-20
C11015 _032_ net18 4.23e-19
C11016 mask\[0\] _315_/a_1108_47# 6.28e-21
C11017 _060_ clk 1.07e-20
C11018 net4 _335_/a_193_47# 0.00102f
C11019 _272_/a_81_21# _272_/a_384_47# 0.00138f
C11020 mask\[5\] _152_/a_150_297# 9.54e-19
C11021 _023_ _310_/a_27_47# 6.27e-19
C11022 _327_/a_639_47# _136_ 3.85e-19
C11023 net12 net54 3.08e-20
C11024 net47 _068_ 3.15e-19
C11025 cal_itt\[0\] _041_ 0.0129f
C11026 _336_/a_543_47# _336_/a_1108_47# 7.99e-20
C11027 _336_/a_193_47# _336_/a_651_413# 0.0346f
C11028 _050_ _028_ 0.182f
C11029 _319_/a_761_289# _319_/a_639_47# 3.16e-19
C11030 _319_/a_27_47# _319_/a_1217_47# 2.56e-19
C11031 output35/a_27_47# _047_ 0.00251f
C11032 _106_ wire42/a_75_212# 1.27e-20
C11033 _237_/a_218_47# _048_ 1.16e-19
C11034 _276_/a_59_75# _032_ 0.0323f
C11035 trim_mask\[0\] _332_/a_1108_47# 0.0462f
C11036 _329_/a_27_47# _329_/a_761_289# 0.0701f
C11037 _327_/a_27_47# _341_/a_27_47# 4.43e-21
C11038 _078_ _086_ 0.00406f
C11039 _286_/a_218_374# _122_ 7.33e-19
C11040 _060_ net4 1.05e-19
C11041 net24 _074_ 0.05f
C11042 _121_ _049_ 0.0172f
C11043 _324_/a_1108_47# _020_ 0.00287f
C11044 _006_ _310_/a_193_47# 1.06e-20
C11045 net54 net44 1.35e-20
C11046 fanout43/a_27_47# _245_/a_27_297# 0.0216f
C11047 net13 net3 0.0105f
C11048 _002_ _202_/a_79_21# 0.107f
C11049 _144_/a_27_47# output40/a_27_47# 2.19e-20
C11050 clknet_2_2__leaf_clk _330_/a_1217_47# 4.62e-19
C11051 _209_/a_27_47# _076_ 0.00552f
C11052 state\[0\] _051_ 0.205f
C11053 _062_ net19 0.248f
C11054 _328_/a_543_47# net46 0.155f
C11055 _064_ _066_ 6.91e-19
C11056 _008_ _218_/a_113_297# 0.15f
C11057 _197_/a_199_47# _069_ 0.00189f
C11058 _259_/a_27_297# _033_ 4.61e-19
C11059 _104_ _336_/a_651_413# 5.97e-19
C11060 _074_ _313_/a_805_47# 1.15e-20
C11061 _334_/a_761_289# clknet_2_2__leaf_clk 5.11e-19
C11062 _088_ _260_/a_93_21# 2.44e-19
C11063 _327_/a_27_47# clknet_2_2__leaf_clk 0.3f
C11064 VPWR _304_/a_805_47# 1.82e-19
C11065 _097_ _232_/a_32_297# 3.18e-20
C11066 net28 _222_/a_113_297# 0.00758f
C11067 _325_/a_543_47# net13 0.00146f
C11068 net44 _068_ 0.0278f
C11069 VPWR _340_/a_652_21# 0.25f
C11070 net54 _263_/a_79_21# 0.00361f
C11071 output21/a_27_47# _156_/a_27_47# 1.13e-19
C11072 _218_/a_113_297# mask\[5\] 9e-21
C11073 _303_/a_1108_47# _001_ 2.64e-20
C11074 _053_ _338_/a_27_47# 1.98e-21
C11075 _249_/a_27_297# _084_ 1.18e-20
C11076 _195_/a_76_199# net19 7.11e-20
C11077 _274_/a_75_212# rebuffer1/a_75_212# 1.32e-20
C11078 trim[2] _056_ 0.00662f
C11079 _107_ _062_ 0.0161f
C11080 net33 net32 1.61e-19
C11081 ctln[5] ctln[6] 0.00305f
C11082 _251_/a_27_297# _022_ 0.11f
C11083 _081_ _039_ 9.79e-21
C11084 net12 net27 0.331f
C11085 net31 trim[0] 0.0191f
C11086 rebuffer3/a_75_212# _278_/a_27_47# 2.1e-20
C11087 net52 _310_/a_1108_47# 9.14e-20
C11088 _308_/a_1108_47# mask\[1\] 1.87e-20
C11089 _335_/a_27_47# clknet_2_2__leaf_clk 0.247f
C11090 _269_/a_299_297# _172_/a_150_297# 8.01e-20
C11091 _328_/a_639_47# _058_ 5.31e-19
C11092 _321_/a_1283_21# _018_ 4.83e-21
C11093 trim_mask\[2\] _335_/a_1108_47# 5.98e-21
C11094 _341_/a_1283_21# net46 0.293f
C11095 _282_/a_68_297# _065_ 0.181f
C11096 _052_ _242_/a_297_47# 0.00891f
C11097 clknet_2_1__leaf_clk _078_ 0.0378f
C11098 _246_/a_27_297# _246_/a_373_47# 0.0134f
C11099 net27 _159_/a_27_47# 0.0334f
C11100 mask\[0\] _319_/a_543_47# 0.036f
C11101 _202_/a_297_47# _070_ 0.0486f
C11102 trimb[1] net37 0.0164f
C11103 _333_/a_27_47# net46 0.665f
C11104 _321_/a_543_47# net26 6.88e-20
C11105 _307_/a_193_47# _137_/a_150_297# 5.99e-20
C11106 _083_ mask\[4\] 0.365f
C11107 _329_/a_1108_47# net48 2.35e-20
C11108 _325_/a_1283_21# _322_/a_27_47# 1.42e-20
C11109 _336_/a_1108_47# _106_ 3.75e-20
C11110 cal_count\[0\] net34 1.94e-19
C11111 en_co_clk _095_ 0.648f
C11112 trim_mask\[2\] rebuffer2/a_75_212# 6.01e-22
C11113 net44 _311_/a_448_47# 8.11e-19
C11114 net43 _080_ 0.00271f
C11115 net27 net44 0.105f
C11116 _322_/a_1108_47# rebuffer5/a_161_47# 2.12e-19
C11117 _267_/a_59_75# _109_ 0.0986f
C11118 _189_/a_408_47# _103_ 2.68e-19
C11119 _329_/a_543_47# _329_/a_805_47# 0.00171f
C11120 _329_/a_761_289# _329_/a_1217_47# 4.2e-19
C11121 _329_/a_1108_47# _329_/a_1270_413# 0.00645f
C11122 _094_ _337_/a_193_47# 0.0221f
C11123 VPWR _321_/a_805_47# 1.18e-19
C11124 _323_/a_27_47# _311_/a_1108_47# 5.58e-19
C11125 _323_/a_193_47# _311_/a_1283_21# 1.72e-19
C11126 _105_ _278_/a_27_47# 8.14e-20
C11127 _188_/a_27_47# _135_ 1.17e-19
C11128 _319_/a_27_47# _282_/a_68_297# 7.58e-19
C11129 clknet_2_1__leaf_clk _313_/a_651_413# 0.00144f
C11130 _306_/a_1108_47# clkbuf_0_clk/a_110_47# 2.75e-19
C11131 _306_/a_193_47# clk 2.25e-19
C11132 mask\[7\] _224_/a_199_47# 0.0106f
C11133 _220_/a_113_297# _084_ 0.0981f
C11134 net13 fanout44/a_27_47# 0.00419f
C11135 VPWR _337_/a_805_47# 1.5e-19
C11136 _247_/a_109_297# _101_ 0.0133f
C11137 _327_/a_1108_47# _265_/a_299_297# 1.68e-20
C11138 _281_/a_253_297# _281_/a_253_47# 0.00137f
C11139 _286_/a_439_47# net18 2.47e-19
C11140 _065_ _204_/a_75_212# 1.15e-19
C11141 net7 net14 3.57e-21
C11142 net12 _306_/a_27_47# 0.0176f
C11143 _110_ net10 1.95e-20
C11144 _317_/a_193_47# net14 5.64e-19
C11145 _014_ _316_/a_651_413# 0.00325f
C11146 net45 _316_/a_448_47# 7.54e-19
C11147 _326_/a_193_47# net14 0.00884f
C11148 _097_ net55 1.31e-20
C11149 _325_/a_543_47# net43 0.161f
C11150 trim_mask\[4\] _027_ 3.06e-19
C11151 _061_ net34 6.04e-19
C11152 _015_ state\[0\] 0.268f
C11153 _305_/a_543_47# _073_ 4.8e-21
C11154 net5 _061_ 0.00366f
C11155 _322_/a_805_47# mask\[2\] 1.81e-19
C11156 net35 _333_/a_1283_21# 1.16e-19
C11157 net15 _245_/a_109_297# 4.09e-19
C11158 _214_/a_113_297# _247_/a_27_297# 5.11e-20
C11159 _182_/a_27_47# _109_ 1.08e-19
C11160 fanout45/a_27_47# _317_/a_1283_21# 0.00344f
C11161 _309_/a_193_47# mask\[3\] 1.96e-19
C11162 _309_/a_761_289# net25 1.47e-19
C11163 _329_/a_1270_413# net9 1.44e-19
C11164 net8 _176_/a_27_47# 2.96e-19
C11165 _050_ _095_ 0.501f
C11166 _026_ _064_ 9.32e-20
C11167 _253_/a_299_297# net26 6.75e-19
C11168 _134_ _332_/a_761_289# 2.32e-19
C11169 trim[2] _173_/a_27_47# 8.78e-19
C11170 VPWR _245_/a_373_47# 6.3e-19
C11171 clknet_0_clk cal_itt\[3\] 0.0237f
C11172 VPWR _338_/a_27_47# 0.697f
C11173 _306_/a_27_47# net44 0.304f
C11174 clk _227_/a_109_93# 0.00819f
C11175 _326_/a_1283_21# _253_/a_299_297# 0.00155f
C11176 _333_/a_761_289# rebuffer2/a_75_212# 7.71e-20
C11177 _291_/a_35_297# _291_/a_117_297# 0.00641f
C11178 VPWR _340_/a_1056_47# 4.86e-19
C11179 _275_/a_384_47# net50 3.6e-19
C11180 _333_/a_651_413# rebuffer1/a_75_212# 4.98e-20
C11181 _333_/a_543_47# _108_ 0.0112f
C11182 _333_/a_193_47# _332_/a_1108_47# 1.42e-21
C11183 _341_/a_543_47# _053_ 3.23e-19
C11184 trim_mask\[0\] _171_/a_27_47# 3.71e-19
C11185 VPWR _102_ 0.508f
C11186 _275_/a_299_297# _057_ 2.45e-19
C11187 _109_ net37 7.01e-21
C11188 trim[2] net48 2.08e-19
C11189 _265_/a_384_47# _108_ 1.18e-19
C11190 _178_/a_68_297# _057_ 0.106f
C11191 clk net7 0.0053f
C11192 _304_/a_27_47# _065_ 0.0109f
C11193 _337_/a_1270_413# _049_ 1.04e-19
C11194 clk _317_/a_193_47# 0.00965f
C11195 _103_ clone1/a_27_47# 0.00696f
C11196 _336_/a_1283_21# _278_/a_27_47# 2.4e-21
C11197 clknet_0_clk _262_/a_205_47# 1.91e-20
C11198 _210_/a_113_297# _078_ 0.0496f
C11199 _210_/a_199_47# mask\[0\] 0.0106f
C11200 net23 _212_/a_199_47# 0.0015f
C11201 _304_/a_543_47# net2 3.56e-20
C11202 output32/a_27_47# net33 0.00242f
C11203 _164_/a_161_47# en_co_clk 9.44e-19
C11204 _321_/a_193_47# _074_ 1.2e-19
C11205 net4 _227_/a_109_93# 1.04e-21
C11206 _306_/a_543_47# _101_ 4.44e-21
C11207 _081_ net15 4.63e-20
C11208 net43 fanout44/a_27_47# 0.0499f
C11209 net14 net30 0.0107f
C11210 _333_/a_1217_47# net46 6.24e-19
C11211 _096_ clone7/a_27_47# 0.00608f
C11212 _307_/a_1108_47# _039_ 0.0336f
C11213 net33 clkc 2.25e-19
C11214 VPWR _331_/a_1270_413# 7.89e-19
C11215 net4 net7 0.0774f
C11216 VPWR _006_ 0.689f
C11217 _322_/a_543_47# mask\[3\] 0.0512f
C11218 _124_ clknet_2_3__leaf_clk 2.19e-19
C11219 _332_/a_805_47# clknet_2_2__leaf_clk 2.34e-19
C11220 net4 _317_/a_193_47# 0.0134f
C11221 _321_/a_761_289# clknet_2_0__leaf_clk 1.49e-20
C11222 _307_/a_1283_21# fanout43/a_27_47# 3.85e-22
C11223 result[0] _039_ 2.93e-19
C11224 VPWR _328_/a_761_289# 0.215f
C11225 _078_ _313_/a_27_47# 0.00921f
C11226 cal_itt\[0\] _303_/a_1108_47# 0.00177f
C11227 cal_itt\[1\] _303_/a_1283_21# 4.77e-20
C11228 _233_/a_373_47# net14 7.15e-19
C11229 VPWR net17 1.33f
C11230 calibrate _013_ 0.0224f
C11231 _300_/a_129_47# clknet_2_3__leaf_clk 0.00307f
C11232 _094_ _337_/a_1462_47# 2.57e-19
C11233 VPWR _089_ 0.255f
C11234 _337_/a_27_47# net45 2.29e-20
C11235 _337_/a_761_289# clknet_2_0__leaf_clk 6.55e-19
C11236 net28 _314_/a_448_47# 0.0037f
C11237 _309_/a_193_47# _310_/a_1283_21# 5.38e-20
C11238 _309_/a_27_47# _310_/a_1108_47# 3.96e-19
C11239 trim_mask\[3\] _330_/a_27_47# 7.85e-20
C11240 _018_ _101_ 0.0498f
C11241 _064_ net40 0.347f
C11242 _257_/a_109_47# _058_ 1.22e-19
C11243 VPWR _312_/a_193_47# 0.574f
C11244 net2 _035_ 4.55e-20
C11245 _090_ net41 0.00615f
C11246 net12 _306_/a_1217_47# 8.28e-20
C11247 _062_ _118_ 0.0742f
C11248 net4 _286_/a_76_199# 7.84e-21
C11249 _110_ _271_/a_75_212# 0.00989f
C11250 net45 _013_ 0.0723f
C11251 _166_/a_161_47# _048_ 7.08e-20
C11252 _050_ _164_/a_161_47# 5.94e-19
C11253 VPWR _323_/a_761_289# 0.215f
C11254 net43 _082_ 0.00876f
C11255 net23 net25 2.16e-22
C11256 _313_/a_27_47# _313_/a_651_413# 9.73e-19
C11257 _313_/a_761_289# _313_/a_1108_47# 0.0512f
C11258 _313_/a_193_47# _313_/a_448_47# 0.0612f
C11259 _336_/a_193_47# clkbuf_2_2__f_clk/a_110_47# 0.0151f
C11260 clk _054_ 0.00996f
C11261 _312_/a_193_47# net53 5.31e-20
C11262 cal_itt\[2\] _190_/a_655_47# 4.48e-19
C11263 cal_itt\[1\] _190_/a_215_47# 7.48e-20
C11264 _041_ net26 5.16e-20
C11265 clk _318_/a_1283_21# 0.031f
C11266 _337_/a_27_47# _065_ 0.0302f
C11267 clk net30 1.03f
C11268 net15 _016_ 0.0382f
C11269 net12 _318_/a_543_47# 7.82e-19
C11270 _326_/a_193_47# net52 0.00214f
C11271 en_co_clk _207_/a_109_297# 0.00235f
C11272 _259_/a_109_297# net18 5.32e-19
C11273 VPWR _301_/a_285_47# 0.0118f
C11274 output35/a_27_47# trim_val\[0\] 6.59e-20
C11275 _169_/a_215_311# _092_ 1.18e-21
C11276 _325_/a_193_47# mask\[2\] 9.95e-20
C11277 _306_/a_1217_47# net44 6.03e-19
C11278 VPWR _341_/a_543_47# 0.204f
C11279 _312_/a_193_47# _009_ 0.234f
C11280 _326_/a_639_47# mask\[7\] 1.47e-19
C11281 _326_/a_1270_413# _102_ 5.01e-20
C11282 _173_/a_27_47# _055_ 0.197f
C11283 _136_ _300_/a_377_297# 6.58e-19
C11284 _309_/a_193_47# fanout43/a_27_47# 3.37e-20
C11285 net4 net30 0.0619f
C11286 _041_ _286_/a_535_374# 3.12e-19
C11287 _208_/a_76_199# _077_ 0.105f
C11288 _330_/a_193_47# _330_/a_543_47# 0.22f
C11289 _330_/a_27_47# _330_/a_1283_21# 0.0436f
C11290 _208_/a_505_21# _076_ 0.254f
C11291 _304_/a_1217_47# _065_ 2.55e-19
C11292 net43 _314_/a_805_47# 0.00316f
C11293 clk _317_/a_1462_47# 2.24e-19
C11294 VPWR _308_/a_193_47# 0.605f
C11295 en_co_clk _226_/a_27_47# 0.00555f
C11296 _264_/a_27_297# net40 1.87e-19
C11297 net55 _240_/a_109_297# 0.00361f
C11298 _315_/a_651_413# net14 0.00176f
C11299 trim_val\[2\] net34 0.0981f
C11300 _116_ fanout46/a_27_47# 9.48e-21
C11301 _104_ clkbuf_2_2__f_clk/a_110_47# 0.0012f
C11302 _288_/a_59_75# cal_count\[2\] 8.42e-19
C11303 _340_/a_1602_47# net2 4.96e-19
C11304 output24/a_27_47# result[2] 0.332f
C11305 _319_/a_1283_21# clknet_0_clk 0.0256f
C11306 VPWR trimb[1] 0.537f
C11307 _222_/a_113_297# _085_ 0.0972f
C11308 _249_/a_27_297# _311_/a_193_47# 3.43e-19
C11309 clk _072_ 0.207f
C11310 VPWR _320_/a_448_47# 0.0828f
C11311 _097_ _316_/a_543_47# 3.7e-19
C11312 clkbuf_2_2__f_clk/a_110_47# net55 3.7e-19
C11313 net16 net34 0.0142f
C11314 net12 cal_itt\[3\] 0.012f
C11315 VPWR _339_/a_193_47# 0.294f
C11316 net5 net16 3.66e-20
C11317 _094_ _090_ 2.67e-20
C11318 net43 _310_/a_448_47# 5.45e-19
C11319 output16/a_27_47# trimb[3] 6.54e-19
C11320 ctlp[2] output39/a_27_47# 0.0101f
C11321 result[5] output28/a_27_47# 6.68e-19
C11322 output27/a_27_47# result[6] 7.93e-20
C11323 _051_ calibrate 0.00542f
C11324 _035_ _123_ 1.21e-19
C11325 _232_/a_32_297# _337_/a_543_47# 5.02e-21
C11326 _303_/a_639_47# _068_ 2.23e-19
C11327 net33 _130_ 0.00557f
C11328 cal_itt\[2\] _000_ 0.00363f
C11329 _263_/a_382_297# _049_ 2.17e-20
C11330 net52 net30 1.74e-20
C11331 ctlp[6] _312_/a_761_289# 0.00104f
C11332 _324_/a_1283_21# net27 0.00397f
C11333 _063_ net30 0.0247f
C11334 _162_/a_27_47# trim_val\[1\] 3.66e-20
C11335 _305_/a_193_47# clk 0.00448f
C11336 _305_/a_1108_47# clkbuf_0_clk/a_110_47# 0.00789f
C11337 _322_/a_193_47# _247_/a_27_297# 1.58e-20
C11338 net31 net35 1.68e-19
C11339 net2 _198_/a_27_47# 3.03e-20
C11340 net12 _305_/a_27_47# 5.89e-19
C11341 trim_mask\[3\] _330_/a_1217_47# 1.1e-19
C11342 _275_/a_81_21# net46 1.21e-19
C11343 _051_ net45 0.00193f
C11344 _325_/a_193_47# _325_/a_1108_47# 0.125f
C11345 _325_/a_27_47# _325_/a_448_47# 0.0919f
C11346 _110_ _269_/a_384_47# 1.12e-19
C11347 _050_ _226_/a_27_47# 6.6e-19
C11348 net4 cal_count\[0\] 2.07e-19
C11349 _255_/a_27_47# _103_ 0.0945f
C11350 net16 _299_/a_298_297# 0.00289f
C11351 VPWR _307_/a_651_413# 0.143f
C11352 _302_/a_109_297# trim_mask\[1\] 2.79e-21
C11353 _090_ _192_/a_505_280# 0.00181f
C11354 _107_ _227_/a_209_311# 0.00952f
C11355 net44 cal_itt\[3\] 0.0612f
C11356 mask\[4\] _311_/a_27_47# 0.228f
C11357 mask\[7\] _086_ 0.0853f
C11358 _185_/a_68_297# _048_ 8.76e-22
C11359 _313_/a_193_47# _010_ 0.217f
C11360 _126_ _122_ 1.19e-19
C11361 _334_/a_27_47# _057_ 9.67e-20
C11362 _337_/a_1217_47# _065_ 9.91e-20
C11363 trim_mask\[3\] _327_/a_27_47# 1.68e-20
C11364 _305_/a_193_47# net4 6.04e-21
C11365 _051_ _065_ 8.6e-23
C11366 net43 _247_/a_27_297# 4.34e-21
C11367 net23 _039_ 1.96e-19
C11368 net3 _062_ 0.0875f
C11369 _321_/a_1108_47# _042_ 0.016f
C11370 _064_ _256_/a_109_47# 0.00344f
C11371 _104_ _256_/a_27_297# 0.226f
C11372 _305_/a_27_47# net44 0.0191f
C11373 output35/a_27_47# _131_ 4.38e-22
C11374 _322_/a_1108_47# net51 3.81e-20
C11375 _028_ _049_ 0.00101f
C11376 _053_ _092_ 0.0183f
C11377 mask\[3\] mask\[2\] 0.0187f
C11378 result[1] net14 5.96e-20
C11379 _321_/a_639_47# clknet_2_1__leaf_clk 0.00108f
C11380 _289_/a_68_297# _129_ 0.00941f
C11381 _126_ _299_/a_27_413# 4.82e-20
C11382 trim_mask\[4\] _171_/a_27_47# 7.91e-20
C11383 _316_/a_27_47# _316_/a_193_47# 0.904f
C11384 net43 result[5] 7.57e-19
C11385 _058_ _193_/a_109_297# 2.5e-19
C11386 VPWR _333_/a_805_47# 4.56e-19
C11387 VPWR _303_/a_193_47# 0.581f
C11388 _340_/a_1602_47# _123_ 0.00883f
C11389 _063_ _072_ 0.00253f
C11390 trim_mask\[3\] _335_/a_27_47# 0.002f
C11391 trim_val\[3\] _335_/a_193_47# 8.29e-19
C11392 output28/a_27_47# net29 2.96e-19
C11393 VPWR _109_ 0.355f
C11394 _008_ _311_/a_543_47# 5.01e-19
C11395 _330_/a_448_47# _330_/a_639_47# 4.61e-19
C11396 _172_/a_68_297# _055_ 0.105f
C11397 _301_/a_47_47# _300_/a_285_47# 1.53e-19
C11398 _301_/a_285_47# _300_/a_47_47# 1.53e-19
C11399 trim_mask\[1\] cal_count\[3\] 2.64e-20
C11400 _037_ cal_count\[0\] 2.17e-20
C11401 _338_/a_193_47# _065_ 1.8e-20
C11402 VPWR _308_/a_1462_47# 4.04e-19
C11403 _337_/a_543_47# net55 0.00186f
C11404 net27 _044_ 0.00619f
C11405 _048_ _088_ 0.283f
C11406 _341_/a_27_47# _300_/a_285_47# 6.92e-21
C11407 state\[2\] _318_/a_448_47# 3.21e-21
C11408 _305_/a_193_47# _063_ 7.72e-20
C11409 _125_ _131_ 3e-21
C11410 _307_/a_543_47# net30 1.21e-19
C11411 _262_/a_465_47# _063_ 2.79e-19
C11412 net2 _297_/a_129_47# 5.79e-19
C11413 _284_/a_68_297# _122_ 0.111f
C11414 _187_/a_27_413# _134_ 6.26e-19
C11415 VPWR _309_/a_1283_21# 0.392f
C11416 VPWR _152_/a_68_297# 0.175f
C11417 net43 rebuffer6/a_27_47# 9.98e-21
C11418 mask\[1\] _076_ 2.4e-19
C11419 net16 _133_ 0.0261f
C11420 net45 _331_/a_639_47# 9.54e-19
C11421 _271_/a_75_212# clknet_2_2__leaf_clk 0.0696f
C11422 _074_ _312_/a_543_47# 3.22e-20
C11423 clkbuf_2_1__f_clk/a_110_47# _101_ 0.0272f
C11424 trim_mask\[0\] net49 5.76e-20
C11425 _200_/a_80_21# _200_/a_209_297# 0.0626f
C11426 VPWR _339_/a_796_47# 1.16e-19
C11427 _015_ calibrate 0.0209f
C11428 net15 _040_ 0.0131f
C11429 _328_/a_1108_47# _030_ 0.00135f
C11430 trim_mask\[0\] _336_/a_543_47# 4.83e-20
C11431 _014_ _090_ 0.00256f
C11432 en_co_clk _195_/a_535_374# 0.00124f
C11433 cal_itt\[1\] en_co_clk 0.133f
C11434 mask\[7\] clknet_2_1__leaf_clk 0.00293f
C11435 net43 _306_/a_761_289# 1.24e-20
C11436 calibrate _242_/a_79_21# 0.00314f
C11437 VPWR _279_/a_490_47# 9.97e-19
C11438 _015_ net45 0.0237f
C11439 net12 _250_/a_109_297# 0.00775f
C11440 VPWR _292_/a_493_297# 0.00253f
C11441 _335_/a_27_47# _330_/a_1283_21# 0.011f
C11442 _064_ _280_/a_75_212# 0.0176f
C11443 _216_/a_113_297# net25 0.021f
C11444 output34/a_27_47# _334_/a_1283_21# 9e-19
C11445 _110_ _336_/a_1270_413# 1.39e-19
C11446 VPWR _324_/a_651_413# 0.144f
C11447 output22/a_27_47# clknet_2_0__leaf_clk 0.0311f
C11448 net43 net29 0.0617f
C11449 VPWR _158_/a_150_297# 0.00213f
C11450 _329_/a_1108_47# _110_ 2.85e-19
C11451 _048_ _108_ 0.00102f
C11452 _302_/a_109_47# _067_ 1.47e-19
C11453 mask\[4\] _311_/a_1217_47# 8.37e-19
C11454 cal_count\[1\] _125_ 0.0748f
C11455 net15 _095_ 0.0835f
C11456 _235_/a_79_21# _095_ 0.111f
C11457 _313_/a_1462_47# _010_ 4.67e-20
C11458 _239_/a_27_297# _051_ 4.51e-19
C11459 net19 _150_/a_27_47# 8.67e-19
C11460 output20/a_27_47# output21/a_27_47# 4.46e-21
C11461 _104_ _331_/a_193_47# 1.36e-22
C11462 _324_/a_651_413# net53 6.01e-19
C11463 _320_/a_27_47# clkbuf_2_1__f_clk/a_110_47# 0.013f
C11464 _237_/a_439_47# _049_ 7.78e-20
C11465 _015_ _065_ 2.22e-19
C11466 _255_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 1.92e-20
C11467 VPWR _322_/a_448_47# 0.0794f
C11468 _259_/a_27_297# trim_mask\[2\] 9.79e-20
C11469 VPWR _092_ 3.61f
C11470 _064_ _258_/a_109_297# 0.0106f
C11471 _083_ _311_/a_1108_47# 1.65e-20
C11472 _001_ _068_ 1.8e-20
C11473 output25/a_27_47# net26 6.71e-20
C11474 _308_/a_543_47# _074_ 0.0157f
C11475 _041_ _123_ 0.0407f
C11476 _030_ _333_/a_761_289# 7.67e-19
C11477 _113_ _333_/a_543_47# 3.51e-20
C11478 _293_/a_81_21# trimb[4] 9.37e-20
C11479 _338_/a_1182_261# _123_ 3.03e-20
C11480 ctln[7] _318_/a_543_47# 1.28e-19
C11481 net13 _318_/a_1108_47# 0.00312f
C11482 _316_/a_543_47# _316_/a_639_47# 0.0138f
C11483 _316_/a_193_47# _316_/a_1217_47# 2.36e-20
C11484 _316_/a_761_289# _316_/a_805_47# 3.69e-19
C11485 _050_ _052_ 0.349f
C11486 _195_/a_76_199# _062_ 0.109f
C11487 _322_/a_448_47# net53 5.51e-21
C11488 net34 net40 0.002f
C11489 net5 net40 1.96e-19
C11490 VPWR _303_/a_1462_47# 2.56e-19
C11491 _040_ _049_ 2.28e-19
C11492 net50 _335_/a_805_47# 2.13e-19
C11493 mask\[3\] mask\[1\] 9.14e-20
C11494 net23 net15 0.00814f
C11495 _090_ _243_/a_27_297# 8.83e-19
C11496 _229_/a_27_297# _100_ 0.0509f
C11497 clknet_2_1__leaf_clk _312_/a_27_47# 0.303f
C11498 net44 _319_/a_1283_21# 1.61e-19
C11499 _110_ net9 0.138f
C11500 en_co_clk _332_/a_1283_21# 3.21e-19
C11501 net22 _138_/a_27_47# 0.0015f
C11502 _308_/a_1283_21# clknet_2_0__leaf_clk 1.65e-19
C11503 net30 _279_/a_396_47# 0.00106f
C11504 _326_/a_761_289# net43 0.175f
C11505 clknet_0_clk clone7/a_27_47# 4.43e-21
C11506 _330_/a_1270_413# net46 8.41e-20
C11507 _336_/a_448_47# _119_ 0.0083f
C11508 _323_/a_193_47# clknet_2_1__leaf_clk 0.00196f
C11509 _338_/a_796_47# _065_ 1.61e-20
C11510 net18 _278_/a_109_297# 1.3e-20
C11511 _267_/a_59_75# net46 2.04e-20
C11512 _341_/a_1283_21# _135_ 1.09e-19
C11513 _337_/a_27_47# _282_/a_68_297# 6.09e-19
C11514 _015_ _243_/a_109_297# 0.00189f
C11515 _198_/a_27_47# _067_ 0.248f
C11516 _251_/a_109_47# _101_ 0.00145f
C11517 _251_/a_27_297# net52 0.245f
C11518 _306_/a_1270_413# _092_ 5.17e-21
C11519 output10/a_27_47# _275_/a_81_21# 8.07e-20
C11520 _198_/a_27_47# _070_ 0.089f
C11521 net27 mask\[2\] 4.53e-21
C11522 VPWR _008_ 0.534f
C11523 _320_/a_639_47# clknet_2_0__leaf_clk 3.68e-19
C11524 trimb[0] net34 0.0659f
C11525 _299_/a_298_297# net40 0.00128f
C11526 _315_/a_27_47# _241_/a_105_352# 2.24e-21
C11527 trim_mask\[2\] net33 0.00626f
C11528 net9 net47 0.131f
C11529 _249_/a_109_47# net26 0.00123f
C11530 _232_/a_220_297# _090_ 0.0146f
C11531 _328_/a_1108_47# trim_mask\[1\] 0.049f
C11532 _102_ mask\[6\] 0.00305f
C11533 trim_mask\[2\] trim_mask\[1\] 0.0266f
C11534 _244_/a_27_297# _076_ 2.71e-19
C11535 _200_/a_209_297# _071_ 4.88e-19
C11536 _319_/a_543_47# _016_ 0.00139f
C11537 VPWR _246_/a_109_297# 0.196f
C11538 net9 _340_/a_1140_413# 1.65e-19
C11539 _253_/a_81_21# _078_ 0.011f
C11540 net4 _066_ 2.22e-19
C11541 _095_ _049_ 0.0214f
C11542 _289_/a_68_297# _297_/a_47_47# 4.35e-19
C11543 trim_mask\[2\] _336_/a_761_289# 1.41e-21
C11544 _008_ net53 0.028f
C11545 _307_/a_639_47# _074_ 0.00166f
C11546 _140_/a_68_297# net45 3.35e-20
C11547 trim_mask\[0\] _106_ 0.152f
C11548 _149_/a_68_297# _149_/a_150_297# 0.00477f
C11549 output26/a_27_47# net25 3.74e-20
C11550 _334_/a_193_47# _334_/a_651_413# 0.0346f
C11551 _334_/a_543_47# _334_/a_1108_47# 7.99e-20
C11552 trim[3] net46 1.66e-19
C11553 _314_/a_193_47# _314_/a_1270_413# 1.46e-19
C11554 _314_/a_27_47# _314_/a_639_47# 0.00188f
C11555 _314_/a_543_47# _314_/a_448_47# 0.0498f
C11556 _314_/a_761_289# _314_/a_651_413# 0.0977f
C11557 _314_/a_1283_21# _314_/a_1108_47# 0.234f
C11558 VPWR _199_/a_109_297# 0.00273f
C11559 VPWR mask\[5\] 1.68f
C11560 _326_/a_639_47# net28 1.7e-19
C11561 _228_/a_297_47# _052_ 0.0542f
C11562 _327_/a_193_47# _327_/a_543_47# 0.23f
C11563 _327_/a_27_47# _327_/a_1283_21# 0.0435f
C11564 _164_/a_161_47# net15 0.00151f
C11565 net12 _021_ 7.98e-19
C11566 ctln[5] _330_/a_448_47# 4.12e-20
C11567 net2 _339_/a_1032_413# 2.56e-20
C11568 _308_/a_193_47# _319_/a_193_47# 0.00148f
C11569 _168_/a_207_413# _331_/a_193_47# 2.79e-21
C11570 _029_ _109_ 7.06e-19
C11571 mask\[5\] net53 0.188f
C11572 _185_/a_68_297# net54 0.167f
C11573 _336_/a_651_413# _266_/a_68_297# 4.89e-21
C11574 _060_ _075_ 0.245f
C11575 _299_/a_215_297# _299_/a_298_297# 0.0718f
C11576 mask\[7\] _313_/a_27_47# 6.7e-19
C11577 _304_/a_193_47# _298_/a_78_199# 4.02e-20
C11578 VPWR _291_/a_35_297# 0.179f
C11579 _327_/a_543_47# _058_ 0.0112f
C11580 clknet_0_clk _073_ 5.34e-22
C11581 net46 net37 1.7e-19
C11582 _259_/a_109_297# trim_mask\[4\] 0.00151f
C11583 _320_/a_1108_47# clknet_2_1__leaf_clk 6.67e-22
C11584 _104_ _260_/a_93_21# 0.0789f
C11585 _041_ _067_ 2.26e-20
C11586 clone1/a_27_47# _242_/a_297_47# 0.0382f
C11587 net3 output41/a_27_47# 9.02e-19
C11588 VPWR _019_ 0.476f
C11589 _304_/a_651_413# _122_ 0.00442f
C11590 _041_ _070_ 6.58e-20
C11591 _034_ net30 0.0547f
C11592 _072_ _201_/a_113_47# 0.0096f
C11593 mask\[5\] _009_ 1.37e-19
C11594 _333_/a_1283_21# _056_ 1.36e-20
C11595 _115_ net33 1.51e-21
C11596 _106_ _191_/a_27_297# 5e-19
C11597 _021_ net44 0.0069f
C11598 mask\[6\] _312_/a_193_47# 3.48e-20
C11599 _112_ _333_/a_27_47# 0.0184f
C11600 trim_val\[1\] _333_/a_543_47# 0.00171f
C11601 net49 _333_/a_193_47# 0.0129f
C11602 trim_mask\[1\] _333_/a_761_289# 7.01e-19
C11603 _115_ trim_mask\[1\] 1.95e-19
C11604 _133_ net40 0.00147f
C11605 _260_/a_93_21# net55 3.94e-21
C11606 net35 _058_ 0.00401f
C11607 _298_/a_78_199# _298_/a_493_297# 3.15e-19
C11608 _310_/a_27_47# _310_/a_193_47# 0.887f
C11609 _042_ net19 0.0106f
C11610 _316_/a_448_47# _013_ 0.167f
C11611 _200_/a_80_21# _053_ 0.0384f
C11612 _019_ net53 0.00889f
C11613 _127_ _297_/a_285_47# 7.44e-21
C11614 _329_/a_1108_47# _274_/a_75_212# 0.00253f
C11615 _064_ net19 4.18e-20
C11616 _327_/a_27_47# _108_ 0.03f
C11617 _306_/a_1283_21# _048_ 3.18e-20
C11618 _323_/a_1270_413# _042_ 3.5e-19
C11619 _309_/a_448_47# _074_ 0.0102f
C11620 _159_/a_27_47# _313_/a_761_289# 0.00138f
C11621 net54 _088_ 6.12e-21
C11622 _335_/a_193_47# _335_/a_543_47# 0.23f
C11623 _335_/a_27_47# _335_/a_1283_21# 0.0436f
C11624 _059_ en_co_clk 0.091f
C11625 _033_ _119_ 0.728f
C11626 _262_/a_27_47# _092_ 8.22e-20
C11627 net10 trim_mask\[3\] 0.00217f
C11628 _074_ _249_/a_27_297# 4.66e-19
C11629 net28 _086_ 0.106f
C11630 net35 _332_/a_27_47# 7.94e-19
C11631 _058_ _332_/a_761_289# 0.00357f
C11632 fanout43/a_27_47# mask\[1\] 0.0536f
C11633 net9 _301_/a_47_47# 4.82e-20
C11634 _303_/a_1108_47# net2 4.77e-21
C11635 _334_/a_805_47# net46 0.0036f
C11636 VPWR _208_/a_218_47# 2.26e-19
C11637 _315_/a_1283_21# _099_ 3e-19
C11638 _315_/a_1108_47# _095_ 7.61e-19
C11639 net27 _314_/a_193_47# 8.02e-20
C11640 _327_/a_1270_413# net46 3.35e-19
C11641 cal_itt\[0\] _068_ 0.0535f
C11642 _129_ _298_/a_78_199# 1.27e-19
C11643 _299_/a_215_297# _133_ 4.06e-19
C11644 net9 _341_/a_27_47# 0.00101f
C11645 _336_/a_543_47# trim_mask\[4\] 0.0358f
C11646 _064_ _107_ 0.00119f
C11647 VPWR _017_ 0.42f
C11648 _329_/a_27_47# trim_mask\[4\] 4.49e-19
C11649 _329_/a_1108_47# clknet_2_2__leaf_clk 0.00393f
C11650 clkbuf_0_clk/a_110_47# fanout47/a_27_47# 2.1e-19
C11651 _304_/a_27_47# _304_/a_1217_47# 2.56e-19
C11652 _304_/a_761_289# _304_/a_639_47# 3.16e-19
C11653 _126_ _297_/a_285_47# 2.58e-20
C11654 net14 sample 8.01e-20
C11655 _047_ _055_ 3.3e-20
C11656 _230_/a_59_75# _091_ 0.128f
C11657 _339_/a_1032_413# _123_ 0.0695f
C11658 _048_ _227_/a_368_53# 3.75e-19
C11659 net43 _305_/a_761_289# 0.203f
C11660 trim[1] _162_/a_27_47# 6.46e-19
C11661 _329_/a_805_47# trim_mask\[2\] 9.76e-20
C11662 clk _316_/a_27_47# 2.74e-19
C11663 _107_ _100_ 0.0129f
C11664 input1/a_75_212# net1 0.11f
C11665 _332_/a_27_47# _332_/a_761_289# 0.0623f
C11666 rebuffer1/a_75_212# _108_ 0.188f
C11667 _059_ _050_ 0.239f
C11668 _327_/a_448_47# _327_/a_639_47# 4.61e-19
C11669 net12 clone7/a_27_47# 1.4e-20
C11670 _264_/a_27_297# net19 2.68e-19
C11671 _335_/a_1270_413# net46 2.76e-19
C11672 _048_ _317_/a_1283_21# 1.69e-19
C11673 VPWR _226_/a_197_47# 2.43e-19
C11674 _093_ _092_ 1.08e-19
C11675 _169_/a_215_311# state\[0\] 0.216f
C11676 _168_/a_207_413# _260_/a_93_21# 0.016f
C11677 ctlp[7] _074_ 0.0518f
C11678 net51 rebuffer4/a_27_47# 0.111f
C11679 net43 clkbuf_2_0__f_clk/a_110_47# 4.53e-20
C11680 output37/a_27_47# _126_ 0.0104f
C11681 _304_/a_543_47# clknet_2_3__leaf_clk 0.00312f
C11682 _082_ _247_/a_27_297# 1.82e-20
C11683 _333_/a_1283_21# _173_/a_27_47# 4.74e-19
C11684 _340_/a_1182_261# _298_/a_78_199# 0.00134f
C11685 net9 clknet_2_2__leaf_clk 0.185f
C11686 _309_/a_543_47# clknet_2_1__leaf_clk 5.3e-20
C11687 _078_ net21 0.427f
C11688 _074_ _220_/a_113_297# 3.15e-19
C11689 _294_/a_150_297# net33 3.68e-19
C11690 net13 _042_ 0.0188f
C11691 VPWR _330_/a_651_413# 0.145f
C11692 net24 _006_ 0.0752f
C11693 result[2] _081_ 5.8e-19
C11694 _257_/a_27_297# _336_/a_27_47# 6.17e-21
C11695 _332_/a_651_413# net46 0.0388f
C11696 _136_ clkc 5.39e-20
C11697 _207_/a_109_297# _049_ 0.00121f
C11698 _237_/a_505_21# _096_ 0.247f
C11699 _304_/a_1270_413# _035_ 1.07e-21
C11700 wire42/a_75_212# _092_ 0.00229f
C11701 net47 _122_ 0.1f
C11702 _048_ _192_/a_174_21# 0.0772f
C11703 output38/a_27_47# net16 0.00105f
C11704 _306_/a_1108_47# _050_ 5.7e-20
C11705 _325_/a_193_47# net26 4.29e-20
C11706 _053_ net46 6.57e-19
C11707 _336_/a_805_47# _107_ 1.48e-19
C11708 _264_/a_27_297# _107_ 0.0841f
C11709 _340_/a_1140_413# _122_ 2.73e-19
C11710 _064_ _279_/a_27_47# 1.42e-20
C11711 VPWR _200_/a_80_21# 0.17f
C11712 _337_/a_1283_21# clknet_0_clk 2.34e-19
C11713 _326_/a_1108_47# _325_/a_27_47# 3.16e-20
C11714 _310_/a_543_47# _310_/a_639_47# 0.0138f
C11715 _310_/a_193_47# _310_/a_1217_47# 2.36e-20
C11716 _310_/a_761_289# _310_/a_805_47# 3.69e-19
C11717 net13 _100_ 0.00763f
C11718 net28 clknet_2_1__leaf_clk 0.242f
C11719 _071_ _053_ 0.00497f
C11720 _116_ clkbuf_2_2__f_clk/a_110_47# 3.83e-19
C11721 _307_/a_193_47# net22 0.21f
C11722 _307_/a_27_47# mask\[0\] 0.0111f
C11723 _059_ _228_/a_297_47# 8.65e-21
C11724 _186_/a_109_297# _088_ 9.11e-21
C11725 _327_/a_1217_47# _108_ 3.22e-20
C11726 VPWR _325_/a_1270_413# 8.1e-19
C11727 net21 _313_/a_651_413# 2.12e-19
C11728 _335_/a_448_47# _335_/a_639_47# 4.61e-19
C11729 net16 _333_/a_448_47# 0.00323f
C11730 _324_/a_448_47# clknet_2_1__leaf_clk 8.22e-19
C11731 _340_/a_652_21# _129_ 2.33e-21
C11732 clknet_2_1__leaf_clk _158_/a_68_297# 0.00905f
C11733 net26 _076_ 0.00189f
C11734 _226_/a_27_47# _049_ 6.98e-19
C11735 _035_ clknet_2_3__leaf_clk 0.107f
C11736 _322_/a_1283_21# _250_/a_27_297# 9.71e-22
C11737 clk _003_ 2.86e-19
C11738 _311_/a_27_47# _311_/a_1108_47# 0.102f
C11739 _311_/a_193_47# _311_/a_1283_21# 0.0424f
C11740 _311_/a_761_289# _311_/a_543_47# 0.21f
C11741 _042_ _248_/a_109_297# 3.94e-19
C11742 _322_/a_193_47# _042_ 7.52e-20
C11743 net12 _073_ 0.00478f
C11744 en_co_clk _192_/a_27_47# 0.00756f
C11745 _304_/a_761_289# _136_ 0.00121f
C11746 _064_ _257_/a_109_297# 0.0165f
C11747 cal_itt\[2\] _306_/a_193_47# 8.89e-21
C11748 _322_/a_1108_47# clknet_2_1__leaf_clk 1.12e-19
C11749 _227_/a_209_311# _062_ 1.75e-20
C11750 _106_ trim_mask\[4\] 1.48e-20
C11751 _304_/a_1283_21# net47 0.286f
C11752 _096_ _241_/a_297_47# 7.33e-19
C11753 _326_/a_27_47# _314_/a_193_47# 3.41e-19
C11754 _326_/a_193_47# _314_/a_27_47# 7.79e-19
C11755 _336_/a_27_47# trim_val\[4\] 6.67e-19
C11756 VPWR _314_/a_1283_21# 0.408f
C11757 _187_/a_297_47# en_co_clk 6.97e-19
C11758 _264_/a_27_297# _279_/a_27_47# 6.6e-19
C11759 result[3] clknet_2_1__leaf_clk 0.0234f
C11760 _308_/a_1108_47# mask\[0\] 0.00229f
C11761 _308_/a_1283_21# _078_ 0.00166f
C11762 _321_/a_27_47# _321_/a_1217_47# 2.56e-19
C11763 _321_/a_761_289# _321_/a_639_47# 3.16e-19
C11764 output15/a_27_47# net28 2.54e-19
C11765 net43 _042_ 0.377f
C11766 _332_/a_805_47# _108_ 6.71e-19
C11767 _340_/a_27_47# _340_/a_1602_47# 4.5e-20
C11768 _340_/a_193_47# _340_/a_1032_413# 0.0573f
C11769 _332_/a_1108_47# _332_/a_1270_413# 0.00645f
C11770 _332_/a_761_289# _332_/a_1217_47# 4.2e-19
C11771 _332_/a_543_47# _332_/a_805_47# 0.00171f
C11772 _074_ _213_/a_109_297# 0.0012f
C11773 _228_/a_297_47# _170_/a_384_47# 2.15e-20
C11774 net44 _073_ 6.49e-20
C11775 _136_ _298_/a_215_47# 0.00109f
C11776 _308_/a_193_47# net24 5.52e-22
C11777 _302_/a_109_47# clknet_2_3__leaf_clk 0.00176f
C11778 _136_ clkbuf_2_3__f_clk/a_110_47# 8.86e-19
C11779 ctlp[0] _314_/a_761_289# 9.95e-19
C11780 _164_/a_161_47# state\[1\] 2.13e-19
C11781 net43 _319_/a_448_47# 2.77e-19
C11782 state\[0\] _053_ 0.0174f
C11783 _063_ net40 4.59e-19
C11784 _074_ _222_/a_113_297# 1.18e-19
C11785 _199_/a_193_297# _065_ 0.00156f
C11786 net31 _056_ 9.97e-20
C11787 _050_ _192_/a_27_47# 8.37e-19
C11788 _337_/a_27_47# _337_/a_1217_47# 2.56e-19
C11789 _337_/a_761_289# _337_/a_639_47# 3.16e-19
C11790 _303_/a_1283_21# _069_ 4.45e-19
C11791 _007_ net26 0.00175f
C11792 _037_ net40 3.14e-19
C11793 VPWR _310_/a_27_47# 0.488f
C11794 net13 _022_ 1.44e-20
C11795 _333_/a_639_47# net32 1.09e-19
C11796 _288_/a_145_75# _125_ 5.76e-19
C11797 _340_/a_193_47# cal_count\[3\] 1.07e-20
C11798 net9 _339_/a_956_413# 2.92e-19
C11799 net50 fanout46/a_27_47# 1.66e-20
C11800 VPWR net46 4.73f
C11801 _333_/a_1283_21# _172_/a_68_297# 2.46e-19
C11802 _287_/a_75_212# _338_/a_476_47# 3.15e-19
C11803 clknet_2_1__leaf_clk _246_/a_27_297# 0.00409f
C11804 _341_/a_27_47# _122_ 5.3e-19
C11805 mask\[3\] net26 0.00358f
C11806 _276_/a_145_75# _117_ 5.76e-19
C11807 VPWR _195_/a_439_47# 0.00127f
C11808 _064_ _118_ 0.0875f
C11809 VPWR _071_ 0.473f
C11810 _303_/a_1108_47# _067_ 5.17e-21
C11811 _306_/a_27_47# _244_/a_27_297# 0.0129f
C11812 _338_/a_27_47# net18 0.016f
C11813 _324_/a_1283_21# _021_ 6.94e-21
C11814 _303_/a_1108_47# _070_ 2.47e-19
C11815 _119_ clkbuf_2_3__f_clk/a_110_47# 2.64e-20
C11816 _321_/a_1108_47# _143_/a_68_297# 5.65e-20
C11817 _239_/a_277_297# _092_ 0.0588f
C11818 VPWR _334_/a_639_47# 0.00447f
C11819 _326_/a_1108_47# net25 8.95e-20
C11820 mask\[6\] _158_/a_150_297# 1.07e-19
C11821 clknet_2_0__leaf_clk en_co_clk 0.0128f
C11822 output23/a_27_47# _213_/a_109_297# 5.98e-20
C11823 _307_/a_1462_47# net22 5.12e-19
C11824 VPWR _327_/a_651_413# 0.144f
C11825 _266_/a_68_297# clkbuf_2_2__f_clk/a_110_47# 1.71e-19
C11826 net13 _313_/a_1283_21# 4.31e-19
C11827 _335_/a_639_47# _032_ 3.71e-19
C11828 _189_/a_218_47# _048_ 0.0814f
C11829 _313_/a_1283_21# _155_/a_68_297# 7.54e-19
C11830 _185_/a_150_297# _049_ 3.24e-20
C11831 _302_/a_109_297# _136_ 0.0131f
C11832 _092_ _206_/a_27_93# 5.28e-20
C11833 cal net41 0.0709f
C11834 _307_/a_193_47# _079_ 4.88e-19
C11835 net15 _141_/a_27_47# 0.109f
C11836 trim[4] comp 6.05e-20
C11837 net28 _313_/a_27_47# 0.209f
C11838 _311_/a_1108_47# _311_/a_1217_47# 0.00742f
C11839 _311_/a_1283_21# _311_/a_1462_47# 0.0074f
C11840 output22/a_27_47# _004_ 0.00117f
C11841 _161_/a_68_297# net46 0.00116f
C11842 clknet_0_clk _101_ 0.00175f
C11843 _074_ _212_/a_113_297# 0.0208f
C11844 _064_ _025_ 1.51e-19
C11845 clkbuf_2_0__f_clk/a_110_47# net3 0.0132f
C11846 VPWR _335_/a_651_413# 0.145f
C11847 _313_/a_27_47# _158_/a_68_297# 4.15e-19
C11848 trim[4] _332_/a_1270_413# 9.46e-21
C11849 VPWR output27/a_27_47# 0.329f
C11850 VPWR _311_/a_761_289# 0.215f
C11851 _304_/a_1108_47# _063_ 0.00103f
C11852 net12 _337_/a_1283_21# 8.78e-19
C11853 _167_/a_161_47# clk 0.00238f
C11854 _341_/a_193_47# _304_/a_543_47# 9.04e-20
C11855 _111_ _267_/a_59_75# 0.109f
C11856 _018_ _310_/a_1108_47# 5.62e-19
C11857 _050_ clknet_2_0__leaf_clk 0.115f
C11858 _328_/a_27_47# _256_/a_27_297# 0.0111f
C11859 net9 _131_ 7.01e-21
C11860 net43 _022_ 0.00451f
C11861 output14/a_27_47# net27 2.42e-20
C11862 net17 net18 0.0821f
C11863 _340_/a_381_47# net47 1.05e-20
C11864 _037_ _304_/a_1108_47# 7.95e-20
C11865 _264_/a_27_297# _118_ 0.0112f
C11866 _065_ _208_/a_439_47# 0.00369f
C11867 clknet_2_1__leaf_clk _084_ 0.277f
C11868 _311_/a_761_289# net53 0.00351f
C11869 _097_ _095_ 9.72e-19
C11870 _005_ net22 0.00141f
C11871 _048_ _232_/a_32_297# 4.6e-19
C11872 VPWR _332_/a_448_47# 0.0829f
C11873 cal_itt\[2\] net30 0.00218f
C11874 net31 _173_/a_27_47# 0.00232f
C11875 _052_ _049_ 0.59f
C11876 net2 _076_ 0.44f
C11877 net8 _333_/a_543_47# 9.56e-21
C11878 _136_ cal_count\[3\] 0.258f
C11879 VPWR state\[0\] 1.13f
C11880 _128_ _127_ 0.0211f
C11881 _008_ mask\[6\] 6.33e-21
C11882 net26 _310_/a_1283_21# 6.96e-20
C11883 _149_/a_150_297# net19 4.36e-19
C11884 _253_/a_81_21# mask\[7\] 0.0581f
C11885 _309_/a_651_413# _078_ 0.00281f
C11886 _187_/a_27_413# _058_ 1.98e-20
C11887 _167_/a_161_47# net4 0.0473f
C11888 _144_/a_27_47# _041_ 0.207f
C11889 _323_/a_193_47# _043_ 7e-20
C11890 _110_ _024_ 1.51e-21
C11891 _326_/a_543_47# _310_/a_1108_47# 1.16e-20
C11892 _326_/a_1283_21# _310_/a_1283_21# 1.51e-20
C11893 _326_/a_651_413# _310_/a_193_47# 2.21e-20
C11894 _320_/a_27_47# clknet_0_clk 3.01e-19
C11895 _337_/a_1283_21# net44 0.289f
C11896 _309_/a_1283_21# net24 0.133f
C11897 _041_ clknet_2_3__leaf_clk 0.011f
C11898 _338_/a_1182_261# clknet_2_3__leaf_clk 0.0623f
C11899 result[4] net26 0.00579f
C11900 VPWR _310_/a_1217_47# 5.52e-20
C11901 calibrate _228_/a_79_21# 0.0432f
C11902 _068_ net26 3.89e-20
C11903 clknet_2_1__leaf_clk _208_/a_535_374# 3.1e-19
C11904 _233_/a_109_297# input1/a_75_212# 7.12e-21
C11905 net54 _192_/a_174_21# 0.0437f
C11906 net30 _137_/a_150_297# 1.66e-19
C11907 state\[2\] _098_ 0.0595f
C11908 _058_ _268_/a_75_212# 0.00368f
C11909 output36/a_27_47# trimb[2] 0.00188f
C11910 trimb[0] output38/a_27_47# 6.66e-20
C11911 net43 _313_/a_1283_21# 0.27f
C11912 mask\[6\] mask\[5\] 0.017f
C11913 net31 _127_ 3.67e-20
C11914 _078_ _045_ 7.44e-19
C11915 _141_/a_27_47# _049_ 4.22e-19
C11916 _078_ _249_/a_109_297# 1.15e-19
C11917 _293_/a_384_47# _126_ 2.2e-20
C11918 result[5] net29 6.48e-20
C11919 _232_/a_114_297# en_co_clk 4.78e-19
C11920 trim[0] net16 3.49e-20
C11921 _189_/a_408_47# _050_ 0.042f
C11922 _306_/a_448_47# net51 6.51e-21
C11923 en_co_clk net33 4.99e-19
C11924 _321_/a_651_413# _101_ 8.49e-19
C11925 _341_/a_27_47# _091_ 0.00191f
C11926 _119_ cal_count\[3\] 3.29e-21
C11927 _128_ _126_ 3.32e-19
C11928 state\[2\] clknet_0_clk 5.82e-21
C11929 _134_ _299_/a_382_47# 5.12e-19
C11930 _306_/a_761_289# rebuffer6/a_27_47# 3.83e-20
C11931 cal_itt\[2\] _072_ 0.145f
C11932 _300_/a_47_47# net46 6.86e-20
C11933 cal_itt\[0\] cal_itt\[3\] 0.00179f
C11934 _268_/a_75_212# _332_/a_27_47# 5.61e-20
C11935 _337_/a_1283_21# _263_/a_79_21# 7.38e-22
C11936 _104_ _048_ 0.0872f
C11937 _136_ _038_ 0.0457f
C11938 state\[0\] _318_/a_27_47# 0.00104f
C11939 _291_/a_285_297# _289_/a_68_297# 6.54e-21
C11940 clk _331_/a_543_47# 0.00889f
C11941 _060_ _318_/a_448_47# 3.19e-20
C11942 _019_ mask\[6\] 1.18e-20
C11943 _258_/a_109_47# _280_/a_75_212# 3.49e-20
C11944 _314_/a_193_47# _011_ 0.26f
C11945 _314_/a_543_47# _086_ 9.06e-19
C11946 _066_ _193_/a_109_297# 0.0125f
C11947 net12 _331_/a_761_289# 7.17e-20
C11948 net28 _313_/a_1217_47# 8.92e-19
C11949 net31 _126_ 0.00137f
C11950 _311_/a_448_47# net26 0.0163f
C11951 _078_ mask\[4\] 0.174f
C11952 net27 net26 1.42e-19
C11953 net4 _280_/a_75_212# 3.38e-19
C11954 _064_ _330_/a_761_289# 1.87e-21
C11955 _104_ _330_/a_27_47# 3.03e-20
C11956 _306_/a_27_47# _306_/a_1283_21# 0.0436f
C11957 _306_/a_193_47# _306_/a_543_47# 0.23f
C11958 _303_/a_1283_21# fanout47/a_27_47# 0.0139f
C11959 cal_itt\[2\] _305_/a_193_47# 0.00182f
C11960 _074_ _314_/a_448_47# 1.14e-19
C11961 _048_ net55 0.907f
C11962 _329_/a_1108_47# trim_mask\[3\] 1.06e-19
C11963 _326_/a_761_289# result[5] 9.44e-20
C11964 net3 _100_ 3.82e-21
C11965 _331_/a_27_47# _331_/a_651_413# 9.73e-19
C11966 _331_/a_761_289# _331_/a_1108_47# 0.0512f
C11967 _331_/a_193_47# _331_/a_448_47# 0.0612f
C11968 _169_/a_215_311# calibrate 1.25e-21
C11969 _097_ _164_/a_161_47# 0.00108f
C11970 _245_/a_27_297# _101_ 0.142f
C11971 _325_/a_1108_47# _250_/a_109_297# 7.36e-20
C11972 net4 _198_/a_181_47# 4.12e-19
C11973 _029_ net46 0.0415f
C11974 clknet_2_1__leaf_clk _085_ 0.196f
C11975 _321_/a_1283_21# _320_/a_543_47# 1.26e-21
C11976 _002_ rebuffer5/a_161_47# 2.85e-20
C11977 _256_/a_109_297# clknet_2_2__leaf_clk 0.00629f
C11978 _078_ _220_/a_199_47# 1.28e-19
C11979 _325_/a_543_47# _042_ 0.00153f
C11980 net25 _146_/a_68_297# 0.12f
C11981 net4 _331_/a_543_47# 1.41e-19
C11982 net47 _338_/a_1032_413# 0.245f
C11983 _338_/a_27_47# _338_/a_652_21# 0.185f
C11984 _258_/a_27_297# _258_/a_373_47# 0.0134f
C11985 output40/a_27_47# trimb[4] 0.337f
C11986 VPWR output10/a_27_47# 0.297f
C11987 cal _315_/a_193_47# 0.00305f
C11988 net1 _315_/a_27_47# 4.25e-19
C11989 _169_/a_215_311# net45 2.97e-19
C11990 net39 net34 0.147f
C11991 _325_/a_651_413# clknet_2_1__leaf_clk 5.87e-19
C11992 _074_ _310_/a_761_289# 0.0091f
C11993 net47 _297_/a_285_47# 1.15e-19
C11994 _340_/a_562_413# _037_ 1.08e-19
C11995 _326_/a_27_47# output14/a_27_47# 4.86e-21
C11996 net23 result[2] 4.23e-19
C11997 _051_ _331_/a_639_47# 2.63e-19
C11998 _050_ clone1/a_27_47# 0.00933f
C11999 _120_ net55 2.09e-21
C12000 net31 _172_/a_68_297# 0.0148f
C12001 trim_mask\[3\] net9 0.0183f
C12002 _061_ net35 0.0122f
C12003 net12 _101_ 0.0151f
C12004 _341_/a_761_289# cal_count\[3\] 0.0186f
C12005 _338_/a_1296_47# clknet_2_3__leaf_clk 3.98e-19
C12006 _135_ net37 1.53e-20
C12007 _341_/a_651_413# clknet_2_3__leaf_clk 0.00499f
C12008 _012_ input1/a_75_212# 5.56e-21
C12009 _074_ cal 0.00431f
C12010 _198_/a_181_47# _063_ 1.28e-19
C12011 _320_/a_193_47# _143_/a_68_297# 0.00162f
C12012 _015_ _051_ 0.0399f
C12013 _078_ _020_ 3.53e-21
C12014 clkbuf_2_2__f_clk/a_110_47# _279_/a_314_297# 1.04e-20
C12015 VPWR _306_/a_651_413# 0.143f
C12016 net31 output5/a_27_47# 0.00676f
C12017 net9 _001_ 0.00129f
C12018 trim_mask\[1\] _334_/a_193_47# 1.13e-20
C12019 trim_mask\[0\] _301_/a_285_47# 1.56e-19
C12020 output15/a_27_47# _085_ 0.0257f
C12021 _272_/a_81_21# _334_/a_27_47# 4.16e-20
C12022 _340_/a_1032_413# _339_/a_27_47# 4.51e-20
C12023 _340_/a_1182_261# _339_/a_193_47# 1.55e-19
C12024 _340_/a_652_21# _339_/a_476_47# 4.14e-22
C12025 _340_/a_476_47# _339_/a_652_21# 4.26e-20
C12026 _340_/a_27_47# _339_/a_1032_413# 2.42e-20
C12027 _168_/a_207_413# _048_ 2.41e-23
C12028 _307_/a_761_289# net14 0.00982f
C12029 clknet_2_1__leaf_clk _314_/a_543_47# 6.19e-19
C12030 cal _014_ 3e-20
C12031 net1 clknet_2_0__leaf_clk 1.47e-19
C12032 _051_ _242_/a_79_21# 2.03e-20
C12033 _307_/a_1283_21# _138_/a_27_47# 0.00116f
C12034 _326_/a_761_289# net29 7.76e-20
C12035 mask\[1\] _319_/a_1283_21# 9.46e-20
C12036 _227_/a_109_93# _227_/a_296_53# 1.84e-19
C12037 _122_ _131_ 0.0065f
C12038 _043_ _303_/a_27_47# 0.00115f
C12039 _064_ _062_ 0.516f
C12040 net44 _101_ 0.158f
C12041 _029_ _332_/a_448_47# 0.158f
C12042 clknet_2_1__leaf_clk rebuffer4/a_27_47# 0.012f
C12043 _059_ _049_ 0.00658f
C12044 _144_/a_27_47# _339_/a_1032_413# 4.27e-19
C12045 clknet_2_0__leaf_clk _039_ 0.00324f
C12046 _169_/a_109_53# _243_/a_27_297# 6.94e-21
C12047 net12 _320_/a_27_47# 1.15e-21
C12048 net2 _068_ 0.00928f
C12049 _047_ _333_/a_1283_21# 0.0012f
C12050 _323_/a_651_413# net47 0.0122f
C12051 trim_mask\[2\] _119_ 0.104f
C12052 _312_/a_1108_47# net20 0.00215f
C12053 _322_/a_27_47# clknet_0_clk 1.13e-19
C12054 _299_/a_27_413# _131_ 0.253f
C12055 _299_/a_382_47# cal_count\[2\] 8.88e-19
C12056 _305_/a_1283_21# _068_ 6.01e-19
C12057 _259_/a_373_47# net46 1.02e-19
C12058 _306_/a_448_47# _306_/a_639_47# 4.61e-19
C12059 _076_ _070_ 2.23e-20
C12060 cal_itt\[2\] _305_/a_1462_47# 8.36e-19
C12061 _326_/a_27_47# net26 0.00144f
C12062 _341_/a_761_289# _038_ 0.00104f
C12063 _341_/a_448_47# _136_ 0.00158f
C12064 _331_/a_761_289# clknet_2_2__leaf_clk 1.82e-19
C12065 _331_/a_193_47# _028_ 0.547f
C12066 _064_ _195_/a_76_199# 1.78e-19
C12067 net7 _317_/a_543_47# 1.06e-19
C12068 net15 _317_/a_1108_47# 0.0035f
C12069 state\[0\] _093_ 0.0554f
C12070 _053_ calibrate 0.145f
C12071 _074_ net51 5.04e-19
C12072 _326_/a_1108_47# net15 2.21e-20
C12073 _325_/a_543_47# _022_ 5.3e-19
C12074 _317_/a_193_47# _317_/a_543_47# 0.217f
C12075 _317_/a_27_47# _317_/a_1283_21# 0.0435f
C12076 _325_/a_1108_47# _021_ 1.91e-20
C12077 clk net19 0.039f
C12078 _233_/a_27_297# net41 2.45e-20
C12079 _258_/a_27_297# clknet_2_2__leaf_clk 0.0569f
C12080 _326_/a_27_47# _326_/a_1283_21# 0.0436f
C12081 _326_/a_193_47# _326_/a_543_47# 0.23f
C12082 VPWR ctlp[6] 0.774f
C12083 _325_/a_27_47# _078_ 0.0104f
C12084 _024_ clknet_2_2__leaf_clk 0.153f
C12085 net54 _232_/a_32_297# 0.172f
C12086 _082_ _042_ 0.00156f
C12087 _308_/a_651_413# net14 0.00291f
C12088 mask\[0\] _120_ 0.00193f
C12089 trim_val\[1\] rebuffer1/a_75_212# 8.86e-20
C12090 _338_/a_27_47# _338_/a_1056_47# 0.00248f
C12091 _328_/a_193_47# _328_/a_1108_47# 0.119f
C12092 _328_/a_27_47# _328_/a_448_47# 0.0902f
C12093 VPWR _317_/a_651_413# 0.133f
C12094 state\[2\] net12 0.261f
C12095 _104_ _327_/a_27_47# 7.3e-20
C12096 VPWR _326_/a_651_413# 0.145f
C12097 _320_/a_27_47# net44 0.296f
C12098 _290_/a_297_47# net37 0.00147f
C12099 _053_ net45 5.85e-20
C12100 cal_count\[1\] _122_ 0.201f
C12101 output29/a_27_47# _314_/a_1283_21# 5.15e-19
C12102 _277_/a_75_212# net19 2.95e-21
C12103 _053_ rebuffer3/a_75_212# 1.3e-19
C12104 _089_ _090_ 0.205f
C12105 _313_/a_27_47# _085_ 0.00843f
C12106 net13 _337_/a_448_47# 0.00342f
C12107 state\[2\] _331_/a_1108_47# 6.44e-20
C12108 net21 _312_/a_27_47# 2.25e-21
C12109 output35/a_27_47# net2 4.69e-19
C12110 _170_/a_81_21# _054_ 0.119f
C12111 _170_/a_384_47# _049_ 0.0101f
C12112 _273_/a_59_75# _273_/a_145_75# 0.00658f
C12113 net30 _170_/a_81_21# 2.4e-19
C12114 _040_ _337_/a_543_47# 8.12e-20
C12115 _250_/a_27_297# _311_/a_27_47# 1.96e-20
C12116 net4 net19 0.346f
C12117 clk _107_ 0.0308f
C12118 VPWR _192_/a_476_47# 1.11e-19
C12119 cal_count\[1\] _299_/a_27_413# 4.98e-21
C12120 _104_ _335_/a_27_47# 1.78e-19
C12121 _272_/a_384_47# net46 1.37e-19
C12122 net44 _312_/a_448_47# 5.97e-19
C12123 _312_/a_193_47# _312_/a_543_47# 0.23f
C12124 _312_/a_27_47# _312_/a_1283_21# 0.0435f
C12125 _168_/a_297_47# _050_ 0.00186f
C12126 _033_ _330_/a_448_47# 6.61e-19
C12127 _336_/a_1108_47# net46 0.223f
C12128 _053_ _065_ 0.352f
C12129 ctlp[6] _009_ 2.05e-20
C12130 _286_/a_76_199# _286_/a_218_374# 0.00557f
C12131 _214_/a_113_297# _214_/a_199_47# 2.42e-19
C12132 _320_/a_193_47# net52 0.00316f
C12133 net24 _017_ 0.00128f
C12134 clknet_2_1__leaf_clk _311_/a_193_47# 0.00421f
C12135 _329_/a_543_47# _027_ 1.42e-20
C12136 _329_/a_761_289# net46 0.166f
C12137 _323_/a_651_413# net44 5.32e-19
C12138 _303_/a_1108_47# clknet_2_3__leaf_clk 0.0604f
C12139 _320_/a_1283_21# _041_ 1.05e-19
C12140 net47 _339_/a_1602_47# 0.00217f
C12141 _305_/a_448_47# net51 0.00158f
C12142 _092_ net18 4.21e-19
C12143 net2 _125_ 0.0333f
C12144 _114_ _334_/a_761_289# 0.00204f
C12145 trim_val\[2\] _334_/a_1108_47# 0.00214f
C12146 _323_/a_193_47# _323_/a_1108_47# 0.119f
C12147 _323_/a_27_47# _323_/a_448_47# 0.0931f
C12148 net13 _143_/a_68_297# 9.7e-19
C12149 _200_/a_209_47# _106_ 1.13e-19
C12150 _053_ _105_ 0.154f
C12151 VPWR _315_/a_761_289# 0.222f
C12152 net4 _107_ 0.0857f
C12153 _306_/a_1283_21# cal_itt\[3\] 0.0644f
C12154 _306_/a_543_47# _072_ 1.35e-19
C12155 _104_ net54 0.00148f
C12156 _337_/a_193_47# _092_ 5.56e-19
C12157 _337_/a_543_47# _095_ 3.65e-19
C12158 net3 _316_/a_193_47# 1.57e-20
C12159 VPWR _111_ 0.369f
C12160 VPWR _318_/a_805_47# 5.1e-19
C12161 net16 _334_/a_1108_47# 2.65e-19
C12162 _063_ net19 0.824f
C12163 _315_/a_761_289# valid 9.39e-19
C12164 _308_/a_543_47# _006_ 8.48e-20
C12165 _308_/a_1108_47# _081_ 3.75e-21
C12166 trim_mask\[0\] _109_ 0.103f
C12167 state\[2\] _263_/a_79_21# 7.14e-20
C12168 _060_ _096_ 0.0589f
C12169 net54 net55 0.395f
C12170 _049_ _203_/a_59_75# 7.54e-22
C12171 _306_/a_543_47# _305_/a_193_47# 0.00115f
C12172 _306_/a_1283_21# _305_/a_27_47# 9.58e-19
C12173 net13 clk 0.015f
C12174 _302_/a_27_297# _092_ 0.0688f
C12175 net43 _321_/a_448_47# 0.0251f
C12176 _324_/a_27_47# net20 0.0134f
C12177 _320_/a_27_47# _320_/a_543_47# 0.11f
C12178 _320_/a_193_47# _320_/a_761_289# 0.181f
C12179 _293_/a_299_297# _144_/a_27_47# 3.09e-19
C12180 _192_/a_27_47# _049_ 0.00826f
C12181 VPWR calibrate 4.54f
C12182 _208_/a_76_199# _003_ 4.11e-20
C12183 output24/a_27_47# _007_ 4.85e-19
C12184 _301_/a_47_47# _134_ 0.0393f
C12185 _048_ _121_ 1.12e-20
C12186 ctlp[0] _225_/a_109_297# 4.39e-19
C12187 output14/a_27_47# _011_ 1.29e-19
C12188 _331_/a_1462_47# _028_ 2.52e-19
C12189 en_co_clk _316_/a_1283_21# 3.25e-21
C12190 clknet_2_2__leaf_clk _260_/a_250_297# 1.54e-21
C12191 _028_ _260_/a_93_21# 0.0854f
C12192 _101_ _209_/a_27_47# 0.0126f
C12193 net15 clknet_2_0__leaf_clk 0.153f
C12194 net35 net16 0.0519f
C12195 _260_/a_250_297# _260_/a_584_47# 2.43e-19
C12196 _317_/a_448_47# _317_/a_639_47# 4.61e-19
C12197 net9 _334_/a_448_47# 3.67e-19
C12198 _341_/a_1108_47# _301_/a_285_47# 3.78e-20
C12199 _328_/a_651_413# clknet_2_2__leaf_clk 0.00165f
C12200 calibrate valid 0.00353f
C12201 _326_/a_448_47# _326_/a_639_47# 4.61e-19
C12202 mask\[3\] mask\[0\] 1.07e-20
C12203 _107_ _063_ 0.019f
C12204 net25 _078_ 0.407f
C12205 _001_ _122_ 0.589f
C12206 _337_/a_1108_47# _034_ 1.97e-19
C12207 _327_/a_1283_21# net9 0.0171f
C12208 net43 net14 2.29f
C12209 VPWR net45 4.53f
C12210 output22/a_27_47# _308_/a_27_47# 0.0131f
C12211 net12 _324_/a_193_47# 3.78e-20
C12212 _341_/a_543_47# _341_/a_1108_47# 7.99e-20
C12213 _341_/a_193_47# _341_/a_651_413# 0.0276f
C12214 VPWR rebuffer3/a_75_212# 0.242f
C12215 net13 net4 0.00859f
C12216 _059_ state\[1\] 0.00785f
C12217 _320_/a_1217_47# net44 6.59e-20
C12218 _053_ _194_/a_113_297# 2.1e-19
C12219 _036_ _035_ 4.23e-21
C12220 net47 _303_/a_448_47# 2.48e-19
C12221 trim_mask\[0\] _279_/a_490_47# 3.36e-19
C12222 _024_ _279_/a_204_297# 6.23e-22
C12223 net4 _279_/a_27_47# 5.29e-20
C12224 net45 valid 3.94e-19
C12225 net47 cal_count\[2\] 0.00129f
C12226 _042_ _247_/a_27_297# 0.0322f
C12227 state\[2\] clknet_2_2__leaf_clk 2.67e-22
C12228 state\[2\] _260_/a_584_47# 0.00134f
C12229 _308_/a_1108_47# _016_ 6.48e-19
C12230 _005_ _245_/a_27_297# 7.7e-20
C12231 net16 _332_/a_761_289# 0.00716f
C12232 _318_/a_193_47# _318_/a_639_47# 2.28e-19
C12233 _318_/a_761_289# _318_/a_1270_413# 2.6e-19
C12234 _318_/a_543_47# _318_/a_651_413# 0.0572f
C12235 _304_/a_1283_21# _231_/a_161_47# 0.00128f
C12236 net12 _322_/a_27_47# 6.71e-21
C12237 _189_/a_27_47# _227_/a_109_93# 2.21e-20
C12238 _125_ _123_ 1.37e-21
C12239 net9 _335_/a_1283_21# 1.72e-19
C12240 _121_ _120_ 0.00179f
C12241 _325_/a_193_47# _010_ 3.98e-19
C12242 VPWR _065_ 3.3f
C12243 _233_/a_109_297# _315_/a_27_47# 1.46e-19
C12244 _233_/a_27_297# _315_/a_193_47# 9.55e-19
C12245 _110_ trim_val\[4\] 0.0123f
C12246 VPWR _135_ 0.394f
C12247 _312_/a_448_47# _312_/a_639_47# 4.61e-19
C12248 _309_/a_193_47# _101_ 2.73e-19
C12249 rstn net6 0.00668f
C12250 _033_ _027_ 2.18e-19
C12251 _324_/a_193_47# net44 0.0485f
C12252 _320_/a_27_47# _209_/a_27_47# 2.73e-21
C12253 _286_/a_218_47# _124_ 2.88e-19
C12254 _286_/a_218_374# cal_count\[0\] 0.00688f
C12255 VPWR _305_/a_651_413# 0.144f
C12256 _068_ _067_ 0.0116f
C12257 _041_ _205_/a_27_47# 0.0753f
C12258 _068_ _070_ 0.0108f
C12259 _308_/a_27_47# _308_/a_1283_21# 0.0436f
C12260 _308_/a_193_47# _308_/a_543_47# 0.23f
C12261 _323_/a_639_47# net19 8.84e-19
C12262 VPWR _105_ 0.27f
C12263 net33 output40/a_27_47# 0.00169f
C12264 _324_/a_27_47# _323_/a_27_47# 8.63e-20
C12265 _065_ net53 1.47e-19
C12266 _291_/a_35_297# _129_ 7.54e-21
C12267 trim_mask\[0\] _092_ 0.00122f
C12268 _002_ net51 0.0071f
C12269 net13 net52 0.0204f
C12270 _107_ _260_/a_346_47# 2.81e-19
C12271 _192_/a_505_280# _192_/a_639_47# 8e-19
C12272 _019_ _321_/a_193_47# 1.38e-19
C12273 net9 _108_ 0.0117f
C12274 net9 _332_/a_543_47# 5.4e-20
C12275 _307_/a_761_289# _307_/a_543_47# 0.21f
C12276 _307_/a_193_47# _307_/a_1283_21# 0.0424f
C12277 _307_/a_27_47# _307_/a_1108_47# 0.102f
C12278 VPWR _259_/a_109_47# 6e-20
C12279 net43 clk 0.00926f
C12280 _037_ _339_/a_381_47# 1.56e-19
C12281 net31 _047_ 0.105f
C12282 result[0] _307_/a_27_47# 0.0108f
C12283 trim[3] _179_/a_27_47# 7.28e-19
C12284 output34/a_27_47# net34 0.22f
C12285 _290_/a_27_413# output40/a_27_47# 0.0126f
C12286 clknet_2_0__leaf_clk _049_ 0.221f
C12287 _041_ _040_ 4.32e-20
C12288 _063_ _279_/a_27_47# 3.67e-19
C12289 VPWR _319_/a_27_47# 0.479f
C12290 _322_/a_27_47# net44 0.301f
C12291 _337_/a_1462_47# _092_ 3.4e-20
C12292 _329_/a_1108_47# _031_ 8.91e-19
C12293 _318_/a_27_47# net45 0.297f
C12294 _233_/a_27_297# _074_ 0.096f
C12295 net3 _316_/a_1462_47# 9.82e-20
C12296 _026_ _327_/a_543_47# 4.33e-20
C12297 net31 _110_ 6.29e-20
C12298 _128_ net47 0.0987f
C12299 net12 _219_/a_109_297# 4.53e-19
C12300 _058_ _172_/a_68_297# 1.31e-19
C12301 VPWR _243_/a_109_297# 0.178f
C12302 _186_/a_109_297# net55 2.48e-19
C12303 clkbuf_2_2__f_clk/a_110_47# _330_/a_1108_47# 0.00167f
C12304 _231_/a_161_47# _091_ 0.222f
C12305 net24 _310_/a_27_47# 2.97e-21
C12306 _303_/a_448_47# net44 4.4e-19
C12307 net43 net4 2.72e-21
C12308 _326_/a_639_47# _074_ 0.00132f
C12309 trim[2] _108_ 4.34e-20
C12310 _309_/a_448_47# _006_ 0.158f
C12311 _309_/a_1270_413# _081_ 2.96e-20
C12312 _323_/a_1283_21# _303_/a_193_47# 3.34e-19
C12313 _323_/a_543_47# _303_/a_761_289# 4.73e-19
C12314 _323_/a_1108_47# _303_/a_27_47# 4.49e-21
C12315 trim_mask\[3\] _256_/a_109_297# 1.18e-20
C12316 net50 _256_/a_27_297# 0.00768f
C12317 _339_/a_27_47# _339_/a_1182_261# 0.0608f
C12318 _339_/a_193_47# _339_/a_476_47# 0.198f
C12319 _248_/a_373_47# _101_ 2.72e-19
C12320 _322_/a_543_47# _101_ 0.00139f
C12321 _322_/a_193_47# net52 5.82e-23
C12322 _088_ clone7/a_27_47# 6.68e-21
C12323 _322_/a_1283_21# _041_ 7.76e-20
C12324 net13 _320_/a_761_289# 0.00446f
C12325 _306_/a_448_47# clknet_2_1__leaf_clk 2.39e-19
C12326 _188_/a_27_47# net37 0.0139f
C12327 VPWR _232_/a_304_297# 0.00452f
C12328 _317_/a_639_47# _014_ 9.32e-19
C12329 _317_/a_1270_413# net45 1.7e-19
C12330 _317_/a_1108_47# state\[1\] 0.00189f
C12331 _187_/a_27_413# _061_ 0.00275f
C12332 net9 _031_ 7.5e-19
C12333 _305_/a_543_47# net30 8.41e-21
C12334 VPWR _194_/a_113_297# 0.235f
C12335 VPWR _112_ 0.709f
C12336 _321_/a_1283_21# mask\[2\] 0.062f
C12337 _271_/a_75_212# _113_ 0.201f
C12338 VPWR _272_/a_299_297# 0.276f
C12339 _315_/a_27_47# _315_/a_1108_47# 0.102f
C12340 _315_/a_193_47# _315_/a_1283_21# 0.0424f
C12341 _315_/a_761_289# _315_/a_543_47# 0.21f
C12342 _189_/a_27_47# _054_ 3.69e-21
C12343 _048_ clknet_2_3__leaf_clk 2.42e-19
C12344 VPWR _336_/a_1283_21# 0.371f
C12345 _189_/a_408_47# _049_ 9.24e-19
C12346 _189_/a_27_47# net30 0.00307f
C12347 _134_ trim_val\[0\] 1.07e-20
C12348 net47 _000_ 0.00829f
C12349 VPWR _329_/a_193_47# 0.612f
C12350 net28 net21 0.0199f
C12351 net8 _334_/a_761_289# 0.00805f
C12352 clkbuf_2_1__f_clk/a_110_47# net30 3.38e-20
C12353 _078_ _039_ 0.2f
C12354 net4 _118_ 0.00759f
C12355 _333_/a_761_289# _333_/a_639_47# 3.16e-19
C12356 _333_/a_27_47# _333_/a_1217_47# 2.56e-19
C12357 _111_ _029_ 0.00664f
C12358 _312_/a_27_47# _045_ 6.75e-19
C12359 net43 net52 0.151f
C12360 fanout43/a_27_47# mask\[0\] 0.00867f
C12361 VPWR _239_/a_27_297# 0.274f
C12362 net43 _063_ 0.00244f
C12363 _249_/a_27_297# _312_/a_193_47# 2.91e-21
C12364 _250_/a_109_297# net26 5.73e-20
C12365 net19 _279_/a_396_47# 0.0147f
C12366 _265_/a_81_21# _109_ 0.125f
C12367 _093_ _315_/a_761_289# 1.4e-19
C12368 calibrate _315_/a_543_47# 0.00737f
C12369 _012_ _315_/a_27_47# 0.17f
C12370 _309_/a_1462_47# _101_ 4.66e-20
C12371 _324_/a_1462_47# net44 0.00323f
C12372 _324_/a_1108_47# _312_/a_1108_47# 4.89e-20
C12373 _334_/a_1283_21# net34 0.0166f
C12374 _257_/a_27_297# clknet_2_2__leaf_clk 0.0282f
C12375 _324_/a_543_47# net19 6.58e-20
C12376 net43 _214_/a_199_47# 1.37e-20
C12377 _308_/a_448_47# _308_/a_639_47# 4.61e-19
C12378 cal_itt\[0\] _122_ 6.25e-20
C12379 net2 cal_itt\[3\] 2.98e-22
C12380 net15 _319_/a_639_47# 7.77e-19
C12381 _232_/a_114_297# _049_ 2.35e-19
C12382 VPWR _289_/a_150_297# 0.00246f
C12383 VPWR output9/a_27_47# 0.268f
C12384 _014_ _315_/a_1283_21# 6.06e-19
C12385 clknet_2_0__leaf_clk _315_/a_1108_47# 0.016f
C12386 _307_/a_1283_21# _307_/a_1462_47# 0.0074f
C12387 _307_/a_1108_47# _307_/a_1217_47# 0.00742f
C12388 net45 _315_/a_543_47# 0.153f
C12389 _192_/a_548_47# _065_ 1.74e-20
C12390 net42 _227_/a_109_93# 2.25e-19
C12391 _090_ _092_ 0.187f
C12392 _326_/a_448_47# clknet_2_1__leaf_clk 0.00313f
C12393 _305_/a_543_47# _072_ 0.00622f
C12394 _305_/a_1283_21# cal_itt\[3\] 1.82e-20
C12395 _074_ _086_ 0.0915f
C12396 _235_/a_382_297# net55 0.00112f
C12397 trim_val\[3\] _280_/a_75_212# 4.87e-21
C12398 net35 net40 0.175f
C12399 _063_ _118_ 0.00299f
C12400 _322_/a_1217_47# net44 0.00148f
C12401 VPWR _319_/a_1217_47# 4.45e-20
C12402 _300_/a_47_47# _135_ 0.149f
C12403 _300_/a_285_47# net2 0.0685f
C12404 _318_/a_1217_47# net45 6.03e-19
C12405 output38/a_27_47# net39 0.0374f
C12406 net3 net14 0.0121f
C12407 _107_ _279_/a_396_47# 0.0111f
C12408 calibrate _093_ 1.41f
C12409 _110_ _330_/a_193_47# 0.00736f
C12410 _336_/a_27_47# net30 6.14e-21
C12411 _189_/a_27_47# _072_ 5.62e-20
C12412 _189_/a_218_47# cal_itt\[3\] 1.94e-19
C12413 _305_/a_27_47# net2 1.9e-19
C12414 net43 _320_/a_761_289# 2.8e-19
C12415 _080_ net14 0.00104f
C12416 output8/a_27_47# _108_ 9.16e-20
C12417 net8 rebuffer1/a_75_212# 4.41e-20
C12418 _036_ _041_ 0.00246f
C12419 trim[4] net32 0.00269f
C12420 _323_/a_193_47# mask\[4\] 0.00152f
C12421 _325_/a_448_47# _321_/a_543_47# 1.3e-20
C12422 _305_/a_27_47# _305_/a_1283_21# 0.0435f
C12423 _305_/a_193_47# _305_/a_543_47# 0.219f
C12424 clone1/a_27_47# _049_ 0.0108f
C12425 _242_/a_297_47# _099_ 4.21e-19
C12426 _000_ net44 0.024f
C12427 _093_ net45 0.0295f
C12428 _012_ clknet_2_0__leaf_clk 0.00553f
C12429 _337_/a_639_47# en_co_clk 4.18e-19
C12430 _262_/a_27_47# _105_ 0.165f
C12431 _303_/a_1270_413# net19 9.48e-20
C12432 _306_/a_27_47# mask\[0\] 4.4e-20
C12433 _332_/a_761_289# net40 3.26e-19
C12434 _033_ _032_ 5.83e-21
C12435 trim_val\[3\] _258_/a_109_297# 3.19e-20
C12436 trim_mask\[3\] _258_/a_27_297# 0.0609f
C12437 _339_/a_652_21# _339_/a_1056_47# 3.94e-19
C12438 _339_/a_476_47# _339_/a_796_47# 0.00184f
C12439 _339_/a_1032_413# _339_/a_1140_413# 0.00523f
C12440 _339_/a_381_47# _339_/a_562_413# 8.75e-19
C12441 _291_/a_35_297# _297_/a_47_47# 1.75e-19
C12442 _055_ _108_ 0.00609f
C12443 _309_/a_1108_47# _140_/a_68_297# 1.48e-19
C12444 _341_/a_1108_47# _092_ 8.65e-22
C12445 clknet_2_0__leaf_clk state\[1\] 0.027f
C12446 _288_/a_59_75# net40 0.00443f
C12447 net43 _307_/a_543_47# 1.29e-20
C12448 _136_ en_co_clk 0.00657f
C12449 _320_/a_805_47# _040_ 0.00239f
C12450 cal_itt\[1\] _304_/a_543_47# 1.58e-19
C12451 net12 _156_/a_27_47# 2.04e-19
C12452 _293_/a_81_21# _339_/a_27_47# 5.65e-20
C12453 _122_ _108_ 4.53e-21
C12454 _315_/a_1108_47# _315_/a_1217_47# 0.00742f
C12455 _315_/a_1283_21# _315_/a_1462_47# 0.0074f
C12456 _337_/a_1270_413# _076_ 3.59e-20
C12457 trim_mask\[4\] _279_/a_490_47# 9.91e-21
C12458 clknet_2_2__leaf_clk trim_val\[4\] 1.6e-19
C12459 _093_ _065_ 0.0062f
C12460 _155_/a_68_297# _155_/a_150_297# 0.00477f
C12461 clk net3 0.00563f
C12462 mask\[7\] _222_/a_199_47# 5.21e-21
C12463 _083_ _041_ 3.53e-21
C12464 _168_/a_27_413# _227_/a_109_93# 1.68e-19
C12465 _134_ _131_ 0.0982f
C12466 _292_/a_78_199# _339_/a_1032_413# 0.00155f
C12467 VPWR _329_/a_1462_47# 2.5e-19
C12468 _288_/a_145_75# _122_ 5.55e-20
C12469 _279_/a_27_47# _279_/a_396_47# 0.00537f
C12470 _303_/a_193_47# _303_/a_543_47# 0.22f
C12471 _303_/a_27_47# _303_/a_1283_21# 0.0436f
C12472 _325_/a_27_47# mask\[7\] 6.45e-19
C12473 _096_ net30 1.8e-20
C12474 _004_ _039_ 1.08e-19
C12475 _237_/a_76_199# _095_ 0.00196f
C12476 net42 _054_ 1.86e-19
C12477 _323_/a_193_47# _020_ 0.227f
C12478 _074_ clknet_2_1__leaf_clk 0.473f
C12479 _331_/a_27_47# _330_/a_448_47# 3.88e-21
C12480 _331_/a_448_47# _330_/a_27_47# 3.88e-21
C12481 _060_ _098_ 3.68e-19
C12482 net42 net30 0.00662f
C12483 _285_/a_113_47# _065_ 8.6e-21
C12484 _320_/a_1108_47# mask\[4\] 8.26e-21
C12485 _337_/a_1108_47# _075_ 0.00231f
C12486 net15 _078_ 0.00631f
C12487 net3 net4 0.416f
C12488 _321_/a_193_47# _310_/a_27_47# 1.77e-21
C12489 _321_/a_27_47# _310_/a_193_47# 1.7e-22
C12490 _300_/a_285_47# _123_ 1.36e-19
C12491 trim_mask\[4\] _092_ 2.7e-22
C12492 _051_ _226_/a_303_47# 7.24e-19
C12493 _093_ _243_/a_109_297# 0.00354f
C12494 _324_/a_761_289# _324_/a_543_47# 0.21f
C12495 _324_/a_193_47# _324_/a_1283_21# 0.0424f
C12496 _324_/a_27_47# _324_/a_1108_47# 0.102f
C12497 net46 net18 0.0539f
C12498 _327_/a_27_47# clknet_2_3__leaf_clk 3.43e-20
C12499 net13 _248_/a_109_47# 6.47e-19
C12500 net13 _322_/a_761_289# 9.37e-19
C12501 net4 _330_/a_761_289# 0.00111f
C12502 mask\[2\] _101_ 0.269f
C12503 _308_/a_1108_47# net23 0.00198f
C12504 _308_/a_1270_413# net43 2.06e-19
C12505 _328_/a_639_47# _025_ 2.82e-19
C12506 _105_ wire42/a_75_212# 8.03e-20
C12507 _316_/a_193_47# output41/a_27_47# 9.62e-20
C12508 _238_/a_75_212# _233_/a_27_297# 5.09e-20
C12509 output21/a_27_47# _155_/a_68_297# 0.005f
C12510 _319_/a_193_47# net45 2.36e-19
C12511 _319_/a_543_47# clknet_2_0__leaf_clk 0.0375f
C12512 _060_ clknet_0_clk 1.05e-20
C12513 cal_itt\[0\] _091_ 0.134f
C12514 _048_ _266_/a_68_297# 0.206f
C12515 _200_/a_80_21# trim_mask\[0\] 1.5e-19
C12516 _338_/a_1032_413# _001_ 2.61e-19
C12517 cal_count\[1\] _134_ 2.26e-21
C12518 net27 _010_ 1.37e-19
C12519 _309_/a_27_47# net43 0.303f
C12520 net21 _084_ 1.92e-20
C12521 _325_/a_761_289# _159_/a_27_47# 0.00118f
C12522 _042_ _150_/a_27_47# 0.0295f
C12523 _187_/a_27_413# net16 0.0078f
C12524 _110_ _330_/a_1462_47# 4.63e-19
C12525 _276_/a_59_75# net46 3.42e-21
C12526 _053_ _304_/a_27_47# 0.0108f
C12527 _323_/a_1462_47# mask\[4\] 0.00237f
C12528 _305_/a_448_47# _305_/a_639_47# 4.61e-19
C12529 _093_ _232_/a_304_297# 5.61e-19
C12530 en_co_clk _087_ 1.01e-24
C12531 net12 _077_ 0.00266f
C12532 VPWR _282_/a_68_297# 0.157f
C12533 _302_/a_27_297# net46 4.03e-20
C12534 net16 _268_/a_75_212# 1.21e-20
C12535 _309_/a_543_47# _309_/a_651_413# 0.0572f
C12536 _309_/a_761_289# _309_/a_1270_413# 2.6e-19
C12537 _309_/a_193_47# _309_/a_639_47# 2.28e-19
C12538 _312_/a_1283_21# _084_ 1.03e-21
C12539 _319_/a_193_47# _065_ 5.84e-19
C12540 output32/a_27_47# trim[4] 0.00125f
C12541 trim[1] output35/a_27_47# 9.24e-19
C12542 _110_ _334_/a_543_47# 3.4e-20
C12543 _050_ _119_ 2.53e-20
C12544 VPWR _278_/a_27_47# 0.00812f
C12545 output15/a_27_47# _074_ 3.47e-20
C12546 _080_ net52 2.07e-22
C12547 _110_ _327_/a_193_47# 6.59e-21
C12548 _024_ _181_/a_68_297# 9.19e-21
C12549 _322_/a_27_47# _322_/a_543_47# 0.114f
C12550 _322_/a_193_47# _322_/a_761_289# 0.173f
C12551 _248_/a_27_297# _248_/a_373_47# 0.0134f
C12552 _176_/a_27_47# net33 0.11f
C12553 _241_/a_105_352# _099_ 0.0595f
C12554 _305_/a_448_47# clknet_2_1__leaf_clk 4.84e-20
C12555 net42 _072_ 1.06e-20
C12556 net13 _034_ 0.00173f
C12557 _257_/a_27_297# _257_/a_373_47# 0.0134f
C12558 _320_/a_27_47# mask\[2\] 0.00131f
C12559 _289_/a_68_297# _132_ 0.00342f
C12560 _168_/a_297_47# _049_ 7.02e-19
C12561 _168_/a_27_413# _054_ 0.00299f
C12562 trim_mask\[2\] _057_ 2.32e-20
C12563 _210_/a_113_297# _315_/a_193_47# 3.16e-20
C12564 _082_ net14 0.00888f
C12565 _269_/a_384_47# trim_val\[1\] 1.99e-19
C12566 _269_/a_81_21# net49 8.25e-19
C12567 _269_/a_299_297# trim_mask\[1\] 0.0595f
C12568 VPWR _179_/a_27_47# 0.244f
C12569 _168_/a_27_413# net30 0.00119f
C12570 VPWR _188_/a_27_47# 0.259f
C12571 _146_/a_150_297# clknet_2_1__leaf_clk 0.00154f
C12572 _239_/a_277_297# calibrate 0.024f
C12573 clk _062_ 0.0102f
C12574 _058_ _047_ 2.25e-19
C12575 trim[4] clkc 0.0371f
C12576 trim_val\[3\] net19 5.82e-23
C12577 _262_/a_205_47# net55 3.16e-19
C12578 _303_/a_27_47# mask\[4\] 9.47e-20
C12579 net44 _077_ 0.00501f
C12580 net22 net30 0.0562f
C12581 net31 trim_val\[0\] 1.55e-19
C12582 clkbuf_2_1__f_clk/a_110_47# _319_/a_1108_47# 0.00376f
C12583 _319_/a_27_47# _319_/a_193_47# 0.582f
C12584 VPWR _204_/a_75_212# 0.263f
C12585 net43 _201_/a_113_47# 3.14e-20
C12586 _110_ _058_ 0.0486f
C12587 _325_/a_1108_47# _101_ 2.63e-19
C12588 _325_/a_543_47# net52 5.95e-20
C12589 mask\[3\] _245_/a_109_297# 2.59e-20
C12590 _237_/a_76_199# _164_/a_161_47# 5.85e-19
C12591 cal_count\[1\] _339_/a_1602_47# 0.0975f
C12592 _036_ _339_/a_1032_413# 2.02e-20
C12593 _091_ _108_ 3.2e-20
C12594 _110_ _335_/a_193_47# 0.0115f
C12595 _116_ _335_/a_27_47# 4.14e-20
C12596 _256_/a_109_297# _108_ 7.11e-19
C12597 en_co_clk _263_/a_297_47# 8.37e-19
C12598 _050_ _087_ 6.6e-20
C12599 net28 _045_ 1.65e-19
C12600 _279_/a_204_297# trim_val\[4\] 0.0098f
C12601 _279_/a_396_47# _118_ 0.052f
C12602 _303_/a_448_47# _303_/a_639_47# 4.61e-19
C12603 _162_/a_27_47# rebuffer2/a_75_212# 3.09e-20
C12604 _048_ _028_ 8.13e-20
C12605 _291_/a_285_297# trimb[1] 5.07e-19
C12606 _065_ _202_/a_79_21# 0.0512f
C12607 _243_/a_27_297# _243_/a_373_47# 0.0134f
C12608 mask\[7\] net25 4.43e-19
C12609 _127_ cal_count\[0\] 0.286f
C12610 _047_ _332_/a_27_47# 1.63e-20
C12611 net4 _062_ 0.34f
C12612 net15 _316_/a_1283_21# 0.0144f
C12613 _103_ _171_/a_27_47# 1.75e-19
C12614 _317_/a_193_47# _316_/a_761_289# 1.78e-20
C12615 _317_/a_27_47# _316_/a_543_47# 1.37e-20
C12616 state\[2\] _166_/a_161_47# 0.26f
C12617 _068_ clknet_2_3__leaf_clk 1.16e-19
C12618 _305_/a_27_47# _067_ 1.18e-20
C12619 cal_count\[2\] _131_ 0.643f
C12620 _305_/a_27_47# _070_ 3.36e-21
C12621 _305_/a_1108_47# _202_/a_297_47# 3.77e-19
C12622 _028_ _330_/a_27_47# 5.1e-19
C12623 _331_/a_27_47# _027_ 4.98e-19
C12624 clknet_2_2__leaf_clk _330_/a_193_47# 0.0446f
C12625 _190_/a_27_47# _092_ 3.77e-20
C12626 _110_ _332_/a_27_47# 0.00426f
C12627 _188_/a_27_47# _161_/a_68_297# 1.06e-20
C12628 _314_/a_805_47# net14 6.71e-19
C12629 _169_/a_215_311# _051_ 0.0381f
C12630 VPWR _316_/a_448_47# 0.0846f
C12631 cal_itt\[1\] _198_/a_27_47# 0.215f
C12632 trim_mask\[0\] net46 0.352f
C12633 _306_/a_543_47# _003_ 3.12e-19
C12634 _324_/a_1283_21# _324_/a_1462_47# 0.0074f
C12635 _324_/a_1108_47# _324_/a_1217_47# 0.00742f
C12636 _306_/a_1283_21# _073_ 0.00125f
C12637 _106_ _262_/a_109_297# 3.99e-19
C12638 _302_/a_373_47# _108_ 8.63e-21
C12639 net9 _113_ 3.21e-20
C12640 output7/a_27_47# net15 0.00137f
C12641 _115_ _057_ 1.61e-20
C12642 net21 _085_ 8.48e-20
C12643 _074_ _313_/a_27_47# 0.0119f
C12644 _257_/a_373_47# trim_val\[4\] 2.41e-20
C12645 net4 _195_/a_76_199# 0.0136f
C12646 mask\[1\] _101_ 0.407f
C12647 _330_/a_193_47# net11 3.59e-19
C12648 _330_/a_543_47# net19 0.0116f
C12649 VPWR _304_/a_27_47# 0.501f
C12650 mask\[3\] _081_ 2.32e-20
C12651 net43 _034_ 0.021f
C12652 _050_ _263_/a_297_47# 2.23e-20
C12653 _309_/a_1217_47# net43 2.95e-19
C12654 _126_ cal_count\[0\] 0.239f
C12655 _327_/a_1283_21# _024_ 2.09e-19
C12656 _327_/a_651_413# trim_mask\[0\] 2.51e-19
C12657 _303_/a_27_47# _020_ 0.00106f
C12658 output33/a_27_47# _176_/a_27_47# 0.00817f
C12659 _097_ clknet_2_0__leaf_clk 1.42e-19
C12660 _063_ _062_ 0.322f
C12661 _305_/a_639_47# _002_ 0.00467f
C12662 fanout44/a_27_47# net52 4.86e-20
C12663 _053_ _340_/a_476_47# 5.85e-20
C12664 _251_/a_27_297# _251_/a_109_47# 0.00393f
C12665 net9 net2 0.0285f
C12666 _320_/a_543_47# _077_ 2.5e-20
C12667 _319_/a_1462_47# _065_ 1.27e-19
C12668 _277_/a_75_212# _335_/a_761_289# 7.23e-19
C12669 _320_/a_1283_21# _076_ 5.33e-20
C12670 cal_count\[1\] cal_count\[2\] 4.34e-19
C12671 _306_/a_193_47# clknet_0_clk 8.12e-20
C12672 net27 _153_/a_27_47# 0.00138f
C12673 _322_/a_1108_47# mask\[4\] 1.63e-20
C12674 VPWR _298_/a_292_297# 0.00802f
C12675 _002_ clknet_2_1__leaf_clk 0.00753f
C12676 _008_ _249_/a_27_297# 1.5e-20
C12677 trim_val\[2\] _056_ 0.228f
C12678 _228_/a_79_21# _242_/a_79_21# 0.0132f
C12679 _194_/a_113_297# _194_/a_199_47# 2.42e-19
C12680 _078_ _315_/a_1108_47# 1.81e-19
C12681 _272_/a_299_297# _272_/a_384_47# 1.48e-19
C12682 _023_ _310_/a_193_47# 4.6e-19
C12683 _327_/a_448_47# _038_ 2.76e-19
C12684 _327_/a_805_47# _136_ 1.89e-19
C12685 _195_/a_76_199# _063_ 5.74e-19
C12686 _144_/a_27_47# _125_ 0.00216f
C12687 net12 _060_ 2.45e-20
C12688 _320_/a_27_47# mask\[1\] 0.00686f
C12689 _329_/a_1283_21# trim_mask\[1\] 1.09e-19
C12690 _336_/a_1283_21# _336_/a_1108_47# 0.234f
C12691 _336_/a_761_289# _336_/a_651_413# 0.0977f
C12692 _336_/a_543_47# _336_/a_448_47# 0.0498f
C12693 _336_/a_27_47# _336_/a_639_47# 3.82e-19
C12694 _336_/a_193_47# _336_/a_1270_413# 1.46e-19
C12695 net31 _131_ 0.0059f
C12696 trim[4] _130_ 2.59e-20
C12697 _281_/a_103_199# _095_ 0.152f
C12698 _314_/a_1108_47# _046_ 3.69e-20
C12699 net16 _056_ 0.00292f
C12700 _319_/a_193_47# _319_/a_1217_47# 2.36e-20
C12701 _319_/a_543_47# _319_/a_639_47# 0.0138f
C12702 _319_/a_761_289# _319_/a_805_47# 3.69e-19
C12703 output10/a_27_47# net18 0.00701f
C12704 _237_/a_439_47# _048_ 0.00406f
C12705 _249_/a_27_297# mask\[5\] 0.112f
C12706 _276_/a_145_75# _032_ 0.00138f
C12707 _024_ _108_ 0.0014f
C12708 trim_mask\[0\] _332_/a_448_47# 5.1e-19
C12709 _329_/a_27_47# _329_/a_543_47# 0.115f
C12710 _329_/a_193_47# _329_/a_761_289# 0.186f
C12711 VPWR _321_/a_27_47# 0.445f
C12712 _079_ net30 0.0937f
C12713 _286_/a_535_374# _122_ 2.48e-19
C12714 _237_/a_535_374# net3 2.81e-19
C12715 clknet_0_clk _227_/a_109_93# 2.5e-19
C12716 _303_/a_639_47# _000_ 9.32e-19
C12717 result[5] net14 8.01e-20
C12718 VPWR _337_/a_27_47# 0.413f
C12719 _309_/a_27_47# _080_ 5.04e-20
C12720 _059_ _337_/a_543_47# 4.42e-20
C12721 trim_mask\[3\] _257_/a_27_297# 3.91e-19
C12722 _324_/a_639_47# mask\[5\] 1.48e-19
C12723 _187_/a_27_413# net40 0.00448f
C12724 _058_ _301_/a_47_47# 2.94e-19
C12725 _006_ _310_/a_761_289# 2.15e-19
C12726 _321_/a_27_47# net53 2.51e-22
C12727 _128_ cal_count\[1\] 0.18f
C12728 _305_/a_1217_47# _067_ 2.25e-21
C12729 net34 _296_/a_113_47# 1.59e-19
C12730 _209_/a_27_47# _077_ 0.326f
C12731 net5 _296_/a_113_47# 1.24e-19
C12732 clknet_2_2__leaf_clk _330_/a_1462_47# 4.64e-19
C12733 _239_/a_27_297# _239_/a_277_297# 0.145f
C12734 _239_/a_694_21# _239_/a_474_297# 0.0922f
C12735 _015_ _169_/a_215_311# 5.91e-19
C12736 _053_ _051_ 0.0391f
C12737 VPWR _013_ 0.491f
C12738 _268_/a_75_212# net40 0.0221f
C12739 _248_/a_27_297# mask\[2\] 0.00222f
C12740 _322_/a_27_47# mask\[2\] 0.0965f
C12741 _328_/a_1283_21# net46 0.347f
C12742 fanout47/a_27_47# _124_ 2.13e-19
C12743 net24 net45 2.76e-20
C12744 result[2] clknet_2_0__leaf_clk 0.00281f
C12745 VPWR net38 0.411f
C12746 _104_ _336_/a_1270_413# 3.05e-19
C12747 net14 output41/a_27_47# 0.00326f
C12748 _013_ valid 6.4e-21
C12749 _064_ _264_/a_27_297# 3.08e-19
C12750 _334_/a_543_47# clknet_2_2__leaf_clk 7.44e-19
C12751 _211_/a_109_297# clknet_2_0__leaf_clk 0.00371f
C12752 net9 _123_ 0.0156f
C12753 _331_/a_1462_47# _052_ 5.97e-20
C12754 net27 net20 0.0479f
C12755 _320_/a_1283_21# mask\[3\] 4.04e-19
C12756 _301_/a_47_47# _332_/a_27_47# 7.08e-21
C12757 _052_ _260_/a_93_21# 0.22f
C12758 _327_/a_193_47# clknet_2_2__leaf_clk 0.115f
C12759 VPWR _304_/a_1217_47# 7.1e-20
C12760 _101_ _244_/a_27_297# 0.17f
C12761 _325_/a_1283_21# net13 0.0175f
C12762 VPWR _340_/a_476_47# 0.296f
C12763 _045_ _084_ 0.0144f
C12764 _060_ _263_/a_79_21# 0.0144f
C12765 net54 _263_/a_382_297# 5.19e-19
C12766 _218_/a_199_47# mask\[5\] 1.96e-20
C12767 _053_ _338_/a_193_47# 1.27e-21
C12768 mask\[5\] _220_/a_113_297# 0.0821f
C12769 _249_/a_109_297# _084_ 5e-20
C12770 _048_ _095_ 0.0407f
C12771 _107_ _075_ 5.06e-19
C12772 net24 _065_ 3.63e-21
C12773 cal_itt\[2\] net19 9.46e-19
C12774 _251_/a_109_297# _022_ 0.00252f
C12775 _325_/a_27_47# net28 9.8e-20
C12776 _323_/a_27_47# _068_ 1.08e-20
C12777 net49 net32 1.42e-20
C12778 _250_/a_27_297# _078_ 0.00401f
C12779 _058_ clknet_2_2__leaf_clk 0.0751f
C12780 state\[2\] _088_ 0.00635f
C12781 _076_ _205_/a_27_47# 3.4e-20
C12782 _335_/a_193_47# clknet_2_2__leaf_clk 0.00249f
C12783 net30 _098_ 8.93e-20
C12784 _321_/a_1108_47# _018_ 2.29e-21
C12785 _328_/a_805_47# _058_ 2.61e-19
C12786 _341_/a_1108_47# net46 0.227f
C12787 net14 net29 0.0335f
C12788 _104_ net9 3.84e-19
C12789 _282_/a_150_297# _065_ 2.58e-19
C12790 mask\[0\] _319_/a_1283_21# 0.109f
C12791 trim_val\[2\] net48 0.0604f
C12792 _333_/a_193_47# net46 0.0553f
C12793 _040_ _076_ 3.91e-20
C12794 clk output41/a_27_47# 1.65e-19
C12795 clknet_0_clk _054_ 3.05e-19
C12796 cal_itt\[2\] _107_ 5.64e-19
C12797 _336_/a_543_47# _033_ 4.76e-19
C12798 _325_/a_1108_47# _248_/a_27_297# 4.4e-20
C12799 _321_/a_639_47# net15 1.49e-19
C12800 _325_/a_1283_21# _322_/a_193_47# 1.15e-20
C12801 clknet_0_clk net30 0.237f
C12802 _265_/a_81_21# net46 0.00127f
C12803 _332_/a_27_47# clknet_2_2__leaf_clk 0.262f
C12804 mask\[4\] _084_ 3.07e-20
C12805 en_co_clk _099_ 0.00304f
C12806 _120_ _095_ 0.0356f
C12807 net44 _311_/a_651_413# 0.0134f
C12808 output11/a_27_47# net19 2.97e-19
C12809 _110_ _227_/a_109_93# 4.49e-21
C12810 net48 net16 0.22f
C12811 _094_ _337_/a_761_289# 0.0133f
C12812 VPWR input4/a_27_47# 0.275f
C12813 VPWR _321_/a_1217_47# 4.26e-20
C12814 _287_/a_75_212# _124_ 0.242f
C12815 _035_ _286_/a_218_47# 6.37e-20
C12816 output28/a_27_47# _314_/a_27_47# 0.0132f
C12817 _323_/a_27_47# net27 4.72e-19
C12818 net3 _034_ 2.54e-21
C12819 _127_ net16 0.00342f
C12820 net13 _075_ 2.54e-20
C12821 _319_/a_193_47# _282_/a_68_297# 4.88e-19
C12822 clknet_2_1__leaf_clk _313_/a_1270_413# 3.05e-19
C12823 state\[0\] _090_ 1.04e-19
C12824 _220_/a_199_47# _084_ 0.00151f
C12825 _306_/a_761_289# clk 6.33e-21
C12826 VPWR _337_/a_1217_47# 1.14e-19
C12827 _247_/a_27_297# net52 0.177f
C12828 _247_/a_109_47# _101_ 0.00172f
C12829 _281_/a_337_297# _281_/a_253_47# 0.00219f
C12830 net2 _122_ 0.244f
C12831 net12 _306_/a_193_47# 0.0173f
C12832 _062_ _279_/a_396_47# 1.82e-19
C12833 VPWR _051_ 2.08f
C12834 _317_/a_761_289# net14 6.77e-20
C12835 _014_ _316_/a_1270_413# 5.82e-20
C12836 net45 _316_/a_651_413# 0.0138f
C12837 fanout43/a_27_47# _016_ 2.63e-19
C12838 _326_/a_761_289# net14 0.00502f
C12839 _012_ _004_ 0.00219f
C12840 _325_/a_1283_21# net43 0.272f
C12841 trim_mask\[4\] net46 0.468f
C12842 net35 _333_/a_1108_47# 3.91e-20
C12843 _322_/a_1217_47# mask\[2\] 3.77e-21
C12844 _058_ _333_/a_651_413# 6.29e-19
C12845 net2 _299_/a_27_413# 9.13e-19
C12846 _058_ trim_val\[0\] 0.0634f
C12847 fanout45/a_27_47# _317_/a_1108_47# 6.5e-20
C12848 _309_/a_761_289# mask\[3\] 9.58e-19
C12849 _309_/a_543_47# net25 3.39e-19
C12850 _309_/a_27_47# _082_ 5.57e-20
C12851 _329_/a_639_47# net9 7.53e-19
C12852 _164_/a_161_47# _048_ 0.315f
C12853 _322_/a_27_47# mask\[1\] 2.06e-20
C12854 _050_ _099_ 2.42e-19
C12855 mask\[3\] _205_/a_27_47# 5.26e-20
C12856 _134_ _108_ 3.3e-20
C12857 _253_/a_384_47# net26 0.00117f
C12858 _134_ _332_/a_543_47# 1.86e-19
C12859 clknet_0_clk _072_ 0.00187f
C12860 net16 _126_ 0.00142f
C12861 VPWR _338_/a_193_47# 0.273f
C12862 _306_/a_193_47# net44 0.0299f
C12863 mask\[7\] net15 0.0158f
C12864 _331_/a_27_47# _171_/a_27_47# 3.56e-21
C12865 clk _227_/a_209_311# 5.87e-19
C12866 _333_/a_543_47# rebuffer2/a_75_212# 0.00125f
C12867 _291_/a_35_297# _291_/a_285_297# 0.025f
C12868 VPWR _340_/a_1224_47# 9.06e-20
C12869 _111_ net18 7.79e-21
C12870 _333_/a_1283_21# _108_ 0.0051f
C12871 VPWR _023_ 0.916f
C12872 mask\[3\] _040_ 3.21e-20
C12873 net47 _286_/a_76_199# 2.22e-19
C12874 trim[2] _114_ 9.22e-20
C12875 trim_val\[0\] _332_/a_27_47# 1.33e-19
C12876 _178_/a_150_297# _057_ 4.96e-19
C12877 net43 _314_/a_27_47# 0.311f
C12878 _304_/a_193_47# _065_ 0.0205f
C12879 _337_/a_639_47# _049_ 7.11e-19
C12880 clk _317_/a_761_289# 0.00393f
C12881 _005_ mask\[1\] 2.2e-19
C12882 _210_/a_199_47# _078_ 0.00106f
C12883 _239_/a_694_21# _103_ 4.25e-20
C12884 _104_ clone7/a_27_47# 2.64e-21
C12885 trim_val\[2\] _172_/a_68_297# 5.43e-19
C12886 trim_val\[1\] _055_ 0.125f
C12887 _051_ _318_/a_27_47# 9.02e-20
C12888 _164_/a_161_47# _120_ 5.12e-20
C12889 net4 _227_/a_209_311# 2.66e-21
C12890 _110_ net30 0.214f
C12891 _181_/a_68_297# trim_val\[4\] 0.187f
C12892 _246_/a_373_47# _017_ 1.97e-19
C12893 _200_/a_209_47# _092_ 0.00314f
C12894 net3 _281_/a_253_47# 2.32e-20
C12895 _333_/a_1462_47# net46 0.00288f
C12896 net55 clone7/a_27_47# 0.0294f
C12897 net16 _172_/a_68_297# 0.00115f
C12898 _307_/a_448_47# _039_ 1.22e-19
C12899 VPWR _331_/a_639_47# 1.22e-19
C12900 _033_ _106_ 6.82e-20
C12901 _322_/a_1283_21# mask\[3\] 0.101f
C12902 rebuffer3/a_75_212# net18 0.0112f
C12903 net4 _317_/a_761_289# 0.00189f
C12904 _123_ _122_ 0.941f
C12905 VPWR _046_ 0.778f
C12906 _307_/a_1108_47# fanout43/a_27_47# 4.94e-22
C12907 output25/a_27_47# output26/a_27_47# 5.69e-19
C12908 VPWR _328_/a_543_47# 0.209f
C12909 _078_ _313_/a_193_47# 8.12e-19
C12910 output20/a_27_47# net44 0.00394f
C12911 cal_itt\[0\] _303_/a_448_47# 7.63e-20
C12912 cal_itt\[1\] _303_/a_1108_47# 1.16e-20
C12913 _093_ _013_ 0.0321f
C12914 _300_/a_285_47# clknet_2_3__leaf_clk 0.0447f
C12915 _337_/a_193_47# net45 2.77e-20
C12916 _337_/a_543_47# clknet_2_0__leaf_clk 0.00278f
C12917 net28 _314_/a_651_413# 0.00362f
C12918 result[6] _314_/a_1108_47# 1.96e-19
C12919 net23 _007_ 3.02e-20
C12920 _309_/a_761_289# _310_/a_1283_21# 3.87e-22
C12921 _309_/a_27_47# _310_/a_448_47# 1.58e-20
C12922 trim_mask\[3\] _330_/a_193_47# 1.89e-19
C12923 _319_/a_1283_21# _121_ 0.00141f
C12924 cal_itt\[2\] net43 0.00853f
C12925 result[3] net25 0.00624f
C12926 VPWR _312_/a_761_289# 0.203f
C12927 _123_ _299_/a_27_413# 5.11e-22
C12928 net12 _306_/a_1462_47# 1.18e-19
C12929 _015_ VPWR 0.564f
C12930 _257_/a_27_297# _335_/a_1283_21# 1.03e-20
C12931 _065_ net18 0.661f
C12932 VPWR _323_/a_543_47# 0.197f
C12933 net23 mask\[3\] 2.04e-20
C12934 _119_ _049_ 1.08e-19
C12935 _302_/a_27_297# rebuffer3/a_75_212# 1.03e-19
C12936 _313_/a_193_47# _313_/a_651_413# 0.0346f
C12937 _313_/a_543_47# _313_/a_1108_47# 7.99e-20
C12938 _101_ net26 0.261f
C12939 _336_/a_761_289# clkbuf_2_2__f_clk/a_110_47# 0.00792f
C12940 clk _318_/a_1108_47# 0.0526f
C12941 cal_itt\[1\] _190_/a_465_47# 0.0111f
C12942 cal_itt\[0\] _190_/a_655_47# 0.102f
C12943 VPWR _242_/a_79_21# 0.236f
C12944 _071_ _190_/a_27_47# 0.00405f
C12945 _236_/a_109_297# en_co_clk 2.11e-19
C12946 _337_/a_193_47# _065_ 0.00349f
C12947 _048_ _226_/a_27_47# 0.0335f
C12948 net28 _310_/a_543_47# 1.51e-20
C12949 net12 _054_ 2.18e-21
C12950 output31/a_27_47# net37 1.08e-19
C12951 _253_/a_81_21# _074_ 0.206f
C12952 _234_/a_109_297# mask\[0\] 4.5e-19
C12953 net12 _318_/a_1283_21# 0.00577f
C12954 _135_ _129_ 7.86e-20
C12955 net12 net30 0.011f
C12956 fanout45/a_27_47# clknet_2_0__leaf_clk 4.69e-20
C12957 _326_/a_761_289# net52 2.03e-19
C12958 _259_/a_109_47# net18 3.1e-19
C12959 _257_/a_27_297# _108_ 1.61e-21
C12960 net54 _095_ 0.173f
C12961 _325_/a_761_289# mask\[2\] 1.27e-19
C12962 _306_/a_1462_47# net44 0.00288f
C12963 VPWR _341_/a_1283_21# 0.36f
C12964 _302_/a_27_297# _065_ 0.0274f
C12965 _326_/a_805_47# mask\[7\] 9e-20
C12966 trim_mask\[0\] _111_ 0.226f
C12967 VPWR _333_/a_27_47# 0.436f
C12968 _136_ _300_/a_129_47# 0.00104f
C12969 _103_ _106_ 0.00163f
C12970 _087_ _049_ 8.72e-19
C12971 trimb[3] net16 3.69e-19
C12972 VPWR ctlp[4] 0.346f
C12973 _041_ _286_/a_218_47# 0.0019f
C12974 net47 cal_count\[0\] 0.268f
C12975 trim_val\[0\] _332_/a_1217_47# 3.85e-20
C12976 _330_/a_27_47# _330_/a_1108_47# 0.102f
C12977 _330_/a_193_47# _330_/a_1283_21# 0.0424f
C12978 _330_/a_761_289# _330_/a_543_47# 0.21f
C12979 _208_/a_218_374# _076_ 0.00733f
C12980 _208_/a_505_21# _077_ 4.91e-20
C12981 _207_/a_109_297# _076_ 0.0142f
C12982 net43 _314_/a_1217_47# 6.03e-19
C12983 _304_/a_1462_47# _065_ 4.06e-19
C12984 VPWR _308_/a_761_289# 0.227f
C12985 _311_/a_1283_21# _152_/a_68_297# 6.2e-22
C12986 net44 net30 0.0123f
C12987 en_co_clk _226_/a_109_47# 1.05e-19
C12988 state\[2\] _170_/a_299_297# 0.00523f
C12989 _127_ net40 1.19e-19
C12990 _315_/a_1270_413# net14 1.25e-19
C12991 _015_ _318_/a_27_47# 0.17f
C12992 result[2] _078_ 4.7e-20
C12993 _051_ _318_/a_1217_47# 5.08e-20
C12994 _117_ fanout46/a_27_47# 5.57e-19
C12995 trim_mask\[0\] calibrate 4.16e-20
C12996 _236_/a_109_297# _050_ 0.00217f
C12997 clkbuf_2_0__f_clk/a_110_47# net14 7.11e-22
C12998 _004_ _210_/a_199_47# 1.84e-21
C12999 _319_/a_1108_47# clknet_0_clk 0.0083f
C13000 _122_ _067_ 1.5e-19
C13001 _222_/a_199_47# _085_ 0.00151f
C13002 VPWR _320_/a_651_413# 0.134f
C13003 _097_ _316_/a_1283_21# 5.84e-19
C13004 _256_/a_27_297# trim_mask\[1\] 0.0717f
C13005 net12 _072_ 0.00247f
C13006 VPWR _339_/a_652_21# 0.247f
C13007 net8 net9 0.00149f
C13008 _327_/a_543_47# _025_ 9.83e-21
C13009 _051_ _093_ 1.44e-20
C13010 net43 _310_/a_651_413# 0.0122f
C13011 _328_/a_27_47# _271_/a_75_212# 1.35e-20
C13012 trim_mask\[0\] rebuffer3/a_75_212# 3.37e-21
C13013 _162_/a_27_47# net33 0.00588f
C13014 _329_/a_193_47# net18 5.13e-20
C13015 cal_itt\[0\] _000_ 1.21e-20
C13016 _107_ _170_/a_81_21# 0.00403f
C13017 ctlp[6] _312_/a_543_47# 9.17e-19
C13018 _324_/a_1108_47# net27 0.00103f
C13019 net22 sample 2.63e-19
C13020 VPWR _140_/a_68_297# 0.196f
C13021 _305_/a_761_289# clk 3.45e-19
C13022 _108_ trim_val\[4\] 0.299f
C13023 _322_/a_193_47# _247_/a_109_297# 1.26e-20
C13024 net12 _305_/a_193_47# 3.97e-19
C13025 _275_/a_299_297# net46 6.39e-20
C13026 trim_mask\[3\] _330_/a_1462_47# 4.97e-19
C13027 _325_/a_193_47# _325_/a_448_47# 0.0642f
C13028 _325_/a_761_289# _325_/a_1108_47# 0.0512f
C13029 _325_/a_27_47# _325_/a_651_413# 9.73e-19
C13030 _083_ mask\[3\] 6.93e-20
C13031 _126_ net40 0.234f
C13032 _305_/a_1108_47# _198_/a_27_47# 5.62e-20
C13033 _051_ wire42/a_75_212# 2.15e-20
C13034 net16 _299_/a_382_47# 4.83e-19
C13035 VPWR _307_/a_1270_413# 6.74e-19
C13036 _107_ _227_/a_296_53# 9.57e-20
C13037 _282_/a_68_297# _282_/a_150_297# 0.00477f
C13038 mask\[4\] _311_/a_193_47# 0.0256f
C13039 fanout46/a_27_47# _119_ 0.0686f
C13040 net44 _072_ 0.477f
C13041 net8 trim[2] 2.25e-19
C13042 trim_mask\[0\] _135_ 2.05e-20
C13043 _313_/a_761_289# _010_ 4.31e-19
C13044 _334_/a_193_47# _057_ 5.45e-20
C13045 net50 _327_/a_27_47# 0.00315f
C13046 _321_/a_27_47# mask\[6\] 6.01e-19
C13047 trim_mask\[0\] _105_ 0.00879f
C13048 net31 _108_ 0.0162f
C13049 _304_/a_1283_21# _067_ 0.013f
C13050 output9/a_27_47# net18 5.56e-21
C13051 _321_/a_448_47# _042_ 2.86e-19
C13052 _041_ clknet_2_0__leaf_clk 4.53e-21
C13053 _339_/a_1032_413# trimb[4] 2.64e-22
C13054 _064_ _256_/a_373_47# 2.84e-19
C13055 _104_ _256_/a_109_297# 0.00732f
C13056 _305_/a_193_47# net44 0.0117f
C13057 net23 fanout43/a_27_47# 0.0294f
C13058 _321_/a_805_47# clknet_2_1__leaf_clk 4.26e-19
C13059 _289_/a_150_297# _129_ 3.83e-19
C13060 _289_/a_68_297# _130_ 3.28e-21
C13061 clknet_2_2__leaf_clk net30 0.00237f
C13062 _328_/a_1283_21# _111_ 2.19e-19
C13063 _316_/a_27_47# _316_/a_761_289# 0.0701f
C13064 trim_mask\[3\] _058_ 4.79e-21
C13065 VPWR _333_/a_1217_47# 3.36e-20
C13066 VPWR _303_/a_761_289# 0.213f
C13067 _340_/a_381_47# _123_ 0.0144f
C13068 trim[1] trim[2] 3.16e-20
C13069 trim_mask\[3\] _335_/a_193_47# 0.00315f
C13070 net50 _335_/a_27_47# 0.00398f
C13071 trim_val\[3\] _335_/a_761_289# 4.26e-20
C13072 _234_/a_109_297# _121_ 3.7e-19
C13073 _042_ net14 1.65e-20
C13074 VPWR _295_/a_113_47# 4.85e-19
C13075 _330_/a_1108_47# _330_/a_1217_47# 0.00742f
C13076 _330_/a_1283_21# _330_/a_1462_47# 0.0074f
C13077 _172_/a_150_297# _055_ 4.96e-19
C13078 _008_ _311_/a_1283_21# 3.61e-20
C13079 _284_/a_68_297# net40 2.83e-21
C13080 _307_/a_27_47# _315_/a_27_47# 2.09e-19
C13081 _338_/a_652_21# _065_ 7.36e-20
C13082 net2 _101_ 3.53e-21
C13083 _048_ _052_ 0.119f
C13084 _074_ net21 0.473f
C13085 _341_/a_1283_21# _300_/a_47_47# 2.14e-19
C13086 state\[2\] _318_/a_651_413# 9.5e-19
C13087 _167_/a_161_47# _096_ 4.21e-21
C13088 _305_/a_761_289# _063_ 4.1e-20
C13089 _106_ clkbuf_2_3__f_clk/a_110_47# 0.00664f
C13090 calibrate _090_ 0.0169f
C13091 _217_/a_109_297# _007_ 0.0154f
C13092 _307_/a_1283_21# net30 6.9e-19
C13093 net2 _297_/a_285_47# 0.00117f
C13094 output33/a_27_47# _162_/a_27_47# 2.14e-20
C13095 _042_ _143_/a_68_297# 7.6e-19
C13096 _284_/a_150_297# _122_ 4.96e-19
C13097 VPWR _309_/a_1108_47# 0.32f
C13098 mask\[1\] _077_ 4.87e-19
C13099 _187_/a_212_413# _134_ 6.6e-19
C13100 _061_ _301_/a_47_47# 5.51e-19
C13101 net45 _331_/a_805_47# 0.00316f
C13102 VPWR _152_/a_150_297# 0.00224f
C13103 mask\[5\] _311_/a_1283_21# 5.66e-20
C13104 _091_ _067_ 0.00473f
C13105 _200_/a_80_21# _200_/a_209_47# 0.0101f
C13106 trim_mask\[0\] _194_/a_113_297# 0.0872f
C13107 clknet_2_1__leaf_clk _245_/a_373_47# 1.69e-19
C13108 trim_mask\[0\] _112_ 1.56e-19
C13109 net9 _340_/a_27_47# 0.019f
C13110 VPWR _339_/a_1056_47# 1.63e-19
C13111 _015_ _093_ 0.0433f
C13112 _211_/a_109_297# _004_ 0.0113f
C13113 trim_mask\[0\] _336_/a_1283_21# 5.37e-20
C13114 _007_ _216_/a_113_297# 2.9e-19
C13115 net45 _090_ 1.49e-20
C13116 net28 net15 0.0994f
C13117 _324_/a_193_47# net26 2.1e-21
C13118 output22/a_27_47# _074_ 0.00596f
C13119 _102_ clknet_2_1__leaf_clk 1.34e-19
C13120 _002_ clkbuf_0_clk/a_110_47# 0.00165f
C13121 calibrate _242_/a_382_297# 4.65e-19
C13122 net43 _306_/a_543_47# 1.25e-19
C13123 _339_/a_27_47# _124_ 2.96e-21
C13124 VPWR result[6] 0.49f
C13125 output8/a_27_47# net8 0.17f
C13126 _029_ _333_/a_27_47# 2.08e-20
C13127 output37/a_27_47# net2 3.29e-20
C13128 VPWR _292_/a_215_47# 0.00846f
C13129 net12 _250_/a_109_47# 3.88e-20
C13130 net15 _158_/a_68_297# 8.23e-19
C13131 _216_/a_113_297# mask\[3\] 0.0523f
C13132 _216_/a_199_47# net25 5.39e-20
C13133 _214_/a_113_297# clkbuf_2_1__f_clk/a_110_47# 1.49e-19
C13134 _335_/a_27_47# _330_/a_1108_47# 8.91e-19
C13135 _335_/a_193_47# _330_/a_1283_21# 0.00203f
C13136 _110_ trim_val\[2\] 2.39e-19
C13137 _307_/a_27_47# clknet_2_0__leaf_clk 0.259f
C13138 net7 net6 0.00138f
C13139 output34/a_27_47# _334_/a_1108_47# 5.37e-19
C13140 _079_ sample 0.00111f
C13141 net9 clknet_2_3__leaf_clk 0.162f
C13142 _111_ _265_/a_81_21# 3.52e-20
C13143 VPWR _324_/a_1270_413# 7.73e-19
C13144 ctlp[0] net28 0.0759f
C13145 _090_ _065_ 1.37e-19
C13146 mask\[4\] _311_/a_1462_47# 0.00185f
C13147 _322_/a_27_47# net26 1.42e-20
C13148 _062_ _075_ 0.442f
C13149 net15 _099_ 0.0134f
C13150 _235_/a_79_21# _099_ 6.65e-20
C13151 _235_/a_382_297# _095_ 1.16e-19
C13152 _239_/a_277_297# _051_ 1.67e-19
C13153 _110_ net16 0.0575f
C13154 VPWR output31/a_27_47# 0.358f
C13155 _320_/a_193_47# clkbuf_2_1__f_clk/a_110_47# 0.00198f
C13156 net43 _018_ 0.193f
C13157 VPWR _322_/a_651_413# 0.138f
C13158 _006_ clknet_2_1__leaf_clk 0.00374f
C13159 _259_/a_109_297# trim_mask\[2\] 8.17e-20
C13160 _064_ _258_/a_109_47# 0.00344f
C13161 _104_ _258_/a_27_297# 0.233f
C13162 _083_ _311_/a_448_47# 4.21e-20
C13163 _104_ _024_ 0.00874f
C13164 net27 _083_ 2.92e-21
C13165 net24 _321_/a_27_47# 1.24e-20
C13166 _273_/a_59_75# _056_ 8.32e-21
C13167 _064_ net4 0.0666f
C13168 _051_ _206_/a_27_93# 0.2f
C13169 _293_/a_299_297# trimb[4] 1.92e-19
C13170 output22/a_27_47# output23/a_27_47# 5.69e-19
C13171 _113_ _333_/a_1283_21# 3.12e-21
C13172 _181_/a_68_297# _058_ 0.107f
C13173 _030_ _333_/a_543_47# 5.3e-19
C13174 _338_/a_1032_413# _123_ 6.77e-19
C13175 net13 _318_/a_448_47# 0.00562f
C13176 _316_/a_1108_47# _316_/a_1270_413# 0.00645f
C13177 _316_/a_761_289# _316_/a_1217_47# 4.2e-19
C13178 _316_/a_543_47# _316_/a_805_47# 0.00171f
C13179 _198_/a_27_47# _069_ 0.044f
C13180 _195_/a_505_21# _062_ 0.0383f
C13181 VPWR _218_/a_113_297# 0.178f
C13182 net47 net16 7.59e-20
C13183 cal_itt\[2\] _062_ 0.00126f
C13184 net50 _335_/a_1217_47# 1.51e-19
C13185 _275_/a_384_47# _032_ 7.95e-20
C13186 clknet_2_1__leaf_clk _312_/a_193_47# 0.0256f
C13187 net44 _319_/a_1108_47# 1.96e-19
C13188 _308_/a_1108_47# clknet_2_0__leaf_clk 0.00133f
C13189 net30 _279_/a_204_297# 1.45e-19
C13190 _326_/a_543_47# net43 0.157f
C13191 _330_/a_639_47# net46 1.79e-19
C13192 _219_/a_109_297# net26 1.97e-19
C13193 net5 net34 0.217f
C13194 _134_ net2 0.501f
C13195 calibrate trim_mask\[4\] 0.0447f
C13196 _323_/a_761_289# clknet_2_1__leaf_clk 2.53e-19
C13197 trim[1] _055_ 0.00585f
C13198 _341_/a_1108_47# _135_ 2.01e-19
C13199 _337_/a_193_47# _282_/a_68_297# 2.71e-19
C13200 _106_ cal_count\[3\] 0.00111f
C13201 _237_/a_76_199# clknet_2_0__leaf_clk 4.11e-20
C13202 _251_/a_109_297# net52 0.0474f
C13203 _251_/a_373_47# _101_ 3.04e-19
C13204 _198_/a_109_47# _067_ 0.00165f
C13205 output10/a_27_47# _275_/a_299_297# 4.68e-19
C13206 VPWR _275_/a_81_21# 0.209f
C13207 _042_ net52 0.0113f
C13208 _334_/a_27_47# net46 0.502f
C13209 output26/a_27_47# _007_ 0.00126f
C13210 net15 _246_/a_27_297# 0.0109f
C13211 _320_/a_805_47# clknet_2_0__leaf_clk 1.55e-19
C13212 _216_/a_113_297# _310_/a_1283_21# 0.00123f
C13213 _299_/a_382_47# net40 2.78e-19
C13214 net45 trim_mask\[4\] 0.103f
C13215 _135_ _265_/a_81_21# 2.87e-21
C13216 _064_ _063_ 0.219f
C13217 output39/a_27_47# net38 4.96e-20
C13218 trim_mask\[4\] rebuffer3/a_75_212# 1.36e-21
C13219 cal_itt\[2\] _195_/a_76_199# 5.23e-21
C13220 _232_/a_304_297# _090_ 0.00148f
C13221 _328_/a_448_47# trim_mask\[1\] 0.0164f
C13222 trim_mask\[2\] net49 1.51e-19
C13223 _189_/a_27_47# _107_ 0.00319f
C13224 _021_ net20 1.25e-19
C13225 trim_mask\[2\] _272_/a_81_21# 0.111f
C13226 _200_/a_209_47# _071_ 9.76e-19
C13227 net51 _208_/a_218_47# 1.68e-19
C13228 net9 _340_/a_586_47# 7.81e-19
C13229 VPWR _246_/a_109_47# 2.99e-19
C13230 _253_/a_299_297# _078_ 0.00324f
C13231 _319_/a_1283_21# _016_ 6.74e-20
C13232 _304_/a_27_47# _304_/a_193_47# 0.827f
C13233 _099_ _049_ 0.0156f
C13234 trim_mask\[2\] _336_/a_543_47# 1.15e-20
C13235 _307_/a_639_47# calibrate 2.23e-20
C13236 _307_/a_805_47# _074_ 6.43e-19
C13237 net4 _336_/a_805_47# 4.25e-19
C13238 _329_/a_27_47# trim_mask\[2\] 2.31e-19
C13239 _334_/a_193_47# _334_/a_1270_413# 1.46e-19
C13240 _334_/a_543_47# _334_/a_448_47# 0.0498f
C13241 _334_/a_761_289# _334_/a_651_413# 0.0977f
C13242 _334_/a_1283_21# _334_/a_1108_47# 0.234f
C13243 _314_/a_193_47# _314_/a_639_47# 2.28e-19
C13244 _314_/a_761_289# _314_/a_1270_413# 2.6e-19
C13245 _314_/a_543_47# _314_/a_651_413# 0.0572f
C13246 clone1/a_27_47# _260_/a_93_21# 2.25e-20
C13247 net4 _264_/a_27_297# 0.00976f
C13248 state\[2\] _232_/a_32_297# 1.3e-19
C13249 VPWR _199_/a_193_297# 0.00241f
C13250 _326_/a_805_47# net28 2.68e-20
C13251 _187_/a_212_413# cal_count\[2\] 3.89e-19
C13252 _327_/a_761_289# _327_/a_543_47# 0.21f
C13253 _327_/a_193_47# _327_/a_1283_21# 0.0424f
C13254 _327_/a_27_47# _327_/a_1108_47# 0.102f
C13255 _336_/a_27_47# net19 0.0145f
C13256 _307_/a_639_47# net45 9.54e-19
C13257 _041_ _069_ 1.36e-19
C13258 net2 _339_/a_1602_47# 3.98e-20
C13259 _185_/a_68_297# _060_ 0.132f
C13260 _299_/a_215_297# _299_/a_382_47# 0.0105f
C13261 mask\[7\] _313_/a_193_47# 2.26e-19
C13262 _304_/a_193_47# _298_/a_292_297# 8.14e-21
C13263 _026_ _110_ 4.25e-20
C13264 _059_ _048_ 0.0919f
C13265 VPWR input3/a_75_212# 0.283f
C13266 mask\[6\] _046_ 0.075f
C13267 VPWR _291_/a_117_297# 0.00849f
C13268 clknet_0_clk _003_ 1.8e-20
C13269 _327_/a_1283_21# _058_ 0.0143f
C13270 ctlp[6] ctlp[7] 0.0358f
C13271 _014_ _241_/a_105_352# 0.171f
C13272 _259_/a_109_47# trim_mask\[4\] 5.34e-19
C13273 _104_ _260_/a_250_297# 0.0126f
C13274 _328_/a_27_47# net9 0.00722f
C13275 _341_/a_27_47# _066_ 0.0126f
C13276 input3/a_75_212# valid 9.25e-19
C13277 _000_ net26 5.23e-20
C13278 _333_/a_1108_47# _056_ 1.92e-19
C13279 _137_/a_68_297# _137_/a_150_297# 0.00477f
C13280 net13 clkbuf_2_1__f_clk/a_110_47# 2.91e-19
C13281 _336_/a_27_47# _107_ 0.00341f
C13282 _264_/a_27_297# _063_ 3.05e-19
C13283 _134_ _123_ 2.37e-20
C13284 _112_ _333_/a_193_47# 0.0105f
C13285 net49 _333_/a_761_289# 0.0106f
C13286 trim_mask\[1\] _333_/a_543_47# 7.04e-19
C13287 trim_val\[1\] _333_/a_1283_21# 0.103f
C13288 _340_/a_27_47# _122_ 0.00249f
C13289 _304_/a_27_47# net18 0.00548f
C13290 _115_ _272_/a_81_21# 0.00215f
C13291 _273_/a_59_75# net48 4.38e-19
C13292 _274_/a_75_212# trim_val\[2\] 1.82e-19
C13293 cal_count\[3\] _278_/a_109_297# 9.2e-19
C13294 _298_/a_78_199# _298_/a_215_47# 0.0907f
C13295 _301_/a_47_47# net16 0.0132f
C13296 _316_/a_193_47# net14 3.78e-20
C13297 _310_/a_27_47# _310_/a_761_289# 0.0701f
C13298 _200_/a_209_297# _053_ 2.12e-19
C13299 net34 _133_ 2.23e-20
C13300 _327_/a_193_47# _108_ 0.00281f
C13301 state\[2\] _104_ 0.0326f
C13302 _309_/a_651_413# _074_ 1.23e-20
C13303 _159_/a_27_47# _313_/a_543_47# 9.58e-20
C13304 net54 _052_ 1.63e-20
C13305 _060_ _088_ 5.91e-21
C13306 _335_/a_27_47# _335_/a_1108_47# 0.102f
C13307 _335_/a_193_47# _335_/a_1283_21# 0.0424f
C13308 _335_/a_761_289# _335_/a_543_47# 0.21f
C13309 _274_/a_75_212# net16 6.84e-19
C13310 _122_ clknet_2_3__leaf_clk 0.15f
C13311 en_co_clk net41 3.57e-19
C13312 fanout45/a_27_47# _316_/a_1283_21# 0.0122f
C13313 trim_mask\[0\] _278_/a_27_47# 6.4e-21
C13314 _262_/a_109_297# _092_ 1.19e-19
C13315 state\[2\] net55 0.0135f
C13316 _074_ _045_ 0.158f
C13317 _022_ net52 0.00375f
C13318 ctln[4] trim_val\[3\] 0.00181f
C13319 net10 net50 0.0105f
C13320 _074_ _249_/a_109_297# 3.35e-20
C13321 _058_ _332_/a_543_47# 0.00456f
C13322 net35 _332_/a_193_47# 8.54e-19
C13323 _058_ _108_ 0.228f
C13324 mask\[0\] _101_ 0.115f
C13325 _304_/a_27_47# _302_/a_27_297# 2.43e-20
C13326 net42 net19 5.45e-21
C13327 _304_/a_1108_47# clknet_0_clk 1.9e-19
C13328 _287_/a_75_212# _035_ 0.12f
C13329 _334_/a_1217_47# net46 6.14e-19
C13330 _041_ _078_ 0.409f
C13331 _194_/a_113_297# trim_mask\[4\] 1.81e-20
C13332 _188_/a_27_47# trim_mask\[0\] 3.43e-20
C13333 _082_ _310_/a_651_413# 9.17e-19
C13334 _066_ clknet_2_2__leaf_clk 6.69e-19
C13335 output26/a_27_47# result[4] 0.158f
C13336 VPWR _208_/a_439_47# 7.04e-19
C13337 _315_/a_1108_47# _099_ 1.31e-19
C13338 _327_/a_639_47# net46 0.00142f
C13339 net2 cal_count\[2\] 0.244f
C13340 net27 _314_/a_761_289# 3.66e-19
C13341 net9 _338_/a_956_413# 1.21e-19
C13342 _129_ _298_/a_292_297# 2.17e-20
C13343 _299_/a_298_297# _133_ 1.4e-21
C13344 net9 _341_/a_193_47# 0.00198f
C13345 _336_/a_1283_21# trim_mask\[4\] 0.052f
C13346 cal_itt\[1\] _068_ 0.171f
C13347 _329_/a_193_47# trim_mask\[4\] 1.26e-19
C13348 _329_/a_448_47# clknet_2_2__leaf_clk 1.12e-19
C13349 _304_/a_761_289# _304_/a_805_47# 3.69e-19
C13350 _304_/a_193_47# _304_/a_1217_47# 2.36e-20
C13351 _304_/a_543_47# _304_/a_639_47# 0.0138f
C13352 _110_ net40 1.8e-20
C13353 _230_/a_145_75# _091_ 5.76e-19
C13354 net43 _305_/a_543_47# 0.187f
C13355 _334_/a_543_47# _031_ 7.35e-20
C13356 _329_/a_1217_47# trim_mask\[2\] 1.33e-19
C13357 _026_ _258_/a_373_47# 2.43e-19
C13358 clk _316_/a_193_47# 6.05e-19
C13359 _336_/a_27_47# _279_/a_27_47# 1.13e-20
C13360 net16 clknet_2_2__leaf_clk 1.2e-19
C13361 _283_/a_75_212# _065_ 0.0287f
C13362 rebuffer1/a_75_212# rebuffer2/a_75_212# 5.35e-19
C13363 fanout47/a_27_47# _198_/a_27_47# 2.81e-20
C13364 _239_/a_27_297# trim_mask\[4\] 1.85e-21
C13365 _107_ _096_ 3.94e-19
C13366 _332_/a_27_47# _108_ 0.445f
C13367 _321_/a_27_47# _321_/a_193_47# 0.586f
C13368 _332_/a_193_47# _332_/a_761_289# 0.175f
C13369 _332_/a_27_47# _332_/a_543_47# 0.112f
C13370 _327_/a_1108_47# _327_/a_1217_47# 0.00742f
C13371 _327_/a_1283_21# _327_/a_1462_47# 0.0074f
C13372 net42 _107_ 0.0111f
C13373 _335_/a_639_47# net46 0.00482f
C13374 _074_ mask\[4\] 0.189f
C13375 VPWR _226_/a_303_47# 3.86e-19
C13376 _286_/a_76_199# _001_ 1.8e-19
C13377 net43 clkbuf_2_1__f_clk/a_110_47# 0.00886f
C13378 _169_/a_109_53# state\[0\] 0.034f
C13379 _169_/a_215_311# _053_ 0.128f
C13380 _050_ net41 1.45e-20
C13381 net47 net40 1.13e-20
C13382 _105_ _190_/a_27_47# 9.22e-20
C13383 _304_/a_448_47# _133_ 8.76e-21
C13384 _337_/a_27_47# _337_/a_193_47# 0.855f
C13385 _304_/a_1283_21# clknet_2_3__leaf_clk 4.73e-20
C13386 cal_count\[1\] cal_count\[0\] 0.112f
C13387 mask\[3\] _247_/a_373_47# 0.00178f
C13388 _333_/a_1108_47# _173_/a_27_47# 4.54e-19
C13389 _231_/a_161_47# net30 7.08e-21
C13390 output26/a_27_47# net27 7.85e-21
C13391 _340_/a_1032_413# _298_/a_78_199# 0.00129f
C13392 _309_/a_1283_21# clknet_2_1__leaf_clk 5.21e-21
C13393 _236_/a_109_297# _049_ 7.62e-20
C13394 net31 _113_ 2.53e-20
C13395 state\[1\] _099_ 6.04e-22
C13396 _048_ _203_/a_59_75# 1.4e-20
C13397 VPWR _330_/a_1270_413# 9.76e-19
C13398 net15 _085_ 0.46f
C13399 _257_/a_27_297# _336_/a_193_47# 1.28e-19
C13400 _332_/a_1270_413# net46 7.94e-19
C13401 _128_ net2 0.0683f
C13402 clkbuf_2_0__f_clk/a_110_47# _034_ 4.34e-20
C13403 _328_/a_1217_47# net9 1.84e-20
C13404 _237_/a_505_21# net55 3.76e-21
C13405 _237_/a_218_374# _096_ 0.00688f
C13406 _048_ _192_/a_27_47# 0.0203f
C13407 VPWR _267_/a_59_75# 0.22f
C13408 net47 _149_/a_68_297# 0.00372f
C13409 _337_/a_1108_47# clknet_0_clk 8.64e-21
C13410 VPWR _200_/a_209_297# 0.191f
C13411 _094_ en_co_clk 0.112f
C13412 _326_/a_1108_47# _325_/a_193_47# 1.29e-20
C13413 clknet_2_0__leaf_clk _281_/a_103_199# 1.79e-19
C13414 _326_/a_27_47# _216_/a_113_297# 5.86e-22
C13415 _310_/a_1108_47# _310_/a_1270_413# 0.00645f
C13416 _310_/a_761_289# _310_/a_1217_47# 4.2e-19
C13417 _310_/a_543_47# _310_/a_805_47# 0.00171f
C13418 net13 _096_ 0.649f
C13419 VPWR _228_/a_79_21# 0.256f
C13420 _324_/a_543_47# _042_ 8.95e-20
C13421 _314_/a_27_47# net29 0.00205f
C13422 _307_/a_27_47# _078_ 0.00861f
C13423 _307_/a_193_47# mask\[0\] 0.00201f
C13424 _307_/a_761_289# net22 0.0371f
C13425 VPWR _325_/a_639_47# 5.51e-19
C13426 _327_/a_1462_47# _108_ 4.2e-20
C13427 net31 net2 0.00231f
C13428 net21 _313_/a_1270_413# 5.17e-20
C13429 _050_ _171_/a_27_47# 0.0108f
C13430 _335_/a_1108_47# _335_/a_1217_47# 0.00742f
C13431 _335_/a_1283_21# _335_/a_1462_47# 0.0074f
C13432 net16 _333_/a_651_413# 0.0056f
C13433 _340_/a_476_47# _129_ 6.87e-21
C13434 _282_/a_68_297# _090_ 3.1e-19
C13435 _041_ fanout47/a_27_47# 0.0425f
C13436 _123_ cal_count\[2\] 0.277f
C13437 _228_/a_297_47# net41 4.1e-20
C13438 clknet_2_1__leaf_clk _158_/a_150_297# 6.18e-21
C13439 result[4] _310_/a_639_47# 3.91e-19
C13440 _062_ _170_/a_81_21# 6.81e-21
C13441 VPWR trim[3] 0.564f
C13442 _322_/a_1283_21# _250_/a_109_297# 1.33e-21
C13443 net16 trim_val\[0\] 0.0338f
C13444 _168_/a_27_413# _107_ 0.00152f
C13445 _311_/a_27_47# _311_/a_448_47# 0.0897f
C13446 _311_/a_193_47# _311_/a_1108_47# 0.119f
C13447 net27 _311_/a_27_47# 1.98e-21
C13448 net12 _003_ 0.181f
C13449 _091_ clknet_2_3__leaf_clk 0.0011f
C13450 VPWR _182_/a_27_47# 0.242f
C13451 _256_/a_109_297# clknet_2_3__leaf_clk 1.28e-20
C13452 en_co_clk _192_/a_505_280# 0.0534f
C13453 _304_/a_543_47# _136_ 0.00126f
C13454 _064_ _257_/a_109_47# 0.00489f
C13455 _104_ _257_/a_27_297# 0.242f
C13456 _000_ net2 9.24e-22
C13457 _319_/a_761_289# _092_ 2.39e-20
C13458 net9 _341_/a_1462_47# 4.41e-20
C13459 _026_ clknet_2_2__leaf_clk 0.0985f
C13460 _304_/a_1108_47# net47 0.254f
C13461 _094_ _050_ 0.00885f
C13462 _326_/a_193_47# _314_/a_193_47# 6.68e-19
C13463 _326_/a_27_47# _314_/a_761_289# 4.89e-21
C13464 output22/a_27_47# output30/a_27_47# 7.06e-19
C13465 net43 _251_/a_109_47# 3.35e-21
C13466 _336_/a_27_47# _118_ 1.22e-19
C13467 _336_/a_193_47# trim_val\[4\] 0.0128f
C13468 VPWR _314_/a_1108_47# 0.325f
C13469 VPWR net37 0.557f
C13470 _308_/a_1108_47# _078_ 0.0125f
C13471 clkbuf_2_2__f_clk/a_110_47# _119_ 0.151f
C13472 _321_/a_761_289# _321_/a_805_47# 3.69e-19
C13473 _321_/a_193_47# _321_/a_1217_47# 2.36e-20
C13474 _321_/a_543_47# _321_/a_639_47# 0.0138f
C13475 _340_/a_27_47# _340_/a_381_47# 0.069f
C13476 _340_/a_193_47# _340_/a_1602_47# 4.25e-19
C13477 _340_/a_652_21# _340_/a_1032_413# 0.00971f
C13478 net44 _003_ 0.00554f
C13479 _308_/a_27_47# result[2] 9.42e-19
C13480 VPWR _169_/a_215_311# 0.268f
C13481 _302_/a_373_47# clknet_2_3__leaf_clk 0.00164f
C13482 output28/a_27_47# result[7] 0.0564f
C13483 _149_/a_68_297# net44 1.91e-19
C13484 _001_ _072_ 1.65e-20
C13485 ctlp[0] _314_/a_543_47# 0.00126f
C13486 _048_ clknet_2_0__leaf_clk 7.83e-20
C13487 _128_ _123_ 0.281f
C13488 _059_ net54 0.318f
C13489 _301_/a_47_47# net40 0.00154f
C13490 clkbuf_2_0__f_clk/a_110_47# _281_/a_253_47# 2.55e-19
C13491 cal_count\[0\] _001_ 4.97e-19
C13492 net43 _319_/a_651_413# 0.0122f
C13493 _229_/a_27_297# _098_ 4.93e-19
C13494 _087_ _240_/a_109_297# 0.00257f
C13495 _341_/a_27_47# net40 4.38e-21
C13496 _050_ _192_/a_505_280# 0.115f
C13497 _337_/a_761_289# _337_/a_805_47# 3.69e-19
C13498 _337_/a_193_47# _337_/a_1217_47# 2.36e-20
C13499 _337_/a_543_47# _337_/a_639_47# 0.0138f
C13500 _213_/a_109_297# net45 5.77e-21
C13501 net31 trim_val\[1\] 0.0297f
C13502 _008_ clknet_2_1__leaf_clk 0.116f
C13503 _303_/a_1108_47# _069_ 0.00103f
C13504 _082_ _018_ 9.07e-20
C13505 _333_/a_805_47# net32 6.64e-20
C13506 VPWR _310_/a_193_47# 0.277f
C13507 net4 _316_/a_1462_47# 4.88e-20
C13508 _088_ _227_/a_109_93# 4e-20
C13509 _340_/a_652_21# cal_count\[3\] 8.19e-20
C13510 _340_/a_381_47# clknet_2_3__leaf_clk 0.00224f
C13511 _325_/a_27_47# _074_ 1.71e-20
C13512 _025_ _336_/a_27_47# 2.56e-21
C13513 _333_/a_1108_47# _172_/a_68_297# 1.43e-19
C13514 _326_/a_27_47# output26/a_27_47# 3.9e-19
C13515 _041_ _287_/a_75_212# 0.0515f
C13516 clknet_2_1__leaf_clk _246_/a_109_297# 0.00544f
C13517 _293_/a_81_21# _289_/a_68_297# 5.27e-19
C13518 _247_/a_27_297# _247_/a_109_297# 0.171f
C13519 _341_/a_193_47# _122_ 5.13e-19
C13520 _161_/a_68_297# net37 0.00916f
C13521 net24 _140_/a_68_297# 1.86e-19
C13522 _306_/a_193_47# _244_/a_27_297# 3.15e-19
C13523 _104_ trim_val\[4\] 0.0488f
C13524 clknet_2_1__leaf_clk mask\[5\] 0.0811f
C13525 _338_/a_193_47# net18 0.0121f
C13526 _324_/a_1108_47# _021_ 7.95e-20
C13527 _320_/a_27_47# _121_ 2.11e-20
C13528 _239_/a_474_297# _092_ 0.0755f
C13529 VPWR _334_/a_805_47# 0.0022f
C13530 _326_/a_1108_47# mask\[3\] 1.09e-21
C13531 clknet_2_0__leaf_clk _120_ 0.0431f
C13532 _314_/a_1217_47# net29 1.37e-19
C13533 net45 rebuffer5/a_161_47# 3.93e-19
C13534 _307_/a_1462_47# mask\[0\] 3.18e-19
C13535 VPWR _327_/a_1270_413# 7.99e-19
C13536 _307_/a_1217_47# _078_ 5.09e-19
C13537 net13 _313_/a_1108_47# 0.00232f
C13538 _335_/a_805_47# _032_ 1.01e-19
C13539 _189_/a_408_47# _048_ 2.21e-19
C13540 _313_/a_1108_47# _155_/a_68_297# 2.65e-19
C13541 trim_mask\[4\] _278_/a_27_47# 2.53e-20
C13542 clknet_2_2__leaf_clk net40 0.0226f
C13543 _302_/a_109_47# _136_ 0.00158f
C13544 _169_/a_215_311# _318_/a_27_47# 2.83e-20
C13545 net1 net41 0.0625f
C13546 _307_/a_761_289# _079_ 3.2e-19
C13547 _307_/a_27_47# _004_ 0.17f
C13548 net16 _131_ 0.0107f
C13549 net28 _313_/a_193_47# 0.0255f
C13550 net43 result[7] 9.52e-20
C13551 _259_/a_27_297# _330_/a_27_47# 1.16e-20
C13552 _161_/a_150_297# net46 1.6e-19
C13553 clknet_2_0__leaf_clk _076_ 0.00551f
C13554 _067_ _190_/a_655_47# 6.58e-21
C13555 _074_ _212_/a_199_47# 4.22e-19
C13556 _306_/a_1108_47# _068_ 9.75e-21
C13557 _065_ rebuffer5/a_161_47# 6.42e-19
C13558 VPWR _335_/a_1270_413# 8.38e-19
C13559 _313_/a_193_47# _158_/a_68_297# 2.04e-19
C13560 _019_ clknet_2_1__leaf_clk 0.00835f
C13561 VPWR _311_/a_543_47# 0.211f
C13562 _218_/a_113_297# mask\[6\] 2.62e-20
C13563 _250_/a_27_297# _084_ 4.16e-19
C13564 net12 _337_/a_1108_47# 2.05e-19
C13565 _110_ _280_/a_75_212# 7.08e-22
C13566 _067_ trim_val\[4\] 0.00182f
C13567 _029_ _267_/a_59_75# 1.07e-19
C13568 _111_ _267_/a_145_75# 7.45e-19
C13569 _212_/a_113_297# net45 0.00109f
C13570 _328_/a_193_47# _256_/a_27_297# 3.43e-19
C13571 _037_ _304_/a_448_47# 2.13e-19
C13572 clk net14 0.0521f
C13573 _195_/a_218_374# net30 8.83e-21
C13574 _097_ _099_ 0.0211f
C13575 _311_/a_543_47# net53 0.00637f
C13576 net43 net22 2.63e-19
C13577 _005_ mask\[0\] 3.99e-20
C13578 VPWR _332_/a_651_413# 0.142f
C13579 cal_itt\[0\] net30 3.6e-20
C13580 _340_/a_1032_413# _340_/a_1056_47# 0.0016f
C13581 _340_/a_381_47# _340_/a_586_47# 3.7e-19
C13582 _088_ _054_ 0.0123f
C13583 net2 _077_ 8.99e-20
C13584 _237_/a_76_199# _316_/a_1283_21# 1.98e-19
C13585 _005_ output24/a_27_47# 7.02e-19
C13586 _186_/a_109_297# _059_ 3.87e-19
C13587 VPWR _053_ 2.55f
C13588 _088_ net30 2.51e-19
C13589 output38/a_27_47# net34 0.0944f
C13590 net26 _310_/a_1108_47# 1.19e-19
C13591 en_co_clk _243_/a_27_297# 0.00177f
C13592 _337_/a_27_47# _090_ 5.41e-22
C13593 _253_/a_81_21# _102_ 7.47e-19
C13594 _253_/a_299_297# mask\[7\] 0.0671f
C13595 trim_mask\[0\] _051_ 0.0111f
C13596 _309_/a_1270_413# _078_ 9.62e-20
C13597 _064_ trim_val\[3\] 4.87e-20
C13598 _187_/a_212_413# _058_ 7.15e-20
C13599 _323_/a_761_289# _043_ 2.03e-21
C13600 cal_count\[1\] net16 0.0384f
C13601 _326_/a_1283_21# _310_/a_1108_47# 3.98e-19
C13602 _326_/a_1108_47# _310_/a_1283_21# 3.09e-21
C13603 _320_/a_193_47# clknet_0_clk 9.18e-19
C13604 _309_/a_1108_47# net24 0.0587f
C13605 _337_/a_1108_47# net44 0.263f
C13606 _338_/a_1032_413# clknet_2_3__leaf_clk 0.0853f
C13607 calibrate _228_/a_382_297# 0.00142f
C13608 _048_ clone1/a_27_47# 0.0259f
C13609 VPWR _310_/a_1462_47# 2.01e-19
C13610 net4 net14 1.54e-19
C13611 _060_ _192_/a_174_21# 2.07e-20
C13612 net54 _192_/a_27_47# 0.142f
C13613 _037_ _133_ 0.0115f
C13614 _051_ _337_/a_1462_47# 3.32e-20
C13615 output20/a_27_47# output19/a_27_47# 3.07e-21
C13616 net43 _313_/a_1108_47# 0.213f
C13617 _074_ net25 0.123f
C13618 trim_val\[0\] net40 3.63e-20
C13619 clknet_2_1__leaf_clk _017_ 6.06e-19
C13620 trim[1] _333_/a_1283_21# 3.74e-20
C13621 _247_/a_27_297# _018_ 0.116f
C13622 _232_/a_220_297# en_co_clk 2.85e-19
C13623 _230_/a_59_75# _107_ 2.31e-19
C13624 _306_/a_651_413# net51 3.67e-19
C13625 _341_/a_193_47# _091_ 2.12e-20
C13626 _321_/a_1270_413# _101_ 3.07e-19
C13627 _321_/a_448_47# net52 6.06e-21
C13628 output32/a_27_47# _109_ 4.83e-20
C13629 _338_/a_796_47# net18 4.63e-19
C13630 _000_ _070_ 6.75e-20
C13631 _036_ net9 0.18f
C13632 clknet_0_clk net19 0.0411f
C13633 mask\[3\] clknet_2_0__leaf_clk 1.61e-20
C13634 output34/a_27_47# _056_ 7.29e-19
C13635 _306_/a_543_47# rebuffer6/a_27_47# 4.26e-21
C13636 _189_/a_27_47# _062_ 0.4f
C13637 VPWR _224_/a_113_297# 0.24f
C13638 _337_/a_1270_413# _101_ 8.97e-21
C13639 _108_ _054_ 1.4e-20
C13640 cal_itt\[0\] _072_ 0.00264f
C13641 cal_itt\[1\] cal_itt\[3\] 0.00338f
C13642 output12/a_27_47# ctln[6] 0.342f
C13643 _337_/a_1108_47# _263_/a_79_21# 3.12e-19
C13644 ctlp[4] net18 0.00798f
C13645 _231_/a_161_47# _066_ 0.00683f
C13646 cal_itt\[0\] cal_count\[0\] 4.18e-21
C13647 _107_ _098_ 0.0442f
C13648 net30 _108_ 0.0409f
C13649 _094_ _039_ 1.23e-20
C13650 _125_ trimb[4] 0.00214f
C13651 clk _331_/a_1283_21# 5.3e-21
C13652 state\[0\] _318_/a_193_47# 4.22e-20
C13653 net52 net14 2.19e-20
C13654 _314_/a_761_289# _011_ 7.65e-19
C13655 net12 _331_/a_543_47# 5.19e-20
C13656 trimb[3] net39 0.0254f
C13657 net28 _313_/a_1462_47# 0.002f
C13658 _311_/a_651_413# net26 0.0265f
C13659 _113_ _058_ 0.00723f
C13660 _064_ _330_/a_543_47# 1.16e-21
C13661 _104_ _330_/a_193_47# 1.8e-20
C13662 _303_/a_1108_47# fanout47/a_27_47# 0.0021f
C13663 _306_/a_761_289# _306_/a_543_47# 0.21f
C13664 _306_/a_193_47# _306_/a_1283_21# 0.0424f
C13665 _306_/a_27_47# _306_/a_1108_47# 0.102f
C13666 cal_itt\[2\] _305_/a_761_289# 6.11e-19
C13667 cal_itt\[0\] _305_/a_193_47# 4.7e-21
C13668 clk net4 0.0808f
C13669 _110_ _273_/a_59_75# 0.084f
C13670 _329_/a_448_47# trim_mask\[3\] 8.81e-19
C13671 clknet_0_clk _107_ 0.039f
C13672 _326_/a_543_47# result[5] 2.17e-19
C13673 _035_ _339_/a_27_47# 2.25e-20
C13674 net3 _096_ 0.027f
C13675 net12 _229_/a_27_297# 0.00101f
C13676 _331_/a_193_47# _331_/a_651_413# 0.0346f
C13677 _331_/a_543_47# _331_/a_1108_47# 7.99e-20
C13678 fanout46/a_27_47# _027_ 2.72e-19
C13679 _215_/a_109_297# _081_ 7.96e-20
C13680 _245_/a_109_297# _101_ 0.0116f
C13681 _143_/a_68_297# net52 0.00329f
C13682 mask\[3\] _146_/a_68_297# 0.173f
C13683 net25 _146_/a_150_297# 2.14e-19
C13684 net47 _338_/a_1602_47# 0.0549f
C13685 _059_ _235_/a_382_297# 5.19e-20
C13686 _338_/a_193_47# _338_/a_652_21# 0.078f
C13687 _338_/a_27_47# _338_/a_476_47# 0.209f
C13688 _328_/a_27_47# _258_/a_27_297# 1.75e-19
C13689 _086_ _310_/a_27_47# 3.93e-22
C13690 result[2] result[3] 0.037f
C13691 _328_/a_27_47# _024_ 0.00115f
C13692 _103_ _092_ 0.0584f
C13693 _113_ _332_/a_27_47# 1.61e-20
C13694 cal _315_/a_761_289# 6.15e-19
C13695 net1 _315_/a_193_47# 0.00824f
C13696 _169_/a_109_53# net45 4.09e-21
C13697 _292_/a_78_199# _122_ 0.0843f
C13698 _074_ _310_/a_543_47# 0.0136f
C13699 net15 net41 0.00739f
C13700 _326_/a_193_47# output14/a_27_47# 3.39e-21
C13701 _214_/a_113_297# _245_/a_27_297# 2.2e-20
C13702 _327_/a_639_47# _111_ 1.76e-19
C13703 net13 _098_ 2.72e-21
C13704 VPWR valid 0.59f
C13705 net43 _079_ 2.56e-19
C13706 VPWR net53 0.629f
C13707 _134_ clknet_2_3__leaf_clk 0.0566f
C13708 clk _063_ 7.88e-20
C13709 _051_ _090_ 0.202f
C13710 _313_/a_193_47# _084_ 3.03e-21
C13711 _259_/a_27_297# _335_/a_27_47# 2.31e-19
C13712 _269_/a_81_21# net46 2.74e-20
C13713 _341_/a_543_47# cal_count\[3\] 0.0299f
C13714 _341_/a_1270_413# clknet_2_3__leaf_clk 8.2e-20
C13715 net2 _332_/a_27_47# 2.97e-19
C13716 calibrate cal 0.0111f
C13717 trim_mask\[0\] _242_/a_79_21# 2.03e-20
C13718 _074_ net1 0.113f
C13719 net13 clknet_0_clk 0.0596f
C13720 _131_ net40 0.0122f
C13721 _110_ net19 0.0477f
C13722 _081_ _101_ 0.024f
C13723 VPWR _306_/a_1270_413# 7.67e-19
C13724 VPWR _009_ 0.35f
C13725 _272_/a_299_297# _334_/a_27_47# 2.64e-20
C13726 _272_/a_81_21# _334_/a_193_47# 4.54e-19
C13727 VPWR _161_/a_68_297# 0.167f
C13728 _053_ _262_/a_27_47# 0.111f
C13729 _340_/a_476_47# _339_/a_476_47# 0.00255f
C13730 _340_/a_1032_413# _339_/a_193_47# 2.36e-20
C13731 _340_/a_193_47# _339_/a_1032_413# 1.02e-20
C13732 _327_/a_27_47# trim_mask\[1\] 6.42e-19
C13733 _074_ _039_ 4.18e-20
C13734 net1 _014_ 1.44e-20
C13735 cal net45 3.14e-19
C13736 _307_/a_543_47# net14 0.00307f
C13737 clknet_2_1__leaf_clk _314_/a_1283_21# 2.14e-20
C13738 _303_/a_27_47# _035_ 1.88e-19
C13739 _307_/a_1108_47# _138_/a_27_47# 8.52e-19
C13740 _051_ _242_/a_382_297# 1.34e-21
C13741 net4 _063_ 0.0356f
C13742 _326_/a_543_47# net29 1.9e-19
C13743 mask\[1\] _319_/a_1108_47# 2.41e-19
C13744 _227_/a_209_311# _227_/a_296_53# 0.0049f
C13745 _099_ _240_/a_109_297# 0.0113f
C13746 trim_mask\[0\] _333_/a_27_47# 4.34e-20
C13747 _043_ _303_/a_193_47# 5.52e-19
C13748 output27/a_27_47# _086_ 8.35e-19
C13749 _009_ net53 1.32e-20
C13750 VPWR _318_/a_27_47# 0.518f
C13751 _280_/a_75_212# clknet_2_2__leaf_clk 0.0284f
C13752 net47 net19 0.152f
C13753 _146_/a_68_297# _310_/a_1283_21# 9.04e-19
C13754 _144_/a_27_47# _339_/a_1602_47# 2.69e-19
C13755 trimb[2] net38 0.0166f
C13756 _058_ trim_val\[1\] 7.73e-19
C13757 _181_/a_68_297# _066_ 1.06e-20
C13758 _049_ net41 0.0018f
C13759 _323_/a_1270_413# net47 1.7e-19
C13760 _110_ _107_ 0.0146f
C13761 _318_/a_761_289# net41 2.4e-20
C13762 _100_ _075_ 1.35e-20
C13763 _312_/a_448_47# net20 0.0146f
C13764 _299_/a_215_297# _131_ 0.0586f
C13765 _305_/a_1108_47# _068_ 1.61e-21
C13766 clknet_2_1__leaf_clk _310_/a_27_47# 0.324f
C13767 _306_/a_1283_21# _306_/a_1462_47# 0.0074f
C13768 _306_/a_1108_47# _306_/a_1217_47# 0.00742f
C13769 net42 _062_ 7.43e-19
C13770 _255_/a_27_47# _048_ 0.00344f
C13771 _341_/a_543_47# _038_ 0.00788f
C13772 _026_ trim_mask\[3\] 0.00645f
C13773 _341_/a_651_413# _136_ 0.00138f
C13774 _326_/a_193_47# net26 1.15e-20
C13775 _235_/a_79_21# _094_ 0.0948f
C13776 _094_ net15 0.00573f
C13777 _331_/a_761_289# _028_ 0.0322f
C13778 _331_/a_543_47# clknet_2_2__leaf_clk 3.85e-19
C13779 cal_count\[1\] net40 0.0105f
C13780 _331_/a_651_413# _260_/a_93_21# 9.66e-21
C13781 _064_ _195_/a_505_21# 1.39e-19
C13782 net15 _317_/a_448_47# 0.00169f
C13783 _281_/a_103_199# _316_/a_1283_21# 4.66e-21
C13784 _325_/a_639_47# mask\[6\] 0.00432f
C13785 _325_/a_1283_21# _022_ 4.61e-20
C13786 _317_/a_27_47# _317_/a_1108_47# 0.102f
C13787 _317_/a_193_47# _317_/a_1283_21# 0.0418f
C13788 _317_/a_761_289# _317_/a_543_47# 0.21f
C13789 _101_ _016_ 0.0162f
C13790 _258_/a_109_297# clknet_2_2__leaf_clk 0.00682f
C13791 _326_/a_761_289# _326_/a_543_47# 0.21f
C13792 _326_/a_193_47# _326_/a_1283_21# 0.0424f
C13793 _326_/a_27_47# _326_/a_1108_47# 0.102f
C13794 net33 rebuffer1/a_75_212# 5.32e-20
C13795 _325_/a_193_47# _078_ 7.8e-19
C13796 _337_/a_27_47# _283_/a_75_212# 1.36e-19
C13797 trim_mask\[1\] rebuffer1/a_75_212# 2.07e-19
C13798 net54 _232_/a_114_297# 0.003f
C13799 _060_ _232_/a_32_297# 0.0107f
C13800 _338_/a_476_47# _338_/a_586_47# 0.00807f
C13801 _338_/a_1032_413# _338_/a_956_413# 0.00212f
C13802 _338_/a_27_47# _338_/a_1224_47# 1.63e-19
C13803 _338_/a_652_21# _338_/a_796_47# 0.00196f
C13804 VPWR _317_/a_1270_413# 5.3e-19
C13805 _104_ _327_/a_193_47# 1.35e-19
C13806 VPWR _326_/a_1270_413# 8.42e-19
C13807 _328_/a_193_47# _328_/a_448_47# 0.0564f
C13808 _328_/a_761_289# _328_/a_1108_47# 0.0512f
C13809 _328_/a_27_47# _328_/a_651_413# 9.73e-19
C13810 _306_/a_1283_21# net30 2.19e-20
C13811 _320_/a_193_47# net44 0.0241f
C13812 _036_ _122_ 0.00237f
C13813 net43 clknet_0_clk 0.152f
C13814 net45 net51 1.03e-19
C13815 output29/a_27_47# _314_/a_1108_47# 7.19e-19
C13816 _065_ _311_/a_1283_21# 2.03e-21
C13817 _313_/a_193_47# _085_ 0.0013f
C13818 net13 _337_/a_651_413# 0.00431f
C13819 net21 _312_/a_193_47# 2.49e-21
C13820 _309_/a_27_47# net14 0.0121f
C13821 _274_/a_75_212# _273_/a_59_75# 0.00216f
C13822 _051_ trim_mask\[4\] 0.266f
C13823 _053_ wire42/a_75_212# 1.84e-20
C13824 _171_/a_27_47# _049_ 0.00707f
C13825 net30 _170_/a_299_297# 8.72e-20
C13826 _340_/a_27_47# cal_count\[2\] 0.00358f
C13827 trim[0] net34 0.105f
C13828 clkbuf_2_3__f_clk/a_110_47# _092_ 0.00248f
C13829 clkbuf_2_1__f_clk/a_110_47# _247_/a_27_297# 1.56e-20
C13830 _104_ _058_ 0.00402f
C13831 _078_ _076_ 0.0104f
C13832 _015_ _090_ 6.44e-20
C13833 net31 trim[1] 0.0412f
C13834 _325_/a_1283_21# _313_/a_1283_21# 9.75e-19
C13835 VPWR _192_/a_548_47# 6.97e-20
C13836 cal_count\[1\] _299_/a_215_297# 1.12e-20
C13837 _104_ _335_/a_193_47# 0.0025f
C13838 net44 _312_/a_651_413# 0.0135f
C13839 net12 _107_ 0.0371f
C13840 _110_ _279_/a_27_47# 0.00639f
C13841 VPWR _300_/a_47_47# 0.389f
C13842 _312_/a_27_47# _312_/a_1108_47# 0.102f
C13843 _312_/a_193_47# _312_/a_1283_21# 0.0424f
C13844 _312_/a_761_289# _312_/a_543_47# 0.21f
C13845 net44 net19 0.0822f
C13846 _336_/a_448_47# net46 2.46e-19
C13847 _065_ net51 0.153f
C13848 _286_/a_76_199# _286_/a_535_374# 6.64e-19
C13849 _306_/a_27_47# clknet_2_0__leaf_clk 0.248f
C13850 _320_/a_761_289# net52 7.52e-19
C13851 _320_/a_1283_21# _101_ 5.34e-21
C13852 clknet_2_1__leaf_clk _311_/a_761_289# 7.33e-21
C13853 _090_ _242_/a_79_21# 1.33e-20
C13854 output27/a_27_47# clknet_2_1__leaf_clk 0.0124f
C13855 _329_/a_543_47# net46 0.153f
C13856 _303_/a_448_47# clknet_2_3__leaf_clk 0.0138f
C13857 VPWR _262_/a_27_47# 0.222f
C13858 _041_ _339_/a_27_47# 0.0381f
C13859 clknet_0_clk _118_ 2.72e-21
C13860 net47 _339_/a_381_47# 1.31e-20
C13861 clknet_2_3__leaf_clk cal_count\[2\] 3.1e-20
C13862 _305_/a_651_413# net51 7.46e-20
C13863 trim_val\[2\] _334_/a_448_47# 7.84e-20
C13864 _323_/a_193_47# _323_/a_448_47# 0.0594f
C13865 _323_/a_761_289# _323_/a_1108_47# 0.0512f
C13866 _323_/a_27_47# _323_/a_651_413# 9.73e-19
C13867 net13 _143_/a_150_297# 5.75e-20
C13868 _231_/a_161_47# net40 4.22e-19
C13869 _094_ _049_ 0.166f
C13870 _273_/a_59_75# clknet_2_2__leaf_clk 0.00184f
C13871 VPWR _315_/a_543_47# 0.228f
C13872 _337_/a_761_289# _092_ 1.3e-19
C13873 _306_/a_1108_47# cal_itt\[3\] 0.00238f
C13874 _306_/a_1283_21# _072_ 0.00214f
C13875 _337_/a_543_47# _099_ 1.53e-21
C13876 _328_/a_1283_21# _333_/a_27_47# 8.44e-21
C13877 net3 _316_/a_761_289# 2.15e-19
C13878 VPWR _029_ 0.411f
C13879 _319_/a_1108_47# _244_/a_27_297# 4.17e-20
C13880 VPWR _318_/a_1217_47# 2.19e-19
C13881 _242_/a_79_21# _242_/a_382_297# 0.00145f
C13882 _315_/a_543_47# valid 0.00124f
C13883 _042_ _310_/a_651_413# 1.29e-20
C13884 _306_/a_193_47# net2 1.04e-20
C13885 state\[0\] _243_/a_373_47# 6.15e-20
C13886 _060_ net55 0.168f
C13887 _074_ net15 0.00832f
C13888 _306_/a_1108_47# _305_/a_27_47# 1.65e-19
C13889 _306_/a_1283_21# _305_/a_193_47# 0.00444f
C13890 _302_/a_109_297# _092_ 0.00303f
C13891 net43 _321_/a_651_413# 0.0122f
C13892 output35/a_27_47# net33 0.0075f
C13893 _324_/a_193_47# net20 5.31e-21
C13894 _320_/a_27_47# _320_/a_1283_21# 0.0436f
C13895 _320_/a_193_47# _320_/a_543_47# 0.217f
C13896 net12 net13 0.0452f
C13897 _007_ _078_ 1.77e-19
C13898 _192_/a_505_280# _049_ 9.03e-19
C13899 VPWR _093_ 1.07f
C13900 _053_ _197_/a_113_297# 3.07e-19
C13901 _275_/a_81_21# net18 0.00275f
C13902 net43 _337_/a_651_413# 1e-19
C13903 _301_/a_377_297# _134_ 0.00106f
C13904 _331_/a_639_47# trim_mask\[4\] 2.12e-19
C13905 net15 _014_ 0.0791f
C13906 _028_ _260_/a_250_297# 9.92e-19
C13907 _128_ _144_/a_27_47# 0.00276f
C13908 _128_ clknet_2_3__leaf_clk 1.4e-20
C13909 net9 _334_/a_651_413# 4.52e-19
C13910 _317_/a_1108_47# _317_/a_1217_47# 0.00742f
C13911 _317_/a_1283_21# _317_/a_1462_47# 0.0074f
C13912 _317_/a_27_47# clknet_2_0__leaf_clk 0.323f
C13913 _308_/a_27_47# _307_/a_27_47# 5.57e-19
C13914 _328_/a_1270_413# clknet_2_2__leaf_clk 2.74e-19
C13915 _093_ valid 9.09e-19
C13916 _012_ net41 9.64e-19
C13917 ctlp[0] _074_ 0.00279f
C13918 _326_/a_1283_21# _326_/a_1462_47# 0.0074f
C13919 _326_/a_1108_47# _326_/a_1217_47# 0.00742f
C13920 mask\[3\] _078_ 0.248f
C13921 _337_/a_448_47# _034_ 0.157f
C13922 net13 _159_/a_27_47# 2.62e-19
C13923 _327_/a_1108_47# net9 0.00184f
C13924 _263_/a_79_21# _107_ 0.112f
C13925 output22/a_27_47# _308_/a_193_47# 2.68e-19
C13926 _066_ _108_ 0.0118f
C13927 trim_val\[2\] _108_ 0.0396f
C13928 _341_/a_1283_21# _341_/a_1108_47# 0.234f
C13929 _341_/a_761_289# _341_/a_651_413# 0.0977f
C13930 _341_/a_543_47# _341_/a_448_47# 0.0498f
C13931 _341_/a_27_47# _341_/a_639_47# 0.00188f
C13932 _341_/a_193_47# _341_/a_1270_413# 1.46e-19
C13933 net26 _072_ 1.07e-20
C13934 _320_/a_1462_47# net44 0.00331f
C13935 _053_ _194_/a_199_47# 0.00139f
C13936 net47 _303_/a_651_413# 0.0129f
C13937 VPWR wire42/a_75_212# 0.205f
C13938 _125_ net33 0.401f
C13939 _303_/a_27_47# _041_ 2.19e-19
C13940 _303_/a_1283_21# _338_/a_27_47# 7.36e-19
C13941 VPWR _285_/a_113_47# 7.03e-20
C13942 clknet_2_2__leaf_clk net19 0.125f
C13943 net46 net32 2.32e-19
C13944 net22 _137_/a_68_297# 0.174f
C13945 state\[1\] net41 0.00658f
C13946 _042_ _247_/a_109_297# 0.0466f
C13947 net4 _279_/a_396_47# 0.0117f
C13948 state\[2\] _028_ 0.00598f
C13949 _333_/a_27_47# _333_/a_193_47# 0.845f
C13950 net13 net44 0.217f
C13951 _069_ _068_ 1.84e-20
C13952 net16 _108_ 0.253f
C13953 _005_ _245_/a_109_297# 5e-20
C13954 net16 _332_/a_543_47# 0.00336f
C13955 clkbuf_0_clk/a_110_47# _092_ 5e-20
C13956 _290_/a_27_413# _125_ 0.243f
C13957 _318_/a_761_289# _318_/a_639_47# 3.16e-19
C13958 _318_/a_27_47# _318_/a_1217_47# 2.56e-19
C13959 cal_count\[3\] _092_ 0.0602f
C13960 _265_/a_81_21# _333_/a_27_47# 8.6e-21
C13961 net12 _322_/a_193_47# 3.45e-20
C13962 _238_/a_75_212# net1 1.02e-19
C13963 _021_ _311_/a_27_47# 7.16e-21
C13964 _189_/a_27_47# _227_/a_209_311# 4.59e-21
C13965 _233_/a_27_297# _315_/a_761_289# 3.84e-19
C13966 _203_/a_59_75# cal_itt\[3\] 0.14f
C13967 _110_ _118_ 0.0398f
C13968 _312_/a_1108_47# _312_/a_1217_47# 0.00742f
C13969 _312_/a_1283_21# _312_/a_1462_47# 0.0074f
C13970 _309_/a_761_289# _101_ 1.29e-19
C13971 _324_/a_761_289# net44 0.177f
C13972 _033_ net46 0.176f
C13973 _324_/a_27_47# _312_/a_27_47# 1.9e-20
C13974 _320_/a_193_47# _209_/a_27_47# 2.58e-19
C13975 _286_/a_535_374# cal_count\[0\] 0.00526f
C13976 net19 net11 0.0983f
C13977 VPWR _305_/a_1270_413# 5.12e-19
C13978 _101_ _205_/a_27_47# 0.0103f
C13979 _000_ clknet_2_3__leaf_clk 0.0294f
C13980 _185_/a_68_297# _316_/a_27_47# 6.01e-22
C13981 _308_/a_761_289# _308_/a_543_47# 0.21f
C13982 _308_/a_193_47# _308_/a_1283_21# 0.0424f
C13983 _308_/a_27_47# _308_/a_1108_47# 0.102f
C13984 _323_/a_805_47# net19 5.15e-19
C13985 _328_/a_27_47# _257_/a_27_297# 2.44e-19
C13986 _324_/a_193_47# _323_/a_27_47# 0.00123f
C13987 _041_ _339_/a_586_47# 0.0018f
C13988 _107_ clknet_2_2__leaf_clk 0.00487f
C13989 _107_ _260_/a_584_47# 7.02e-20
C13990 net2 _286_/a_76_199# 2.09e-21
C13991 _307_/a_193_47# _307_/a_1108_47# 0.125f
C13992 _307_/a_27_47# _307_/a_448_47# 0.0931f
C13993 trim_val\[2\] _031_ 1.29e-19
C13994 _305_/a_27_47# _203_/a_59_75# 1.32e-21
C13995 VPWR _259_/a_373_47# 2.07e-19
C13996 _333_/a_1108_47# clknet_2_2__leaf_clk 2.36e-21
C13997 _304_/a_1108_47# _001_ 6.56e-21
C13998 result[0] _307_/a_193_47# 0.001f
C13999 _040_ _101_ 0.0781f
C14000 net12 net43 0.00841f
C14001 _235_/a_79_21# _243_/a_27_297# 9.24e-21
C14002 _290_/a_207_413# output40/a_27_47# 9.59e-19
C14003 _014_ _049_ 1.21e-21
C14004 _063_ _279_/a_396_47# 2.43e-20
C14005 _181_/a_68_297# net40 4.36e-20
C14006 VPWR _319_/a_193_47# 0.561f
C14007 _322_/a_193_47# net44 0.0319f
C14008 _329_/a_448_47# _031_ 3.97e-20
C14009 _318_/a_193_47# net45 0.026f
C14010 _233_/a_27_297# calibrate 0.129f
C14011 _233_/a_109_297# _074_ 0.0159f
C14012 _058_ _172_/a_150_297# 5.6e-20
C14013 VPWR _243_/a_109_47# 1.97e-19
C14014 output29/a_27_47# _224_/a_113_297# 1.79e-20
C14015 net16 _031_ 2.98e-19
C14016 net3 clknet_0_clk 8.51e-19
C14017 _078_ _310_/a_1283_21# 0.00703f
C14018 net43 _159_/a_27_47# 0.00878f
C14019 clkbuf_2_2__f_clk/a_110_47# _330_/a_448_47# 8.5e-19
C14020 net24 _310_/a_193_47# 2.6e-21
C14021 _303_/a_651_413# net44 3.05e-19
C14022 _233_/a_27_297# net45 2.35e-19
C14023 _038_ _092_ 0.00841f
C14024 VPWR _197_/a_113_297# 0.208f
C14025 _326_/a_805_47# _074_ 5.87e-19
C14026 _320_/a_448_47# _320_/a_639_47# 4.61e-19
C14027 result[4] _078_ 5.53e-20
C14028 _323_/a_1283_21# _303_/a_761_289# 2.87e-20
C14029 _323_/a_543_47# _303_/a_543_47# 1.15e-19
C14030 _323_/a_1108_47# _303_/a_193_47# 0.00107f
C14031 _323_/a_448_47# _303_/a_27_47# 1.6e-20
C14032 net50 _256_/a_109_297# 0.0024f
C14033 net43 net44 0.0814f
C14034 _322_/a_1283_21# _101_ 1.38e-19
C14035 _322_/a_761_289# net52 3.59e-21
C14036 _339_/a_27_47# _339_/a_1032_413# 0.178f
C14037 _339_/a_193_47# _339_/a_1182_261# 0.0728f
C14038 _339_/a_652_21# _339_/a_476_47# 0.26f
C14039 _052_ clone7/a_27_47# 2.83e-37
C14040 net13 _320_/a_543_47# 0.00303f
C14041 _094_ state\[1\] 3.09e-22
C14042 _306_/a_651_413# clknet_2_1__leaf_clk 7.92e-19
C14043 _317_/a_805_47# _014_ 3.81e-19
C14044 _317_/a_448_47# state\[1\] 7.84e-20
C14045 _187_/a_212_413# _061_ 0.16f
C14046 _317_/a_639_47# net45 9.54e-19
C14047 result[5] result[7] 7.15e-19
C14048 _320_/a_27_47# _040_ 0.359f
C14049 VPWR _194_/a_199_47# 2.07e-19
C14050 VPWR _272_/a_384_47# 3.03e-19
C14051 _321_/a_1108_47# mask\[2\] 0.00219f
C14052 _271_/a_75_212# _030_ 0.109f
C14053 _315_/a_27_47# _315_/a_448_47# 0.0931f
C14054 _315_/a_193_47# _315_/a_1108_47# 0.119f
C14055 VPWR _202_/a_79_21# 0.266f
C14056 VPWR _336_/a_1108_47# 0.323f
C14057 _312_/a_1283_21# _152_/a_68_297# 3.24e-19
C14058 _328_/a_27_47# trim_val\[4\] 3.04e-21
C14059 VPWR _329_/a_761_289# 0.224f
C14060 net8 _334_/a_543_47# 0.00525f
C14061 VPWR output29/a_27_47# 0.294f
C14062 _140_/a_68_297# _140_/a_150_297# 0.00477f
C14063 _042_ _018_ 0.172f
C14064 _333_/a_543_47# _333_/a_639_47# 0.0138f
C14065 _333_/a_193_47# _333_/a_1217_47# 2.36e-20
C14066 _333_/a_761_289# _333_/a_805_47# 3.69e-19
C14067 _312_/a_193_47# _045_ 3.32e-19
C14068 fanout43/a_27_47# _078_ 0.053f
C14069 net23 _101_ 0.0393f
C14070 _230_/a_59_75# _062_ 0.00845f
C14071 _243_/a_27_297# _049_ 6.11e-19
C14072 VPWR _239_/a_277_297# 0.183f
C14073 trim_val\[0\] _333_/a_1108_47# 2.64e-21
C14074 net12 _322_/a_1462_47# 3.73e-19
C14075 _104_ _227_/a_109_93# 0.00139f
C14076 cal_itt\[0\] net40 5.38e-21
C14077 net19 _279_/a_204_297# 3.29e-19
C14078 _286_/a_76_199# _123_ 0.202f
C14079 net27 _078_ 0.445f
C14080 _078_ _311_/a_448_47# 1.55e-20
C14081 _093_ _315_/a_543_47# 1.44e-19
C14082 _265_/a_299_297# _109_ 0.00133f
C14083 calibrate _315_/a_1283_21# 0.0914f
C14084 _012_ _315_/a_193_47# 0.263f
C14085 _200_/a_80_21# clkbuf_2_3__f_clk/a_110_47# 0.00682f
C14086 _322_/a_27_47# _320_/a_1283_21# 0.00137f
C14087 _337_/a_1283_21# _226_/a_27_47# 0.00132f
C14088 _327_/a_1283_21# net40 5.37e-20
C14089 _062_ _098_ 3.97e-19
C14090 VPWR _206_/a_27_93# 0.137f
C14091 _257_/a_109_297# clknet_2_2__leaf_clk 2.86e-20
C14092 _334_/a_1108_47# net34 0.00409f
C14093 _324_/a_1283_21# net19 0.00291f
C14094 VPWR mask\[6\] 0.717f
C14095 _227_/a_109_93# net55 0.0976f
C14096 net54 _316_/a_1283_21# 6.52e-20
C14097 _262_/a_27_47# wire42/a_75_212# 3.51e-19
C14098 _308_/a_1283_21# _308_/a_1462_47# 0.0074f
C14099 _308_/a_1108_47# _308_/a_1217_47# 0.00742f
C14100 cal_itt\[1\] _122_ 1.33e-20
C14101 net2 _072_ 0.234f
C14102 _225_/a_109_297# _011_ 0.0157f
C14103 net15 _319_/a_805_47# 3.43e-19
C14104 _232_/a_220_297# _049_ 0.00703f
C14105 net2 cal_count\[0\] 1.05e-19
C14106 _230_/a_59_75# _195_/a_76_199# 1.86e-19
C14107 clknet_2_0__leaf_clk _315_/a_448_47# 0.00154f
C14108 _014_ _315_/a_1108_47# 3.11e-19
C14109 net42 _227_/a_209_311# 7.88e-20
C14110 net45 _315_/a_1283_21# 0.344f
C14111 cal_itt\[1\] _073_ 4.66e-20
C14112 _305_/a_1283_21# _072_ 0.0404f
C14113 _305_/a_1108_47# cal_itt\[3\] 4.63e-19
C14114 _321_/a_543_47# _085_ 3.19e-20
C14115 clknet_0_clk _062_ 0.142f
C14116 mask\[6\] net53 0.0795f
C14117 _235_/a_297_47# net55 0.0563f
C14118 trim_mask\[3\] _280_/a_75_212# 6.83e-19
C14119 _300_/a_377_297# _135_ 0.00232f
C14120 _322_/a_1462_47# net44 0.00384f
C14121 VPWR _319_/a_1462_47# 1.14e-19
C14122 _026_ _031_ 1.79e-20
C14123 _107_ _279_/a_204_297# 0.00129f
C14124 _318_/a_1462_47# net45 0.00288f
C14125 _309_/a_1283_21# _308_/a_1283_21# 4.89e-20
C14126 _309_/a_193_47# _308_/a_651_413# 4.01e-21
C14127 fanout44/a_27_47# clknet_0_clk 1.96e-21
C14128 _309_/a_651_413# _308_/a_193_47# 2.17e-21
C14129 _074_ _012_ 0.0814f
C14130 _110_ _330_/a_761_289# 2.26e-19
C14131 _336_/a_193_47# net30 5.93e-22
C14132 _238_/a_75_212# net15 4.65e-20
C14133 net43 _320_/a_543_47# 1.01e-19
C14134 net23 _320_/a_27_47# 1.89e-20
C14135 _305_/a_193_47# net2 1.92e-19
C14136 net35 net34 0.00132f
C14137 result[7] net29 0.00528f
C14138 _323_/a_761_289# mask\[4\] 0.00101f
C14139 _305_/a_761_289# _305_/a_543_47# 0.21f
C14140 _305_/a_193_47# _305_/a_1283_21# 0.0424f
C14141 _305_/a_27_47# _305_/a_1108_47# 0.102f
C14142 fanout47/a_27_47# _068_ 3.24e-19
C14143 trim[1] _058_ 0.00145f
C14144 clkbuf_2_2__f_clk/a_110_47# _027_ 0.0137f
C14145 _277_/a_75_212# trim_val\[3\] 4.8e-19
C14146 _239_/a_694_21# _049_ 0.00157f
C14147 _242_/a_297_47# _092_ 2.32e-20
C14148 _061_ net2 1.78e-19
C14149 _012_ _014_ 1.56e-20
C14150 _337_/a_805_47# en_co_clk 2.38e-19
C14151 _303_/a_639_47# net19 0.00129f
C14152 _262_/a_109_297# _105_ 0.00736f
C14153 net20 _156_/a_27_47# 0.111f
C14154 mask\[6\] _009_ 4.05e-19
C14155 _306_/a_193_47# mask\[0\] 7.13e-21
C14156 _108_ net40 1.01f
C14157 _332_/a_543_47# net40 7.76e-19
C14158 clknet_0_clk _195_/a_76_199# 1.29e-19
C14159 net50 _258_/a_27_297# 0.00128f
C14160 trim_mask\[3\] _258_/a_109_297# 0.00299f
C14161 _323_/a_27_47# _000_ 4.43e-20
C14162 net50 _024_ 2.32e-20
C14163 _097_ net41 3.65e-19
C14164 cal _316_/a_448_47# 3.68e-20
C14165 _339_/a_652_21# _339_/a_1224_47# 1.57e-19
C14166 _341_/a_448_47# _092_ 5.82e-21
C14167 _014_ state\[1\] 1.65e-20
C14168 _271_/a_75_212# trim_mask\[1\] 0.118f
C14169 net43 _307_/a_1283_21# 2.34e-20
C14170 _048_ _119_ 6.77e-19
C14171 _320_/a_1217_47# _040_ 0.00102f
C14172 cal_itt\[1\] _304_/a_1283_21# 0.0627f
C14173 net13 ctln[7] 0.101f
C14174 _293_/a_299_297# _339_/a_27_47# 3.38e-20
C14175 clknet_2_2__leaf_clk _118_ 2.09e-19
C14176 _104_ _054_ 0.0343f
C14177 net19 _044_ 0.00813f
C14178 _083_ _101_ 0.0013f
C14179 _104_ net30 0.677f
C14180 _168_/a_27_413# _227_/a_209_311# 6.04e-21
C14181 _168_/a_207_413# _227_/a_109_93# 2.38e-20
C14182 _119_ _330_/a_27_47# 8.06e-19
C14183 _319_/a_805_47# _049_ 2.4e-20
C14184 _244_/a_27_297# _003_ 9.28e-20
C14185 clk _330_/a_543_47# 1.65e-19
C14186 _250_/a_27_297# _074_ 3.55e-20
C14187 _279_/a_27_47# _279_/a_204_297# 0.0153f
C14188 net43 _209_/a_27_47# 3.21e-20
C14189 _303_/a_761_289# _303_/a_543_47# 0.21f
C14190 _303_/a_193_47# _303_/a_1283_21# 0.0425f
C14191 _303_/a_27_47# _303_/a_1108_47# 0.102f
C14192 net37 _129_ 1.3e-19
C14193 net55 _054_ 4.54e-20
C14194 _325_/a_193_47# mask\[7\] 1.79e-19
C14195 _325_/a_27_47# _102_ 3.99e-21
C14196 mask\[5\] _312_/a_1283_21# 5.46e-20
C14197 net55 net30 0.0559f
C14198 _237_/a_505_21# _095_ 0.00165f
C14199 _237_/a_76_199# _099_ 0.0546f
C14200 cal_count\[0\] _123_ 0.293f
C14201 _200_/a_80_21# clkbuf_0_clk/a_110_47# 1.35e-20
C14202 _048_ _087_ 0.463f
C14203 _071_ clkbuf_2_3__f_clk/a_110_47# 0.00225f
C14204 _314_/a_27_47# net14 0.00552f
C14205 _322_/a_27_47# _205_/a_27_47# 0.0117f
C14206 net52 _208_/a_76_199# 0.00104f
C14207 fanout44/a_27_47# _337_/a_651_413# 5.72e-20
C14208 _025_ clknet_2_2__leaf_clk 0.149f
C14209 _326_/a_27_47# _078_ 0.00936f
C14210 _324_/a_193_47# _324_/a_1108_47# 0.125f
C14211 _324_/a_27_47# _324_/a_448_47# 0.0931f
C14212 _327_/a_193_47# clknet_2_3__leaf_clk 4.14e-19
C14213 calibrate _243_/a_373_47# 1.78e-19
C14214 net13 _248_/a_373_47# 5.63e-19
C14215 net13 _322_/a_543_47# 0.00836f
C14216 state\[0\] _316_/a_1270_413# 8.89e-21
C14217 net4 _330_/a_543_47# 3.94e-19
C14218 _059_ clone7/a_27_47# 0.00398f
C14219 _110_ _062_ 3.13e-19
C14220 _308_/a_639_47# net43 0.00168f
C14221 _308_/a_448_47# net23 5e-20
C14222 _328_/a_805_47# _025_ 1.11e-19
C14223 net3 net44 1.09e-20
C14224 _046_ _222_/a_113_297# 0.0555f
C14225 trim_mask\[0\] _267_/a_59_75# 0.0743f
C14226 clknet_2_1__leaf_clk net45 0.266f
C14227 VPWR net24 1.61f
C14228 _322_/a_27_47# _040_ 1.61e-20
C14229 _319_/a_1283_21# clknet_2_0__leaf_clk 0.0582f
C14230 _319_/a_761_289# net45 7.31e-20
C14231 cal_itt\[1\] _091_ 0.00111f
C14232 _048_ _266_/a_150_297# 5.59e-19
C14233 output6/a_27_47# ctln[0] 0.156f
C14234 state\[1\] _243_/a_27_297# 3.97e-19
C14235 _309_/a_193_47# net43 0.031f
C14236 _325_/a_543_47# _159_/a_27_47# 1.05e-19
C14237 VPWR output39/a_27_47# 0.407f
C14238 _106_ _049_ 2e-20
C14239 _187_/a_212_413# net16 0.00604f
C14240 _058_ clknet_2_3__leaf_clk 6.52e-19
C14241 _327_/a_448_47# _256_/a_27_297# 6.81e-19
C14242 _053_ _304_/a_193_47# 0.00902f
C14243 _214_/a_113_297# mask\[2\] 0.0502f
C14244 _305_/a_1283_21# _305_/a_1462_47# 0.0074f
C14245 _305_/a_1108_47# _305_/a_1217_47# 0.00742f
C14246 VPWR _282_/a_150_297# 0.00193f
C14247 VPWR _313_/a_805_47# 3.71e-20
C14248 _309_/a_27_47# _309_/a_1217_47# 2.56e-19
C14249 _309_/a_761_289# _309_/a_639_47# 3.16e-19
C14250 _048_ _263_/a_297_47# 0.00665f
C14251 clknet_2_1__leaf_clk _065_ 0.0218f
C14252 _312_/a_1108_47# _084_ 1.83e-20
C14253 _292_/a_78_199# cal_count\[2\] 1.5e-19
C14254 trim_mask\[0\] _182_/a_27_47# 2.95e-19
C14255 _322_/a_27_47# _322_/a_1283_21# 0.0436f
C14256 _322_/a_193_47# _322_/a_543_47# 0.212f
C14257 _241_/a_105_352# _092_ 9.7e-21
C14258 _110_ _327_/a_761_289# 1.61e-20
C14259 _241_/a_388_297# _099_ 0.00421f
C14260 _241_/a_297_47# _095_ 0.00346f
C14261 _320_/a_193_47# mask\[2\] 5.9e-19
C14262 cal _013_ 4.03e-19
C14263 _168_/a_207_413# _054_ 3.69e-20
C14264 _269_/a_384_47# trim_mask\[1\] 0.0103f
C14265 _269_/a_299_297# net49 0.0484f
C14266 _269_/a_81_21# _112_ 0.115f
C14267 _253_/a_81_21# _310_/a_27_47# 0.0015f
C14268 _327_/a_27_47# _136_ 0.00263f
C14269 _239_/a_474_297# calibrate 0.0297f
C14270 _262_/a_465_47# net55 2.93e-19
C14271 net12 _062_ 0.00931f
C14272 _303_/a_193_47# mask\[4\] 2.28e-19
C14273 mask\[0\] net30 0.228f
C14274 clknet_2_1__leaf_clk _319_/a_27_47# 0.00309f
C14275 clkbuf_2_1__f_clk/a_110_47# _319_/a_448_47# 6.83e-19
C14276 _319_/a_27_47# _319_/a_761_289# 0.0535f
C14277 _325_/a_448_47# _101_ 2e-19
C14278 trim_mask\[0\] net37 0.00301f
C14279 _237_/a_505_21# _164_/a_161_47# 0.00601f
C14280 _036_ _339_/a_1602_47# 1.37e-20
C14281 _116_ _335_/a_193_47# 3.56e-20
C14282 _117_ _335_/a_27_47# 0.00205f
C14283 _110_ _335_/a_761_289# 1.39e-20
C14284 _256_/a_109_47# _108_ 1.46e-20
C14285 _067_ _072_ 0.0964f
C14286 _072_ _070_ 0.0703f
C14287 net43 _248_/a_373_47# 3.4e-20
C14288 net43 _322_/a_543_47# 2.97e-20
C14289 _050_ _089_ 5.45e-21
C14290 _113_ net16 0.00136f
C14291 cal_count\[3\] net46 0.0794f
C14292 _053_ net18 0.829f
C14293 _279_/a_204_297# _118_ 0.0147f
C14294 _279_/a_314_297# trim_val\[4\] 0.0263f
C14295 _303_/a_1108_47# _303_/a_1217_47# 0.00742f
C14296 _303_/a_1283_21# _303_/a_1462_47# 0.0074f
C14297 _065_ _202_/a_382_297# 0.00191f
C14298 clkbuf_2_0__f_clk/a_110_47# _096_ 0.0044f
C14299 output25/a_27_47# result[3] 0.159f
C14300 _032_ clkbuf_2_2__f_clk/a_110_47# 1.45e-19
C14301 _102_ net25 2.7e-20
C14302 mask\[7\] mask\[3\] 5.1e-19
C14303 _001_ net19 2.07e-19
C14304 _231_/a_161_47# _107_ 4.94e-19
C14305 net15 _316_/a_1108_47# 0.00642f
C14306 cal_itt\[2\] clk 0.0131f
C14307 _071_ clkbuf_0_clk/a_110_47# 0.0217f
C14308 _317_/a_27_47# _316_/a_1283_21# 4.57e-20
C14309 _317_/a_193_47# _316_/a_543_47# 2.29e-20
C14310 _292_/a_78_199# _128_ 0.233f
C14311 _305_/a_193_47# _067_ 6.85e-20
C14312 _305_/a_193_47# _070_ 2.92e-20
C14313 _028_ _330_/a_193_47# 2e-19
C14314 clknet_2_2__leaf_clk _330_/a_761_289# 0.0325f
C14315 _331_/a_193_47# _027_ 1.93e-19
C14316 _110_ _332_/a_193_47# 0.00146f
C14317 _314_/a_1217_47# net14 1.84e-19
C14318 net44 _062_ 5.01e-19
C14319 _169_/a_109_53# _051_ 0.0198f
C14320 VPWR _316_/a_651_413# 0.142f
C14321 _210_/a_113_297# net45 0.00159f
C14322 cal_itt\[1\] _198_/a_109_47# 0.00108f
C14323 fanout44/a_27_47# net44 0.156f
C14324 cal_itt\[0\] _198_/a_181_47# 4.2e-20
C14325 _326_/a_1217_47# _078_ 2.97e-20
C14326 _106_ _262_/a_193_297# 0.00367f
C14327 _306_/a_1108_47# _073_ 1.09e-19
C14328 _306_/a_1283_21# _003_ 1.29e-20
C14329 net2 net16 0.203f
C14330 net9 _030_ 3.65e-20
C14331 _005_ net23 0.0439f
C14332 _064_ _336_/a_27_47# 8.59e-21
C14333 _328_/a_1283_21# _267_/a_59_75# 3.41e-19
C14334 _316_/a_639_47# net41 0.0043f
C14335 _238_/a_75_212# _012_ 1.22e-19
C14336 _074_ _313_/a_193_47# 6.67e-19
C14337 _053_ _302_/a_27_297# 0.0625f
C14338 _331_/a_543_47# _088_ 1.96e-21
C14339 net4 _195_/a_505_21# 7.28e-19
C14340 cal_itt\[2\] net4 1.64e-21
C14341 VPWR _304_/a_193_47# 0.597f
C14342 _166_/a_161_47# _107_ 1.77e-19
C14343 net25 _006_ 1.92e-19
C14344 _335_/a_27_47# _119_ 1.68e-19
C14345 _309_/a_1462_47# net43 0.00196f
C14346 _328_/a_27_47# _327_/a_193_47# 2.53e-20
C14347 _328_/a_193_47# _327_/a_27_47# 2.52e-20
C14348 net14 _310_/a_651_413# 0.00145f
C14349 _327_/a_1108_47# _024_ 0.00102f
C14350 _327_/a_1270_413# trim_mask\[0\] 7.89e-20
C14351 _090_ _228_/a_79_21# 1.96e-20
C14352 _229_/a_27_297# _088_ 1.01e-19
C14353 _023_ _314_/a_448_47# 1.94e-20
C14354 _097_ _014_ 0.0205f
C14355 _263_/a_79_21# _062_ 3.44e-19
C14356 _305_/a_805_47# _002_ 0.0023f
C14357 _251_/a_27_297# _251_/a_373_47# 0.0134f
C14358 _038_ net46 0.0265f
C14359 _214_/a_113_297# mask\[1\] 0.0423f
C14360 _320_/a_1283_21# _077_ 2.48e-19
C14361 _277_/a_75_212# _335_/a_543_47# 6.3e-19
C14362 _320_/a_1108_47# _076_ 0.00196f
C14363 _308_/a_761_289# _212_/a_113_297# 0.00133f
C14364 _328_/a_27_47# _058_ 0.00513f
C14365 _322_/a_448_47# _322_/a_639_47# 4.61e-19
C14366 _322_/a_448_47# mask\[4\] 8.95e-19
C14367 VPWR _298_/a_493_297# 0.00254f
C14368 _257_/a_373_47# _025_ 1.8e-19
C14369 _258_/a_27_297# _335_/a_1108_47# 3.02e-20
C14370 net4 _335_/a_543_47# 3.88e-20
C14371 trim_val\[2\] trim_val\[1\] 0.0161f
C14372 _149_/a_68_297# net26 0.104f
C14373 _020_ _152_/a_68_297# 0.00129f
C14374 mask\[7\] _310_/a_1283_21# 0.00273f
C14375 _327_/a_1217_47# _136_ 7.17e-20
C14376 trim_mask\[1\] _336_/a_1270_413# 1.19e-20
C14377 net13 mask\[2\] 0.0636f
C14378 _195_/a_505_21# _063_ 1.54e-19
C14379 _320_/a_193_47# mask\[1\] 0.402f
C14380 cal_itt\[2\] _063_ 0.36f
C14381 clkbuf_2_0__f_clk/a_110_47# net22 1.84e-20
C14382 _227_/a_209_311# _098_ 7.16e-19
C14383 _329_/a_1108_47# trim_mask\[1\] 2.78e-20
C14384 _336_/a_543_47# _336_/a_651_413# 0.0572f
C14385 _336_/a_761_289# _336_/a_1270_413# 2.6e-19
C14386 _336_/a_193_47# _336_/a_639_47# 2.28e-19
C14387 _234_/a_109_297# clknet_2_0__leaf_clk 1.76e-21
C14388 _336_/a_27_47# _264_/a_27_297# 1.96e-20
C14389 _281_/a_103_199# _099_ 7.1e-21
C14390 _281_/a_253_297# _095_ 0.00135f
C14391 _319_/a_1108_47# _319_/a_1270_413# 0.00645f
C14392 _319_/a_761_289# _319_/a_1217_47# 4.2e-19
C14393 _319_/a_543_47# _319_/a_805_47# 0.00171f
C14394 net13 _166_/a_161_47# 1.58e-19
C14395 mask\[5\] _045_ 3.91e-21
C14396 result[4] mask\[7\] 5.8e-20
C14397 net16 trim_val\[1\] 0.0116f
C14398 _058_ _266_/a_68_297# 3.24e-19
C14399 _267_/a_59_75# _265_/a_81_21# 0.00147f
C14400 VPWR net18 1.45f
C14401 _249_/a_109_297# mask\[5\] 0.0146f
C14402 trim_mask\[0\] _332_/a_651_413# 1.2e-19
C14403 _329_/a_27_47# _329_/a_1283_21# 0.0423f
C14404 _329_/a_193_47# _329_/a_543_47# 0.23f
C14405 VPWR _321_/a_193_47# 0.585f
C14406 _273_/a_59_75# _334_/a_448_47# 2.34e-19
C14407 _073_ _203_/a_59_75# 0.111f
C14408 trim_mask\[0\] _053_ 0.396f
C14409 _218_/a_113_297# _218_/a_199_47# 2.42e-19
C14410 _169_/a_215_311# _090_ 2.65e-21
C14411 _303_/a_805_47# _000_ 3.81e-19
C14412 net54 _087_ 9.32e-20
C14413 VPWR _129_ 0.627f
C14414 VPWR _337_/a_193_47# 0.528f
C14415 net16 _123_ 0.036f
C14416 _100_ _096_ 0.0909f
C14417 _008_ mask\[4\] 0.0966f
C14418 _187_/a_212_413# net40 0.0142f
C14419 result[2] _074_ 0.00705f
C14420 output35/a_27_47# _136_ 4.5e-19
C14421 _059_ _337_/a_1283_21# 4.91e-20
C14422 trim_mask\[3\] _257_/a_109_297# 1.15e-19
C14423 net50 _257_/a_27_297# 0.00549f
C14424 _324_/a_805_47# mask\[5\] 9.25e-20
C14425 _321_/a_193_47# net53 7.04e-20
C14426 _006_ _310_/a_543_47# 2.82e-20
C14427 _128_ _036_ 0.0109f
C14428 _305_/a_1462_47# _067_ 1.46e-21
C14429 fanout43/a_27_47# _245_/a_109_47# 5.73e-20
C14430 _121_ net30 0.0346f
C14431 _181_/a_68_297# _107_ 2.75e-20
C14432 _074_ _211_/a_109_297# 0.00107f
C14433 _002_ _202_/a_297_47# 0.00166f
C14434 _239_/a_27_297# _239_/a_474_297# 0.0551f
C14435 VPWR _276_/a_59_75# 0.237f
C14436 _188_/a_27_47# _132_ 4.11e-22
C14437 _015_ _169_/a_109_53# 0.00193f
C14438 _051_ net51 3.7e-20
C14439 net5 _187_/a_27_413# 1.94e-19
C14440 _293_/a_81_21# _291_/a_35_297# 6.66e-19
C14441 _322_/a_193_47# mask\[2\] 0.0128f
C14442 _101_ _311_/a_27_47# 6.71e-21
C14443 net9 trim_mask\[1\] 0.00869f
C14444 _328_/a_1108_47# net46 0.262f
C14445 trim_mask\[2\] net46 0.25f
C14446 _033_ _105_ 1.58e-21
C14447 VPWR _302_/a_27_297# 0.216f
C14448 _219_/a_109_297# _083_ 3.99e-21
C14449 _103_ calibrate 0.00146f
C14450 _104_ _336_/a_639_47# 0.00118f
C14451 mask\[5\] mask\[4\] 0.071f
C14452 _334_/a_1283_21# clknet_2_2__leaf_clk 1.24e-20
C14453 input2/a_27_47# _297_/a_285_47# 7.66e-20
C14454 _301_/a_47_47# _332_/a_193_47# 9.75e-21
C14455 _052_ _260_/a_250_297# 0.00804f
C14456 mask\[7\] net27 0.0419f
C14457 _012_ output30/a_27_47# 1.46e-19
C14458 _327_/a_761_289# clknet_2_2__leaf_clk 5.58e-19
C14459 _325_/a_1108_47# net13 0.0152f
C14460 VPWR _340_/a_1182_261# 0.234f
C14461 _060_ _263_/a_382_297# 2.06e-19
C14462 net54 _263_/a_297_47# 0.0492f
C14463 _053_ _338_/a_652_21# 9.89e-22
C14464 _275_/a_81_21# _275_/a_299_297# 0.0821f
C14465 mask\[5\] _220_/a_199_47# 0.0103f
C14466 fanout45/a_27_47# net41 5.27e-20
C14467 _048_ _099_ 0.0926f
C14468 trim[2] net33 0.11f
C14469 net43 mask\[2\] 0.00171f
C14470 _275_/a_81_21# _178_/a_68_297# 0.00128f
C14471 cal_itt\[0\] net19 0.0181f
C14472 _323_/a_193_47# _068_ 2.08e-22
C14473 output23/a_27_47# result[2] 7.83e-19
C14474 result[1] output24/a_27_47# 0.00235f
C14475 _250_/a_109_297# _078_ 7.17e-19
C14476 _320_/a_27_47# _141_/a_27_47# 3.45e-19
C14477 state\[2\] _052_ 0.346f
C14478 _308_/a_651_413# mask\[1\] 2.4e-19
C14479 _335_/a_761_289# clknet_2_2__leaf_clk 2.9e-19
C14480 _328_/a_1217_47# _058_ 1e-20
C14481 _321_/a_448_47# _018_ 0.158f
C14482 _231_/a_161_47# _118_ 3.89e-19
C14483 _019_ mask\[4\] 0.00537f
C14484 _030_ _055_ 1.99e-20
C14485 _008_ _020_ 3.4e-20
C14486 _181_/a_68_297# _279_/a_27_47# 0.0158f
C14487 _341_/a_448_47# net46 2.46e-19
C14488 _066_ _067_ 0.155f
C14489 net50 trim_val\[4\] 7.69e-20
C14490 mask\[0\] _319_/a_1108_47# 0.0388f
C14491 trim_val\[2\] _114_ 0.0134f
C14492 _040_ _077_ 8.91e-20
C14493 _333_/a_761_289# net46 0.167f
C14494 _115_ net46 0.241f
C14495 _307_/a_1283_21# _137_/a_68_297# 0.0135f
C14496 _336_/a_1283_21# _033_ 2.48e-20
C14497 cal_itt\[0\] _107_ 3.22e-19
C14498 _265_/a_299_297# net46 3.28e-19
C14499 _325_/a_1108_47# _322_/a_193_47# 2.21e-19
C14500 _325_/a_1108_47# _248_/a_109_297# 5.3e-21
C14501 _286_/a_76_199# clknet_2_3__leaf_clk 0.00387f
C14502 _332_/a_193_47# clknet_2_2__leaf_clk 0.00303f
C14503 _018_ net14 9.06e-21
C14504 en_co_clk _092_ 0.274f
C14505 net44 _311_/a_1270_413# 3.41e-19
C14506 _107_ _088_ 0.0421f
C14507 net2 net40 0.0254f
C14508 net13 mask\[1\] 0.0277f
C14509 net27 _312_/a_27_47# 2.6e-19
C14510 VPWR trim_mask\[0\] 3.23f
C14511 _114_ net16 8.85e-19
C14512 mask\[5\] _020_ 0.00752f
C14513 clkbuf_2_0__f_clk/a_110_47# _079_ 8.04e-21
C14514 _233_/a_27_297# _013_ 2.65e-19
C14515 _329_/a_448_47# _329_/a_639_47# 4.61e-19
C14516 _094_ _337_/a_543_47# 0.038f
C14517 VPWR _321_/a_1462_47# 2.24e-19
C14518 _273_/a_59_75# _031_ 0.00952f
C14519 net13 _185_/a_68_297# 0.00304f
C14520 _035_ _286_/a_439_47# 3.12e-20
C14521 _323_/a_193_47# net27 1.6e-19
C14522 _053_ _090_ 2.67e-20
C14523 _306_/a_543_47# clk 3.57e-21
C14524 VPWR _337_/a_1462_47# 2.55e-19
C14525 _247_/a_109_297# net52 0.0105f
C14526 _247_/a_373_47# _101_ 0.00199f
C14527 net12 _306_/a_761_289# 0.00389f
C14528 _108_ net19 8.39e-19
C14529 _110_ ctln[4] 1.91e-19
C14530 _317_/a_543_47# net14 1.93e-19
C14531 _321_/a_1462_47# net53 2.16e-19
C14532 _322_/a_1283_21# _077_ 4.15e-20
C14533 _014_ _316_/a_639_47# 8.45e-19
C14534 net45 _316_/a_1270_413# 3.67e-19
C14535 _326_/a_543_47# net14 0.00717f
C14536 net2 _003_ 4.96e-20
C14537 _325_/a_1108_47# net43 0.222f
C14538 net44 rebuffer6/a_27_47# 0.00106f
C14539 _238_/a_75_212# _097_ 0.183f
C14540 trim[1] _061_ 6.73e-21
C14541 _058_ _333_/a_1270_413# 3.76e-21
C14542 _135_ clkc 2.25e-19
C14543 _330_/a_1283_21# _118_ 3.87e-22
C14544 clknet_2_3__leaf_clk net30 3.13e-21
C14545 net2 _299_/a_215_297# 0.0259f
C14546 _308_/a_193_47# _039_ 4.38e-19
C14547 ctln[1] clknet_2_0__leaf_clk 4.53e-21
C14548 _322_/a_193_47# mask\[1\] 2e-21
C14549 _309_/a_543_47# mask\[3\] 0.00691f
C14550 _329_/a_805_47# net9 4.44e-19
C14551 trim_mask\[0\] _161_/a_68_297# 0.102f
C14552 output33/a_27_47# trim[2] 0.337f
C14553 _050_ _092_ 0.882f
C14554 _026_ _104_ 0.00621f
C14555 _308_/a_27_47# fanout43/a_27_47# 0.00358f
C14556 _294_/a_68_297# net37 8.7e-20
C14557 output20/a_27_47# net20 0.238f
C14558 VPWR _191_/a_27_297# 0.459f
C14559 VPWR _338_/a_652_21# 0.242f
C14560 _102_ net15 7.88e-20
C14561 _306_/a_761_289# net44 0.168f
C14562 _107_ _108_ 0.412f
C14563 _331_/a_193_47# _171_/a_27_47# 1.18e-21
C14564 _326_/a_27_47# mask\[7\] 0.0132f
C14565 _326_/a_651_413# _253_/a_81_21# 6.67e-19
C14566 _291_/a_35_297# _291_/a_285_47# 0.00723f
C14567 VPWR _340_/a_1296_47# 5.16e-19
C14568 output19/a_27_47# net19 0.172f
C14569 _333_/a_1108_47# _108_ 0.0171f
C14570 _325_/a_27_47# mask\[5\] 2.2e-21
C14571 VPWR _297_/a_47_47# 0.376f
C14572 net47 _286_/a_505_21# 0.0104f
C14573 _265_/a_81_21# _332_/a_651_413# 2.18e-21
C14574 trim_val\[0\] _332_/a_193_47# 1.93e-19
C14575 _021_ _078_ 5.51e-21
C14576 _304_/a_761_289# _065_ 0.00475f
C14577 _337_/a_805_47# _049_ 3.28e-19
C14578 net43 _314_/a_193_47# 0.0393f
C14579 clk _317_/a_543_47# 0.00437f
C14580 _340_/a_27_47# cal_count\[0\] 3.14e-19
C14581 net34 _056_ 0.0887f
C14582 net33 _055_ 0.0246f
C14583 net43 mask\[1\] 0.144f
C14584 _239_/a_27_297# _103_ 7.91e-19
C14585 trim_mask\[1\] _055_ 0.00218f
C14586 _051_ _318_/a_193_47# 2.52e-19
C14587 cal_itt\[2\] _201_/a_113_47# 2.46e-19
C14588 _123_ net40 1.12e-20
C14589 _321_/a_543_47# _074_ 4.42e-20
C14590 _122_ net33 9.06e-21
C14591 _181_/a_150_297# trim_val\[4\] 8.47e-19
C14592 _181_/a_68_297# _118_ 0.0224f
C14593 _200_/a_303_47# _092_ 0.00324f
C14594 clkbuf_2_0__f_clk/a_110_47# clknet_0_clk 0.346f
C14595 _144_/a_27_47# cal_count\[0\] 0.0451f
C14596 _307_/a_651_413# _039_ 6.5e-19
C14597 VPWR _331_/a_805_47# 5.66e-20
C14598 _322_/a_1108_47# mask\[3\] 0.058f
C14599 cal_count\[0\] clknet_2_3__leaf_clk 0.36f
C14600 net4 _317_/a_543_47# 3.81e-19
C14601 result[3] _007_ 0.00262f
C14602 _303_/a_27_47# _068_ 0.00323f
C14603 VPWR _328_/a_1283_21# 0.353f
C14604 net33 _299_/a_27_413# 1.21e-19
C14605 _078_ _313_/a_761_289# 6.56e-20
C14606 _053_ trim_mask\[4\] 0.0186f
C14607 _329_/a_639_47# _026_ 7.96e-19
C14608 VPWR _090_ 1.24f
C14609 _125_ _339_/a_27_47# 2.29e-20
C14610 _337_/a_761_289# net45 4.08e-19
C14611 result[6] _314_/a_448_47# 9.22e-19
C14612 _108_ _279_/a_27_47# 0.235f
C14613 _309_/a_651_413# _310_/a_27_47# 6.14e-21
C14614 _309_/a_543_47# _310_/a_1283_21# 9.43e-19
C14615 _319_/a_1108_47# _121_ 1.8e-19
C14616 trim_mask\[3\] _330_/a_761_289# 8.58e-21
C14617 result[3] mask\[3\] 1.45e-19
C14618 _105_ clkbuf_2_3__f_clk/a_110_47# 0.00233f
C14619 _018_ net52 0.19f
C14620 VPWR _312_/a_543_47# 0.195f
C14621 _257_/a_109_297# _335_/a_1283_21# 8.88e-21
C14622 _257_/a_27_297# _335_/a_1108_47# 4.52e-21
C14623 state\[2\] _059_ 3.46e-20
C14624 _061_ clknet_2_3__leaf_clk 0.00543f
C14625 VPWR _323_/a_1283_21# 0.364f
C14626 _302_/a_109_297# rebuffer3/a_75_212# 1.6e-19
C14627 _166_/a_161_47# net3 3.74e-21
C14628 _313_/a_193_47# _313_/a_1270_413# 1.46e-19
C14629 _313_/a_27_47# _313_/a_639_47# 3.82e-19
C14630 _313_/a_543_47# _313_/a_448_47# 0.0498f
C14631 _313_/a_761_289# _313_/a_651_413# 0.0977f
C14632 _313_/a_1283_21# _313_/a_1108_47# 0.234f
C14633 _336_/a_543_47# clkbuf_2_2__f_clk/a_110_47# 0.00882f
C14634 cal_itt\[1\] _190_/a_655_47# 0.134f
C14635 VPWR _242_/a_382_297# 0.00464f
C14636 _071_ _190_/a_215_47# 0.00714f
C14637 clk _318_/a_448_47# 0.0164f
C14638 _111_ cal_count\[3\] 0.00281f
C14639 _337_/a_761_289# _065_ 8.96e-21
C14640 _048_ _226_/a_109_47# 0.00218f
C14641 _253_/a_299_297# _074_ 0.0564f
C14642 output37/a_27_47# trimb[4] 2.97e-20
C14643 trimb[1] output40/a_27_47# 0.00214f
C14644 trim_mask\[0\] _262_/a_27_47# 0.00833f
C14645 net12 _318_/a_1108_47# 0.00278f
C14646 _083_ _077_ 5.66e-20
C14647 _326_/a_1108_47# _101_ 6.61e-20
C14648 _326_/a_543_47# net52 1.38e-19
C14649 _064_ _230_/a_59_75# 0.00158f
C14650 net8 trim_val\[2\] 0.179f
C14651 input2/a_27_47# cal_count\[2\] 9.26e-21
C14652 _060_ _095_ 3.3e-20
C14653 net54 _099_ 0.0742f
C14654 _321_/a_27_47# clknet_2_1__leaf_clk 0.423f
C14655 VPWR _341_/a_1108_47# 0.297f
C14656 cal_itt\[0\] _118_ 0.0023f
C14657 _331_/a_448_47# net30 5.29e-20
C14658 _312_/a_543_47# _009_ 2.71e-19
C14659 _326_/a_1217_47# mask\[7\] 7.28e-19
C14660 _302_/a_109_297# _065_ 3.33e-21
C14661 VPWR _175_/a_68_297# 0.147f
C14662 trim_mask\[0\] _029_ 0.00237f
C14663 net34 _173_/a_27_47# 0.0121f
C14664 VPWR _333_/a_193_47# 0.623f
C14665 _136_ _300_/a_285_47# 0.00637f
C14666 _089_ _049_ 0.00246f
C14667 net4 _318_/a_448_47# 1.7e-19
C14668 _041_ _286_/a_439_47# 0.00175f
C14669 VPWR _265_/a_81_21# 0.245f
C14670 _124_ _338_/a_27_47# 2.26e-20
C14671 _067_ net40 3.32e-19
C14672 net8 net16 0.103f
C14673 net47 _150_/a_27_47# 6.57e-19
C14674 _208_/a_218_374# _077_ 1.1e-19
C14675 trim_val\[0\] _332_/a_1462_47# 1.25e-19
C14676 _330_/a_27_47# _330_/a_448_47# 0.0867f
C14677 _330_/a_193_47# _330_/a_1108_47# 0.125f
C14678 _208_/a_535_374# _076_ 0.00551f
C14679 calibrate _331_/a_27_47# 6.64e-20
C14680 net43 _314_/a_1462_47# 0.00288f
C14681 VPWR _308_/a_543_47# 0.23f
C14682 _194_/a_113_297# clkbuf_2_3__f_clk/a_110_47# 5.57e-19
C14683 state\[2\] _170_/a_384_47# 8.2e-20
C14684 _100_ _098_ 0.048f
C14685 cal_count\[3\] rebuffer3/a_75_212# 0.012f
C14686 _315_/a_639_47# net14 7.18e-19
C14687 _015_ _318_/a_193_47# 0.255f
C14688 _064_ clknet_0_clk 1.04e-19
C14689 net43 _244_/a_27_297# 0.00135f
C14690 _127_ net34 1.73e-19
C14691 _231_/a_161_47# _062_ 7.77e-21
C14692 _266_/a_68_297# net30 0.0328f
C14693 _059_ _237_/a_505_21# 7.37e-21
C14694 net45 _331_/a_27_47# 0.298f
C14695 ctlp[6] net21 3.56e-20
C14696 VPWR _320_/a_1270_413# 5.58e-19
C14697 _097_ _316_/a_1108_47# 9.37e-19
C14698 _256_/a_109_297# trim_mask\[1\] 0.00342f
C14699 VPWR _339_/a_476_47# 0.285f
C14700 VPWR trim_mask\[4\] 1.13f
C14701 _143_/a_68_297# clkbuf_2_1__f_clk/a_110_47# 5.14e-19
C14702 net43 _310_/a_1270_413# 1.09e-19
C14703 net27 net28 0.41f
C14704 _328_/a_193_47# _271_/a_75_212# 1.96e-19
C14705 clkbuf_0_clk/a_110_47# _065_ 1.79e-20
C14706 trim[1] net16 5.53e-20
C14707 _336_/a_1108_47# net18 1.3e-20
C14708 _065_ cal_count\[3\] 0.0151f
C14709 VPWR output13/a_27_47# 0.472f
C14710 result[3] result[4] 0.0472f
C14711 _329_/a_27_47# _256_/a_27_297# 1.23e-19
C14712 trim_mask\[0\] wire42/a_75_212# 4.51e-19
C14713 net26 net19 0.0105f
C14714 _107_ _170_/a_299_297# 0.00161f
C14715 _135_ cal_count\[3\] 0.00333f
C14716 _016_ net30 1.45e-19
C14717 _200_/a_80_21# en_co_clk 0.0268f
C14718 _162_/a_27_47# net49 5.55e-21
C14719 mask\[0\] sample 1.96e-19
C14720 VPWR _140_/a_150_297# 0.00335f
C14721 _108_ _118_ 0.445f
C14722 net12 _305_/a_761_289# 7.74e-20
C14723 _325_/a_543_47# _325_/a_1108_47# 7.99e-20
C14724 _325_/a_193_47# _325_/a_651_413# 0.0346f
C14725 _105_ cal_count\[3\] 0.0584f
C14726 _189_/a_27_47# clk 0.0122f
C14727 output14/a_27_47# output28/a_27_47# 0.00151f
C14728 _126_ net34 0.00327f
C14729 net31 input2/a_27_47# 0.00901f
C14730 VPWR _307_/a_639_47# 4.04e-19
C14731 _074_ _041_ 0.0864f
C14732 _090_ _192_/a_548_47# 6.74e-20
C14733 _107_ _227_/a_368_53# 2.25e-19
C14734 mask\[4\] _311_/a_761_289# 0.0219f
C14735 mask\[7\] _011_ 2.81e-19
C14736 _313_/a_543_47# _010_ 0.00139f
C14737 clkbuf_2_2__f_clk/a_110_47# _106_ 5.96e-21
C14738 _080_ mask\[1\] 0.0845f
C14739 VPWR trimb[2] 0.581f
C14740 net31 rebuffer2/a_75_212# 6.95e-19
C14741 _321_/a_193_47# mask\[6\] 7.54e-20
C14742 _185_/a_68_297# net3 7.88e-22
C14743 clknet_2_0__leaf_clk _101_ 0.137f
C14744 _304_/a_1108_47# _067_ 0.0051f
C14745 _321_/a_651_413# _042_ 0.00176f
C14746 _104_ _256_/a_109_47# 0.00354f
C14747 _305_/a_761_289# net44 0.0065f
C14748 _294_/a_68_297# VPWR 0.156f
C14749 _320_/a_1283_21# net30 4.43e-21
C14750 _321_/a_1217_47# clknet_2_1__leaf_clk 8.36e-20
C14751 _028_ net30 6.27e-21
C14752 _316_/a_193_47# _316_/a_761_289# 0.186f
C14753 _316_/a_27_47# _316_/a_543_47# 0.111f
C14754 _038_ _065_ 0.243f
C14755 _328_/a_1283_21# _029_ 5.83e-21
C14756 net50 _058_ 0.0378f
C14757 VPWR _333_/a_1462_47# 8.45e-20
C14758 VPWR _303_/a_543_47# 0.222f
C14759 _340_/a_562_413# _123_ 0.00221f
C14760 net50 _335_/a_193_47# 0.00563f
C14761 trim_mask\[3\] _335_/a_761_289# 5.63e-20
C14762 trim_val\[3\] _335_/a_543_47# 1.48e-20
C14763 _110_ _064_ 0.00401f
C14764 _008_ _311_/a_1108_47# 1.09e-19
C14765 _330_/a_27_47# _027_ 0.617f
C14766 _194_/a_113_297# cal_count\[3\] 1.5e-19
C14767 calibrate _331_/a_1217_47# 6.96e-20
C14768 _338_/a_476_47# _065_ 4.08e-20
C14769 output32/a_27_47# _188_/a_27_47# 2.58e-19
C14770 _066_ clknet_2_3__leaf_clk 0.29f
C14771 clk _336_/a_27_47# 2.69e-21
C14772 state\[2\] _318_/a_1270_413# 8.41e-20
C14773 _341_/a_1108_47# _300_/a_47_47# 3.89e-19
C14774 _305_/a_543_47# _063_ 1.33e-20
C14775 cal input3/a_75_212# 0.00459f
C14776 _093_ _090_ 0.0849f
C14777 _307_/a_1108_47# net30 1.86e-19
C14778 _267_/a_59_75# _267_/a_145_75# 0.00658f
C14779 _320_/a_27_47# clknet_2_0__leaf_clk 0.264f
C14780 net43 output14/a_27_47# 0.0031f
C14781 net13 net26 0.0114f
C14782 VPWR _283_/a_75_212# 0.224f
C14783 net16 _144_/a_27_47# 0.118f
C14784 net47 _042_ 0.0705f
C14785 VPWR _309_/a_448_47# 0.0791f
C14786 net45 _331_/a_1217_47# 6.03e-19
C14787 VPWR _190_/a_27_47# 0.31f
C14788 net34 output5/a_27_47# 0.00396f
C14789 net16 clknet_2_3__leaf_clk 0.016f
C14790 net5 output5/a_27_47# 0.197f
C14791 _188_/a_27_47# clkc 7.28e-19
C14792 _181_/a_68_297# _062_ 3.02e-20
C14793 _258_/a_27_297# trim_mask\[1\] 2.65e-19
C14794 _024_ trim_mask\[1\] 1.13e-19
C14795 _200_/a_209_297# _200_/a_209_47# 6.96e-20
C14796 _200_/a_80_21# _200_/a_303_47# 0.0115f
C14797 trim_mask\[0\] _194_/a_199_47# 0.00917f
C14798 clkbuf_2_1__f_clk/a_110_47# net52 0.241f
C14799 net9 _340_/a_193_47# 0.0212f
C14800 VPWR _339_/a_1224_47# 8.97e-20
C14801 _076_ rebuffer4/a_27_47# 0.246f
C14802 trim_mask\[0\] _336_/a_1108_47# 5.1e-20
C14803 state\[1\] _089_ 3.47e-20
C14804 _307_/a_27_47# _074_ 0.0166f
C14805 net4 _336_/a_27_47# 0.00723f
C14806 VPWR _249_/a_27_297# 0.226f
C14807 _326_/a_27_47# net28 9.15e-20
C14808 _228_/a_79_21# _228_/a_382_297# 0.00145f
C14809 _071_ en_co_clk 0.125f
C14810 _023_ clknet_2_1__leaf_clk 0.184f
C14811 net43 _306_/a_1283_21# 0.00135f
C14812 calibrate _242_/a_297_47# 0.0509f
C14813 _339_/a_193_47# _124_ 1.29e-20
C14814 net12 _250_/a_373_47# 0.00129f
C14815 _335_/a_193_47# _330_/a_1108_47# 1.74e-20
C14816 _104_ _280_/a_75_212# 0.0245f
C14817 _216_/a_199_47# mask\[3\] 0.0105f
C14818 _051_ _336_/a_448_47# 8.21e-21
C14819 _307_/a_193_47# clknet_2_0__leaf_clk 0.00805f
C14820 net12 _042_ 0.00452f
C14821 trim[3] _334_/a_27_47# 4.94e-20
C14822 _249_/a_27_297# net53 0.242f
C14823 VPWR _324_/a_639_47# 8.07e-19
C14824 fanout44/a_27_47# mask\[1\] 9.97e-21
C14825 _110_ _264_/a_27_297# 0.109f
C14826 _060_ _226_/a_27_47# 0.127f
C14827 _322_/a_193_47# net26 2.09e-20
C14828 net15 _092_ 0.167f
C14829 _235_/a_79_21# _092_ 0.0527f
C14830 _239_/a_474_297# _051_ 0.00417f
C14831 result[7] net14 0.0254f
C14832 trimb[3] net34 0.00164f
C14833 _104_ _331_/a_543_47# 1.29e-21
C14834 net12 _100_ 0.0959f
C14835 _321_/a_1283_21# _078_ 1.24e-21
C14836 VPWR _322_/a_1270_413# 7.93e-19
C14837 net2 net19 0.00927f
C14838 _064_ _258_/a_373_47# 6.38e-21
C14839 net42 clk 0.0128f
C14840 _104_ _258_/a_109_297# 0.0601f
C14841 _336_/a_27_47# _063_ 9.79e-21
C14842 _303_/a_651_413# net26 1.01e-19
C14843 _249_/a_27_297# _009_ 4.03e-20
C14844 net27 _084_ 0.14f
C14845 clknet_2_1__leaf_clk _046_ 0.0278f
C14846 VPWR ctlp[7] 0.639f
C14847 _051_ _206_/a_206_47# 5.53e-21
C14848 _269_/a_81_21# _333_/a_27_47# 0.00145f
C14849 _042_ net44 0.0115f
C14850 _030_ _333_/a_1283_21# 4.61e-20
C14851 _113_ _333_/a_1108_47# 3.38e-21
C14852 _338_/a_1602_47# _123_ 4.3e-20
C14853 _181_/a_150_297# _058_ 9.62e-19
C14854 net13 _318_/a_651_413# 0.00247f
C14855 _198_/a_109_47# _069_ 6.92e-19
C14856 net43 net26 0.0143f
C14857 _195_/a_218_374# _062_ 2.49e-20
C14858 VPWR _218_/a_199_47# 5.72e-19
C14859 VPWR _220_/a_113_297# 0.254f
C14860 net50 _335_/a_1462_47# 1.92e-19
C14861 cal_itt\[0\] _062_ 0.266f
C14862 _049_ _279_/a_490_47# 5.81e-20
C14863 net4 _096_ 3.61e-21
C14864 _229_/a_27_297# net55 6.38e-20
C14865 clknet_2_1__leaf_clk _312_/a_761_289# 4.98e-19
C14866 _110_ ctln[3] 1.44e-20
C14867 net22 net14 0.467f
C14868 _040_ net30 1.71e-20
C14869 _247_/a_27_297# mask\[2\] 0.0574f
C14870 _078_ _138_/a_27_47# 0.0117f
C14871 _308_/a_1283_21# net45 0.0158f
C14872 _308_/a_448_47# clknet_2_0__leaf_clk 0.00154f
C14873 net30 _279_/a_314_297# 2.29e-19
C14874 _326_/a_1283_21# net43 0.278f
C14875 _088_ _062_ 1.38e-19
C14876 _330_/a_805_47# net46 0.0019f
C14877 state\[0\] en_co_clk 0.00123f
C14878 _323_/a_543_47# clknet_2_1__leaf_clk 1.49e-19
C14879 _341_/a_448_47# _065_ 0.00802f
C14880 net9 _136_ 0.0501f
C14881 _218_/a_199_47# net53 4.92e-21
C14882 output37/a_27_47# net33 0.0101f
C14883 _337_/a_193_47# _282_/a_150_297# 1.24e-19
C14884 _015_ _243_/a_373_47# 7.21e-19
C14885 _237_/a_76_199# _014_ 7.24e-19
C14886 _237_/a_505_21# clknet_2_0__leaf_clk 7.15e-20
C14887 _198_/a_181_47# _067_ 0.00258f
C14888 _002_ _041_ 3.63e-20
C14889 _198_/a_181_47# _070_ 2.89e-20
C14890 VPWR _275_/a_299_297# 0.236f
C14891 _320_/a_1217_47# clknet_2_0__leaf_clk 1.2e-21
C14892 _334_/a_193_47# net46 0.042f
C14893 net15 _246_/a_109_297# 0.00523f
C14894 net25 _310_/a_27_47# 0.00131f
C14895 _216_/a_113_297# _310_/a_1108_47# 0.00151f
C14896 net31 trimb[4] 0.109f
C14897 _287_/a_75_212# _122_ 8.88e-21
C14898 _195_/a_76_199# _195_/a_218_374# 0.00557f
C14899 VPWR _178_/a_68_297# 0.171f
C14900 _315_/a_27_47# _241_/a_297_47# 1.52e-21
C14901 _290_/a_27_413# output37/a_27_47# 0.011f
C14902 cal_itt\[0\] _195_/a_76_199# 0.379f
C14903 ctlp[6] _045_ 6.87e-19
C14904 cal_itt\[2\] _195_/a_505_21# 3.68e-21
C14905 _328_/a_651_413# trim_mask\[1\] 0.0265f
C14906 _328_/a_1108_47# _112_ 1.1e-20
C14907 _189_/a_218_47# _107_ 6.77e-19
C14908 trim_mask\[2\] _112_ 6.44e-20
C14909 net51 _208_/a_439_47# 4.69e-19
C14910 trim_mask\[2\] _272_/a_299_297# 0.0586f
C14911 output7/a_27_47# ctln[1] 0.159f
C14912 _200_/a_303_47# _071_ 6.01e-19
C14913 VPWR _246_/a_373_47# 5.57e-19
C14914 net9 _340_/a_796_47# 5.14e-19
C14915 _319_/a_651_413# net52 3.39e-19
C14916 _319_/a_1108_47# _016_ 1.93e-19
C14917 _253_/a_384_47# _078_ 5.45e-19
C14918 _092_ _049_ 0.291f
C14919 _304_/a_27_47# _304_/a_761_289# 0.0701f
C14920 output15/a_27_47# _046_ 0.00266f
C14921 _188_/a_27_47# _130_ 5.13e-22
C14922 trim_mask\[2\] _336_/a_1283_21# 0.00755f
C14923 _095_ net30 1.44e-19
C14924 _307_/a_805_47# calibrate 3.52e-21
C14925 _334_/a_193_47# _334_/a_639_47# 2.28e-19
C14926 _334_/a_761_289# _334_/a_1270_413# 2.6e-19
C14927 _334_/a_543_47# _334_/a_651_413# 0.0572f
C14928 _168_/a_27_413# clk 0.00939f
C14929 _329_/a_193_47# trim_mask\[2\] 4.46e-19
C14930 _314_/a_761_289# _314_/a_639_47# 3.16e-19
C14931 _314_/a_27_47# _314_/a_1217_47# 2.56e-19
C14932 clone1/a_27_47# _260_/a_250_297# 7.24e-21
C14933 _296_/a_113_47# _131_ 7.51e-19
C14934 state\[2\] _232_/a_114_297# 2.02e-19
C14935 _263_/a_79_21# _100_ 2.66e-19
C14936 _339_/a_1140_413# cal_count\[0\] 1.36e-19
C14937 _320_/a_639_47# _065_ 2.56e-20
C14938 _327_/a_27_47# _327_/a_448_47# 0.0894f
C14939 _327_/a_193_47# _327_/a_1108_47# 0.125f
C14940 net42 _063_ 0.00633f
C14941 state\[0\] _050_ 5.44e-19
C14942 _336_/a_193_47# net19 0.014f
C14943 _335_/a_27_47# _027_ 6.08e-20
C14944 _051_ _033_ 4.8e-20
C14945 calibrate _241_/a_105_352# 9.55e-20
C14946 _307_/a_805_47# net45 0.00316f
C14947 _062_ _108_ 0.0054f
C14948 _308_/a_1283_21# _319_/a_27_47# 2.4e-19
C14949 _168_/a_207_413# _331_/a_543_47# 3.65e-21
C14950 _169_/a_215_311# _169_/a_109_53# 0.179f
C14951 _185_/a_150_297# _060_ 4.96e-19
C14952 _306_/a_761_289# _208_/a_505_21# 8.62e-21
C14953 _262_/a_27_47# _190_/a_27_47# 2.9e-21
C14954 _299_/a_298_297# _299_/a_382_47# 1.58e-20
C14955 state\[2\] clone1/a_27_47# 0.166f
C14956 fanout44/a_27_47# _244_/a_27_297# 2.31e-19
C14957 _292_/a_78_199# cal_count\[0\] 1.96e-20
C14958 _036_ _286_/a_76_199# 8.26e-20
C14959 _168_/a_27_413# net4 3.44e-21
C14960 VPWR _291_/a_285_297# 0.26f
C14961 _134_ net33 3.12e-20
C14962 net27 _085_ 0.0174f
C14963 _327_/a_1108_47# _058_ 0.0142f
C14964 VPWR _213_/a_109_297# 0.00725f
C14965 net45 _241_/a_105_352# 9.84e-19
C14966 _232_/a_32_297# _107_ 6.74e-19
C14967 _014_ _241_/a_388_297# 0.00855f
C14968 _048_ net41 2.36e-19
C14969 _064_ clknet_2_2__leaf_clk 0.246f
C14970 output25/a_27_47# _074_ 4.25e-19
C14971 _104_ _260_/a_256_47# 4.85e-19
C14972 _328_/a_193_47# net9 0.00793f
C14973 _304_/a_639_47# _122_ 0.00166f
C14974 _341_/a_193_47# _066_ 1.06e-20
C14975 _239_/a_474_297# _242_/a_79_21# 1.54e-19
C14976 _333_/a_1283_21# net33 0.00975f
C14977 _336_/a_193_47# _107_ 0.00241f
C14978 VPWR _222_/a_113_297# 0.261f
C14979 _021_ _312_/a_27_47# 3.92e-20
C14980 _340_/a_193_47# _122_ 0.00197f
C14981 _112_ _333_/a_761_289# 4.82e-19
C14982 net49 _333_/a_543_47# 0.00704f
C14983 _272_/a_299_297# _333_/a_761_289# 9.29e-21
C14984 trim_val\[1\] _333_/a_1108_47# 0.0209f
C14985 _115_ _112_ 0.00388f
C14986 _144_/a_27_47# net40 2.09e-19
C14987 _304_/a_193_47# net18 0.0092f
C14988 _115_ _272_/a_299_297# 5.06e-19
C14989 _273_/a_59_75# _114_ 0.18f
C14990 cal_count\[3\] _278_/a_27_47# 1.1e-19
C14991 result[0] result[1] 0.0489f
C14992 clknet_2_3__leaf_clk net40 0.00271f
C14993 _334_/a_1283_21# _108_ 4.38e-19
C14994 _310_/a_193_47# _310_/a_761_289# 0.181f
C14995 _310_/a_27_47# _310_/a_543_47# 0.115f
C14996 _104_ net19 0.122f
C14997 _329_/a_193_47# _115_ 7.12e-20
C14998 _327_/a_761_289# _108_ 2.33e-19
C14999 _046_ _313_/a_27_47# 0.0294f
C15000 _335_/a_27_47# _335_/a_448_47# 0.0931f
C15001 _335_/a_193_47# _335_/a_1108_47# 0.125f
C15002 VPWR rebuffer5/a_161_47# 0.595f
C15003 _005_ clknet_2_0__leaf_clk 0.00317f
C15004 fanout45/a_27_47# _316_/a_1108_47# 0.00133f
C15005 net55 net19 1.79e-20
C15006 mask\[1\] _247_/a_27_297# 4.05e-20
C15007 _079_ net14 0.0167f
C15008 _262_/a_193_297# _092_ 9.77e-20
C15009 _058_ rebuffer2/a_75_212# 0.005f
C15010 _303_/a_1283_21# _065_ 2.22e-20
C15011 ctln[4] trim_mask\[3\] 1.69e-19
C15012 net28 _011_ 0.0751f
C15013 _149_/a_68_297# clknet_2_3__leaf_clk 6.28e-21
C15014 _281_/a_103_199# _192_/a_505_280# 0.00113f
C15015 _103_ _051_ 0.0432f
C15016 _048_ _171_/a_27_47# 0.00273f
C15017 _058_ _332_/a_1283_21# 0.00241f
C15018 _078_ _101_ 1.01f
C15019 _304_/a_27_47# _302_/a_109_297# 4.56e-21
C15020 _304_/a_193_47# _302_/a_27_297# 3.45e-21
C15021 net9 _301_/a_129_47# 9.57e-21
C15022 net10 _057_ 8.16e-19
C15023 net13 _232_/a_32_297# 0.00856f
C15024 _334_/a_1462_47# net46 0.00288f
C15025 net15 _017_ 6.48e-20
C15026 _195_/a_218_47# _068_ 2.88e-19
C15027 net27 _314_/a_543_47# 9.2e-20
C15028 net9 _338_/a_1140_413# 1.04e-19
C15029 comp net37 8.58e-19
C15030 _327_/a_805_47# net46 0.00343f
C15031 _129_ _298_/a_493_297# 1.98e-20
C15032 net9 _341_/a_761_289# 7.52e-19
C15033 _336_/a_1108_47# trim_mask\[4\] 0.0389f
C15034 _104_ _107_ 0.0234f
C15035 _264_/a_27_297# clknet_2_2__leaf_clk 7.38e-19
C15036 net43 net2 3.18e-20
C15037 _304_/a_543_47# _304_/a_805_47# 0.00171f
C15038 _304_/a_761_289# _304_/a_1217_47# 4.2e-19
C15039 _304_/a_1108_47# _304_/a_1270_413# 0.00645f
C15040 _047_ net34 0.103f
C15041 _339_/a_381_47# _123_ 0.0146f
C15042 net5 _047_ 4.5e-19
C15043 net43 _305_/a_1283_21# 0.285f
C15044 _026_ _328_/a_27_47# 8.37e-20
C15045 _329_/a_1462_47# trim_mask\[2\] 5.43e-19
C15046 clk _316_/a_761_289# 2.77e-19
C15047 _336_/a_27_47# _279_/a_396_47# 0.00922f
C15048 _336_/a_193_47# _279_/a_27_47# 0.0013f
C15049 VPWR _212_/a_113_297# 0.241f
C15050 _235_/a_297_47# _226_/a_27_47# 0.0143f
C15051 _107_ net55 0.116f
C15052 _321_/a_27_47# _321_/a_761_289# 0.0535f
C15053 _332_/a_193_47# _108_ 0.397f
C15054 _332_/a_193_47# _332_/a_543_47# 0.21f
C15055 _332_/a_27_47# _332_/a_1283_21# 0.0427f
C15056 _067_ net19 0.0106f
C15057 net19 _070_ 0.0709f
C15058 _094_ _048_ 0.00253f
C15059 _335_/a_805_47# net46 0.00447f
C15060 _286_/a_505_21# _001_ 1.03e-19
C15061 _169_/a_301_53# state\[0\] 1.53e-19
C15062 net3 _317_/a_1283_21# 4.42e-20
C15063 _306_/a_448_47# _076_ 2.94e-20
C15064 clkbuf_0_clk/a_110_47# _304_/a_27_47# 8.33e-21
C15065 _276_/a_59_75# net18 4.1e-19
C15066 _320_/a_27_47# _078_ 3.44e-19
C15067 _304_/a_27_47# cal_count\[3\] 8.79e-21
C15068 _337_/a_27_47# _337_/a_761_289# 0.0701f
C15069 _136_ _122_ 0.00727f
C15070 output33/a_27_47# _333_/a_1283_21# 9.71e-21
C15071 _304_/a_1108_47# clknet_2_3__leaf_clk 1.68e-19
C15072 _036_ cal_count\[0\] 0.083f
C15073 _333_/a_27_47# net32 7.72e-20
C15074 net31 _030_ 1.25e-20
C15075 _257_/a_27_297# trim_mask\[1\] 0.18f
C15076 net9 _339_/a_27_47# 0.0159f
C15077 _309_/a_1108_47# clknet_2_1__leaf_clk 3.88e-21
C15078 state\[1\] _092_ 0.00946f
C15079 _302_/a_27_297# net18 0.0108f
C15080 VPWR _330_/a_639_47# 4.33e-19
C15081 result[2] _006_ 8.61e-19
C15082 _257_/a_109_297# _336_/a_193_47# 1.7e-19
C15083 _332_/a_639_47# net46 9.54e-19
C15084 _328_/a_1462_47# net9 2.57e-19
C15085 net50 net30 3.8e-20
C15086 _237_/a_535_374# _096_ 0.00526f
C15087 _048_ _192_/a_505_280# 0.155f
C15088 VPWR _267_/a_145_75# 3.29e-19
C15089 _104_ _279_/a_27_47# 1.94e-19
C15090 VPWR _200_/a_209_47# 2.27e-19
C15091 net3 _192_/a_174_21# 0.0689f
C15092 net47 _149_/a_150_297# 2.47e-19
C15093 _337_/a_448_47# clknet_0_clk 6.06e-21
C15094 net33 cal_count\[2\] 3.22e-19
C15095 _306_/a_27_47# rebuffer4/a_27_47# 7.75e-22
C15096 _094_ _120_ 0.0625f
C15097 VPWR _334_/a_27_47# 0.51f
C15098 _326_/a_193_47# _216_/a_113_297# 7.22e-21
C15099 VPWR _228_/a_382_297# 0.00468f
C15100 _324_/a_1283_21# _042_ 2.73e-20
C15101 net13 net55 0.314f
C15102 _314_/a_193_47# net29 0.00662f
C15103 result[6] clknet_2_1__leaf_clk 0.0373f
C15104 _307_/a_193_47# _078_ 0.0115f
C15105 _307_/a_543_47# net22 0.015f
C15106 _307_/a_761_289# mask\[0\] 7.07e-20
C15107 VPWR _325_/a_805_47# 3.44e-19
C15108 net21 _313_/a_639_47# 1.32e-19
C15109 _335_/a_27_47# _032_ 0.169f
C15110 _340_/a_1182_261# _129_ 5.56e-20
C15111 _282_/a_150_297# _090_ 2.4e-20
C15112 result[4] _310_/a_805_47# 1.99e-19
C15113 _226_/a_197_47# _049_ 7.09e-20
C15114 _311_/a_27_47# _311_/a_651_413# 9.73e-19
C15115 _311_/a_761_289# _311_/a_1108_47# 0.0512f
C15116 _311_/a_193_47# _311_/a_448_47# 0.0594f
C15117 _168_/a_207_413# _107_ 0.0022f
C15118 en _315_/a_27_47# 1.21e-19
C15119 _094_ _076_ 5.86e-20
C15120 _322_/a_543_47# _042_ 3.29e-20
C15121 state\[2\] _255_/a_27_47# 3.59e-21
C15122 _120_ _192_/a_505_280# 0.183f
C15123 en_co_clk _192_/a_476_47# 1.07e-19
C15124 _304_/a_27_47# _038_ 1.35e-20
C15125 _064_ _257_/a_373_47# 1.56e-20
C15126 _104_ _257_/a_109_297# 0.0322f
C15127 clk _098_ 3.92e-19
C15128 _103_ _242_/a_79_21# 7.62e-20
C15129 _307_/a_27_47# output30/a_27_47# 0.0123f
C15130 result[1] net23 0.00612f
C15131 _304_/a_448_47# net47 1.1e-20
C15132 _326_/a_27_47# _314_/a_543_47# 1.17e-20
C15133 _326_/a_193_47# _314_/a_761_289# 5.38e-22
C15134 _326_/a_761_289# _314_/a_193_47# 5.17e-21
C15135 _326_/a_543_47# _314_/a_27_47# 8.69e-21
C15136 trim_mask\[1\] trim_val\[4\] 0.00357f
C15137 _051_ clkbuf_2_3__f_clk/a_110_47# 0.00607f
C15138 _128_ net33 0.00162f
C15139 net43 _251_/a_373_47# 6.22e-20
C15140 trim_mask\[0\] net18 0.0149f
C15141 _230_/a_59_75# net4 0.012f
C15142 _336_/a_193_47# _118_ 3.81e-21
C15143 VPWR _314_/a_448_47# 0.0836f
C15144 _218_/a_113_297# clknet_2_1__leaf_clk 5.24e-19
C15145 _254_/a_109_297# _092_ 0.00184f
C15146 _321_/a_543_47# _321_/a_805_47# 0.00171f
C15147 _321_/a_761_289# _321_/a_1217_47# 4.2e-19
C15148 _321_/a_1108_47# _321_/a_1270_413# 0.00645f
C15149 _340_/a_27_47# _340_/a_562_413# 6.02e-19
C15150 _340_/a_193_47# _340_/a_381_47# 0.157f
C15151 _340_/a_476_47# _340_/a_1032_413# 0.00329f
C15152 _332_/a_448_47# _332_/a_639_47# 4.61e-19
C15153 clk clknet_0_clk 0.191f
C15154 _308_/a_543_47# net24 7.21e-21
C15155 net8 _273_/a_59_75# 7.89e-20
C15156 VPWR _169_/a_109_53# 0.138f
C15157 _008_ _250_/a_27_297# 2.07e-21
C15158 _059_ _060_ 0.654f
C15159 _048_ _014_ 1.92e-19
C15160 _292_/a_78_199# net16 5.04e-19
C15161 en clknet_2_0__leaf_clk 6.3e-20
C15162 _323_/a_27_47# _149_/a_68_297# 7.54e-19
C15163 net31 net33 0.485f
C15164 net54 net41 0.407f
C15165 net47 _133_ 1.57e-19
C15166 _337_/a_543_47# _337_/a_805_47# 0.00171f
C15167 _337_/a_761_289# _337_/a_1217_47# 4.2e-19
C15168 _337_/a_1108_47# _337_/a_1270_413# 0.00645f
C15169 net5 _301_/a_47_47# 7.27e-20
C15170 net31 trim_mask\[1\] 4.83e-19
C15171 net43 net55 0.00162f
C15172 VPWR _310_/a_761_289# 0.22f
C15173 _333_/a_1217_47# net32 7.32e-20
C15174 _088_ _227_/a_209_311# 0.0915f
C15175 _340_/a_476_47# cal_count\[3\] 1.54e-19
C15176 net9 _339_/a_586_47# 2.06e-19
C15177 net13 mask\[0\] 0.00197f
C15178 mask\[6\] _249_/a_27_297# 6.45e-20
C15179 _325_/a_193_47# _074_ 9.03e-20
C15180 trim_mask\[0\] _302_/a_27_297# 4.91e-21
C15181 _250_/a_27_297# mask\[5\] 0.101f
C15182 net31 _290_/a_27_413# 0.00589f
C15183 calibrate en_co_clk 0.00117f
C15184 _025_ _336_/a_193_47# 1.26e-20
C15185 net4 clknet_0_clk 0.12f
C15186 _035_ _338_/a_27_47# 0.114f
C15187 clknet_2_1__leaf_clk _246_/a_109_47# 0.0012f
C15188 _293_/a_299_297# _289_/a_68_297# 0.00117f
C15189 _247_/a_27_297# _247_/a_109_47# 0.00393f
C15190 _161_/a_150_297# net37 3.96e-19
C15191 _230_/a_59_75# _063_ 0.185f
C15192 _191_/a_27_297# net18 1.36e-19
C15193 _104_ _118_ 0.00748f
C15194 _338_/a_652_21# net18 0.0113f
C15195 _324_/a_448_47# _021_ 0.158f
C15196 _320_/a_193_47# _121_ 1.99e-19
C15197 VPWR _334_/a_1217_47# 1.01e-19
C15198 _324_/a_193_47# _078_ 1.08e-20
C15199 net45 en_co_clk 2.3e-20
C15200 en_co_clk rebuffer3/a_75_212# 1.38e-21
C15201 VPWR cal 0.226f
C15202 _314_/a_1462_47# net29 4.31e-19
C15203 VPWR _327_/a_639_47# 5.1e-19
C15204 net43 _067_ 0.00265f
C15205 net43 _070_ 6.25e-20
C15206 _335_/a_1217_47# _032_ 1.04e-20
C15207 _302_/a_373_47# _136_ 3.16e-19
C15208 _169_/a_215_311# _318_/a_193_47# 2.81e-20
C15209 cal valid 0.0947f
C15210 _307_/a_543_47# _079_ 4.49e-19
C15211 _307_/a_193_47# _004_ 0.223f
C15212 _129_ _297_/a_47_47# 0.0732f
C15213 output35/a_27_47# trim[4] 0.337f
C15214 net28 _313_/a_761_289# 0.022f
C15215 ctlp[7] mask\[6\] 5.34e-19
C15216 _078_ _248_/a_27_297# 4.2e-21
C15217 _322_/a_27_47# _078_ 0.0041f
C15218 _048_ _243_/a_27_297# 1.73e-20
C15219 clknet_0_clk net52 0.119f
C15220 en_co_clk _065_ 0.198f
C15221 _050_ calibrate 0.573f
C15222 clknet_0_clk _063_ 0.0459f
C15223 _104_ _025_ 0.00198f
C15224 trimb[2] output39/a_27_47# 0.00275f
C15225 output38/a_27_47# trimb[3] 9.86e-19
C15226 VPWR _335_/a_639_47# 7.26e-19
C15227 _339_/a_27_47# _122_ 6.27e-21
C15228 _135_ en_co_clk 0.00293f
C15229 VPWR ctln[5] 0.195f
C15230 _313_/a_193_47# _158_/a_150_297# 9.72e-20
C15231 VPWR comp 0.245f
C15232 VPWR _311_/a_1283_21# 0.362f
C15233 mask\[6\] _220_/a_113_297# 0.00553f
C15234 _250_/a_109_297# _084_ 1.14e-19
C15235 _143_/a_68_297# _143_/a_150_297# 0.00477f
C15236 _051_ clkbuf_0_clk/a_110_47# 4.12e-20
C15237 _051_ cal_count\[3\] 1.48e-20
C15238 result[0] sample 0.0473f
C15239 _050_ net45 4.41e-19
C15240 state\[0\] net15 0.0042f
C15241 net54 _094_ 0.0691f
C15242 _037_ _304_/a_651_413# 2.26e-19
C15243 _311_/a_1283_21# net53 2.38e-20
C15244 _097_ _092_ 0.0631f
C15245 net43 mask\[0\] 0.601f
C15246 _005_ _078_ 2.11e-19
C15247 net31 output33/a_27_47# 0.00225f
C15248 VPWR _332_/a_1270_413# 5.43e-19
C15249 cal_itt\[1\] net30 0.00168f
C15250 _340_/a_1182_261# _340_/a_1296_47# 1.84e-19
C15251 _340_/a_1032_413# _340_/a_1224_47# 0.00536f
C15252 _052_ _054_ 3.87e-19
C15253 trim[0] _173_/a_27_47# 2.73e-19
C15254 output31/a_27_47# net32 0.00155f
C15255 _051_ _331_/a_27_47# 0.0011f
C15256 VPWR net51 0.641f
C15257 _224_/a_113_297# _224_/a_199_47# 2.42e-19
C15258 _052_ net30 1.34e-20
C15259 _277_/a_75_212# _110_ 0.0273f
C15260 _232_/a_32_297# net3 0.00234f
C15261 _064_ _231_/a_161_47# 7e-19
C15262 _219_/a_109_297# _078_ 0.00526f
C15263 _308_/a_448_47# _004_ 1.79e-20
C15264 _281_/a_253_47# _096_ 2.32e-19
C15265 en_co_clk _243_/a_109_297# 7.06e-19
C15266 _337_/a_193_47# _090_ 2.84e-21
C15267 _007_ _074_ 0.117f
C15268 _253_/a_384_47# mask\[7\] 0.00918f
C15269 _253_/a_299_297# _102_ 0.0476f
C15270 _253_/a_81_21# _023_ 0.114f
C15271 _186_/a_109_297# net41 0.0113f
C15272 _309_/a_639_47# _078_ 9.62e-19
C15273 _187_/a_297_47# _058_ 1.5e-19
C15274 _064_ trim_mask\[3\] 0.394f
C15275 _323_/a_543_47# _043_ 1.57e-20
C15276 _323_/a_1283_21# net18 3.42e-19
C15277 _326_/a_651_413# _310_/a_543_47# 3.01e-20
C15278 _326_/a_1108_47# _310_/a_1108_47# 8.34e-21
C15279 _320_/a_761_289# clknet_0_clk 0.00358f
C15280 _337_/a_448_47# net44 2.85e-19
C15281 _309_/a_448_47# net24 0.0164f
C15282 _050_ _065_ 0.0226f
C15283 _110_ net4 0.326f
C15284 _338_/a_1602_47# clknet_2_3__leaf_clk 0.0097f
C15285 calibrate _228_/a_297_47# 6.83e-19
C15286 _042_ mask\[2\] 0.0316f
C15287 clknet_2_1__leaf_clk _208_/a_439_47# 5.61e-19
C15288 _060_ _192_/a_27_47# 1.36e-20
C15289 _239_/a_694_21# _048_ 0.111f
C15290 net43 _313_/a_448_47# 0.00219f
C15291 _074_ mask\[3\] 0.116f
C15292 _024_ _136_ 7.49e-19
C15293 net2 _062_ 1.3e-20
C15294 _035_ _338_/a_586_47# 3.33e-19
C15295 _247_/a_109_297# _018_ 0.00249f
C15296 net37 _132_ 0.00591f
C15297 _232_/a_304_297# en_co_clk 1.27e-19
C15298 _305_/a_27_47# rebuffer4/a_27_47# 8.38e-19
C15299 trim_val\[0\] net34 8.77e-19
C15300 _230_/a_145_75# _107_ 8.43e-20
C15301 _338_/a_1056_47# net18 4e-19
C15302 net47 net4 0.0335f
C15303 _050_ _319_/a_27_47# 1.58e-21
C15304 net12 clk 0.0267f
C15305 VPWR _224_/a_199_47# 3.34e-19
C15306 _189_/a_27_47# _075_ 4.85e-20
C15307 net13 _121_ 3.21e-20
C15308 cal_itt\[1\] _072_ 2.1e-20
C15309 _337_/a_1283_21# _263_/a_297_47# 1.43e-21
C15310 cal_itt\[0\] _150_/a_27_47# 4.47e-22
C15311 state\[0\] _049_ 4.22e-19
C15312 output23/a_27_47# _007_ 4.13e-20
C15313 _316_/a_27_47# _095_ 1.61e-19
C15314 _110_ _063_ 6.44e-20
C15315 clk _331_/a_1108_47# 9.3e-19
C15316 output14/a_27_47# net29 0.00225f
C15317 _231_/a_161_47# _264_/a_27_297# 3.44e-21
C15318 _258_/a_27_297# _119_ 9.01e-19
C15319 _099_ clone7/a_27_47# 7.04e-20
C15320 _314_/a_543_47# _011_ 0.00291f
C15321 net12 _331_/a_1283_21# 0.00486f
C15322 _311_/a_1270_413# net26 4.38e-19
C15323 _030_ _058_ 0.00101f
C15324 _322_/a_1217_47# _078_ 1.61e-19
C15325 _064_ _330_/a_1283_21# 1.96e-19
C15326 _104_ _330_/a_761_289# 3.01e-20
C15327 _306_/a_193_47# _306_/a_1108_47# 0.125f
C15328 _306_/a_27_47# _306_/a_448_47# 0.0931f
C15329 mask\[6\] _222_/a_113_297# 0.0504f
C15330 cal_itt\[2\] _305_/a_543_47# 9.12e-20
C15331 _329_/a_651_413# trim_mask\[3\] 6.01e-19
C15332 _326_/a_1283_21# result[5] 1.47e-19
C15333 net12 net4 0.00967f
C15334 _035_ _339_/a_193_47# 7.63e-21
C15335 _331_/a_193_47# _331_/a_1270_413# 1.46e-19
C15336 _331_/a_27_47# _331_/a_639_47# 0.00188f
C15337 _331_/a_543_47# _331_/a_448_47# 0.0498f
C15338 _331_/a_761_289# _331_/a_651_413# 0.0977f
C15339 _331_/a_1283_21# _331_/a_1108_47# 0.234f
C15340 net3 net55 0.134f
C15341 fanout46/a_27_47# net46 0.347f
C15342 clk net44 0.00764f
C15343 _245_/a_27_297# net52 0.192f
C15344 _245_/a_109_47# _101_ 0.00145f
C15345 _143_/a_150_297# net52 1.32e-19
C15346 trim_mask\[4\] net18 0.366f
C15347 _256_/a_373_47# clknet_2_2__leaf_clk 0.00102f
C15348 _325_/a_1108_47# _042_ 1.08e-19
C15349 net47 _063_ 0.0107f
C15350 mask\[3\] _146_/a_150_297# 2.27e-19
C15351 _041_ _338_/a_27_47# 4.85e-19
C15352 clknet_2_3__leaf_clk net19 0.0276f
C15353 net47 _338_/a_381_47# 0.0215f
C15354 _308_/a_27_47# _138_/a_27_47# 0.0116f
C15355 _059_ _235_/a_297_47# 1.17e-19
C15356 _338_/a_27_47# _338_/a_1182_261# 0.0608f
C15357 _338_/a_193_47# _338_/a_476_47# 0.196f
C15358 _328_/a_193_47# _258_/a_27_297# 8.11e-20
C15359 _328_/a_27_47# _258_/a_109_297# 3.66e-19
C15360 _328_/a_1283_21# trim_mask\[0\] 4.74e-19
C15361 cal _315_/a_543_47# 0.00152f
C15362 _113_ _332_/a_193_47# 1.3e-20
C15363 _037_ net47 0.00229f
C15364 mask\[7\] _101_ 0.132f
C15365 _292_/a_292_297# _122_ 4.41e-20
C15366 net19 _153_/a_27_47# 0.118f
C15367 _325_/a_639_47# clknet_2_1__leaf_clk 3.39e-19
C15368 _074_ _310_/a_1283_21# 0.0107f
C15369 _317_/a_27_47# net41 1.11e-20
C15370 _326_/a_761_289# output14/a_27_47# 2.73e-21
C15371 _327_/a_805_47# _111_ 1.11e-19
C15372 _002_ _076_ 1.23e-19
C15373 _239_/a_27_297# _050_ 0.148f
C15374 _005_ _004_ 0.00243f
C15375 net31 _270_/a_59_75# 2.36e-20
C15376 trim[0] _172_/a_68_297# 5.41e-20
C15377 _259_/a_27_297# _058_ 1.34e-20
C15378 _064_ _181_/a_68_297# 0.00196f
C15379 result[4] _074_ 2.42e-19
C15380 _048_ _106_ 0.275f
C15381 output31/a_27_47# output32/a_27_47# 1.88e-19
C15382 net9 _057_ 0.0755f
C15383 _259_/a_109_297# _335_/a_27_47# 8.28e-19
C15384 _259_/a_27_297# _335_/a_193_47# 3.27e-19
C15385 _022_ mask\[2\] 9.54e-25
C15386 net12 net52 4.96e-20
C15387 _269_/a_299_297# net46 0.00155f
C15388 _302_/a_27_297# trim_mask\[4\] 1.27e-19
C15389 _341_/a_1283_21# cal_count\[3\] 0.108f
C15390 _107_ clknet_2_3__leaf_clk 0.00643f
C15391 _341_/a_639_47# clknet_2_3__leaf_clk 0.00133f
C15392 net2 _332_/a_193_47# 2.47e-19
C15393 calibrate net1 0.00394f
C15394 net43 _121_ 0.0321f
C15395 ctlp[6] ctlp[5] 1.96e-20
C15396 net43 _010_ 0.015f
C15397 fanout46/a_27_47# _335_/a_651_413# 1.44e-19
C15398 _116_ net19 0.00268f
C15399 clknet_0_clk _279_/a_396_47# 1.14e-20
C15400 _042_ mask\[1\] 0.00296f
C15401 net26 net29 2.24e-20
C15402 trim_mask\[1\] _334_/a_543_47# 8.39e-22
C15403 _272_/a_81_21# _334_/a_761_289# 6.84e-20
C15404 _272_/a_299_297# _334_/a_193_47# 4.55e-20
C15405 net34 _131_ 0.0115f
C15406 VPWR _161_/a_150_297# 0.00225f
C15407 _053_ _262_/a_109_297# 0.00481f
C15408 net5 _131_ 0.00988f
C15409 net17 _041_ 1.18e-20
C15410 _327_/a_193_47# trim_mask\[1\] 9.96e-21
C15411 clknet_2_1__leaf_clk _314_/a_1108_47# 4.87e-19
C15412 _303_/a_193_47# _035_ 1.09e-21
C15413 net1 net45 1.51e-20
C15414 _051_ _242_/a_297_47# 1.36e-20
C15415 _074_ fanout43/a_27_47# 1.42e-19
C15416 _227_/a_209_311# _227_/a_368_53# 0.0026f
C15417 trim_mask\[0\] _333_/a_193_47# 1.91e-19
C15418 _104_ _062_ 4.39e-20
C15419 net44 net52 0.0125f
C15420 _294_/a_68_297# _129_ 4.36e-19
C15421 net44 _063_ 1.71e-20
C15422 _081_ _214_/a_113_297# 0.0913f
C15423 VPWR _318_/a_193_47# 0.291f
C15424 trim_mask\[0\] _265_/a_81_21# 0.112f
C15425 net27 _074_ 0.119f
C15426 _059_ net30 1.8e-20
C15427 _058_ net33 0.0312f
C15428 _146_/a_68_297# _310_/a_1108_47# 3.64e-19
C15429 net45 _039_ 0.214f
C15430 clk clknet_2_2__leaf_clk 0.0052f
C15431 net54 _243_/a_27_297# 0.00149f
C15432 _058_ trim_mask\[1\] 0.00544f
C15433 _323_/a_639_47# net47 9.54e-19
C15434 _339_/a_381_47# clknet_2_3__leaf_clk 6.75e-19
C15435 output24/a_27_47# _080_ 8.56e-20
C15436 net55 _062_ 0.00671f
C15437 _312_/a_651_413# net20 0.00219f
C15438 _096_ _075_ 5.91e-20
C15439 clknet_2_1__leaf_clk _310_/a_193_47# 0.596f
C15440 _299_/a_298_297# _131_ 8.44e-19
C15441 _136_ _134_ 0.00622f
C15442 _000_ fanout47/a_27_47# 1.13e-19
C15443 fanout44/a_27_47# net55 4.46e-19
C15444 VPWR _233_/a_27_297# 0.242f
C15445 _326_/a_761_289# net26 7.11e-20
C15446 _341_/a_1270_413# _136_ 8.32e-20
C15447 _341_/a_1283_21# _038_ 1.39e-19
C15448 _235_/a_382_297# _094_ 0.0159f
C15449 cal_itt\[0\] _042_ 1.18e-20
C15450 _331_/a_1283_21# clknet_2_2__leaf_clk 5.33e-20
C15451 _161_/a_68_297# _161_/a_150_297# 0.00477f
C15452 _331_/a_543_47# _028_ 0.0336f
C15453 net15 _317_/a_651_413# 0.00245f
C15454 _317_/a_27_47# _317_/a_448_47# 0.0931f
C15455 _317_/a_193_47# _317_/a_1108_47# 0.119f
C15456 _325_/a_805_47# mask\[6\] 0.00211f
C15457 _325_/a_1108_47# _022_ 1.61e-19
C15458 cal_itt\[0\] _064_ 2.64e-19
C15459 _233_/a_27_297# valid 0.00378f
C15460 _258_/a_109_47# clknet_2_2__leaf_clk 0.00309f
C15461 _332_/a_27_47# net33 7.1e-21
C15462 _326_/a_193_47# _326_/a_1108_47# 0.125f
C15463 _326_/a_27_47# _326_/a_448_47# 0.0931f
C15464 _325_/a_761_289# _078_ 1.14e-21
C15465 trim_mask\[0\] trim_mask\[4\] 0.115f
C15466 _046_ net21 0.0115f
C15467 cal_count\[1\] net34 1.15e-20
C15468 _306_/a_651_413# _049_ 5.46e-20
C15469 net54 _232_/a_220_297# 0.00188f
C15470 _308_/a_639_47# net14 7.18e-19
C15471 _341_/a_27_47# _063_ 2.69e-20
C15472 net49 rebuffer1/a_75_212# 2.47e-19
C15473 net4 clknet_2_2__leaf_clk 0.744f
C15474 VPWR _317_/a_639_47# 1.75e-20
C15475 _338_/a_652_21# _338_/a_1056_47# 3.94e-19
C15476 _338_/a_476_47# _338_/a_796_47# 0.00184f
C15477 _338_/a_1032_413# _338_/a_1140_413# 0.00523f
C15478 _338_/a_381_47# _338_/a_562_413# 8.75e-19
C15479 _328_/a_543_47# _328_/a_1108_47# 7.99e-20
C15480 _328_/a_193_47# _328_/a_651_413# 0.0276f
C15481 VPWR _326_/a_639_47# 0.00132f
C15482 _306_/a_1108_47# net30 6.43e-20
C15483 _320_/a_761_289# net44 0.159f
C15484 output23/a_27_47# fanout43/a_27_47# 1.78e-20
C15485 state\[0\] state\[1\] 0.215f
C15486 result[7] _314_/a_27_47# 0.00352f
C15487 _277_/a_75_212# net11 4.84e-20
C15488 _067_ _062_ 0.302f
C15489 _062_ _070_ 3.11e-20
C15490 _331_/a_448_47# net19 5.77e-19
C15491 net13 _337_/a_1270_413# 6.96e-20
C15492 _088_ _100_ 3.2e-19
C15493 _309_/a_193_47# net14 0.0121f
C15494 _170_/a_384_47# _054_ 1.88e-20
C15495 _340_/a_193_47# cal_count\[2\] 1.45e-19
C15496 _318_/a_27_47# _318_/a_193_47# 0.887f
C15497 _034_ clknet_0_clk 0.127f
C15498 _078_ _077_ 0.015f
C15499 _282_/a_68_297# en_co_clk 2.2e-21
C15500 state\[2\] _087_ 0.00261f
C15501 _325_/a_1283_21# _313_/a_1108_47# 8.78e-21
C15502 VPWR _192_/a_639_47# 6.94e-20
C15503 cal_count\[1\] _299_/a_298_297# 6.02e-20
C15504 _104_ _335_/a_761_289# 0.00234f
C15505 _064_ _335_/a_1283_21# 0.00209f
C15506 _086_ _224_/a_113_297# 0.0985f
C15507 net44 _312_/a_1270_413# 3.47e-19
C15508 _110_ _279_/a_396_47# 0.00346f
C15509 VPWR _300_/a_377_297# 0.00591f
C15510 _312_/a_27_47# _312_/a_448_47# 0.0931f
C15511 _312_/a_193_47# _312_/a_1108_47# 0.125f
C15512 _336_/a_651_413# net46 0.0122f
C15513 _286_/a_76_199# _286_/a_218_47# 0.00783f
C15514 _306_/a_193_47# clknet_2_0__leaf_clk 0.00196f
C15515 _320_/a_1108_47# _101_ 1.13e-19
C15516 _320_/a_543_47# net52 4.37e-19
C15517 _195_/a_76_199# _067_ 0.187f
C15518 clknet_2_1__leaf_clk _311_/a_543_47# 3.51e-20
C15519 _329_/a_1283_21# net46 0.35f
C15520 _323_/a_639_47# net44 4.2e-19
C15521 _303_/a_651_413# clknet_2_3__leaf_clk 8.49e-19
C15522 output8/a_27_47# _057_ 0.0648f
C15523 VPWR _262_/a_109_297# 0.16f
C15524 _323_/a_27_47# net19 0.0156f
C15525 _133_ _131_ 0.00247f
C15526 cal_itt\[1\] _066_ 9.54e-25
C15527 _041_ _339_/a_193_47# 0.275f
C15528 net47 _339_/a_562_413# 2.38e-19
C15529 _266_/a_68_297# net19 0.00778f
C15530 net48 _334_/a_1108_47# 4.81e-19
C15531 VPWR _132_ 0.778f
C15532 _188_/a_27_47# en_co_clk 0.00106f
C15533 _323_/a_543_47# _323_/a_1108_47# 7.99e-20
C15534 _323_/a_193_47# _323_/a_651_413# 0.0276f
C15535 net2 rebuffer6/a_27_47# 4.99e-20
C15536 _064_ _108_ 0.06f
C15537 _336_/a_639_47# _052_ 4.96e-21
C15538 _182_/a_27_47# net32 1.88e-19
C15539 VPWR _315_/a_1283_21# 0.404f
C15540 _306_/a_448_47# cal_itt\[3\] 1.38e-19
C15541 _306_/a_1108_47# _072_ 4.11e-19
C15542 _337_/a_1283_21# _099_ 1.09e-21
C15543 _337_/a_543_47# _092_ 3.51e-19
C15544 net50 net40 0.0315f
C15545 net14 net6 0.0989f
C15546 _328_/a_1108_47# _333_/a_27_47# 1.39e-19
C15547 fanout44/a_27_47# mask\[0\] 4.45e-19
C15548 net20 _155_/a_68_297# 2.23e-19
C15549 VPWR _318_/a_1462_47# 0.00178f
C15550 _242_/a_79_21# _242_/a_297_47# 0.0326f
C15551 _315_/a_448_47# net41 5.39e-20
C15552 _110_ _257_/a_109_47# 2.49e-21
C15553 _315_/a_1283_21# valid 1.44e-19
C15554 _306_/a_761_289# net2 3.19e-21
C15555 state\[2\] _263_/a_297_47# 1.72e-20
C15556 _292_/a_215_47# _340_/a_1032_413# 8.4e-19
C15557 _314_/a_1108_47# _313_/a_27_47# 1.43e-20
C15558 cal_count\[0\] trimb[4] 5.67e-20
C15559 _050_ _282_/a_68_297# 1.25e-19
C15560 calibrate net15 0.00828f
C15561 _235_/a_79_21# calibrate 1.35e-20
C15562 _306_/a_1283_21# _305_/a_761_289# 0.00118f
C15563 _306_/a_1108_47# _305_/a_193_47# 2.86e-19
C15564 ctln[7] clk 1.18e-20
C15565 _302_/a_109_47# _092_ 0.00216f
C15566 net30 _203_/a_59_75# 0.0435f
C15567 _266_/a_68_297# _107_ 0.00884f
C15568 VPWR _086_ 0.158f
C15569 _326_/a_27_47# _074_ 0.019f
C15570 _002_ _068_ 6.92e-19
C15571 _320_/a_761_289# _320_/a_543_47# 0.21f
C15572 _320_/a_193_47# _320_/a_1283_21# 0.0424f
C15573 _320_/a_27_47# _320_/a_1108_47# 0.102f
C15574 net37 net32 0.129f
C15575 _192_/a_476_47# _049_ 1.44e-19
C15576 _275_/a_299_297# net18 0.00664f
C15577 _311_/a_1283_21# _202_/a_79_21# 5.95e-21
C15578 _178_/a_68_297# net18 0.00254f
C15579 clknet_2_3__leaf_clk _118_ 5.75e-20
C15580 _331_/a_805_47# trim_mask\[4\] 1.36e-19
C15581 net7 clknet_2_0__leaf_clk 2.04e-20
C15582 net15 net45 1.2f
C15583 cal_count\[1\] _133_ 0.00162f
C15584 net52 _209_/a_27_47# 8.83e-19
C15585 _317_/a_27_47# _014_ 0.17f
C15586 _317_/a_193_47# clknet_2_0__leaf_clk 0.584f
C15587 net3 _121_ 1.77e-21
C15588 _308_/a_27_47# _307_/a_193_47# 1.21e-19
C15589 _308_/a_193_47# _307_/a_27_47# 6.5e-21
C15590 _328_/a_639_47# clknet_2_2__leaf_clk 5.75e-19
C15591 VPWR _269_/a_81_21# 0.27f
C15592 _337_/a_651_413# _034_ 7.15e-19
C15593 _136_ cal_count\[2\] 9.64e-19
C15594 _341_/a_543_47# _341_/a_651_413# 0.0572f
C15595 _341_/a_761_289# _341_/a_1270_413# 2.6e-19
C15596 _341_/a_193_47# _341_/a_639_47# 2.28e-19
C15597 _189_/a_27_47# _170_/a_81_21# 1.01e-20
C15598 clk net6 0.00704f
C15599 _264_/a_27_297# _108_ 0.258f
C15600 _303_/a_193_47# _041_ 1.89e-19
C15601 net47 _303_/a_1270_413# 1.81e-19
C15602 _303_/a_1108_47# _338_/a_27_47# 3.5e-19
C15603 _303_/a_1283_21# _338_/a_193_47# 1.98e-19
C15604 _304_/a_27_47# en_co_clk 7.65e-20
C15605 _315_/a_27_47# net30 8.1e-21
C15606 mask\[0\] _137_/a_68_297# 0.163f
C15607 net22 _137_/a_150_297# 1.11e-20
C15608 _028_ net19 0.00127f
C15609 _333_/a_193_47# _175_/a_68_297# 8.23e-20
C15610 net4 _279_/a_204_297# 0.00404f
C15611 net16 rebuffer2/a_75_212# 0.00604f
C15612 _333_/a_27_47# _333_/a_761_289# 0.0701f
C15613 _257_/a_27_297# _119_ 1.41e-19
C15614 net15 _065_ 0.00704f
C15615 net16 _332_/a_1283_21# 0.00684f
C15616 _318_/a_543_47# _318_/a_639_47# 0.0138f
C15617 _318_/a_193_47# _318_/a_1217_47# 2.36e-20
C15618 _318_/a_761_289# _318_/a_805_47# 3.69e-19
C15619 _290_/a_207_413# _125_ 0.0677f
C15620 _265_/a_81_21# _333_/a_193_47# 2.14e-21
C15621 net8 output34/a_27_47# 0.00119f
C15622 _233_/a_109_297# _315_/a_761_289# 3.22e-19
C15623 _233_/a_27_297# _315_/a_543_47# 0.00338f
C15624 _203_/a_59_75# _072_ 0.149f
C15625 _203_/a_145_75# cal_itt\[3\] 0.00121f
C15626 _309_/a_543_47# _101_ 3.1e-20
C15627 rstn ctln[0] 2.27e-19
C15628 net4 net6 0.0663f
C15629 _324_/a_543_47# net44 0.164f
C15630 _324_/a_193_47# _312_/a_27_47# 1.15e-19
C15631 _324_/a_27_47# _312_/a_193_47# 2.78e-21
C15632 calibrate _049_ 0.236f
C15633 VPWR _305_/a_639_47# 3.35e-19
C15634 _185_/a_68_297# _316_/a_193_47# 2.13e-20
C15635 _308_/a_193_47# _308_/a_1108_47# 0.125f
C15636 _308_/a_27_47# _308_/a_448_47# 0.0894f
C15637 net51 _206_/a_27_93# 8.31e-21
C15638 _323_/a_1217_47# net19 2.55e-19
C15639 _041_ _339_/a_796_47# 0.00181f
C15640 _107_ _028_ 7.9e-19
C15641 net15 _319_/a_27_47# 0.0217f
C15642 _307_/a_193_47# _307_/a_448_47# 0.0642f
C15643 _307_/a_761_289# _307_/a_1108_47# 0.0512f
C15644 _307_/a_27_47# _307_/a_651_413# 9.73e-19
C15645 _305_/a_193_47# _203_/a_59_75# 6.15e-20
C15646 _333_/a_448_47# clknet_2_2__leaf_clk 1.96e-20
C15647 trim[0] _047_ 5.54e-19
C15648 _304_/a_448_47# _001_ 0.177f
C15649 _235_/a_79_21# _243_/a_109_297# 2.02e-20
C15650 result[0] _307_/a_761_289# 5.27e-19
C15651 VPWR clknet_2_1__leaf_clk 6.38f
C15652 net45 _049_ 0.00196f
C15653 VPWR _319_/a_761_289# 0.225f
C15654 _322_/a_761_289# net44 0.186f
C15655 net28 _101_ 5.23e-20
C15656 _329_/a_651_413# _031_ 1.38e-19
C15657 _300_/a_47_47# _300_/a_377_297# 0.00899f
C15658 _318_/a_761_289# net45 0.166f
C15659 _233_/a_109_297# calibrate 0.0387f
C15660 _233_/a_109_47# _074_ 0.00145f
C15661 _233_/a_27_297# _093_ 0.205f
C15662 _289_/a_68_297# _125_ 0.00518f
C15663 _126_ _288_/a_59_75# 0.0258f
C15664 clknet_2_0__leaf_clk net30 1.38f
C15665 _270_/a_59_75# _058_ 0.00281f
C15666 _321_/a_1108_47# _083_ 4.68e-23
C15667 VPWR _243_/a_373_47# 2.85e-19
C15668 _325_/a_27_47# _321_/a_27_47# 1.3e-21
C15669 _324_/a_448_47# _101_ 4.94e-21
C15670 net43 _081_ 0.00795f
C15671 output32/a_27_47# _182_/a_27_47# 0.0126f
C15672 _078_ _310_/a_1108_47# 0.0108f
C15673 clknet_2_1__leaf_clk net53 0.87f
C15674 _326_/a_448_47# _011_ 2.6e-20
C15675 clkbuf_2_2__f_clk/a_110_47# _330_/a_651_413# 2.2e-19
C15676 result[2] _310_/a_27_47# 7.53e-20
C15677 _306_/a_27_47# _002_ 0.00358f
C15678 _233_/a_109_297# net45 0.00122f
C15679 _337_/a_27_47# en_co_clk 0.00754f
C15680 VPWR _197_/a_199_47# 9.94e-19
C15681 _262_/a_27_47# _262_/a_109_297# 0.0961f
C15682 state\[0\] _097_ 4.23e-21
C15683 _320_/a_1283_21# _320_/a_1462_47# 0.0074f
C15684 _320_/a_1108_47# _320_/a_1217_47# 0.00742f
C15685 _119_ trim_val\[4\] 5.48e-20
C15686 _001_ _133_ 5.05e-20
C15687 _065_ _049_ 0.339f
C15688 clkbuf_2_0__f_clk/a_110_47# _192_/a_174_21# 4.98e-19
C15689 _323_/a_1283_21# _303_/a_543_47# 3.62e-19
C15690 _323_/a_27_47# _303_/a_651_413# 4.77e-20
C15691 _323_/a_651_413# _303_/a_27_47# 2.28e-20
C15692 net50 _256_/a_109_47# 2.29e-19
C15693 input1/a_75_212# _316_/a_27_47# 4.41e-21
C15694 _322_/a_1108_47# _101_ 0.0104f
C15695 _339_/a_27_47# _339_/a_1602_47# 2.39e-19
C15696 _339_/a_193_47# _339_/a_1032_413# 0.0573f
C15697 net13 _320_/a_1283_21# 0.0124f
C15698 _270_/a_59_75# _332_/a_27_47# 7.88e-19
C15699 output32/a_27_47# net37 0.00802f
C15700 clknet_2_1__leaf_clk _009_ 0.113f
C15701 _187_/a_297_47# _061_ 0.001f
C15702 _317_/a_805_47# net45 0.00316f
C15703 _305_/a_1108_47# net30 8.45e-20
C15704 _105_ _049_ 0.00221f
C15705 _320_/a_193_47# _040_ 0.0371f
C15706 net44 _034_ 7.88e-19
C15707 VPWR _202_/a_382_297# 0.00587f
C15708 _321_/a_448_47# mask\[2\] 6.41e-20
C15709 _315_/a_27_47# _315_/a_651_413# 9.73e-19
C15710 _315_/a_761_289# _315_/a_1108_47# 0.0512f
C15711 _315_/a_193_47# _315_/a_448_47# 0.0642f
C15712 clknet_2_2__leaf_clk _279_/a_396_47# 5.22e-19
C15713 VPWR _336_/a_448_47# 0.0833f
C15714 VPWR output15/a_27_47# 0.242f
C15715 _110_ trim_val\[3\] 0.211f
C15716 _303_/a_639_47# _063_ 3.94e-20
C15717 VPWR _329_/a_543_47# 0.229f
C15718 net8 _334_/a_1283_21# 0.0111f
C15719 _319_/a_27_47# _049_ 0.0011f
C15720 _323_/a_448_47# _152_/a_68_297# 1.63e-20
C15721 net37 clkc 5.01e-19
C15722 _333_/a_1108_47# _333_/a_1270_413# 0.00645f
C15723 _333_/a_761_289# _333_/a_1217_47# 4.2e-19
C15724 _333_/a_543_47# _333_/a_805_47# 0.00171f
C15725 _100_ _170_/a_299_297# 8.93e-20
C15726 _243_/a_109_297# _049_ 0.00162f
C15727 net43 _016_ 8.35e-19
C15728 _312_/a_761_289# _045_ 6.66e-20
C15729 VPWR _239_/a_474_297# 0.136f
C15730 _037_ _131_ 1.12e-19
C15731 _050_ _337_/a_27_47# 1.51e-19
C15732 trim_val\[0\] _333_/a_448_47# 5.91e-20
C15733 _104_ _227_/a_209_311# 1.02e-19
C15734 _286_/a_505_21# _123_ 0.136f
C15735 net19 _279_/a_314_297# 0.00139f
C15736 net42 _170_/a_81_21# 7.65e-19
C15737 _042_ net26 0.0409f
C15738 _012_ _315_/a_761_289# 8.16e-19
C15739 _074_ _315_/a_448_47# 0.00471f
C15740 calibrate _315_/a_1108_47# 0.0542f
C15741 _200_/a_209_297# clkbuf_2_3__f_clk/a_110_47# 2.65e-19
C15742 _320_/a_1283_21# _248_/a_109_297# 1.26e-21
C15743 _337_/a_1108_47# _226_/a_27_47# 9.99e-20
C15744 _322_/a_193_47# _320_/a_1283_21# 1.65e-20
C15745 _322_/a_27_47# _320_/a_1108_47# 3.32e-20
C15746 _326_/a_1108_47# _251_/a_27_297# 2.95e-19
C15747 VPWR _206_/a_206_47# 1.43e-19
C15748 _260_/a_93_21# _092_ 1.12e-20
C15749 _324_/a_1108_47# net19 0.00166f
C15750 _227_/a_209_311# net55 0.0971f
C15751 _246_/a_27_297# _101_ 0.147f
C15752 _124_ _065_ 5.23e-20
C15753 _060_ _316_/a_1283_21# 6.36e-21
C15754 net54 _316_/a_1108_47# 2.02e-20
C15755 _308_/a_27_47# _005_ 0.213f
C15756 VPWR _210_/a_113_297# 0.252f
C15757 _328_/a_27_47# _025_ 0.389f
C15758 _143_/a_68_297# mask\[2\] 0.201f
C15759 _232_/a_304_297# _049_ 0.014f
C15760 _094_ _319_/a_1283_21# 1.33e-20
C15761 net15 _319_/a_1217_47# 6.04e-20
C15762 _014_ _315_/a_448_47# 1.1e-21
C15763 net45 _315_/a_1108_47# 0.245f
C15764 _305_/a_1108_47# _072_ 0.059f
C15765 _074_ _011_ 0.1f
C15766 clknet_0_clk _075_ 0.261f
C15767 net50 _280_/a_75_212# 6.72e-19
C15768 _107_ _279_/a_314_297# 0.00207f
C15769 ctlp[1] net29 5.91e-19
C15770 calibrate _012_ 0.189f
C15771 _336_/a_761_289# net30 2.25e-21
C15772 state\[2\] _099_ 1.26e-19
C15773 net23 _320_/a_193_47# 6.01e-21
C15774 net43 _320_/a_1283_21# 3.85e-19
C15775 net16 trimb[4] 3e-20
C15776 _323_/a_543_47# mask\[4\] 8.93e-19
C15777 _321_/a_27_47# net25 9.67e-20
C15778 input2/a_27_47# net40 2.19e-20
C15779 _305_/a_193_47# _305_/a_1108_47# 0.119f
C15780 _305_/a_27_47# _305_/a_448_47# 0.0867f
C15781 net12 _208_/a_76_199# 0.0113f
C15782 clkbuf_2_2__f_clk/a_110_47# net46 0.0262f
C15783 VPWR _313_/a_27_47# 0.441f
C15784 clone1/a_27_47# net30 5.12e-21
C15785 _309_/a_27_47# _309_/a_193_47# 0.887f
C15786 _239_/a_27_297# _049_ 0.012f
C15787 _277_/a_75_212# trim_mask\[3\] 3.63e-19
C15788 _103_ _053_ 9.49e-19
C15789 calibrate state\[1\] 0.00217f
C15790 _012_ net45 6.1e-19
C15791 _337_/a_1217_47# en_co_clk 3.92e-19
C15792 _262_/a_193_297# _105_ 0.00869f
C15793 _303_/a_805_47# net19 6.71e-19
C15794 _231_/a_161_47# net4 0.005f
C15795 VPWR net32 0.552f
C15796 _332_/a_1283_21# net40 1.44e-20
C15797 _051_ en_co_clk 0.00346f
C15798 _275_/a_81_21# trim_mask\[2\] 2.87e-21
C15799 trim_mask\[3\] _258_/a_109_47# 0.00216f
C15800 _323_/a_193_47# _000_ 2.54e-19
C15801 _320_/a_27_47# _246_/a_27_297# 2.32e-20
C15802 net1 _316_/a_448_47# 1.29e-20
C15803 cal_itt\[2\] clknet_0_clk 0.186f
C15804 trim_mask\[3\] net4 9.76e-21
C15805 _019_ _041_ 8.1e-20
C15806 net34 _108_ 0.00839f
C15807 _149_/a_68_297# _311_/a_27_47# 1.72e-21
C15808 net45 state\[1\] 0.105f
C15809 net43 _307_/a_1108_47# 1.76e-19
C15810 _005_ _307_/a_448_47# 2.65e-19
C15811 _320_/a_1462_47# _040_ 6.28e-19
C15812 cal_itt\[1\] _304_/a_1108_47# 0.00177f
C15813 _062_ clknet_2_3__leaf_clk 0.177f
C15814 net44 _208_/a_76_199# 2.12e-20
C15815 result[0] net43 6.17e-20
C15816 VPWR _033_ 0.844f
C15817 _101_ _084_ 1.37e-19
C15818 net13 _040_ 0.171f
C15819 _168_/a_207_413# _227_/a_209_311# 3.67e-21
C15820 _128_ _339_/a_27_47# 6.99e-19
C15821 _119_ _330_/a_193_47# 2.15e-19
C15822 cal_count\[0\] net33 0.00507f
C15823 net4 _001_ 0.0163f
C15824 _313_/a_27_47# _009_ 1.71e-21
C15825 _319_/a_1217_47# _049_ 5.28e-20
C15826 _166_/a_161_47# net4 0.0367f
C15827 _250_/a_109_297# _074_ 9.52e-21
C15828 _279_/a_396_47# _279_/a_204_297# 0.0127f
C15829 _279_/a_27_47# _279_/a_314_297# 7.66e-19
C15830 _303_/a_27_47# _303_/a_448_47# 0.0902f
C15831 _303_/a_193_47# _303_/a_1108_47# 0.125f
C15832 net37 _130_ 0.0221f
C15833 mask\[5\] _312_/a_1108_47# 2.34e-20
C15834 _231_/a_161_47# _063_ 0.00133f
C15835 _290_/a_27_413# cal_count\[0\] 7.71e-19
C15836 _229_/a_27_297# _226_/a_27_47# 1.02e-19
C15837 _022_ net26 8.91e-20
C15838 result[1] clknet_2_0__leaf_clk 0.0172f
C15839 _313_/a_448_47# net29 1.76e-20
C15840 _237_/a_505_21# _099_ 0.0337f
C15841 _237_/a_76_199# _092_ 0.0622f
C15842 _200_/a_209_297# clkbuf_0_clk/a_110_47# 6.87e-20
C15843 _051_ _050_ 0.567f
C15844 _277_/a_75_212# _330_/a_1283_21# 1.37e-19
C15845 _323_/a_543_47# _020_ 2.71e-19
C15846 _048_ _089_ 0.164f
C15847 _322_/a_193_47# _205_/a_27_47# 0.0108f
C15848 _314_/a_193_47# net14 0.0067f
C15849 mask\[1\] net14 0.00984f
C15850 _326_/a_193_47# _078_ 0.0225f
C15851 _031_ net34 7.71e-23
C15852 _256_/a_27_297# net46 7.71e-19
C15853 _061_ net33 0.0164f
C15854 _324_/a_193_47# _324_/a_448_47# 0.0642f
C15855 _324_/a_761_289# _324_/a_1108_47# 0.0512f
C15856 _324_/a_27_47# _324_/a_651_413# 9.73e-19
C15857 _327_/a_761_289# clknet_2_3__leaf_clk 3e-20
C15858 net4 _330_/a_1283_21# 4.47e-19
C15859 mask\[2\] net52 0.407f
C15860 net13 _095_ 0.00928f
C15861 _308_/a_805_47# net43 0.00368f
C15862 _308_/a_651_413# net23 9.76e-19
C15863 _328_/a_1217_47# _025_ 2.82e-21
C15864 _255_/a_27_47# _227_/a_109_93# 2.21e-19
C15865 trim_mask\[0\] _267_/a_145_75# 0.0029f
C15866 _040_ _248_/a_109_297# 4.45e-20
C15867 _322_/a_193_47# _040_ 1.3e-20
C15868 _002_ cal_itt\[3\] 1.29e-19
C15869 _319_/a_543_47# net45 6.88e-20
C15870 _319_/a_1108_47# clknet_2_0__leaf_clk 0.061f
C15871 clone7/a_27_47# net41 0.00163f
C15872 _143_/a_68_297# mask\[1\] 0.00832f
C15873 state\[1\] _243_/a_109_297# 9.96e-21
C15874 fanout46/a_27_47# _336_/a_1283_21# 0.0114f
C15875 _309_/a_761_289# net43 0.166f
C15876 _325_/a_27_47# _046_ 7.78e-20
C15877 net15 _282_/a_68_297# 0.00169f
C15878 _037_ _001_ 7.89e-19
C15879 _187_/a_297_47# net16 4.92e-19
C15880 _340_/a_1032_413# net37 9.31e-37
C15881 _327_/a_639_47# net18 6.77e-19
C15882 _053_ _304_/a_761_289# 0.00917f
C15883 _214_/a_199_47# mask\[2\] 0.0105f
C15884 _305_/a_27_47# _002_ 0.284f
C15885 VPWR _103_ 0.255f
C15886 VPWR _313_/a_1217_47# 3.99e-20
C15887 _309_/a_761_289# _309_/a_805_47# 3.69e-19
C15888 _309_/a_193_47# _309_/a_1217_47# 2.36e-20
C15889 _309_/a_543_47# _309_/a_639_47# 0.0138f
C15890 _312_/a_448_47# _084_ 4.93e-20
C15891 trim_val\[3\] clknet_2_2__leaf_clk 0.00266f
C15892 net43 _040_ 8.69e-20
C15893 _178_/a_68_297# trim_mask\[4\] 2.49e-20
C15894 _080_ _016_ 8.64e-21
C15895 _015_ en_co_clk 6.27e-19
C15896 _110_ _327_/a_543_47# 1.92e-20
C15897 _322_/a_761_289# _322_/a_543_47# 0.21f
C15898 _322_/a_193_47# _322_/a_1283_21# 0.0424f
C15899 _322_/a_27_47# _322_/a_1108_47# 0.102f
C15900 _241_/a_297_47# _099_ 0.114f
C15901 _320_/a_761_289# mask\[2\] 1.96e-19
C15902 net1 _013_ 0.00186f
C15903 _069_ _072_ 4.94e-20
C15904 _269_/a_299_297# _112_ 0.00116f
C15905 _253_/a_81_21# _310_/a_193_47# 0.00844f
C15906 _327_/a_193_47# _136_ 0.0014f
C15907 _053_ clkbuf_2_3__f_clk/a_110_47# 0.133f
C15908 VPWR output32/a_27_47# 0.499f
C15909 net35 _047_ 2.85e-19
C15910 _094_ _234_/a_109_297# 0.0129f
C15911 _303_/a_761_289# mask\[4\] 5.88e-19
C15912 net12 _075_ 0.057f
C15913 _078_ net30 0.0868f
C15914 _324_/a_27_47# _008_ 2.16e-20
C15915 clkbuf_2_1__f_clk/a_110_47# _319_/a_651_413# 9.92e-19
C15916 clknet_2_1__leaf_clk _319_/a_193_47# 8.29e-19
C15917 _319_/a_27_47# _319_/a_543_47# 0.106f
C15918 _319_/a_193_47# _319_/a_761_289# 0.174f
C15919 comp _129_ 0.00337f
C15920 _325_/a_651_413# _101_ 2.38e-19
C15921 _325_/a_1108_47# net52 2.36e-21
C15922 _216_/a_199_47# _101_ 1.55e-20
C15923 mask\[3\] _245_/a_373_47# 7.06e-20
C15924 _036_ _339_/a_381_47# 0.148f
C15925 _110_ _335_/a_543_47# 0.00158f
C15926 _117_ _335_/a_193_47# 8.94e-20
C15927 _116_ _335_/a_761_289# 1.75e-20
C15928 _030_ net16 0.00367f
C15929 VPWR clkc 0.367f
C15930 _189_/a_27_47# net42 1.7e-19
C15931 _058_ _136_ 0.153f
C15932 _279_/a_206_47# trim_val\[4\] 0.00235f
C15933 _279_/a_314_297# _118_ 0.0157f
C15934 _303_/a_27_47# _000_ 0.162f
C15935 _185_/a_68_297# net4 5.8e-20
C15936 clkbuf_2_0__f_clk/a_110_47# net55 6.68e-20
C15937 _065_ _202_/a_297_47# 2.28e-19
C15938 _102_ mask\[3\] 1.05e-19
C15939 _023_ net25 1.3e-20
C15940 net13 _164_/a_161_47# 4.35e-19
C15941 _324_/a_27_47# mask\[5\] 2.68e-19
C15942 _282_/a_68_297# _049_ 0.0134f
C15943 _255_/a_27_47# net30 0.0396f
C15944 _010_ net29 8.13e-20
C15945 _015_ _050_ 6.2e-21
C15946 cal_itt\[0\] clk 7.41e-21
C15947 _317_/a_27_47# _316_/a_1108_47# 1.69e-20
C15948 _317_/a_193_47# _316_/a_1283_21# 1.12e-20
C15949 _292_/a_292_297# _128_ 0.00566f
C15950 trimb[4] net40 0.0167f
C15951 _209_/a_27_47# _208_/a_76_199# 5.06e-20
C15952 _028_ _330_/a_761_289# 5.82e-23
C15953 clknet_2_2__leaf_clk _330_/a_543_47# 0.0413f
C15954 net50 _107_ 4.2e-20
C15955 _110_ _332_/a_761_289# 7.59e-20
C15956 net44 _075_ 0.0155f
C15957 _314_/a_1462_47# net14 2.52e-19
C15958 clk _088_ 8.97e-20
C15959 _169_/a_301_53# _051_ 3.97e-19
C15960 output32/a_27_47# _161_/a_68_297# 0.00593f
C15961 VPWR _316_/a_1270_413# 7.19e-19
C15962 _210_/a_199_47# net45 1.19e-19
C15963 _071_ _198_/a_27_47# 1.22e-20
C15964 _007_ _006_ 0.00117f
C15965 _306_/a_1108_47# _003_ 5.47e-21
C15966 _106_ _262_/a_205_47# 6.6e-20
C15967 _136_ _332_/a_27_47# 0.00475f
C15968 net43 net23 0.0439f
C15969 output7/a_27_47# net7 0.173f
C15970 _064_ _336_/a_193_47# 3.71e-20
C15971 _266_/a_68_297# _062_ 3.65e-20
C15972 _197_/a_113_297# _197_/a_199_47# 2.42e-19
C15973 trim_mask\[2\] _267_/a_59_75# 3.93e-21
C15974 _316_/a_805_47# net41 0.00208f
C15975 _097_ calibrate 0.0132f
C15976 _074_ _313_/a_761_289# 2.01e-20
C15977 _232_/a_32_297# _100_ 1.42e-20
C15978 _331_/a_543_47# _052_ 2.78e-21
C15979 net4 _195_/a_218_374# 7.36e-19
C15980 mask\[1\] net52 0.114f
C15981 _330_/a_1108_47# net19 9.02e-20
C15982 _058_ _119_ 4.32e-19
C15983 VPWR _304_/a_761_289# 0.207f
C15984 cal_itt\[0\] net4 0.122f
C15985 _335_/a_193_47# _119_ 1.36e-20
C15986 _328_/a_193_47# _327_/a_193_47# 4e-20
C15987 state\[0\] fanout45/a_27_47# 4.75e-21
C15988 _327_/a_639_47# trim_mask\[0\] 5.51e-21
C15989 _327_/a_448_47# _024_ 0.168f
C15990 _229_/a_27_297# _052_ 3.29e-20
C15991 cal_itt\[2\] net44 4.51e-19
C15992 _097_ net45 0.235f
C15993 _107_ _226_/a_27_47# 0.00327f
C15994 _263_/a_79_21# _075_ 0.00358f
C15995 _305_/a_1217_47# _002_ 0.00102f
C15996 _320_/a_1108_47# _077_ 2.9e-19
C15997 _098_ _170_/a_81_21# 1.2e-21
C15998 _308_/a_543_47# _212_/a_113_297# 4.65e-19
C15999 _328_/a_193_47# _058_ 0.00399f
C16000 _309_/a_27_47# mask\[2\] 7.45e-21
C16001 _322_/a_1283_21# _322_/a_1462_47# 0.0074f
C16002 _322_/a_1108_47# _322_/a_1217_47# 0.00742f
C16003 clk _108_ 2.39e-21
C16004 VPWR _298_/a_215_47# 0.0103f
C16005 mask\[6\] clknet_2_1__leaf_clk 0.125f
C16006 VPWR clkbuf_2_3__f_clk/a_110_47# 1.25f
C16007 net48 _056_ 0.0137f
C16008 trim_val\[2\] net33 0.00704f
C16009 trim_mask\[1\] _066_ 1.32e-21
C16010 _053_ clkbuf_0_clk/a_110_47# 8.73e-19
C16011 _064_ _104_ 0.671f
C16012 mask\[7\] _310_/a_1108_47# 1.79e-19
C16013 _023_ _310_/a_543_47# 7.13e-19
C16014 _102_ _310_/a_1283_21# 4.63e-19
C16015 _202_/a_79_21# _202_/a_382_297# 0.00145f
C16016 _149_/a_150_297# net26 1.05e-19
C16017 _053_ cal_count\[3\] 0.0162f
C16018 _327_/a_1462_47# _136_ 1.06e-19
C16019 cal_itt\[0\] _063_ 0.357f
C16020 _320_/a_761_289# mask\[1\] 0.0192f
C16021 clkbuf_2_0__f_clk/a_110_47# mask\[0\] 0.00815f
C16022 _071_ _041_ 1.8e-20
C16023 _336_/a_27_47# _336_/a_1217_47# 2.56e-19
C16024 _336_/a_761_289# _336_/a_639_47# 3.16e-19
C16025 _218_/a_113_297# mask\[4\] 0.0526f
C16026 _321_/a_27_47# net15 0.0128f
C16027 cal_itt\[0\] _338_/a_381_47# 4.41e-19
C16028 _336_/a_193_47# _264_/a_27_297# 1.49e-21
C16029 _103_ _262_/a_27_47# 2.31e-19
C16030 _281_/a_337_297# _095_ 0.00915f
C16031 _281_/a_103_199# _092_ 0.0974f
C16032 net16 net33 0.11f
C16033 VPWR _043_ 0.484f
C16034 result[4] _102_ 2.99e-20
C16035 net16 trim_mask\[1\] 0.0189f
C16036 _058_ _266_/a_150_297# 4.73e-20
C16037 _249_/a_109_47# mask\[5\] 9.26e-19
C16038 _235_/a_79_21# _337_/a_27_47# 5.73e-21
C16039 _329_/a_761_289# _329_/a_543_47# 0.21f
C16040 _329_/a_193_47# _329_/a_1283_21# 0.0424f
C16041 _329_/a_27_47# _329_/a_1108_47# 0.102f
C16042 net15 _337_/a_27_47# 2.65e-20
C16043 VPWR _321_/a_761_289# 0.218f
C16044 _320_/a_1283_21# fanout44/a_27_47# 2.76e-20
C16045 _004_ net30 0.125f
C16046 net4 _108_ 0.0253f
C16047 _286_/a_439_47# _122_ 0.00369f
C16048 _073_ _203_/a_145_75# 5.76e-19
C16049 _003_ _203_/a_59_75# 4.94e-20
C16050 net54 _089_ 4.07e-20
C16051 VPWR _130_ 0.543f
C16052 _060_ _087_ 0.00815f
C16053 _253_/a_81_21# _224_/a_113_297# 1.29e-21
C16054 VPWR _337_/a_761_289# 0.206f
C16055 _100_ net55 0.253f
C16056 _059_ _337_/a_1108_47# 4.98e-19
C16057 _315_/a_27_47# sample 0.00261f
C16058 _058_ _301_/a_129_47# 7.04e-20
C16059 _324_/a_1217_47# mask\[5\] 1.52e-19
C16060 _187_/a_297_47# net40 7.44e-19
C16061 net50 _257_/a_109_297# 0.00363f
C16062 clknet_2_0__leaf_clk _316_/a_27_47# 0.268f
C16063 _168_/a_27_413# _336_/a_27_47# 4.62e-21
C16064 calibrate _211_/a_109_297# 2.18e-19
C16065 VPWR _276_/a_145_75# 0.00228f
C16066 _239_/a_277_297# _239_/a_474_297# 0.149f
C16067 _015_ _169_/a_301_53# 2.51e-20
C16068 net5 _187_/a_212_413# 6.96e-19
C16069 output15/a_27_47# mask\[6\] 5.65e-21
C16070 _101_ _311_/a_193_47# 4.59e-21
C16071 _293_/a_299_297# _291_/a_35_297# 6.34e-20
C16072 _322_/a_761_289# mask\[2\] 1.89e-19
C16073 _328_/a_448_47# net46 6.55e-19
C16074 VPWR _302_/a_109_297# 0.192f
C16075 _064_ _067_ 0.0254f
C16076 fanout47/a_27_47# cal_count\[0\] 1.46e-20
C16077 _330_/a_1108_47# _279_/a_27_47# 5.98e-21
C16078 _104_ _336_/a_805_47# 4.96e-19
C16079 output14/a_27_47# net14 0.201f
C16080 _329_/a_27_47# net9 0.0128f
C16081 _104_ _264_/a_27_297# 6.77e-21
C16082 _334_/a_1108_47# clknet_2_2__leaf_clk 8.02e-20
C16083 _053_ _038_ 0.0563f
C16084 comp _297_/a_47_47# 1.17e-19
C16085 _026_ _259_/a_27_297# 3.79e-20
C16086 _301_/a_47_47# _332_/a_761_289# 2.67e-19
C16087 _052_ _260_/a_256_47# 0.00371f
C16088 _327_/a_543_47# clknet_2_2__leaf_clk 0.00175f
C16089 _063_ _108_ 6.65e-19
C16090 VPWR _340_/a_1032_413# 0.427f
C16091 _206_/a_27_93# _206_/a_206_47# 0.00698f
C16092 _060_ _263_/a_297_47# 0.00436f
C16093 _053_ _338_/a_476_47# 9.6e-21
C16094 _275_/a_81_21# _275_/a_384_47# 0.00138f
C16095 result[1] _078_ 4.11e-20
C16096 _048_ _092_ 0.273f
C16097 VPWR _253_/a_81_21# 0.226f
C16098 cal_itt\[1\] net19 0.215f
C16099 _275_/a_299_297# _178_/a_68_297# 0.00615f
C16100 _103_ wire42/a_75_212# 0.0649f
C16101 trim[2] _272_/a_81_21# 2e-19
C16102 output33/a_27_47# trim_val\[2\] 0.00947f
C16103 clknet_2_0__leaf_clk sample 0.236f
C16104 _251_/a_373_47# _022_ 1.97e-19
C16105 _323_/a_761_289# _068_ 1.5e-21
C16106 net3 _095_ 0.193f
C16107 _320_/a_193_47# _141_/a_27_47# 0.00913f
C16108 _052_ net19 2.02e-21
C16109 _250_/a_109_47# _078_ 1.96e-19
C16110 _337_/a_27_47# _049_ 0.0504f
C16111 _179_/a_27_47# _176_/a_27_47# 1.77e-20
C16112 _056_ _172_/a_68_297# 3.39e-19
C16113 _335_/a_543_47# clknet_2_2__leaf_clk 1.7e-19
C16114 _328_/a_1462_47# _058_ 1.06e-19
C16115 VPWR clkbuf_0_clk/a_110_47# 1.33f
C16116 VPWR cal_count\[3\] 2.99f
C16117 output33/a_27_47# net16 7.09e-19
C16118 _181_/a_150_297# _279_/a_27_47# 1.25e-19
C16119 _341_/a_651_413# net46 0.0122f
C16120 net50 _118_ 0.00284f
C16121 mask\[0\] _319_/a_448_47# 0.0264f
C16122 _309_/a_27_47# mask\[1\] 5.17e-20
C16123 _333_/a_543_47# net46 0.174f
C16124 net24 clknet_2_1__leaf_clk 0.0488f
C16125 _243_/a_27_297# clone7/a_27_47# 0.0806f
C16126 net42 _168_/a_27_413# 3.84e-21
C16127 clknet_2_0__leaf_clk _003_ 0.00196f
C16128 calibrate _240_/a_109_297# 1.7e-21
C16129 cal_itt\[1\] _107_ 3.8e-19
C16130 _307_/a_1108_47# _137_/a_68_297# 3.43e-19
C16131 _026_ trim_mask\[1\] 1.47e-19
C16132 _336_/a_1108_47# _033_ 1.94e-21
C16133 VPWR _331_/a_27_47# 0.449f
C16134 _286_/a_505_21# clknet_2_3__leaf_clk 0.0797f
C16135 _332_/a_761_289# clknet_2_2__leaf_clk 2.34e-19
C16136 _120_ _092_ 0.0763f
C16137 mask\[6\] _313_/a_27_47# 4.14e-19
C16138 net23 _080_ 0.299f
C16139 output11/a_27_47# net11 0.178f
C16140 net44 _311_/a_639_47# 5.93e-19
C16141 _107_ _052_ 0.0314f
C16142 net27 _312_/a_193_47# 2.95e-19
C16143 _311_/a_27_47# net19 7.96e-22
C16144 _300_/a_47_47# _298_/a_215_47# 1.54e-20
C16145 _329_/a_1283_21# _329_/a_1462_47# 0.0074f
C16146 _329_/a_1108_47# _329_/a_1217_47# 0.00742f
C16147 _094_ _337_/a_1283_21# 6.51e-19
C16148 _273_/a_145_75# _031_ 6.16e-19
C16149 net13 _185_/a_150_297# 3.34e-19
C16150 _287_/a_75_212# cal_count\[0\] 4.82e-19
C16151 net2 net34 0.0237f
C16152 net5 net2 9.9e-19
C16153 _051_ net15 2.07e-20
C16154 _051_ _235_/a_79_21# 1.18e-20
C16155 net26 net14 0.00702f
C16156 _306_/a_1283_21# clk 0.0142f
C16157 _262_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.00344f
C16158 _247_/a_109_47# net52 0.00475f
C16159 _327_/a_27_47# _109_ 2.68e-21
C16160 net50 _025_ 9.84e-20
C16161 net12 _306_/a_543_47# 0.00752f
C16162 clkbuf_2_0__f_clk/a_110_47# _121_ 0.00357f
C16163 _014_ _316_/a_805_47# 3.89e-19
C16164 net45 _316_/a_639_47# 5.93e-19
C16165 _322_/a_1108_47# _077_ 5.29e-19
C16166 _092_ _076_ 4.94e-20
C16167 _325_/a_448_47# net43 0.00323f
C16168 net43 _216_/a_113_297# 3.67e-19
C16169 _058_ _333_/a_639_47# 4.87e-19
C16170 VPWR _038_ 0.377f
C16171 net2 _299_/a_298_297# 3.72e-20
C16172 net35 trim_val\[0\] 0.138f
C16173 _127_ _126_ 0.0402f
C16174 _309_/a_761_289# _082_ 5.07e-21
C16175 _329_/a_1217_47# net9 4.37e-19
C16176 _322_/a_761_289# mask\[1\] 2.24e-20
C16177 _308_/a_193_47# fanout43/a_27_47# 0.00553f
C16178 _164_/a_161_47# net3 0.0238f
C16179 VPWR _338_/a_476_47# 0.267f
C16180 _306_/a_543_47# net44 0.154f
C16181 _062_ _095_ 4.99e-20
C16182 _129_ _132_ 0.319f
C16183 _326_/a_193_47# mask\[7\] 0.0143f
C16184 _326_/a_27_47# _102_ 7.75e-20
C16185 _189_/a_27_47# _098_ 1.09e-19
C16186 trim_val\[3\] trim_mask\[3\] 0.57f
C16187 VPWR _297_/a_377_297# 0.00559f
C16188 _325_/a_193_47# mask\[5\] 3.3e-20
C16189 _341_/a_448_47# _053_ 2.94e-20
C16190 net33 net40 0.994f
C16191 trim_mask\[1\] net40 8.96e-22
C16192 trim_val\[0\] _332_/a_761_289# 0.00308f
C16193 _304_/a_543_47# _065_ 0.00211f
C16194 _337_/a_1217_47# _049_ 1.93e-19
C16195 clk _317_/a_1283_21# 0.00588f
C16196 net43 _314_/a_761_289# 0.176f
C16197 _340_/a_193_47# cal_count\[0\] 4.99e-21
C16198 _156_/a_27_47# _084_ 0.00229f
C16199 _290_/a_27_413# net40 1.87e-20
C16200 trim_val\[1\] net34 0.00267f
C16201 _051_ _049_ 0.0328f
C16202 net49 _055_ 1.29e-20
C16203 _051_ _318_/a_761_289# 4.03e-21
C16204 net13 _141_/a_27_47# 0.00464f
C16205 _189_/a_27_47# clknet_0_clk 0.0512f
C16206 _181_/a_150_297# _118_ 8.55e-19
C16207 clkbuf_2_1__f_clk/a_110_47# clknet_0_clk 0.345f
C16208 _306_/a_448_47# _101_ 8.21e-21
C16209 output25/a_27_47# _310_/a_27_47# 0.0112f
C16210 output16/a_27_47# ctlp[2] 0.158f
C16211 net15 _046_ 0.135f
C16212 trimb[0] net33 0.00141f
C16213 _270_/a_59_75# net16 0.00339f
C16214 _307_/a_1270_413# _039_ 3.69e-19
C16215 VPWR _331_/a_1217_47# 6.18e-20
C16216 _340_/a_1182_261# _132_ 5.78e-20
C16217 clknet_2_3__leaf_clk _150_/a_27_47# 6.4e-22
C16218 _322_/a_448_47# mask\[3\] 0.0168f
C16219 _256_/a_27_297# rebuffer3/a_75_212# 4.76e-21
C16220 net4 _317_/a_1283_21# 0.0129f
C16221 VPWR net21 0.803f
C16222 _303_/a_193_47# _068_ 0.00885f
C16223 VPWR _328_/a_1108_47# 0.294f
C16224 _078_ _313_/a_543_47# 0.0015f
C16225 VPWR trim_mask\[2\] 1.14f
C16226 trimb[1] _125_ 0.00521f
C16227 _300_/a_47_47# cal_count\[3\] 0.0717f
C16228 net2 _133_ 0.00134f
C16229 _012_ _013_ 1.91e-19
C16230 _329_/a_805_47# _026_ 3.24e-19
C16231 output20/a_27_47# _312_/a_27_47# 4.41e-19
C16232 _337_/a_543_47# net45 3.42e-20
C16233 _337_/a_1108_47# clknet_2_0__leaf_clk 7.25e-20
C16234 _108_ _279_/a_396_47# 0.333f
C16235 net28 _314_/a_639_47# 0.00177f
C16236 _309_/a_543_47# _310_/a_1108_47# 2.66e-20
C16237 _035_ _065_ 5.27e-20
C16238 trim_mask\[3\] _330_/a_543_47# 5.37e-21
C16239 _167_/a_161_47# clknet_2_0__leaf_clk 1.92e-20
C16240 _262_/a_27_47# cal_count\[3\] 4.56e-19
C16241 net21 net53 1.58e-20
C16242 cal_itt\[1\] net43 6.61e-21
C16243 VPWR _312_/a_1283_21# 0.392f
C16244 _257_/a_109_297# _335_/a_1108_47# 1.11e-20
C16245 calibrate fanout45/a_27_47# 1.6e-20
C16246 VPWR _323_/a_1108_47# 0.28f
C16247 _119_ _054_ 0.00224f
C16248 VPWR output22/a_27_47# 0.311f
C16249 _119_ net30 6.18e-19
C16250 _313_/a_193_47# _313_/a_639_47# 2.28e-19
C16251 _313_/a_761_289# _313_/a_1270_413# 2.6e-19
C16252 _313_/a_543_47# _313_/a_651_413# 0.0572f
C16253 net52 net26 0.0105f
C16254 state\[2\] net41 2.15e-19
C16255 _336_/a_27_47# clknet_0_clk 0.0028f
C16256 _336_/a_1283_21# clkbuf_2_2__f_clk/a_110_47# 0.0067f
C16257 _294_/a_68_297# comp 1.28e-19
C16258 _289_/a_68_297# _122_ 1.55e-19
C16259 clk _318_/a_651_413# 0.0263f
C16260 VPWR _242_/a_297_47# 0.00429f
C16261 _071_ _190_/a_465_47# 0.00198f
C16262 _337_/a_543_47# _065_ 1.69e-19
C16263 _048_ _226_/a_197_47# 0.00231f
C16264 net21 _009_ 5.24e-21
C16265 fanout45/a_27_47# net45 0.181f
C16266 net3 _226_/a_27_47# 0.155f
C16267 _326_/a_1283_21# net52 0.0128f
C16268 net23 _137_/a_68_297# 2.59e-19
C16269 _060_ _099_ 0.00621f
C16270 net54 _092_ 0.204f
C16271 _321_/a_193_47# clknet_2_1__leaf_clk 0.131f
C16272 VPWR _341_/a_448_47# 0.0776f
C16273 _289_/a_68_297# _299_/a_27_413# 6.12e-19
C16274 _059_ _107_ 9.45e-19
C16275 _306_/a_1108_47# net19 2.19e-21
C16276 VPWR _175_/a_150_297# 0.00208f
C16277 _326_/a_1462_47# mask\[7\] 0.00136f
C16278 VPWR _333_/a_761_289# 0.215f
C16279 VPWR _115_ 0.452f
C16280 mask\[3\] mask\[5\] 7.12e-22
C16281 net31 net36 0.152f
C16282 VPWR _265_/a_299_297# 0.292f
C16283 _124_ _338_/a_193_47# 1.13e-19
C16284 _330_/a_27_47# _330_/a_651_413# 9.73e-19
C16285 _330_/a_761_289# _330_/a_1108_47# 0.0512f
C16286 _330_/a_193_47# _330_/a_448_47# 0.0612f
C16287 _208_/a_218_47# _076_ 0.00129f
C16288 _208_/a_535_374# _077_ 2.83e-20
C16289 calibrate _331_/a_193_47# 1.61e-19
C16290 _028_ _227_/a_209_311# 6.9e-20
C16291 VPWR _308_/a_1283_21# 0.42f
C16292 _074_ _215_/a_109_297# 0.00107f
C16293 net27 _152_/a_68_297# 0.107f
C16294 _096_ _098_ 4.83e-19
C16295 output12/a_27_47# net45 5.09e-20
C16296 _315_/a_805_47# net14 5.85e-19
C16297 _015_ _318_/a_761_289# 6.55e-19
C16298 _040_ _247_/a_27_297# 4.86e-21
C16299 _061_ _136_ 0.00202f
C16300 cal_count\[3\] wire42/a_75_212# 2.12e-20
C16301 _123_ _133_ 0.143f
C16302 net42 _098_ 0.174f
C16303 _079_ net22 0.265f
C16304 _319_/a_651_413# clknet_0_clk 3.18e-19
C16305 _266_/a_150_297# net30 0.00133f
C16306 _242_/a_79_21# _049_ 0.0147f
C16307 mask\[1\] _208_/a_76_199# 3.42e-19
C16308 _187_/a_27_413# _301_/a_47_47# 0.0264f
C16309 net45 _331_/a_193_47# 0.0314f
C16310 VPWR _320_/a_639_47# 8.7e-19
C16311 clkbuf_2_1__f_clk/a_110_47# _245_/a_27_297# 0.0172f
C16312 net50 _062_ 1.8e-19
C16313 trim_mask\[0\] _269_/a_81_21# 3.76e-20
C16314 _256_/a_109_47# trim_mask\[1\] 0.00217f
C16315 clknet_0_clk _096_ 0.0288f
C16316 VPWR _339_/a_1182_261# 0.248f
C16317 net8 ctln[3] 2.28e-19
C16318 _019_ mask\[3\] 0.0341f
C16319 net43 _310_/a_639_47# 0.00168f
C16320 _297_/a_47_47# _132_ 0.372f
C16321 _022_ _010_ 5.28e-19
C16322 clk net2 2.48e-20
C16323 net42 clknet_0_clk 0.104f
C16324 net13 _059_ 0.00434f
C16325 _107_ _170_/a_384_47# 8.79e-20
C16326 _200_/a_209_297# en_co_clk 0.0454f
C16327 _078_ sample 1.76e-19
C16328 _205_/a_27_47# rebuffer6/a_27_47# 2.19e-20
C16329 _198_/a_27_47# _065_ 2.44e-19
C16330 _305_/a_1283_21# clk 0.00454f
C16331 _339_/a_27_47# _286_/a_76_199# 5.71e-21
C16332 net12 _305_/a_543_47# 3.3e-19
C16333 _325_/a_1283_21# _325_/a_1108_47# 0.234f
C16334 _325_/a_761_289# _325_/a_651_413# 0.0977f
C16335 _325_/a_543_47# _325_/a_448_47# 0.0498f
C16336 _325_/a_27_47# _325_/a_639_47# 0.00188f
C16337 _325_/a_193_47# _325_/a_1270_413# 1.46e-19
C16338 _231_/a_161_47# _195_/a_505_21# 0.0015f
C16339 _259_/a_27_297# _280_/a_75_212# 6.15e-20
C16340 _051_ state\[1\] 0.355f
C16341 net9 _298_/a_78_199# 0.00188f
C16342 _042_ clknet_2_3__leaf_clk 1.61e-20
C16343 _189_/a_218_47# clk 0.00292f
C16344 _110_ _336_/a_27_47# 0.0106f
C16345 _074_ _101_ 0.969f
C16346 _064_ clknet_2_3__leaf_clk 0.211f
C16347 VPWR _307_/a_805_47# 2.38e-19
C16348 _090_ _192_/a_639_47# 1.09e-19
C16349 mask\[4\] _311_/a_543_47# 0.0356f
C16350 cal_count\[1\] _288_/a_59_75# 0.17f
C16351 _292_/a_493_297# _125_ 2.04e-21
C16352 _226_/a_27_47# _062_ 0.14f
C16353 net2 net4 0.00902f
C16354 _313_/a_1283_21# _010_ 2.58e-19
C16355 _334_/a_543_47# _057_ 1.22e-19
C16356 _182_/a_27_47# en_co_clk 6.91e-20
C16357 trim[0] _108_ 9.39e-20
C16358 _323_/a_27_47# _150_/a_27_47# 1.06e-20
C16359 VPWR _241_/a_105_352# 0.155f
C16360 _321_/a_1270_413# _042_ 2.02e-19
C16361 _041_ net45 1.44e-20
C16362 _104_ _256_/a_373_47# 0.00411f
C16363 _305_/a_543_47# net44 0.00943f
C16364 cal_itt\[2\] _001_ 2.07e-20
C16365 _294_/a_150_297# VPWR 0.00127f
C16366 _268_/a_75_212# clknet_2_2__leaf_clk 0.0215f
C16367 _316_/a_193_47# _316_/a_543_47# 0.23f
C16368 _316_/a_27_47# _316_/a_1283_21# 0.0436f
C16369 _189_/a_27_47# net44 3.35e-21
C16370 _340_/a_956_413# _123_ 0.00237f
C16371 VPWR _303_/a_1283_21# 0.453f
C16372 clkbuf_2_1__f_clk/a_110_47# net44 0.00139f
C16373 trim_mask\[3\] _335_/a_543_47# 4.03e-20
C16374 net50 _335_/a_761_289# 0.00471f
C16375 _168_/a_27_413# clknet_0_clk 0.00165f
C16376 trim_val\[3\] _335_/a_1283_21# 0.0618f
C16377 _214_/a_113_297# clknet_2_0__leaf_clk 1.88e-20
C16378 en_co_clk net37 1.95e-19
C16379 _340_/a_193_47# net16 1.08e-20
C16380 _330_/a_27_47# net46 0.296f
C16381 _330_/a_193_47# _027_ 0.74f
C16382 _008_ _311_/a_448_47# 0.158f
C16383 _008_ net27 9.66e-23
C16384 _041_ _065_ 0.204f
C16385 _301_/a_285_47# _300_/a_285_47# 0.00178f
C16386 _307_/a_193_47# _315_/a_193_47# 2.34e-19
C16387 calibrate _260_/a_93_21# 0.0711f
C16388 _309_/a_27_47# net26 4.53e-21
C16389 net2 _063_ 1.05e-19
C16390 net43 _059_ 1.7e-19
C16391 state\[2\] _318_/a_639_47# 2.38e-19
C16392 _305_/a_1283_21# _063_ 3.38e-19
C16393 _037_ net2 1.05e-19
C16394 _307_/a_448_47# net30 4.57e-19
C16395 _320_/a_193_47# clknet_2_0__leaf_clk 0.00308f
C16396 VPWR _309_/a_651_413# 0.134f
C16397 _061_ _301_/a_129_47# 2.39e-19
C16398 net45 _331_/a_1462_47# 0.00288f
C16399 net45 _260_/a_93_21# 2.59e-20
C16400 VPWR _190_/a_215_47# 0.00277f
C16401 _232_/a_32_297# net4 2.27e-21
C16402 net27 mask\[5\] 0.816f
C16403 mask\[7\] _251_/a_27_297# 0.0953f
C16404 _074_ _312_/a_448_47# 2.76e-20
C16405 net13 _317_/a_1108_47# 2.3e-20
C16406 _200_/a_209_297# _200_/a_303_47# 1.26e-19
C16407 _097_ _013_ 0.00171f
C16408 VPWR _339_/a_1296_47# 1.86e-19
C16409 net9 _340_/a_652_21# 0.00712f
C16410 _042_ net20 1.83e-22
C16411 _077_ rebuffer4/a_27_47# 2.14e-20
C16412 _033_ net18 1.37e-20
C16413 _217_/a_109_297# _082_ 3.1e-19
C16414 _307_/a_193_47# _074_ 0.0168f
C16415 net4 _336_/a_193_47# 0.0115f
C16416 _314_/a_27_47# _314_/a_193_47# 0.883f
C16417 VPWR _045_ 0.513f
C16418 _329_/a_27_47# _258_/a_27_297# 0.0111f
C16419 _329_/a_27_47# _024_ 1.74e-20
C16420 _237_/a_505_21# _192_/a_505_280# 9.76e-19
C16421 VPWR _249_/a_109_297# 0.178f
C16422 _326_/a_193_47# net28 4.64e-20
C16423 VPWR _293_/a_81_21# 0.211f
C16424 _228_/a_79_21# _228_/a_297_47# 0.0326f
C16425 net43 _306_/a_1108_47# 1.11e-19
C16426 _187_/a_27_413# trim_val\[0\] 9.02e-21
C16427 _339_/a_27_47# cal_count\[0\] 0.491f
C16428 output8/a_27_47# ctln[2] 0.16f
C16429 _015_ state\[1\] 0.0493f
C16430 _169_/a_215_311# _050_ 3.11e-19
C16431 _216_/a_113_297# _082_ 0.1f
C16432 _335_/a_543_47# _330_/a_1283_21# 4.14e-19
C16433 _110_ net48 0.00265f
C16434 _051_ _336_/a_651_413# 7.37e-21
C16435 _307_/a_761_289# clknet_2_0__leaf_clk 2.62e-19
C16436 _307_/a_27_47# net45 0.298f
C16437 _045_ net53 1.02e-19
C16438 _104_ clk 0.00692f
C16439 _004_ sample 0.0175f
C16440 trim[3] _334_/a_193_47# 1.78e-19
C16441 VPWR _324_/a_805_47# 4.08e-19
C16442 net31 trim[4] 0.109f
C16443 _110_ _336_/a_1217_47# 1.59e-19
C16444 _249_/a_109_297# net53 0.0573f
C16445 ctlp[0] result[6] 4.71e-19
C16446 _060_ _226_/a_109_47# 8.38e-19
C16447 _136_ _066_ 0.0391f
C16448 _019_ net27 4.53e-21
C16449 state\[0\] _048_ 0.0117f
C16450 _235_/a_382_297# _092_ 0.00169f
C16451 _277_/a_75_212# _104_ 3.86e-19
C16452 clk net55 0.00591f
C16453 _320_/a_543_47# clkbuf_2_1__f_clk/a_110_47# 4.44e-19
C16454 net8 net34 0.0332f
C16455 _321_/a_1108_47# _078_ 1.62e-20
C16456 _045_ _009_ 0.00719f
C16457 _064_ _328_/a_27_47# 3.82e-21
C16458 VPWR mask\[4\] 0.488f
C16459 VPWR _322_/a_639_47# 4.88e-19
C16460 _304_/a_651_413# _284_/a_68_297# 3e-20
C16461 _259_/a_373_47# trim_mask\[2\] 2.72e-20
C16462 _336_/a_193_47# _063_ 1.36e-19
C16463 _291_/a_35_297# _125_ 0.023f
C16464 _136_ net16 0.0255f
C16465 net12 net42 2.81e-20
C16466 _104_ net4 0.166f
C16467 _308_/a_448_47# _074_ 0.00411f
C16468 _269_/a_81_21# _333_/a_193_47# 0.00164f
C16469 _127_ net47 1.52e-20
C16470 _123_ _063_ 0.0556f
C16471 _030_ _333_/a_1108_47# 1.61e-19
C16472 _113_ _333_/a_448_47# 1.68e-20
C16473 ctln[7] _318_/a_448_47# 5.95e-20
C16474 net13 _318_/a_1270_413# 5.91e-20
C16475 _316_/a_448_47# _316_/a_639_47# 4.61e-19
C16476 _198_/a_181_47# _069_ 2.15e-19
C16477 mask\[4\] net53 0.646f
C16478 _037_ _123_ 0.0116f
C16479 VPWR _220_/a_199_47# 9e-19
C16480 cal_itt\[1\] _062_ 0.363f
C16481 _323_/a_27_47# _042_ 0.05f
C16482 net4 net55 1.05e-20
C16483 clknet_2_1__leaf_clk _312_/a_543_47# 2.56e-19
C16484 net44 _319_/a_651_413# 2.61e-20
C16485 _247_/a_109_297# mask\[2\] 0.00166f
C16486 _308_/a_1108_47# net45 0.012f
C16487 mask\[0\] net14 0.00272f
C16488 _326_/a_1108_47# net43 0.237f
C16489 _330_/a_1217_47# net46 6.54e-19
C16490 _052_ _062_ 2.54e-20
C16491 _007_ _310_/a_27_47# 0.169f
C16492 _053_ en_co_clk 0.014f
C16493 trim[1] net34 0.0403f
C16494 _122_ _298_/a_78_199# 0.0898f
C16495 _323_/a_1283_21# clknet_2_1__leaf_clk 1.09e-20
C16496 net51 rebuffer5/a_161_47# 0.293f
C16497 _341_/a_651_413# _065_ 9.16e-19
C16498 state\[2\] _243_/a_27_297# 5.29e-21
C16499 _237_/a_76_199# net45 3.57e-21
C16500 _237_/a_505_21# _014_ 2.65e-20
C16501 _251_/a_373_47# net52 0.00135f
C16502 VPWR _275_/a_384_47# 1.33e-19
C16503 net43 _203_/a_59_75# 1.14e-20
C16504 _334_/a_761_289# net46 0.168f
C16505 net15 _246_/a_109_47# 5.78e-20
C16506 net25 _310_/a_193_47# 0.0081f
C16507 VPWR _178_/a_150_297# 0.00204f
C16508 _195_/a_76_199# _195_/a_535_374# 6.64e-19
C16509 _290_/a_207_413# output37/a_27_47# 0.00114f
C16510 _294_/a_68_297# _132_ 0.0139f
C16511 _104_ _063_ 4.99e-20
C16512 _327_/a_27_47# net46 0.3f
C16513 net9 _338_/a_27_47# 2.21e-19
C16514 _299_/a_27_413# _298_/a_78_199# 4.16e-20
C16515 cal_itt\[0\] _195_/a_505_21# 0.265f
C16516 cal_itt\[1\] _195_/a_76_199# 0.0366f
C16517 _200_/a_80_21# _068_ 4.85e-19
C16518 _336_/a_27_47# clknet_2_2__leaf_clk 0.252f
C16519 _328_/a_1270_413# trim_mask\[1\] 4.1e-19
C16520 _189_/a_408_47# _107_ 0.00102f
C16521 net13 clknet_2_0__leaf_clk 0.164f
C16522 trim_mask\[2\] _272_/a_384_47# 0.0101f
C16523 cal_itt\[2\] cal_itt\[0\] 0.136f
C16524 net9 _340_/a_1056_47# 3.98e-19
C16525 result[1] _308_/a_27_47# 0.0203f
C16526 _319_/a_448_47# _016_ 0.157f
C16527 _324_/a_193_47# _074_ 8.1e-21
C16528 _304_/a_27_47# _304_/a_543_47# 0.113f
C16529 _304_/a_193_47# _304_/a_761_289# 0.186f
C16530 net4 _067_ 0.0556f
C16531 trim_mask\[2\] _336_/a_1108_47# 1.12e-19
C16532 _289_/a_68_297# _297_/a_285_47# 2.98e-19
C16533 net4 _070_ 0.138f
C16534 trim_mask\[0\] _033_ 0.00407f
C16535 _024_ _106_ 7.33e-22
C16536 _099_ net30 7.54e-20
C16537 _329_/a_761_289# trim_mask\[2\] 2.59e-19
C16538 _168_/a_207_413# clk 0.0154f
C16539 _334_/a_761_289# _334_/a_639_47# 3.16e-19
C16540 _334_/a_27_47# _334_/a_1217_47# 2.56e-19
C16541 _314_/a_543_47# _314_/a_639_47# 0.0138f
C16542 _314_/a_193_47# _314_/a_1217_47# 2.36e-20
C16543 _314_/a_761_289# _314_/a_805_47# 3.69e-19
C16544 _034_ _192_/a_174_21# 6.52e-19
C16545 _063_ net55 5.98e-19
C16546 VPWR _020_ 0.452f
C16547 _263_/a_79_21# _096_ 5.63e-20
C16548 _327_/a_193_47# _327_/a_448_47# 0.0604f
C16549 _327_/a_761_289# _327_/a_1108_47# 0.0512f
C16550 _327_/a_27_47# _327_/a_651_413# 9.73e-19
C16551 _336_/a_761_289# net19 6.83e-19
C16552 _053_ _050_ 0.183f
C16553 _335_/a_193_47# _027_ 9.9e-20
C16554 _335_/a_27_47# net46 0.345f
C16555 _322_/a_27_47# _074_ 0.00841f
C16556 _074_ _248_/a_27_297# 0.00126f
C16557 calibrate _241_/a_388_297# 9.09e-20
C16558 _307_/a_1217_47# net45 6.92e-19
C16559 _308_/a_1283_21# _319_/a_193_47# 1.03e-19
C16560 _308_/a_1108_47# _319_/a_27_47# 1.09e-19
C16561 _169_/a_215_311# _169_/a_301_53# 0.0049f
C16562 _020_ net53 0.156f
C16563 _262_/a_109_297# _190_/a_27_47# 8.03e-21
C16564 _266_/a_68_297# _264_/a_27_297# 7.02e-20
C16565 _036_ _286_/a_505_21# 0.00106f
C16566 output27/a_27_47# _007_ 8.94e-20
C16567 mask\[6\] net21 0.00186f
C16568 _168_/a_207_413# net4 8.59e-22
C16569 VPWR _291_/a_285_47# 8.6e-19
C16570 _059_ net3 0.0264f
C16571 _327_/a_448_47# _058_ 0.00438f
C16572 net45 _241_/a_388_297# 0.00113f
C16573 _014_ _241_/a_297_47# 0.0476f
C16574 _104_ _260_/a_346_47# 5.22e-19
C16575 net46 rebuffer1/a_75_212# 3.52e-20
C16576 _067_ _063_ 0.54f
C16577 _328_/a_761_289# net9 0.00368f
C16578 _063_ _070_ 0.0225f
C16579 net9 net17 0.111f
C16580 net47 _284_/a_68_297# 0.00446f
C16581 _304_/a_805_47# _122_ 6.43e-19
C16582 _020_ _009_ 1.89e-20
C16583 _333_/a_1108_47# net33 0.00671f
C16584 _336_/a_761_289# _107_ 0.00133f
C16585 _005_ _074_ 0.124f
C16586 VPWR _222_/a_199_47# 3.71e-19
C16587 _112_ _333_/a_543_47# 0.00315f
C16588 net49 _333_/a_1283_21# 1.09e-19
C16589 trim_mask\[1\] _333_/a_1108_47# 4.23e-19
C16590 trim_val\[1\] _333_/a_448_47# 9.97e-20
C16591 _021_ _312_/a_193_47# 1.23e-20
C16592 _340_/a_652_21# _122_ 0.00191f
C16593 _304_/a_761_289# net18 0.01f
C16594 _274_/a_75_212# net48 1.93e-19
C16595 clknet_0_clk _098_ 4.99e-20
C16596 _246_/a_27_297# net30 7.56e-21
C16597 _092_ cal_itt\[3\] 4.32e-20
C16598 _301_/a_129_47# net16 0.00162f
C16599 _298_/a_493_297# _298_/a_215_47# 3.25e-19
C16600 _310_/a_193_47# _310_/a_543_47# 0.217f
C16601 _310_/a_27_47# _310_/a_1283_21# 0.0436f
C16602 _107_ clone1/a_27_47# 0.00977f
C16603 _144_/a_27_47# net34 3.57e-21
C16604 VPWR _325_/a_27_47# 0.43f
C16605 _327_/a_543_47# _108_ 5.7e-19
C16606 VPWR en_co_clk 6.66f
C16607 _309_/a_639_47# _074_ 2.64e-19
C16608 trim_mask\[0\] _103_ 0.232f
C16609 _046_ _313_/a_193_47# 9.45e-19
C16610 net43 clknet_2_0__leaf_clk 0.373f
C16611 _335_/a_27_47# _335_/a_651_413# 9.73e-19
C16612 _335_/a_761_289# _335_/a_1108_47# 0.0512f
C16613 _335_/a_193_47# _335_/a_448_47# 0.0642f
C16614 _018_ mask\[2\] 4.03e-19
C16615 net5 clknet_2_3__leaf_clk 7.24e-20
C16616 net26 _208_/a_76_199# 1.14e-21
C16617 result[4] _310_/a_27_47# 0.0131f
C16618 _026_ _119_ 2.56e-20
C16619 mask\[1\] _247_/a_109_297# 1.12e-20
C16620 net35 _108_ 0.00122f
C16621 _058_ _332_/a_1108_47# 0.00185f
C16622 mask\[0\] net52 6.74e-19
C16623 _304_/a_761_289# _302_/a_27_297# 4.37e-21
C16624 net9 _301_/a_285_47# 9.99e-20
C16625 net13 _232_/a_114_297# 0.00141f
C16626 net48 clknet_2_2__leaf_clk 2.26e-20
C16627 _069_ net19 2.78e-20
C16628 output32/a_27_47# trim_mask\[0\] 7.18e-21
C16629 _327_/a_1217_47# net46 8.19e-19
C16630 net9 _341_/a_543_47# 1.97e-19
C16631 _336_/a_448_47# trim_mask\[4\] 0.025f
C16632 _071_ _068_ 0.319f
C16633 output23/a_27_47# _005_ 0.0668f
C16634 clkbuf_2_0__f_clk/a_110_47# _095_ 0.117f
C16635 _339_/a_562_413# _123_ 0.00224f
C16636 net43 _305_/a_1108_47# 0.258f
C16637 _026_ _328_/a_193_47# 1.18e-19
C16638 _043_ net18 0.0211f
C16639 clk _316_/a_543_47# 4.67e-19
C16640 _336_/a_193_47# _279_/a_396_47# 0.0116f
C16641 _336_/a_27_47# _279_/a_204_297# 1.34e-19
C16642 _214_/a_113_297# _078_ 0.129f
C16643 net16 _339_/a_27_47# 6.15e-20
C16644 VPWR _212_/a_199_47# 3.44e-19
C16645 VPWR _050_ 1.82f
C16646 net43 _146_/a_68_297# 0.0294f
C16647 _332_/a_761_289# _108_ 0.0315f
C16648 _321_/a_27_47# _321_/a_543_47# 0.106f
C16649 _321_/a_193_47# _321_/a_761_289# 0.176f
C16650 _332_/a_27_47# _332_/a_1108_47# 0.102f
C16651 _332_/a_193_47# _332_/a_1283_21# 0.0418f
C16652 _332_/a_761_289# _332_/a_543_47# 0.21f
C16653 _136_ net40 0.0317f
C16654 net39 net33 1.61e-20
C16655 _302_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 2.93e-20
C16656 output14/a_27_47# _314_/a_27_47# 0.0023f
C16657 _335_/a_1217_47# net46 0.0013f
C16658 _168_/a_27_413# clknet_2_2__leaf_clk 6.96e-20
C16659 _059_ _062_ 0.102f
C16660 state\[0\] net54 0.126f
C16661 _169_/a_373_53# state\[0\] 0.00443f
C16662 net3 _317_/a_1108_47# 1.46e-20
C16663 output31/a_27_47# _176_/a_27_47# 8.27e-21
C16664 clkbuf_0_clk/a_110_47# _304_/a_193_47# 1.02e-19
C16665 _059_ fanout44/a_27_47# 1.22e-21
C16666 _129_ _130_ 0.292f
C16667 _320_/a_193_47# _078_ 3.94e-19
C16668 _337_/a_27_47# _337_/a_543_47# 0.111f
C16669 _337_/a_193_47# _337_/a_761_289# 0.186f
C16670 _304_/a_448_47# clknet_2_3__leaf_clk 0.0162f
C16671 _333_/a_193_47# net32 1.66e-19
C16672 result[4] output27/a_27_47# 1.02e-19
C16673 output26/a_27_47# result[5] 0.00311f
C16674 _340_/a_27_47# _133_ 2.33e-22
C16675 _288_/a_59_75# _288_/a_145_75# 0.00658f
C16676 net9 _339_/a_193_47# 0.0164f
C16677 _309_/a_448_47# clknet_2_1__leaf_clk 2.63e-20
C16678 _257_/a_109_297# trim_mask\[1\] 0.0163f
C16679 _302_/a_109_297# net18 0.0044f
C16680 VPWR _330_/a_805_47# 2.28e-19
C16681 _089_ clone7/a_27_47# 8.68e-20
C16682 _332_/a_805_47# net46 0.00316f
C16683 net28 _251_/a_27_297# 0.00115f
C16684 _338_/a_27_47# _122_ 0.00155f
C16685 _048_ _192_/a_476_47# 0.00275f
C16686 _341_/a_27_47# _284_/a_68_297# 3.15e-19
C16687 _276_/a_59_75# _276_/a_145_75# 0.00658f
C16688 net48 _333_/a_651_413# 6.72e-21
C16689 _104_ _279_/a_396_47# 0.0821f
C16690 net3 _192_/a_27_47# 0.0394f
C16691 VPWR _200_/a_303_47# 1.45e-19
C16692 clknet_2_1__leaf_clk _249_/a_27_297# 0.058f
C16693 net37 output40/a_27_47# 0.00597f
C16694 _306_/a_193_47# rebuffer4/a_27_47# 3.29e-21
C16695 VPWR _334_/a_193_47# 0.601f
C16696 _051_ clkbuf_2_2__f_clk/a_110_47# 6.84e-19
C16697 net45 _281_/a_103_199# 4.61e-20
C16698 _310_/a_448_47# _310_/a_639_47# 4.61e-19
C16699 VPWR _228_/a_297_47# 0.00397f
C16700 _324_/a_1108_47# _042_ 1.03e-19
C16701 clknet_2_3__leaf_clk _133_ 0.00197f
C16702 _314_/a_761_289# net29 0.00218f
C16703 _110_ clknet_0_clk 1.84e-21
C16704 _307_/a_761_289# _078_ 0.00235f
C16705 _307_/a_543_47# mask\[0\] 2.09e-20
C16706 _307_/a_1283_21# net22 0.136f
C16707 VPWR _325_/a_1217_47# 1.19e-19
C16708 VPWR net25 0.637f
C16709 net21 _313_/a_805_47# 7.65e-20
C16710 _335_/a_193_47# _032_ 0.224f
C16711 _324_/a_639_47# clknet_2_1__leaf_clk 3.14e-19
C16712 net16 _333_/a_639_47# 0.0015f
C16713 _302_/a_27_297# _302_/a_109_297# 0.171f
C16714 _340_/a_1032_413# _129_ 4.17e-19
C16715 _232_/a_32_297# _034_ 1.16e-19
C16716 input1/a_75_212# output41/a_27_47# 0.00329f
C16717 result[4] _310_/a_1217_47# 6.14e-21
C16718 _226_/a_303_47# _049_ 1.13e-19
C16719 _311_/a_193_47# _311_/a_651_413# 0.0276f
C16720 _311_/a_543_47# _311_/a_1108_47# 7.99e-20
C16721 _168_/a_297_47# _107_ 2.5e-19
C16722 output27/a_27_47# net27 0.18f
C16723 clkbuf_2_0__f_clk/a_110_47# _164_/a_161_47# 5.09e-19
C16724 cal_count\[3\] net18 0.423f
C16725 trim_mask\[0\] clkbuf_2_3__f_clk/a_110_47# 0.127f
C16726 output10/a_27_47# _335_/a_27_47# 3.61e-19
C16727 en_co_clk _192_/a_548_47# 9.46e-20
C16728 _304_/a_193_47# _038_ 7.11e-21
C16729 _304_/a_1108_47# _136_ 5.64e-19
C16730 _104_ _257_/a_109_47# 5.15e-20
C16731 result[1] result[3] 0.00269f
C16732 net47 clknet_0_clk 5.33e-19
C16733 _071_ _306_/a_27_47# 1.97e-21
C16734 _300_/a_47_47# en_co_clk 1.4e-19
C16735 trim[4] _332_/a_27_47# 6.64e-20
C16736 output36/a_27_47# output37/a_27_47# 0.00254f
C16737 _033_ trim_mask\[4\] 0.0193f
C16738 ctlp[7] clknet_2_1__leaf_clk 1.53e-19
C16739 _307_/a_193_47# output30/a_27_47# 6.7e-19
C16740 _074_ _156_/a_27_47# 2.4e-19
C16741 net15 _314_/a_1108_47# 1.64e-20
C16742 _304_/a_651_413# net47 0.0122f
C16743 net12 _098_ 0.0253f
C16744 _326_/a_543_47# _314_/a_193_47# 1.97e-20
C16745 _326_/a_193_47# _314_/a_543_47# 2.28e-19
C16746 _326_/a_761_289# _314_/a_761_289# 0.00117f
C16747 trim_mask\[1\] _118_ 4.41e-20
C16748 _048_ calibrate 0.262f
C16749 _336_/a_761_289# _118_ 3.01e-19
C16750 _336_/a_543_47# trim_val\[4\] 1.05e-19
C16751 VPWR _314_/a_651_413# 0.143f
C16752 _230_/a_145_75# net4 7.2e-19
C16753 clknet_2_1__leaf_clk _220_/a_113_297# 0.00345f
C16754 _308_/a_651_413# _078_ 8.7e-19
C16755 _340_/a_652_21# _340_/a_381_47# 7.79e-20
C16756 _340_/a_193_47# _340_/a_562_413# 4.45e-20
C16757 _340_/a_1182_261# _340_/a_1032_413# 0.344f
C16758 _340_/a_27_47# _340_/a_956_413# 0.00159f
C16759 _332_/a_1108_47# _332_/a_1217_47# 0.00742f
C16760 _332_/a_1283_21# _332_/a_1462_47# 0.0074f
C16761 _121_ net52 2.08e-20
C16762 _228_/a_79_21# _049_ 0.025f
C16763 _088_ _170_/a_81_21# 0.0285f
C16764 net2 _208_/a_76_199# 0.188f
C16765 _255_/a_27_47# _107_ 0.00512f
C16766 _302_/a_27_297# cal_count\[3\] 0.0968f
C16767 net8 _273_/a_145_75# 1.62e-20
C16768 VPWR _169_/a_301_53# 1.46e-20
C16769 _128_ _290_/a_207_413# 3.1e-21
C16770 net12 clknet_0_clk 0.0103f
C16771 _048_ net45 4.74e-19
C16772 net43 _319_/a_639_47# 4.36e-19
C16773 net3 clknet_2_0__leaf_clk 0.0115f
C16774 _323_/a_193_47# _149_/a_68_297# 1.55e-20
C16775 _292_/a_292_297# net16 1.54e-20
C16776 _067_ _201_/a_113_47# 2.18e-20
C16777 _326_/a_27_47# _310_/a_27_47# 9.43e-22
C16778 _070_ _201_/a_113_47# 3.03e-20
C16779 _060_ net41 0.161f
C16780 _191_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 0.00122f
C16781 _309_/a_27_47# output24/a_27_47# 8.25e-19
C16782 net5 _301_/a_377_297# 5.38e-20
C16783 trim[0] trim_val\[1\] 0.00247f
C16784 net31 net49 0.00371f
C16785 net45 _330_/a_27_47# 7.48e-21
C16786 _062_ _203_/a_59_75# 6.02e-20
C16787 _333_/a_1462_47# net32 2.91e-19
C16788 VPWR _310_/a_543_47# 0.197f
C16789 _052_ _227_/a_209_311# 2.19e-20
C16790 _088_ _227_/a_296_53# 1.25e-20
C16791 mask\[6\] _045_ 0.0215f
C16792 net9 _339_/a_796_47# 2.99e-19
C16793 net10 net46 3.81e-20
C16794 _025_ trim_mask\[1\] 0.12f
C16795 net13 _078_ 0.0381f
C16796 _250_/a_109_297# mask\[5\] 0.0136f
C16797 net31 _290_/a_207_413# 7.34e-19
C16798 mask\[6\] _249_/a_109_297# 1.44e-19
C16799 _038_ net18 0.0268f
C16800 _093_ en_co_clk 0.00338f
C16801 _078_ _155_/a_68_297# 0.00101f
C16802 fanout47/a_27_47# net19 0.00323f
C16803 _110_ _047_ 2.45e-20
C16804 net43 _069_ 7.84e-21
C16805 clkbuf_2_1__f_clk/a_110_47# mask\[2\] 0.014f
C16806 _035_ _338_/a_193_47# 0.173f
C16807 _048_ _065_ 0.0175f
C16808 _247_/a_27_297# _247_/a_373_47# 0.0134f
C16809 _230_/a_145_75# _063_ 6.66e-19
C16810 net44 clknet_0_clk 0.00545f
C16811 output32/a_27_47# _265_/a_81_21# 2.75e-20
C16812 _338_/a_476_47# net18 0.00994f
C16813 _128_ _289_/a_68_297# 2.16e-20
C16814 net45 _120_ 4.53e-21
C16815 VPWR net1 0.177f
C16816 VPWR _327_/a_805_47# 2.51e-19
C16817 _048_ _105_ 0.237f
C16818 _263_/a_79_21# _098_ 4.91e-19
C16819 _051_ fanout45/a_27_47# 3.53e-19
C16820 _169_/a_215_311# _049_ 6.23e-21
C16821 _302_/a_27_297# _038_ 0.111f
C16822 _169_/a_215_311# _318_/a_761_289# 0.00109f
C16823 net1 valid 0.0364f
C16824 _130_ _297_/a_47_47# 5.4e-20
C16825 _129_ _297_/a_377_297# 0.00335f
C16826 _307_/a_761_289# _004_ 0.00175f
C16827 mask\[6\] mask\[4\] 5.62e-20
C16828 net28 _313_/a_543_47# 0.0358f
C16829 VPWR _039_ 0.68f
C16830 _322_/a_193_47# _078_ 0.0036f
C16831 trim_mask\[0\] cal_count\[3\] 2.78e-19
C16832 net45 _076_ 1.28e-20
C16833 _050_ _093_ 2.32e-20
C16834 ctln[4] _335_/a_1108_47# 2.83e-19
C16835 _120_ _065_ 0.123f
C16836 clknet_0_clk _263_/a_79_21# 4.48e-22
C16837 net4 clknet_2_3__leaf_clk 0.0256f
C16838 VPWR _335_/a_805_47# 3.65e-19
C16839 _326_/a_27_47# output27/a_27_47# 3.72e-19
C16840 _339_/a_193_47# _122_ 6.01e-21
C16841 VPWR _311_/a_1108_47# 0.285f
C16842 clknet_2_1__leaf_clk _222_/a_113_297# 0.0129f
C16843 _083_ _042_ 8.1e-20
C16844 trim_mask\[2\] net18 0.00588f
C16845 _060_ _094_ 1.56e-20
C16846 _340_/a_1140_413# net47 9.26e-20
C16847 _037_ _304_/a_1270_413# 8.96e-21
C16848 _106_ trim_val\[4\] 0.0101f
C16849 _065_ _076_ 0.669f
C16850 net43 _078_ 2.58f
C16851 _311_/a_1108_47# net53 0.00102f
C16852 VPWR _332_/a_639_47# 0.00379f
C16853 _050_ wire42/a_75_212# 3.15e-19
C16854 _340_/a_27_47# _037_ 0.151f
C16855 _340_/a_1032_413# _340_/a_1296_47# 0.00384f
C16856 clknet_2_1__leaf_clk rebuffer5/a_161_47# 0.011f
C16857 _319_/a_27_47# _120_ 1.8e-20
C16858 _340_/a_1032_413# _297_/a_47_47# 6.74e-20
C16859 _051_ _331_/a_193_47# 0.00143f
C16860 cal_count\[1\] _127_ 1.22e-19
C16861 _277_/a_75_212# _116_ 0.0372f
C16862 _327_/a_1283_21# _268_/a_75_212# 0.01f
C16863 _327_/a_27_47# _111_ 1.77e-19
C16864 fanout44/a_27_47# clknet_2_0__leaf_clk 0.0446f
C16865 en_co_clk _243_/a_109_47# 4.69e-20
C16866 _253_/a_299_297# _023_ 9.1e-19
C16867 mask\[0\] _034_ 8.14e-22
C16868 _134_ _298_/a_78_199# 2.16e-19
C16869 _081_ net14 0.0112f
C16870 _309_/a_805_47# _078_ 0.00136f
C16871 _187_/a_212_413# net35 0.025f
C16872 _323_/a_1283_21# _043_ 0.0167f
C16873 _104_ trim_val\[3\] 5.05e-20
C16874 _064_ net50 0.465f
C16875 cal_count\[3\] _191_/a_27_297# 0.0689f
C16876 _323_/a_1108_47# net18 2.68e-19
C16877 _320_/a_543_47# clknet_0_clk 0.00449f
C16878 _063_ clknet_2_3__leaf_clk 0.0185f
C16879 _337_/a_651_413# net44 0.0129f
C16880 rebuffer4/a_27_47# _072_ 8.44e-21
C16881 _309_/a_651_413# net24 0.0265f
C16882 clknet_0_clk clknet_2_2__leaf_clk 0.0836f
C16883 _338_/a_381_47# clknet_2_3__leaf_clk 0.0159f
C16884 output17/a_27_47# ctlp[3] 0.157f
C16885 _233_/a_27_297# cal 0.00651f
C16886 _271_/a_75_212# net46 0.0424f
C16887 _037_ clknet_2_3__leaf_clk 0.0387f
C16888 trim_mask\[0\] _038_ 3.83e-20
C16889 _239_/a_27_297# _048_ 2.69e-19
C16890 _021_ mask\[5\] 9.18e-20
C16891 net43 _313_/a_651_413# 0.0154f
C16892 _234_/a_109_297# _092_ 3.9e-19
C16893 VPWR ctlp[5] 0.353f
C16894 _280_/a_75_212# _119_ 0.207f
C16895 _338_/a_1224_47# net18 1.57e-19
C16896 cal_count\[1\] _126_ 0.095f
C16897 mask\[1\] clkbuf_2_1__f_clk/a_110_47# 0.0121f
C16898 _327_/a_27_47# rebuffer3/a_75_212# 3.91e-19
C16899 VPWR output40/a_27_47# 0.499f
C16900 mask\[3\] net45 4.53e-21
C16901 _050_ _319_/a_193_47# 5.42e-21
C16902 output34/a_27_47# net33 0.00131f
C16903 _149_/a_68_297# _303_/a_27_47# 5.08e-21
C16904 _189_/a_408_47# _062_ 0.0985f
C16905 _189_/a_218_47# _075_ 4.95e-20
C16906 _071_ cal_itt\[3\] 1.65e-19
C16907 _268_/a_75_212# _108_ 0.0365f
C16908 net47 net44 6.3e-19
C16909 _015_ fanout45/a_27_47# 6.02e-20
C16910 _053_ _049_ 0.402f
C16911 _316_/a_193_47# _095_ 1.18e-19
C16912 _053_ _318_/a_761_289# 8.36e-20
C16913 clk _331_/a_448_47# 0.00869f
C16914 state\[0\] _318_/a_543_47# 4.69e-20
C16915 output5/a_27_47# _131_ 0.00106f
C16916 _016_ net14 1.04e-20
C16917 _092_ clone7/a_27_47# 2.66e-19
C16918 _100_ _226_/a_27_47# 1.35e-20
C16919 _314_/a_1283_21# _011_ 4.1e-20
C16920 net12 _331_/a_1108_47# 0.00143f
C16921 _067_ _193_/a_109_297# 4.22e-21
C16922 cal_itt\[2\] net2 0.0512f
C16923 _322_/a_1462_47# _078_ 5.11e-19
C16924 _064_ _330_/a_1108_47# 8.48e-20
C16925 _104_ _330_/a_543_47# 3.39e-20
C16926 trim_val\[2\] _057_ 5.23e-20
C16927 _306_/a_193_47# _306_/a_448_47# 0.0642f
C16928 _306_/a_761_289# _306_/a_1108_47# 0.0512f
C16929 _306_/a_27_47# _306_/a_651_413# 9.73e-19
C16930 mask\[6\] _222_/a_199_47# 0.00965f
C16931 _251_/a_27_297# _085_ 1.1e-19
C16932 _327_/a_27_47# _065_ 2.04e-20
C16933 cal_itt\[2\] _305_/a_1283_21# 0.0914f
C16934 _110_ _274_/a_75_212# 0.0044f
C16935 mask\[3\] _065_ 2.22e-20
C16936 _217_/a_109_297# _042_ 4.64e-22
C16937 _326_/a_1108_47# result[5] 1.11e-19
C16938 _331_/a_193_47# _331_/a_639_47# 2.28e-19
C16939 _331_/a_761_289# _331_/a_1270_413# 2.6e-19
C16940 _331_/a_543_47# _331_/a_651_413# 0.0572f
C16941 net54 calibrate 0.0341f
C16942 en_co_clk _206_/a_27_93# 0.00658f
C16943 _215_/a_109_297# _006_ 0.0155f
C16944 _325_/a_27_47# mask\[6\] 0.151f
C16945 _245_/a_109_297# net52 0.00625f
C16946 _245_/a_373_47# _101_ 8.5e-19
C16947 _261_/a_113_47# net19 1.68e-19
C16948 net16 _057_ 1.4e-20
C16949 VPWR _235_/a_79_21# 0.254f
C16950 VPWR net15 2.08f
C16951 net12 net44 0.0433f
C16952 _216_/a_113_297# _042_ 4.09e-19
C16953 _041_ _338_/a_193_47# 1.06e-19
C16954 _189_/a_27_47# _088_ 8.22e-20
C16955 _338_/a_27_47# _338_/a_1032_413# 0.183f
C16956 _338_/a_193_47# _338_/a_1182_261# 0.0728f
C16957 _338_/a_652_21# _338_/a_476_47# 0.26f
C16958 net47 _338_/a_562_413# 1.12e-19
C16959 _308_/a_193_47# _138_/a_27_47# 7.99e-20
C16960 _341_/a_27_47# net47 3.98e-21
C16961 _086_ _310_/a_761_289# 1.59e-22
C16962 output10/a_27_47# net10 0.184f
C16963 trim_mask\[2\] trim_mask\[0\] 2.63e-20
C16964 _328_/a_1108_47# trim_mask\[0\] 5.76e-19
C16965 _030_ _332_/a_193_47# 6.47e-22
C16966 net1 _315_/a_543_47# 0.00105f
C16967 _147_/a_27_47# net17 0.112f
C16968 net35 net2 1.98e-20
C16969 _102_ _101_ 0.00317f
C16970 _074_ _310_/a_1108_47# 5.17e-19
C16971 net54 net45 0.00148f
C16972 _169_/a_215_311# state\[1\] 0.0651f
C16973 _292_/a_493_297# _122_ 0.0107f
C16974 _317_/a_193_47# net41 6.96e-21
C16975 _229_/a_27_297# _087_ 0.0965f
C16976 _326_/a_543_47# output14/a_27_47# 1.43e-20
C16977 _313_/a_27_47# _222_/a_113_297# 2.2e-19
C16978 _170_/a_81_21# _170_/a_299_297# 0.0821f
C16979 _051_ _260_/a_93_21# 0.00143f
C16980 _327_/a_1217_47# _111_ 1.58e-19
C16981 _297_/a_47_47# _297_/a_377_297# 0.00899f
C16982 _110_ clknet_2_2__leaf_clk 1.01f
C16983 VPWR ctlp[0] 0.42f
C16984 _239_/a_277_297# _050_ 7.3e-19
C16985 net31 _270_/a_145_75# 2.11e-20
C16986 _064_ _181_/a_150_297# 4.36e-20
C16987 clone1/a_27_47# _062_ 1.74e-19
C16988 _259_/a_27_297# _335_/a_761_289# 2.67e-19
C16989 _259_/a_109_297# _335_/a_193_47# 4.56e-19
C16990 _107_ _261_/a_113_47# 1.17e-19
C16991 _302_/a_109_297# trim_mask\[4\] 2.67e-20
C16992 _053_ _124_ 1.67e-20
C16993 _341_/a_1108_47# cal_count\[3\] 0.055f
C16994 comp _132_ 0.00448f
C16995 _341_/a_805_47# clknet_2_3__leaf_clk 8.08e-19
C16996 net4 _266_/a_68_297# 0.00574f
C16997 net2 _332_/a_761_289# 1.86e-20
C16998 trim_mask\[0\] _242_/a_297_47# 2.27e-21
C16999 net54 _065_ 0.0165f
C17000 _093_ net1 0.00112f
C17001 _050_ _206_/a_27_93# 0.137f
C17002 _092_ _073_ 4.32e-20
C17003 net31 output36/a_27_47# 0.00817f
C17004 _110_ net11 2.59e-19
C17005 _117_ net19 5.71e-21
C17006 _298_/a_78_199# cal_count\[2\] 0.0138f
C17007 _081_ net52 1.28e-19
C17008 output33/a_27_47# output34/a_27_47# 0.00243f
C17009 VPWR _306_/a_805_47# 6.92e-20
C17010 net2 _288_/a_59_75# 0.138f
C17011 _272_/a_81_21# _334_/a_543_47# 6.99e-19
C17012 _034_ _121_ 0.0165f
C17013 _053_ _262_/a_193_297# 0.018f
C17014 clknet_2_1__leaf_clk _314_/a_448_47# 0.00142f
C17015 _303_/a_761_289# _035_ 7.91e-22
C17016 _307_/a_1108_47# net14 0.00335f
C17017 net15 _318_/a_27_47# 7.97e-21
C17018 _341_/a_193_47# net4 1.23e-21
C17019 result[0] net14 0.00258f
C17020 _043_ _303_/a_543_47# 7.66e-19
C17021 VPWR _049_ 1.51f
C17022 _294_/a_68_297# _130_ 0.175f
C17023 output27/a_27_47# _011_ 0.00178f
C17024 _303_/a_1283_21# net18 6.47e-19
C17025 _294_/a_150_297# _129_ 1.39e-19
C17026 _081_ _214_/a_199_47# 0.00151f
C17027 VPWR _318_/a_761_289# 0.217f
C17028 _029_ _332_/a_639_47# 2.29e-19
C17029 net44 _263_/a_79_21# 9.65e-21
C17030 _315_/a_27_47# output41/a_27_47# 3.29e-20
C17031 trim_mask\[0\] _265_/a_299_297# 0.0595f
C17032 _068_ _065_ 0.00939f
C17033 _190_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.00108f
C17034 _080_ _078_ 0.0018f
C17035 _185_/a_68_297# _096_ 0.00131f
C17036 clk _028_ 0.0679f
C17037 net54 _243_/a_109_297# 4.43e-19
C17038 _060_ _243_/a_27_297# 0.233f
C17039 net35 trim_val\[1\] 0.00225f
C17040 trim_mask\[4\] cal_count\[3\] 1.55e-20
C17041 _058_ net49 0.00402f
C17042 _323_/a_805_47# net47 0.00316f
C17043 _323_/a_543_47# _041_ 7.81e-21
C17044 _266_/a_68_297# _063_ 1.54e-20
C17045 _312_/a_1270_413# net20 4.33e-20
C17046 net55 _075_ 2.15e-19
C17047 fanout43/a_27_47# net45 0.275f
C17048 _299_/a_382_47# _131_ 0.00298f
C17049 clknet_2_1__leaf_clk _310_/a_761_289# 0.0198f
C17050 _047_ trim_val\[0\] 0.039f
C17051 _336_/a_1283_21# _335_/a_27_47# 6.38e-21
C17052 VPWR _233_/a_109_297# 0.179f
C17053 _186_/a_109_297# calibrate 0.00292f
C17054 _341_/a_639_47# _136_ 9.98e-19
C17055 _341_/a_1108_47# _038_ 3.1e-19
C17056 _326_/a_543_47# net26 2.32e-20
C17057 _235_/a_297_47# _094_ 0.0481f
C17058 _331_/a_1283_21# _028_ 0.00204f
C17059 _331_/a_1108_47# clknet_2_2__leaf_clk 1.1e-19
C17060 clknet_2_3__leaf_clk _279_/a_396_47# 4.93e-20
C17061 _110_ trim_val\[0\] 0.00507f
C17062 _331_/a_27_47# trim_mask\[4\] 2.7e-19
C17063 _026_ _057_ 0.00227f
C17064 _304_/a_1283_21# _092_ 4.48e-20
C17065 _119_ net19 0.442f
C17066 _292_/a_78_199# _133_ 1.09e-20
C17067 _128_ _298_/a_78_199# 1.32e-20
C17068 cal_itt\[1\] _064_ 0.00142f
C17069 _325_/a_448_47# _022_ 0.158f
C17070 _325_/a_1217_47# mask\[6\] 8.65e-19
C17071 _317_/a_27_47# _317_/a_651_413# 9.73e-19
C17072 _317_/a_761_289# _317_/a_1108_47# 0.0512f
C17073 _317_/a_193_47# _317_/a_448_47# 0.0594f
C17074 net52 _016_ 0.0278f
C17075 _233_/a_109_297# valid 0.00145f
C17076 _258_/a_373_47# clknet_2_2__leaf_clk 0.00199f
C17077 _326_/a_193_47# _326_/a_448_47# 0.0642f
C17078 _326_/a_761_289# _326_/a_1108_47# 0.0512f
C17079 _326_/a_27_47# _326_/a_651_413# 9.73e-19
C17080 _056_ _108_ 0.00425f
C17081 _325_/a_543_47# _078_ 0.00122f
C17082 _341_/a_193_47# _063_ 1.35e-20
C17083 net12 net11 0.00123f
C17084 net4 _028_ 0.0109f
C17085 net49 _332_/a_27_47# 5.23e-20
C17086 net54 _232_/a_304_297# 0.00231f
C17087 _308_/a_805_47# net14 5.85e-19
C17088 VPWR _317_/a_805_47# 5.66e-20
C17089 _338_/a_652_21# _338_/a_1224_47# 1.57e-19
C17090 _328_/a_1283_21# trim_mask\[2\] 6.44e-20
C17091 _328_/a_1283_21# _328_/a_1108_47# 0.234f
C17092 _328_/a_761_289# _328_/a_651_413# 0.0977f
C17093 _328_/a_543_47# _328_/a_448_47# 0.0498f
C17094 _328_/a_27_47# _328_/a_639_47# 0.00188f
C17095 _328_/a_193_47# _328_/a_1270_413# 1.46e-19
C17096 VPWR _326_/a_805_47# 6.77e-19
C17097 _336_/a_27_47# _108_ 6.55e-19
C17098 _320_/a_543_47# net44 0.152f
C17099 _053_ state\[1\] 0.0276f
C17100 cal_itt\[2\] net55 1.23e-20
C17101 result[7] _314_/a_193_47# 0.0012f
C17102 clknet_2_0__leaf_clk output41/a_27_47# 1.81e-20
C17103 _313_/a_543_47# _085_ 1.84e-19
C17104 net13 _337_/a_639_47# 0.00101f
C17105 _052_ _100_ 0.00194f
C17106 _309_/a_761_289# net14 6.88e-19
C17107 _069_ _195_/a_76_199# 5.64e-21
C17108 _293_/a_81_21# _129_ 0.115f
C17109 _318_/a_27_47# _318_/a_761_289# 0.0701f
C17110 _171_/a_27_47# _054_ 0.23f
C17111 _340_/a_652_21# cal_count\[2\] 1.56e-19
C17112 net42 _088_ 0.00164f
C17113 VPWR _124_ 0.308f
C17114 _119_ _107_ 0.0048f
C17115 _171_/a_27_47# net30 0.185f
C17116 _288_/a_59_75# _123_ 2.1e-21
C17117 state\[2\] _089_ 3.47e-21
C17118 trim[0] trim[1] 0.0363f
C17119 _282_/a_68_297# _120_ 0.103f
C17120 _239_/a_694_21# _060_ 1.71e-19
C17121 net12 _209_/a_27_47# 0.0021f
C17122 _104_ _335_/a_543_47# 1.71e-19
C17123 _064_ _335_/a_1108_47# 0.00192f
C17124 _042_ _311_/a_27_47# 3.4e-21
C17125 _038_ trim_mask\[4\] 1.02e-19
C17126 _086_ _224_/a_199_47# 0.00151f
C17127 net44 _312_/a_639_47# 9.54e-19
C17128 _110_ _279_/a_204_297# 0.00536f
C17129 VPWR _300_/a_129_47# 3.57e-19
C17130 _312_/a_27_47# _312_/a_651_413# 9.73e-19
C17131 _312_/a_761_289# _312_/a_1108_47# 0.0512f
C17132 _312_/a_193_47# _312_/a_448_47# 0.0642f
C17133 input4/a_27_47# output6/a_27_47# 1.74e-20
C17134 _312_/a_27_47# net19 6.86e-20
C17135 _336_/a_1270_413# net46 9.87e-20
C17136 _306_/a_761_289# clknet_2_0__leaf_clk 2.53e-19
C17137 _320_/a_1283_21# net52 2.4e-19
C17138 _306_/a_27_47# net45 1.56e-20
C17139 clknet_2_1__leaf_clk _311_/a_1283_21# 0.00123f
C17140 _195_/a_505_21# _067_ 0.138f
C17141 _323_/a_805_47# net44 1.74e-19
C17142 _329_/a_448_47# _027_ 2e-20
C17143 _329_/a_1108_47# net46 0.266f
C17144 _303_/a_1270_413# clknet_2_3__leaf_clk 3.05e-19
C17145 _091_ _092_ 0.115f
C17146 _323_/a_193_47# net19 0.0188f
C17147 cal_itt\[2\] _067_ 3.46e-19
C17148 mask\[1\] net22 1.8e-20
C17149 VPWR _262_/a_193_297# 0.18f
C17150 _041_ _339_/a_652_21# 0.0173f
C17151 cal_itt\[2\] _070_ 0.166f
C17152 net36 net16 2.74e-19
C17153 mask\[4\] net18 0.00596f
C17154 net47 _339_/a_956_413# 4.53e-19
C17155 _305_/a_639_47# net51 3.68e-19
C17156 _266_/a_150_297# net19 2.11e-19
C17157 _321_/a_193_47# mask\[4\] 2.97e-20
C17158 _341_/a_27_47# clknet_2_2__leaf_clk 1.33e-19
C17159 _323_/a_1283_21# _323_/a_1108_47# 0.234f
C17160 _323_/a_761_289# _323_/a_651_413# 0.0977f
C17161 _323_/a_543_47# _323_/a_448_47# 0.0498f
C17162 _323_/a_27_47# _323_/a_639_47# 0.00188f
C17163 _323_/a_193_47# _323_/a_1270_413# 1.46e-19
C17164 _274_/a_75_212# clknet_2_2__leaf_clk 3.4e-20
C17165 output31/a_27_47# _162_/a_27_47# 8.1e-20
C17166 VPWR _315_/a_1108_47# 0.299f
C17167 _107_ _087_ 0.0797f
C17168 _143_/a_68_297# _040_ 6.46e-21
C17169 _306_/a_448_47# _072_ 1.94e-20
C17170 _337_/a_1283_21# _092_ 7.91e-20
C17171 _337_/a_1108_47# _099_ 2.94e-21
C17172 _094_ net30 2.27e-19
C17173 trim_mask\[2\] _175_/a_68_297# 0.101f
C17174 _328_/a_27_47# _333_/a_448_47# 1.96e-21
C17175 _328_/a_1108_47# _333_/a_193_47# 6.92e-20
C17176 fanout44/a_27_47# _078_ 5.71e-21
C17177 net3 _316_/a_1283_21# 0.00391f
C17178 trim_mask\[2\] _333_/a_193_47# 2.63e-20
C17179 net44 _209_/a_27_47# 0.00315f
C17180 VPWR fanout46/a_27_47# 0.418f
C17181 clknet_2_1__leaf_clk net51 0.331f
C17182 _167_/a_161_47# _099_ 4.06e-21
C17183 _306_/a_27_47# _065_ 9.37e-21
C17184 net16 _334_/a_1270_413# 1.15e-20
C17185 _242_/a_382_297# _242_/a_297_47# 8.13e-19
C17186 clkbuf_0_clk/a_110_47# _190_/a_27_47# 0.012f
C17187 _315_/a_1108_47# valid 5.38e-19
C17188 _292_/a_215_47# _340_/a_1602_47# 6.57e-19
C17189 _306_/a_543_47# net2 2.27e-20
C17190 net14 _095_ 1.78e-20
C17191 _314_/a_1108_47# _313_/a_193_47# 7.01e-21
C17192 _093_ net15 0.00808f
C17193 _306_/a_193_47# _305_/a_448_47# 2.4e-19
C17194 _306_/a_1283_21# _305_/a_543_47# 1.1e-19
C17195 calibrate _317_/a_27_47# 4.43e-22
C17196 net43 _321_/a_639_47# 0.00449f
C17197 output37/a_27_47# trimb[1] 0.337f
C17198 _326_/a_193_47# _074_ 0.0206f
C17199 net9 net46 1.8f
C17200 _266_/a_150_297# _107_ 1.6e-19
C17201 _058_ _106_ 5.05e-19
C17202 _192_/a_548_47# _049_ 4.47e-20
C17203 _320_/a_193_47# _320_/a_1108_47# 0.119f
C17204 _320_/a_27_47# _320_/a_448_47# 0.0864f
C17205 _119_ _279_/a_27_47# 3.79e-19
C17206 net12 ctln[7] 0.00247f
C17207 _309_/a_27_47# _081_ 0.00169f
C17208 VPWR _012_ 0.981f
C17209 _076_ _204_/a_75_212# 7.8e-20
C17210 _189_/a_27_47# _306_/a_1283_21# 5.38e-22
C17211 _261_/a_113_47# _118_ 1.73e-20
C17212 _301_/a_285_47# _134_ 0.0353f
C17213 _178_/a_150_297# net18 3.05e-19
C17214 _331_/a_1217_47# trim_mask\[4\] 2.58e-19
C17215 _187_/a_27_413# _187_/a_212_413# 0.183f
C17216 _317_/a_761_289# clknet_2_0__leaf_clk 0.0196f
C17217 _317_/a_27_47# net45 0.299f
C17218 _317_/a_193_47# _014_ 0.217f
C17219 _308_/a_193_47# _307_/a_193_47# 0.0016f
C17220 _012_ valid 0.0086f
C17221 VPWR _176_/a_27_47# 0.28f
C17222 trim_mask\[2\] trim_mask\[4\] 0.014f
C17223 _328_/a_805_47# clknet_2_2__leaf_clk 2.34e-19
C17224 _262_/a_27_47# _049_ 0.00201f
C17225 _082_ _078_ 0.055f
C17226 _146_/a_68_297# net29 1.71e-20
C17227 VPWR _269_/a_299_297# 0.237f
C17228 _337_/a_1270_413# _034_ 1.66e-20
C17229 net49 _332_/a_1217_47# 3.38e-20
C17230 _263_/a_297_47# _107_ 2.06e-19
C17231 net23 net14 0.00709f
C17232 VPWR state\[1\] 0.552f
C17233 net48 _108_ 0.00244f
C17234 _341_/a_27_47# _341_/a_1217_47# 2.56e-19
C17235 _341_/a_761_289# _341_/a_639_47# 3.16e-19
C17236 net24 net25 1.32e-20
C17237 output21/a_27_47# net20 6.94e-19
C17238 net47 _303_/a_639_47# 9.59e-19
C17239 _301_/a_47_47# trim_val\[0\] 2.33e-21
C17240 _303_/a_1108_47# _338_/a_193_47# 9.13e-19
C17241 _175_/a_68_297# _175_/a_150_297# 0.00477f
C17242 _304_/a_193_47# en_co_clk 2.08e-20
C17243 _315_/a_193_47# net30 1.98e-21
C17244 mask\[0\] _137_/a_150_297# 0.00141f
C17245 clknet_2_2__leaf_clk net11 3.85e-20
C17246 net4 _279_/a_314_297# 0.00558f
C17247 _333_/a_193_47# _333_/a_761_289# 0.186f
C17248 _333_/a_27_47# _333_/a_543_47# 0.107f
C17249 _257_/a_109_297# _119_ 1.08e-19
C17250 _312_/a_27_47# _155_/a_68_297# 2.1e-21
C17251 net16 _332_/a_1108_47# 0.0106f
C17252 _318_/a_1108_47# _318_/a_1270_413# 0.00645f
C17253 _318_/a_761_289# _318_/a_1217_47# 4.2e-19
C17254 _318_/a_543_47# _318_/a_805_47# 0.00171f
C17255 _290_/a_297_47# _125_ 0.00172f
C17256 trim_mask\[4\] _242_/a_297_47# 4.81e-21
C17257 _265_/a_81_21# _265_/a_299_297# 0.0821f
C17258 _203_/a_145_75# _072_ 6.42e-19
C17259 clknet_0_clk mask\[2\] 1.5e-19
C17260 net43 mask\[7\] 0.0343f
C17261 _309_/a_1283_21# _101_ 8.96e-19
C17262 _324_/a_1283_21# net44 0.284f
C17263 _312_/a_1217_47# net19 3.38e-20
C17264 _266_/a_68_297# _279_/a_396_47# 0.00121f
C17265 _324_/a_193_47# _312_/a_193_47# 7.32e-21
C17266 _093_ _049_ 0.0979f
C17267 net52 _205_/a_27_47# 6.74e-22
C17268 VPWR _305_/a_805_47# 1.7e-19
C17269 _048_ _337_/a_27_47# 1.76e-20
C17270 VPWR _250_/a_27_297# 0.313f
C17271 _026_ _027_ 1.14e-19
C17272 _074_ net30 0.0754f
C17273 _185_/a_150_297# _316_/a_193_47# 1.56e-20
C17274 _308_/a_193_47# _308_/a_448_47# 0.0604f
C17275 _308_/a_761_289# _308_/a_1108_47# 0.0512f
C17276 _308_/a_27_47# _308_/a_651_413# 9.73e-19
C17277 _041_ _339_/a_1056_47# 0.00208f
C17278 cal_itt\[0\] _284_/a_68_297# 1.11e-19
C17279 net15 _319_/a_193_47# 0.0179f
C17280 _019_ _321_/a_1283_21# 0.002f
C17281 _090_ _241_/a_105_352# 1.71e-19
C17282 _307_/a_543_47# _307_/a_1108_47# 7.99e-20
C17283 _307_/a_193_47# _307_/a_651_413# 0.0346f
C17284 net48 _031_ 0.00259f
C17285 net9 _332_/a_448_47# 7.31e-20
C17286 _305_/a_761_289# _203_/a_59_75# 1.9e-20
C17287 result[0] _307_/a_543_47# 0.00117f
C17288 _040_ net52 0.153f
C17289 _304_/a_651_413# _001_ 1.44e-20
C17290 _250_/a_27_297# net53 0.185f
C17291 VPWR _319_/a_543_47# 0.223f
C17292 _300_/a_47_47# _300_/a_129_47# 0.00369f
C17293 _322_/a_543_47# net44 0.159f
C17294 _318_/a_27_47# state\[1\] 4.72e-21
C17295 _329_/a_1270_413# _031_ 3.59e-20
C17296 _318_/a_543_47# net45 0.153f
C17297 _233_/a_109_297# _093_ 0.00717f
C17298 _014_ net30 1.8e-20
C17299 trim_val\[0\] clknet_2_2__leaf_clk 2.4e-19
C17300 _289_/a_150_297# _125_ 2.24e-19
C17301 wire42/a_75_212# _049_ 0.00225f
C17302 cal_count\[1\] net47 4.73e-19
C17303 en_co_clk net18 0.00801f
C17304 _270_/a_145_75# _058_ 3.85e-20
C17305 _325_/a_27_47# _321_/a_193_47# 2.01e-19
C17306 _325_/a_193_47# _321_/a_27_47# 5.65e-19
C17307 _293_/a_81_21# _297_/a_47_47# 2.03e-20
C17308 _059_ _100_ 0.0368f
C17309 net12 _044_ 4.19e-20
C17310 VPWR _254_/a_109_297# 0.0075f
C17311 _306_/a_193_47# _002_ 0.00792f
C17312 en_co_clk _129_ 4.52e-19
C17313 _187_/a_27_413# net2 5.73e-21
C17314 _337_/a_193_47# en_co_clk 0.0293f
C17315 _303_/a_27_47# net19 0.015f
C17316 _337_/a_27_47# _120_ 6.92e-19
C17317 _262_/a_27_47# _262_/a_193_297# 0.144f
C17318 output17/a_27_47# net16 5.69e-19
C17319 clkbuf_2_0__f_clk/a_110_47# _192_/a_27_47# 4.09e-20
C17320 _119_ _118_ 3.49e-19
C17321 _323_/a_1108_47# _303_/a_543_47# 3.42e-20
C17322 _323_/a_651_413# _303_/a_193_47# 1.92e-21
C17323 input1/a_75_212# _316_/a_193_47# 1.11e-19
C17324 _339_/a_27_47# _339_/a_381_47# 0.0675f
C17325 _339_/a_193_47# _339_/a_1602_47# 4.25e-19
C17326 _339_/a_652_21# _339_/a_1032_413# 0.00971f
C17327 net13 _320_/a_1108_47# 0.014f
C17328 clone1/a_27_47# _227_/a_209_311# 0.011f
C17329 _172_/a_68_297# _108_ 0.0102f
C17330 _270_/a_59_75# _332_/a_193_47# 1.72e-20
C17331 output8/a_27_47# net46 8.79e-19
C17332 _317_/a_1217_47# net45 6.92e-19
C17333 _320_/a_761_289# _040_ 0.0236f
C17334 trim[4] net16 4.7e-20
C17335 _315_/a_193_47# _315_/a_651_413# 0.0311f
C17336 _315_/a_543_47# _315_/a_1108_47# 7.99e-20
C17337 VPWR _202_/a_297_47# 0.00785f
C17338 output29/a_27_47# net15 1.16e-20
C17339 _321_/a_651_413# mask\[2\] 1.94e-19
C17340 _337_/a_27_47# _076_ 8.74e-20
C17341 net44 _044_ 9.19e-19
C17342 _284_/a_68_297# _108_ 1.4e-20
C17343 clknet_2_2__leaf_clk _279_/a_204_297# 5.17e-20
C17344 _104_ _170_/a_81_21# 0.0544f
C17345 VPWR _336_/a_651_413# 0.144f
C17346 _110_ trim_mask\[3\] 0.121f
C17347 _116_ trim_val\[3\] 0.00305f
C17348 _303_/a_805_47# _063_ 6.23e-21
C17349 VPWR _329_/a_1283_21# 0.375f
C17350 _319_/a_193_47# _049_ 0.00111f
C17351 net8 _334_/a_1108_47# 0.0184f
C17352 _078_ _247_/a_27_297# 0.0114f
C17353 _312_/a_543_47# _045_ 1.35e-19
C17354 net55 _170_/a_81_21# 1.88e-19
C17355 net23 net52 0.00459f
C17356 net46 _055_ 0.00649f
C17357 _050_ _337_/a_193_47# 1.33e-19
C17358 output14/a_27_47# result[7] 0.0905f
C17359 ctlp[0] output29/a_27_47# 6.9e-19
C17360 _286_/a_218_374# _123_ 0.00109f
C17361 result[5] _078_ 4.73e-20
C17362 mask\[6\] net15 0.0927f
C17363 _008_ _101_ 0.00877f
C17364 _164_/a_161_47# net4 3.57e-20
C17365 calibrate _315_/a_448_47# 8.06e-19
C17366 _074_ _315_/a_651_413# 0.00346f
C17367 _012_ _315_/a_543_47# 0.00484f
C17368 _122_ net46 1.07e-20
C17369 _322_/a_761_289# _320_/a_1283_21# 1.22e-19
C17370 _322_/a_193_47# _320_/a_1108_47# 5.87e-21
C17371 _326_/a_1108_47# _251_/a_109_297# 1.24e-19
C17372 trimb[0] net36 0.0182f
C17373 _260_/a_250_297# _092_ 4.55e-21
C17374 _060_ _316_/a_1108_47# 1.92e-20
C17375 _246_/a_109_297# _101_ 0.0301f
C17376 VPWR _210_/a_199_47# 1.43e-19
C17377 _308_/a_193_47# _005_ 0.308f
C17378 _308_/a_27_47# net43 0.313f
C17379 mask\[1\] clknet_0_clk 1.17e-19
C17380 net10 output9/a_27_47# 3.69e-20
C17381 _328_/a_193_47# _025_ 0.219f
C17382 _143_/a_150_297# mask\[2\] 3.43e-19
C17383 _051_ _048_ 0.486f
C17384 ctlp[7] net21 0.0401f
C17385 net15 _319_/a_1462_47# 6.83e-20
C17386 clknet_2_0__leaf_clk _315_/a_1270_413# 1.67e-19
C17387 _014_ _315_/a_651_413# 7.28e-21
C17388 net45 _315_/a_448_47# 2.47e-19
C17389 _305_/a_448_47# _072_ 2.59e-19
C17390 cal_itt\[0\] _230_/a_59_75# 0.0479f
C17391 mask\[5\] _101_ 0.382f
C17392 net47 _001_ 0.0228f
C17393 clkbuf_2_0__f_clk/a_110_47# clknet_2_0__leaf_clk 1.83f
C17394 _300_/a_285_47# _135_ 0.0439f
C17395 _305_/a_27_47# _065_ 8.53e-20
C17396 _309_/a_1108_47# _308_/a_1108_47# 2.99e-21
C17397 _093_ _012_ 0.0256f
C17398 _078_ rebuffer6/a_27_47# 9.27e-20
C17399 _110_ _330_/a_1283_21# 0.0103f
C17400 state\[2\] _092_ 2.44e-20
C17401 _336_/a_543_47# net30 3.34e-21
C17402 _305_/a_543_47# net2 1.86e-19
C17403 net43 _320_/a_1108_47# 5.92e-19
C17404 trim_mask\[0\] en_co_clk 4.6e-20
C17405 _323_/a_1283_21# mask\[4\] 0.122f
C17406 _321_/a_27_47# mask\[3\] 0.00649f
C17407 _321_/a_193_47# net25 6.82e-20
C17408 _305_/a_193_47# _305_/a_448_47# 0.0612f
C17409 _305_/a_761_289# _305_/a_1108_47# 0.0512f
C17410 _305_/a_27_47# _305_/a_651_413# 9.73e-19
C17411 trim[1] net35 0.0359f
C17412 _036_ _037_ 2.57e-20
C17413 VPWR _097_ 0.461f
C17414 _309_/a_27_47# _309_/a_761_289# 0.0701f
C17415 VPWR _313_/a_193_47# 0.593f
C17416 _088_ _098_ 2.83e-19
C17417 input2/a_27_47# net34 0.00866f
C17418 _188_/a_27_47# output35/a_27_47# 0.00787f
C17419 _239_/a_277_297# _049_ 0.0076f
C17420 _277_/a_75_212# net50 0.00108f
C17421 net5 input2/a_27_47# 0.00102f
C17422 _093_ state\[1\] 3.64e-20
C17423 _303_/a_1217_47# net19 1.84e-19
C17424 _337_/a_1462_47# en_co_clk 5.11e-19
C17425 _262_/a_205_47# _105_ 1.74e-20
C17426 _106_ _227_/a_109_93# 3.64e-19
C17427 _328_/a_27_47# trim_val\[3\] 8.55e-21
C17428 _332_/a_1108_47# net40 7.08e-20
C17429 _192_/a_174_21# _096_ 2.5e-20
C17430 cal_itt\[0\] clknet_0_clk 0.00304f
C17431 trim_mask\[2\] _178_/a_68_297# 4.08e-20
C17432 _019_ _101_ 0.0725f
C17433 net12 _166_/a_161_47# 0.00737f
C17434 _339_/a_1032_413# _339_/a_1056_47# 0.0016f
C17435 _339_/a_381_47# _339_/a_586_47# 3.7e-19
C17436 _206_/a_27_93# _049_ 0.00282f
C17437 _107_ _099_ 0.0643f
C17438 _189_/a_27_47# _189_/a_218_47# 0.00788f
C17439 clknet_0_clk _088_ 5.9e-20
C17440 _271_/a_75_212# _112_ 7.61e-19
C17441 _002_ net30 0.00184f
C17442 _294_/a_68_297# _294_/a_150_297# 0.00477f
C17443 _078_ net29 0.109f
C17444 comp clkc 0.0375f
C17445 cal_itt\[1\] _304_/a_448_47# 7.03e-20
C17446 net44 _208_/a_505_21# 2.17e-19
C17447 _128_ trimb[1] 1.84e-19
C17448 _110_ _181_/a_68_297# 3.09e-19
C17449 result[1] _074_ 0.00166f
C17450 _051_ _076_ 8.68e-19
C17451 _128_ _339_/a_193_47# 8.08e-20
C17452 _292_/a_215_47# _339_/a_1032_413# 1.16e-19
C17453 trim_mask\[0\] _050_ 3.24e-20
C17454 net13 net28 3.54e-20
C17455 net44 mask\[2\] 0.00622f
C17456 _319_/a_1462_47# _049_ 9.02e-20
C17457 ctlp[2] ctlp[3] 0.00303f
C17458 net28 _155_/a_68_297# 0.105f
C17459 _279_/a_27_47# _279_/a_206_47# 0.00106f
C17460 _279_/a_396_47# _279_/a_314_297# 0.12f
C17461 _303_/a_193_47# _303_/a_448_47# 0.0612f
C17462 _303_/a_761_289# _303_/a_1108_47# 0.0512f
C17463 _303_/a_27_47# _303_/a_651_413# 9.73e-19
C17464 _325_/a_543_47# mask\[7\] 2.6e-20
C17465 _162_/a_27_47# net37 0.0246f
C17466 output28/a_27_47# net28 0.225f
C17467 en_co_clk _297_/a_47_47# 2.85e-20
C17468 _290_/a_207_413# cal_count\[0\] 0.00352f
C17469 clknet_2_1__leaf_clk _086_ 0.00107f
C17470 _341_/a_27_47# _231_/a_161_47# 4.77e-19
C17471 _237_/a_505_21# _092_ 3.2e-21
C17472 _237_/a_218_374# _099_ 2.1e-19
C17473 net31 trimb[1] 0.109f
C17474 net54 _337_/a_27_47# 0.00143f
C17475 net50 _063_ 2.42e-20
C17476 cal_itt\[2\] clknet_2_3__leaf_clk 2.4e-19
C17477 _314_/a_761_289# net14 0.00489f
C17478 _019_ _320_/a_27_47# 1.79e-19
C17479 _322_/a_761_289# _205_/a_27_47# 0.00152f
C17480 _326_/a_805_47# mask\[6\] 1.94e-21
C17481 _326_/a_1108_47# _022_ 4.8e-20
C17482 _321_/a_27_47# _310_/a_1283_21# 5.37e-21
C17483 _042_ clknet_2_0__leaf_clk 1.44e-20
C17484 _326_/a_761_289# _078_ 0.0108f
C17485 net24 net15 0.00618f
C17486 _256_/a_109_297# net46 2.51e-20
C17487 _324_/a_543_47# _324_/a_1108_47# 7.99e-20
C17488 _324_/a_193_47# _324_/a_651_413# 0.0346f
C17489 _327_/a_543_47# clknet_2_3__leaf_clk 1.94e-19
C17490 _306_/a_27_47# _204_/a_75_212# 0.00414f
C17491 net13 _099_ 0.00749f
C17492 net4 _330_/a_1108_47# 9.85e-20
C17493 _017_ _101_ 8.39e-20
C17494 net12 _325_/a_1108_47# 7.56e-21
C17495 clknet_0_clk _108_ 1.25e-20
C17496 _308_/a_1217_47# net43 0.00157f
C17497 _308_/a_1270_413# net23 5.16e-20
C17498 _015_ _048_ 2.39e-20
C17499 net21 _222_/a_113_297# 4.04e-19
C17500 _316_/a_27_47# net41 0.19f
C17501 VPWR result[2] 0.514f
C17502 _053_ clkbuf_2_2__f_clk/a_110_47# 4.79e-19
C17503 _002_ _072_ 0.0998f
C17504 _319_/a_1283_21# net45 6.73e-19
C17505 _319_/a_448_47# clknet_2_0__leaf_clk 0.0139f
C17506 mask\[1\] _245_/a_27_297# 0.0982f
C17507 output23/a_27_47# result[1] 0.157f
C17508 VPWR _211_/a_109_297# 0.00632f
C17509 _341_/a_27_47# _001_ 5.83e-20
C17510 _048_ _242_/a_79_21# 0.124f
C17511 fanout46/a_27_47# _336_/a_1108_47# 0.00191f
C17512 state\[1\] _243_/a_109_47# 1.67e-19
C17513 _309_/a_543_47# net43 0.157f
C17514 _325_/a_193_47# _046_ 6.44e-20
C17515 _309_/a_27_47# net23 3.7e-20
C17516 net15 _282_/a_150_297# 1.95e-19
C17517 _289_/a_68_297# cal_count\[0\] 4.41e-19
C17518 _327_/a_805_47# net18 2.75e-19
C17519 _053_ _304_/a_543_47# 0.0172f
C17520 _106_ net30 0.084f
C17521 trim[4] net40 0.00188f
C17522 _305_/a_193_47# _002_ 0.23f
C17523 en_co_clk _090_ 0.00578f
C17524 input2/a_27_47# _133_ 1.69e-19
C17525 VPWR _313_/a_1462_47# 8.13e-20
C17526 _254_/a_109_297# wire42/a_75_212# 6.01e-20
C17527 _309_/a_543_47# _309_/a_805_47# 0.00171f
C17528 _309_/a_761_289# _309_/a_1217_47# 4.2e-19
C17529 _309_/a_1108_47# _309_/a_1270_413# 0.00645f
C17530 _319_/a_1283_21# _065_ 8.51e-19
C17531 trim_mask\[3\] clknet_2_2__leaf_clk 0.0111f
C17532 _110_ _334_/a_448_47# 1.14e-20
C17533 _190_/a_27_47# _190_/a_215_47# 0.0716f
C17534 net3 _263_/a_297_47# 2.03e-19
C17535 _146_/a_68_297# _042_ 0.106f
C17536 _322_/a_193_47# _322_/a_1108_47# 0.125f
C17537 _322_/a_27_47# _322_/a_448_47# 0.0931f
C17538 net43 net28 0.435f
C17539 _110_ _327_/a_1283_21# 4.67e-19
C17540 _241_/a_297_47# _092_ 0.0603f
C17541 _305_/a_639_47# clknet_2_1__leaf_clk 1.98e-20
C17542 _320_/a_27_47# _017_ 0.383f
C17543 _320_/a_543_47# mask\[2\] 3.55e-19
C17544 input1/a_75_212# net14 0.00531f
C17545 trim_val\[1\] _056_ 5.31e-19
C17546 net12 mask\[1\] 1.8e-20
C17547 _332_/a_761_289# clknet_2_3__leaf_clk 1.75e-20
C17548 _259_/a_27_297# _064_ 0.0954f
C17549 _104_ _189_/a_27_47# 6.3e-22
C17550 _119_ _062_ 1.74e-19
C17551 _327_/a_761_289# _136_ 9.25e-19
C17552 net13 _246_/a_27_297# 1.03e-19
C17553 net43 _158_/a_68_297# 3.83e-20
C17554 _336_/a_27_47# _336_/a_193_47# 0.735f
C17555 cal_itt\[0\] net47 0.28f
C17556 _303_/a_543_47# mask\[4\] 0.0017f
C17557 net9 _111_ 0.174f
C17558 clknet_2_1__leaf_clk _319_/a_761_289# 1.4e-19
C17559 _023_ _007_ 2.04e-20
C17560 _319_/a_193_47# _319_/a_543_47# 0.22f
C17561 _319_/a_27_47# _319_/a_1283_21# 0.0436f
C17562 comp _130_ 9.2e-19
C17563 _308_/a_27_47# _080_ 1.26e-19
C17564 _189_/a_27_47# net55 8.85e-21
C17565 _325_/a_1270_413# _101_ 1.05e-20
C17566 _325_/a_448_47# net52 1.96e-20
C17567 _324_/a_1283_21# _044_ 5.4e-19
C17568 _116_ _335_/a_543_47# 0.00144f
C17569 _117_ _335_/a_761_289# 0.00241f
C17570 _110_ _335_/a_1283_21# 3.09e-19
C17571 _249_/a_27_297# _249_/a_109_297# 0.171f
C17572 _050_ _090_ 0.0666f
C17573 _341_/a_1108_47# en_co_clk 1.08e-19
C17574 _279_/a_206_47# _118_ 3.03e-20
C17575 _303_/a_193_47# _000_ 0.214f
C17576 mask\[1\] net44 0.145f
C17577 _047_ _108_ 0.00591f
C17578 VPWR _240_/a_109_297# 0.00584f
C17579 _282_/a_150_297# _049_ 2.91e-19
C17580 _324_/a_193_47# mask\[5\] 5.97e-19
C17581 _034_ _095_ 4.95e-20
C17582 _317_/a_193_47# _316_/a_1108_47# 9.92e-21
C17583 _317_/a_543_47# _316_/a_543_47# 9.85e-20
C17584 _292_/a_493_297# _128_ 6.9e-20
C17585 cal_itt\[1\] clk 1.25e-20
C17586 net43 result[3] 6.6e-20
C17587 _028_ _330_/a_543_47# 1.48e-21
C17588 clknet_2_2__leaf_clk _330_/a_1283_21# 0.00182f
C17589 _110_ _332_/a_543_47# 1.5e-20
C17590 _110_ _108_ 0.0421f
C17591 _169_/a_373_53# _051_ 0.00165f
C17592 clk _052_ 0.0283f
C17593 clk input1/a_75_212# 5.57e-20
C17594 VPWR _316_/a_639_47# 1.96e-19
C17595 net54 _051_ 0.00909f
C17596 net30 output30/a_27_47# 0.246f
C17597 net34 trimb[4] 0.0785f
C17598 net12 _088_ 3.71e-19
C17599 net30 _278_/a_109_297# 8.41e-21
C17600 _024_ net46 0.0203f
C17601 _306_/a_448_47# _003_ 0.158f
C17602 _064_ trim_mask\[1\] 0.273f
C17603 _106_ _262_/a_465_47# 5.46e-19
C17604 VPWR clkbuf_2_2__f_clk/a_110_47# 1.25f
C17605 _136_ _332_/a_193_47# 0.00381f
C17606 _104_ _336_/a_27_47# 0.267f
C17607 _249_/a_27_297# mask\[4\] 0.0611f
C17608 _316_/a_1217_47# net41 8.27e-19
C17609 _097_ _093_ 0.507f
C17610 ctlp[7] _045_ 0.0227f
C17611 _074_ _313_/a_543_47# 2.34e-20
C17612 _053_ _302_/a_109_47# 0.00306f
C17613 _232_/a_32_297# _096_ 0.0796f
C17614 _331_/a_1283_21# _052_ 2.16e-19
C17615 net4 _195_/a_535_374# 2.01e-19
C17616 _330_/a_448_47# net19 0.00495f
C17617 trim_mask\[2\] _334_/a_27_47# 0.00247f
C17618 VPWR _304_/a_543_47# 0.207f
C17619 cal_itt\[1\] net4 0.407f
C17620 _125_ net38 1.01e-19
C17621 net13 _084_ 5.3e-20
C17622 net4 _052_ 8.16e-20
C17623 _327_/a_651_413# _024_ 0.00219f
C17624 _327_/a_805_47# trim_mask\[0\] 3.21e-21
C17625 _155_/a_68_297# _084_ 8.19e-19
C17626 _219_/a_109_297# _008_ 0.0125f
C17627 net9 _065_ 3.57e-20
C17628 _129_ output40/a_27_47# 2.28e-19
C17629 _305_/a_1462_47# _002_ 7.49e-19
C17630 net2 _126_ 0.0842f
C17631 mask\[6\] _250_/a_27_297# 0.121f
C17632 net9 _135_ 4.07e-19
C17633 trim_val\[1\] _173_/a_27_47# 0.1f
C17634 _101_ _310_/a_27_47# 5.73e-22
C17635 net13 _236_/a_109_297# 1.33e-19
C17636 _110_ _031_ 0.188f
C17637 cal_count\[1\] _131_ 1.02e-20
C17638 _328_/a_761_289# _058_ 0.0021f
C17639 _322_/a_27_47# _019_ 0.167f
C17640 _019_ _248_/a_27_297# 0.117f
C17641 _114_ _056_ 1.67e-19
C17642 clkbuf_2_1__f_clk/a_110_47# mask\[0\] 3.73e-19
C17643 net48 trim_val\[1\] 9.98e-21
C17644 _272_/a_81_21# trim_val\[2\] 0.189f
C17645 _102_ _310_/a_1108_47# 0.00168f
C17646 _202_/a_79_21# _202_/a_297_47# 0.0326f
C17647 _040_ _208_/a_76_199# 1.12e-19
C17648 _320_/a_543_47# mask\[1\] 0.0346f
C17649 cal_itt\[1\] _063_ 0.39f
C17650 clkbuf_2_0__f_clk/a_110_47# _078_ 1.16e-19
C17651 _336_/a_761_289# _336_/a_805_47# 3.69e-19
C17652 _336_/a_193_47# _336_/a_1217_47# 2.36e-20
C17653 _336_/a_543_47# _336_/a_639_47# 0.0138f
C17654 VPWR _035_ 0.222f
C17655 _218_/a_199_47# mask\[4\] 0.0106f
C17656 _053_ _198_/a_27_47# 3.78e-20
C17657 mask\[4\] _220_/a_113_297# 1.03e-20
C17658 _321_/a_193_47# net15 0.0117f
C17659 cal_itt\[0\] _341_/a_27_47# 1.88e-19
C17660 _050_ trim_mask\[4\] 0.228f
C17661 _103_ _262_/a_109_297# 1.2e-19
C17662 _281_/a_253_297# _092_ 0.00575f
C17663 _281_/a_253_47# _095_ 0.0543f
C17664 _319_/a_448_47# _319_/a_639_47# 4.61e-19
C17665 result[4] _023_ 5.22e-19
C17666 _053_ _331_/a_193_47# 1.48e-22
C17667 net16 net49 0.433f
C17668 _272_/a_81_21# net16 0.00258f
C17669 VPWR _256_/a_27_297# 0.259f
C17670 _249_/a_27_297# _020_ 0.119f
C17671 _249_/a_373_47# mask\[5\] 9.23e-19
C17672 trim_mask\[0\] _332_/a_639_47# 0.00131f
C17673 _329_/a_193_47# _329_/a_1108_47# 0.125f
C17674 _329_/a_27_47# _329_/a_448_47# 0.0931f
C17675 _235_/a_79_21# _337_/a_193_47# 4.82e-19
C17676 net15 _337_/a_193_47# 1.08e-20
C17677 VPWR _321_/a_543_47# 0.216f
C17678 _115_ _334_/a_27_47# 0.00138f
C17679 calibrate clone7/a_27_47# 0.0232f
C17680 _104_ net42 1.36e-20
C17681 _204_/a_75_212# cal_itt\[3\] 5.57e-19
C17682 _003_ _203_/a_145_75# 5.24e-20
C17683 clknet_2_1__leaf_clk _313_/a_27_47# 0.851f
C17684 _060_ _089_ 3.49e-19
C17685 _220_/a_113_297# _220_/a_199_47# 2.42e-19
C17686 VPWR _337_/a_543_47# 0.211f
C17687 VPWR _162_/a_27_47# 0.279f
C17688 _096_ net55 0.13f
C17689 _058_ _301_/a_285_47# 1.75e-19
C17690 _324_/a_1462_47# mask\[5\] 6.42e-19
C17691 _234_/a_109_297# _065_ 2.4e-19
C17692 _317_/a_27_47# _013_ 2.38e-19
C17693 _014_ _316_/a_27_47# 0.0202f
C17694 clknet_2_0__leaf_clk _316_/a_193_47# 0.00439f
C17695 net44 _244_/a_27_297# 0.0642f
C17696 _168_/a_207_413# _336_/a_27_47# 3.37e-21
C17697 net42 net55 0.163f
C17698 _141_/a_27_47# net52 0.0406f
C17699 net45 clone7/a_27_47# 1.48e-20
C17700 _015_ net54 0.00246f
C17701 _322_/a_543_47# mask\[2\] 7.1e-19
C17702 net9 _112_ 1.19e-20
C17703 _328_/a_651_413# net46 0.0122f
C17704 net2 output5/a_27_47# 9.38e-19
C17705 _167_/a_161_47# net41 1.11e-19
C17706 _128_ _291_/a_35_297# 0.167f
C17707 net54 _242_/a_79_21# 1.39e-19
C17708 net13 _085_ 6.8e-21
C17709 _309_/a_27_47# _216_/a_113_297# 2.65e-20
C17710 _329_/a_193_47# net9 0.0159f
C17711 _334_/a_448_47# clknet_2_2__leaf_clk 5.24e-19
C17712 _126_ _123_ 2.34e-21
C17713 _026_ _259_/a_109_297# 1.11e-19
C17714 trim_mask\[4\] _228_/a_297_47# 1.96e-19
C17715 mask\[1\] _209_/a_27_47# 0.00518f
C17716 _301_/a_47_47# _332_/a_543_47# 1.61e-20
C17717 _301_/a_47_47# _108_ 1.67e-20
C17718 en_co_clk _190_/a_27_47# 1.15e-19
C17719 _052_ _260_/a_346_47# 0.00403f
C17720 mask\[7\] result[5] 0.00214f
C17721 _023_ net27 2.27e-19
C17722 _074_ sample 0.0136f
C17723 _327_/a_1283_21# clknet_2_2__leaf_clk 0.00475f
C17724 VPWR fanout45/a_27_47# 0.289f
C17725 _027_ net19 0.0148f
C17726 net16 _289_/a_68_297# 5.02e-19
C17727 _325_/a_651_413# net13 5.88e-19
C17728 _341_/a_27_47# _108_ 5.19e-20
C17729 VPWR _340_/a_1602_47# 0.181f
C17730 _053_ _041_ 2.62e-20
C17731 clknet_0_clk _192_/a_174_21# 0.013f
C17732 _275_/a_299_297# _275_/a_384_47# 1.48e-19
C17733 _000_ mask\[5\] 1.37e-19
C17734 _333_/a_27_47# rebuffer1/a_75_212# 6.92e-21
C17735 VPWR _253_/a_299_297# 0.286f
C17736 _275_/a_299_297# _178_/a_150_297# 8.01e-20
C17737 trim[2] _272_/a_299_297# 1.59e-19
C17738 _304_/a_193_47# _124_ 5.74e-22
C17739 _323_/a_543_47# _068_ 6.22e-19
C17740 net3 _099_ 0.0116f
C17741 _178_/a_68_297# _178_/a_150_297# 0.00477f
C17742 _337_/a_193_47# _049_ 0.0219f
C17743 _104_ _168_/a_27_413# 7.15e-20
C17744 _042_ _078_ 0.0121f
C17745 _335_/a_1283_21# clknet_2_2__leaf_clk 4.35e-20
C17746 trim_val\[1\] _172_/a_68_297# 0.239f
C17747 _134_ net46 6.57e-20
C17748 output9/a_27_47# net9 0.172f
C17749 _341_/a_1270_413# net46 1.7e-19
C17750 VPWR output12/a_27_47# 0.487f
C17751 _168_/a_27_413# net55 2.98e-20
C17752 net27 _046_ 0.0365f
C17753 net48 _114_ 0.00155f
C17754 VPWR _198_/a_27_47# 0.222f
C17755 _309_/a_193_47# mask\[1\] 9.34e-20
C17756 _333_/a_1283_21# net46 0.277f
C17757 net42 _168_/a_207_413# 2.09e-21
C17758 _336_/a_448_47# _033_ 0.158f
C17759 VPWR _331_/a_193_47# 0.602f
C17760 _339_/a_1032_413# net37 4.63e-21
C17761 clknet_2_2__leaf_clk _108_ 0.124f
C17762 _332_/a_543_47# clknet_2_2__leaf_clk 0.00121f
C17763 mask\[6\] _313_/a_193_47# 1.19e-20
C17764 net44 _311_/a_805_47# 0.00215f
C17765 net27 _312_/a_761_289# 3.47e-19
C17766 _053_ _260_/a_93_21# 0.00615f
C17767 ctlp[1] result[7] 8.79e-20
C17768 _329_/a_27_47# _026_ 0.174f
C17769 _094_ _337_/a_1108_47# 0.004f
C17770 _274_/a_75_212# _031_ 0.11f
C17771 _059_ net4 3.63e-20
C17772 clkbuf_2_1__f_clk/a_110_47# _121_ 5.11e-19
C17773 net43 _085_ 0.00429f
C17774 _306_/a_1108_47# clk 0.00192f
C17775 _122_ _065_ 0.0791f
C17776 mask\[7\] net29 1.16f
C17777 _262_/a_109_297# clkbuf_2_3__f_clk/a_110_47# 9e-20
C17778 _247_/a_373_47# net52 7e-19
C17779 mask\[5\] _156_/a_27_47# 2.11e-21
C17780 _124_ net18 0.022f
C17781 _065_ _073_ 3.23e-20
C17782 _327_/a_1283_21# trim_val\[0\] 2.3e-20
C17783 net12 _306_/a_1283_21# 0.00158f
C17784 _135_ _122_ 2.59e-19
C17785 _014_ _316_/a_1217_47# 7.1e-20
C17786 net45 _316_/a_805_47# 0.00215f
C17787 _187_/a_27_413# clknet_2_3__leaf_clk 0.2f
C17788 _325_/a_651_413# net43 0.0154f
C17789 state\[2\] state\[0\] 0.0763f
C17790 _058_ _333_/a_805_47# 2.61e-19
C17791 net47 net26 0.00334f
C17792 _058_ _109_ 0.0221f
C17793 _218_/a_113_297# _076_ 5.93e-20
C17794 _309_/a_543_47# _082_ 9.95e-19
C17795 _322_/a_543_47# mask\[1\] 1.91e-19
C17796 _031_ clknet_2_2__leaf_clk 0.0711f
C17797 net8 _056_ 0.00123f
C17798 _308_/a_761_289# fanout43/a_27_47# 0.00118f
C17799 VPWR _041_ 1.69f
C17800 VPWR _338_/a_1182_261# 0.231f
C17801 _306_/a_1283_21# net44 0.341f
C17802 _244_/a_27_297# _209_/a_27_47# 7.42e-20
C17803 _168_/a_27_413# _168_/a_207_413# 0.185f
C17804 _062_ _099_ 2.25e-21
C17805 ctlp[2] net16 0.00725f
C17806 _130_ _132_ 0.345f
C17807 _075_ _095_ 8.5e-20
C17808 _312_/a_27_47# _221_/a_109_297# 5.89e-20
C17809 _326_/a_27_47# _023_ 0.166f
C17810 _326_/a_761_289# mask\[7\] 0.00354f
C17811 _326_/a_193_47# _102_ 0.00182f
C17812 trim_mask\[0\] _049_ 0.00997f
C17813 trim_val\[3\] net50 0.0617f
C17814 _189_/a_218_47# _098_ 9.31e-21
C17815 VPWR _297_/a_129_47# 2.02e-19
C17816 net2 clknet_0_clk 1.8e-20
C17817 _008_ _077_ 1.23e-20
C17818 _286_/a_76_199# _338_/a_27_47# 1.64e-19
C17819 ctlp[3] net17 0.00723f
C17820 _208_/a_76_199# _208_/a_218_374# 0.00557f
C17821 _041_ net53 0.106f
C17822 _305_/a_1283_21# clknet_0_clk 0.00155f
R0 VGND.n7338 VGND.n877 6.95552e+06
R1 VGND.n7339 VGND.n876 6.95552e+06
R2 VGND.n7341 VGND.n875 6.95552e+06
R3 VGND.n7342 VGND.n874 6.95552e+06
R4 VGND.n7344 VGND.n873 6.95552e+06
R5 VGND.n7345 VGND.n872 6.95552e+06
R6 VGND.n7347 VGND.n871 6.95552e+06
R7 VGND.n7348 VGND.n870 6.95552e+06
R8 VGND.n7350 VGND.n869 6.95552e+06
R9 VGND.n7351 VGND.n868 6.95552e+06
R10 VGND.n7353 VGND.n867 6.95552e+06
R11 VGND.n7354 VGND.n866 6.95552e+06
R12 VGND.n7356 VGND.n865 6.95552e+06
R13 VGND.n7357 VGND.n864 6.95552e+06
R14 VGND.n7359 VGND.n863 6.95552e+06
R15 VGND.n7360 VGND.n862 6.95552e+06
R16 VGND.n7362 VGND.n861 6.95552e+06
R17 VGND.n7363 VGND.n860 6.95552e+06
R18 VGND.n7365 VGND.n858 6.95552e+06
R19 VGND.n7366 VGND.n857 6.95552e+06
R20 VGND.n855 VGND.n850 6.95552e+06
R21 VGND.n854 VGND.n851 6.95552e+06
R22 VGND.n853 VGND.n852 113628
R23 VGND.n7338 VGND 52758.8
R24 VGND.n7367 VGND.n850 40822.2
R25 VGND.n7367 VGND.n7366 40822.2
R26 VGND.n7365 VGND.n7364 40822.2
R27 VGND.n7364 VGND.n7363 40822.2
R28 VGND.n7362 VGND.n7361 40822.2
R29 VGND.n7361 VGND.n7360 40822.2
R30 VGND.n7359 VGND.n7358 40822.2
R31 VGND.n7358 VGND.n7357 40822.2
R32 VGND.n7356 VGND.n7355 40822.2
R33 VGND.n7355 VGND.n7354 40822.2
R34 VGND.n7353 VGND.n7352 40822.2
R35 VGND.n7352 VGND.n7351 40822.2
R36 VGND.n7350 VGND.n7349 40822.2
R37 VGND.n7349 VGND.n7348 40822.2
R38 VGND.n7347 VGND.n7346 40822.2
R39 VGND.n7346 VGND.n7345 40822.2
R40 VGND.n7344 VGND.n7343 40822.2
R41 VGND.n7343 VGND.n7342 40822.2
R42 VGND.n7341 VGND.n7340 40822.2
R43 VGND.n7340 VGND.n7339 40822.2
R44 VGND.n852 VGND.n851 19555.6
R45 VGND VGND.n71 9449.04
R46 VGND VGND.n877 8581.37
R47 VGND.n854 VGND.n853 7652.17
R48 VGND.n856 VGND.n855 7652.17
R49 VGND.n857 VGND.n856 7652.17
R50 VGND.n859 VGND.n858 7652.17
R51 VGND.n860 VGND.n859 7652.17
R52 VGND.n3147 VGND.n861 7652.17
R53 VGND.n3147 VGND.n862 7652.17
R54 VGND.n4244 VGND.n863 7652.17
R55 VGND.n4244 VGND.n864 7652.17
R56 VGND.n2734 VGND.n865 7652.17
R57 VGND.n2734 VGND.n866 7652.17
R58 VGND.n2420 VGND.n867 7652.17
R59 VGND.n2420 VGND.n868 7652.17
R60 VGND.n1828 VGND.n869 7652.17
R61 VGND.n1828 VGND.n870 7652.17
R62 VGND.n1370 VGND.n871 7652.17
R63 VGND.n1370 VGND.n872 7652.17
R64 VGND.n1986 VGND.n873 7652.17
R65 VGND.n1986 VGND.n874 7652.17
R66 VGND.n1040 VGND.n875 7652.17
R67 VGND.n1040 VGND.n876 7652.17
R68 VGND.n851 VGND.n850 7007.41
R69 VGND.n7366 VGND.n7365 7007.41
R70 VGND.n7363 VGND.n7362 7007.41
R71 VGND.n7360 VGND.n7359 7007.41
R72 VGND.n7357 VGND.n7356 7007.41
R73 VGND.n7354 VGND.n7353 7007.41
R74 VGND.n7351 VGND.n7350 7007.41
R75 VGND.n7348 VGND.n7347 7007.41
R76 VGND.n7345 VGND.n7344 7007.41
R77 VGND.n7342 VGND.n7341 7007.41
R78 VGND.n7339 VGND.n7338 7007.41
R79 VGND.n4684 VGND 6347.13
R80 VGND.n7327 VGND.n7326 4831.8
R81 VGND VGND.n4132 4509.58
R82 VGND.n941 VGND 4115.78
R83 VGND.n3254 VGND 3245.21
R84 VGND.n4683 VGND 3245.21
R85 VGND.n2663 VGND 3245.21
R86 VGND.n7969 VGND 3245.21
R87 VGND.n5064 VGND 3228.35
R88 VGND.n6287 VGND 2958.62
R89 VGND.n855 VGND.n854 2742.03
R90 VGND.n858 VGND.n857 2742.03
R91 VGND.n861 VGND.n860 2742.03
R92 VGND.n863 VGND.n862 2742.03
R93 VGND.n865 VGND.n864 2742.03
R94 VGND.n867 VGND.n866 2742.03
R95 VGND.n869 VGND.n868 2742.03
R96 VGND.n871 VGND.n870 2742.03
R97 VGND.n873 VGND.n872 2742.03
R98 VGND.n875 VGND.n874 2742.03
R99 VGND.n877 VGND.n876 2742.03
R100 VGND.n7371 VGND 2469.73
R101 VGND.n112 VGND 2469.73
R102 VGND.n111 VGND 2469.73
R103 VGND.n4132 VGND 2469.73
R104 VGND VGND.n5306 2469.73
R105 VGND.n1830 VGND 2469.73
R106 VGND VGND.n1406 2469.73
R107 VGND VGND.n5788 2469.73
R108 VGND.n5789 VGND 2469.73
R109 VGND.n1363 VGND 2469.73
R110 VGND.n6286 VGND 2469.73
R111 VGND.n7971 VGND 2469.73
R112 VGND.n7967 VGND 2469.73
R113 VGND VGND.n4131 2183.14
R114 VGND.n1012 VGND 2104.35
R115 VGND.n969 VGND 2104.35
R116 VGND.n7369 VGND 1694.25
R117 VGND VGND.n5985 1694.25
R118 VGND.n4685 VGND 1677.39
R119 VGND.n4682 VGND 1677.39
R120 VGND.n5065 VGND 1677.39
R121 VGND.n2665 VGND 1677.39
R122 VGND.n5986 VGND 1677.39
R123 VGND.n1987 VGND 1677.39
R124 VGND VGND.n6107 1677.39
R125 VGND.n6108 VGND 1677.39
R126 VGND.n6763 VGND 1677.39
R127 VGND.n7970 VGND 1677.39
R128 VGND.n856 VGND 1432.95
R129 VGND.n859 VGND 1432.95
R130 VGND VGND.n3147 1432.95
R131 VGND VGND.n4244 1432.95
R132 VGND VGND.n2734 1432.95
R133 VGND VGND.n2420 1432.95
R134 VGND VGND.n1828 1432.95
R135 VGND VGND.n1370 1432.95
R136 VGND VGND.n1986 1432.95
R137 VGND VGND.n1040 1432.95
R138 VGND.n853 VGND 1432.95
R139 VGND.n977 VGND 1087.7
R140 VGND.n7579 VGND.n7578 1010.52
R141 VGND.n7372 VGND 927.203
R142 VGND.n7370 VGND 927.203
R143 VGND.n4135 VGND 927.203
R144 VGND.n4134 VGND 927.203
R145 VGND.n4133 VGND 927.203
R146 VGND.n4245 VGND 927.203
R147 VGND.n5066 VGND 927.203
R148 VGND.n5063 VGND 927.203
R149 VGND.n5062 VGND 927.203
R150 VGND.n5336 VGND 927.203
R151 VGND.n6287 VGND 927.203
R152 VGND.n6766 VGND 927.203
R153 VGND.n6764 VGND 927.203
R154 VGND.n7968 VGND 927.203
R155 VGND VGND.n3253 918.774
R156 VGND.n4131 VGND 918.774
R157 VGND.n2664 VGND 918.774
R158 VGND.n5307 VGND 918.774
R159 VGND.n6765 VGND 918.774
R160 VGND.n6762 VGND 918.774
R161 VGND VGND.n7337 912.795
R162 VGND VGND.n5335 910.346
R163 VGND.n852 VGND 792.337
R164 VGND.n6044 VGND.n6043 671.989
R165 VGND VGND.n4134 649.043
R166 VGND VGND.n4682 649.043
R167 VGND VGND.n2664 649.043
R168 VGND.n5306 VGND 649.043
R169 VGND.n5789 VGND 649.043
R170 VGND.n7372 VGND 632.184
R171 VGND VGND.n7371 632.184
R172 VGND VGND.n7369 632.184
R173 VGND VGND.n7368 632.184
R174 VGND VGND.n112 632.184
R175 VGND VGND.n111 632.184
R176 VGND VGND.n71 632.184
R177 VGND.n3253 VGND 632.184
R178 VGND.n3254 VGND 632.184
R179 VGND.n4135 VGND 632.184
R180 VGND VGND.n4133 632.184
R181 VGND.n4245 VGND 632.184
R182 VGND.n4685 VGND 632.184
R183 VGND VGND.n4683 632.184
R184 VGND.n5066 VGND 632.184
R185 VGND VGND.n5065 632.184
R186 VGND VGND.n5064 632.184
R187 VGND VGND.n5063 632.184
R188 VGND VGND.n5062 632.184
R189 VGND.n2665 VGND 632.184
R190 VGND.n5307 VGND 632.184
R191 VGND.n1830 VGND 632.184
R192 VGND VGND.n1829 632.184
R193 VGND.n5336 VGND 632.184
R194 VGND.n5788 VGND 632.184
R195 VGND VGND.n1363 632.184
R196 VGND.n5985 VGND 632.184
R197 VGND.n5986 VGND 632.184
R198 VGND.n1987 VGND 632.184
R199 VGND VGND.n6286 632.184
R200 VGND.n6107 VGND 632.184
R201 VGND.n6108 VGND 632.184
R202 VGND.n6766 VGND 632.184
R203 VGND VGND.n6765 632.184
R204 VGND VGND.n6764 632.184
R205 VGND VGND.n6763 632.184
R206 VGND VGND.n6762 632.184
R207 VGND.n7971 VGND 632.184
R208 VGND VGND.n7970 632.184
R209 VGND VGND.n7969 632.184
R210 VGND VGND.n7967 632.184
R211 VGND VGND.n7370 623.755
R212 VGND VGND.n4684 623.755
R213 VGND VGND.n2663 623.755
R214 VGND VGND.n1406 623.755
R215 VGND.n5335 VGND 623.755
R216 VGND VGND.n7968 623.755
R217 VGND.n6288 VGND.n6287 613.249
R218 VGND.n6107 VGND.n1224 613.249
R219 VGND.n6109 VGND.n6108 613.249
R220 VGND.n2071 VGND.n1987 613.249
R221 VGND.n7370 VGND.n847 613.249
R222 VGND.n7368 VGND.n849 613.249
R223 VGND.n7794 VGND.n71 613.249
R224 VGND.n3255 VGND.n3254 613.249
R225 VGND.n4134 VGND.n3148 613.249
R226 VGND.n4136 VGND.n4135 613.249
R227 VGND.n4131 VGND.n4130 613.249
R228 VGND.n4246 VGND.n4245 613.249
R229 VGND.n4684 VGND.n2897 613.249
R230 VGND.n4682 VGND.n4681 613.249
R231 VGND.n5063 VGND.n2737 613.249
R232 VGND.n5306 VGND.n5305 613.249
R233 VGND.n5335 VGND.n1450 613.249
R234 VGND.n1831 VGND.n1830 613.249
R235 VGND.n5582 VGND.n1406 613.249
R236 VGND.n5790 VGND.n5789 613.249
R237 VGND.n5985 VGND.n5984 613.249
R238 VGND.n5839 VGND.n1363 613.249
R239 VGND.n6286 VGND.n6285 613.249
R240 VGND.n7037 VGND.n977 613.249
R241 VGND.n7198 VGND.n941 613.249
R242 VGND.n7326 VGND.n7325 613.249
R243 VGND.n7092 VGND.n969 613.249
R244 VGND.n6934 VGND.n1012 613.249
R245 VGND.n7969 VGND.n15 613.249
R246 VGND.n1829 VGND.n1396 611.862
R247 VGND.n7967 VGND.n7966 611.862
R248 VGND.n7371 VGND.n178 611.225
R249 VGND.n111 VGND.n80 611.225
R250 VGND.n7643 VGND.n112 611.225
R251 VGND.n6762 VGND.n6761 610.679
R252 VGND.n7972 VGND.n7971 609.497
R253 VGND.n6763 VGND.n1043 609.497
R254 VGND.n6765 VGND.n1041 609.497
R255 VGND.n7369 VGND.n848 609.497
R256 VGND.n7373 VGND.n7372 609.497
R257 VGND.n3253 VGND.n3252 609.497
R258 VGND.n4132 VGND.n3150 609.497
R259 VGND.n4133 VGND.n3149 609.497
R260 VGND.n4683 VGND.n2898 609.497
R261 VGND.n4686 VGND.n4685 609.497
R262 VGND.n5065 VGND.n2735 609.497
R263 VGND.n5067 VGND.n5066 609.497
R264 VGND.n5064 VGND.n2736 609.497
R265 VGND.n5062 VGND.n5061 609.497
R266 VGND.n2664 VGND.n2421 609.497
R267 VGND.n2666 VGND.n2665 609.497
R268 VGND.n5308 VGND.n5307 609.497
R269 VGND.n2663 VGND.n2662 609.497
R270 VGND.n5337 VGND.n5336 609.497
R271 VGND.n5788 VGND.n5787 609.497
R272 VGND.n5987 VGND.n5986 609.497
R273 VGND.n6767 VGND.n6766 609.497
R274 VGND.n6764 VGND.n1042 609.497
R275 VGND VGND.n7367 564.751
R276 VGND.n7364 VGND 564.751
R277 VGND.n7361 VGND 564.751
R278 VGND.n7358 VGND 564.751
R279 VGND.n7355 VGND 564.751
R280 VGND.n7352 VGND 564.751
R281 VGND.n7349 VGND 564.751
R282 VGND.n7346 VGND 564.751
R283 VGND.n7343 VGND 564.751
R284 VGND.n7340 VGND 564.751
R285 VGND.n7332 VGND.n7331 513.789
R286 VGND.n7329 VGND.n7328 497.392
R287 VGND.n7335 VGND.n7334 480.995
R288 VGND.n7333 VGND.n7332 442.733
R289 VGND.n7334 VGND.n7333 431.801
R290 VGND VGND.n977 420.87
R291 VGND.n1012 VGND 409.938
R292 VGND VGND.n969 409.938
R293 VGND VGND.n941 409.938
R294 VGND.n7326 VGND 409.938
R295 VGND.n7328 VGND.n7327 409.938
R296 VGND.n7336 VGND.n7335 371.678
R297 VGND.n7337 VGND 340.524
R298 VGND VGND.n7329 338.882
R299 VGND.n7968 VGND.n16 306.625
R300 VGND.n7970 VGND.n14 306.625
R301 VGND.n7330 VGND 251.429
R302 VGND VGND.n7330 251.429
R303 VGND.n7337 VGND.n7336 251.429
R304 VGND.n9 VGND.n8 232.784
R305 VGND.n7615 VGND.t174 200.476
R306 VGND.n213 VGND.t93 200.149
R307 VGND.n3654 VGND.t191 200.114
R308 VGND.n740 VGND.t155 193.488
R309 VGND.n7714 VGND.t123 193.488
R310 VGND.n7641 VGND.t164 193.44
R311 VGND.n180 VGND.t141 192.531
R312 VGND.n6352 VGND.t63 192.089
R313 VGND.n7429 VGND.t201 191.915
R314 VGND.n7429 VGND.t9 191.915
R315 VGND.n3 VGND.t181 191.915
R316 VGND.n6662 VGND.t137 191.915
R317 VGND.n6662 VGND.t205 191.915
R318 VGND.n2181 VGND.t243 191.915
R319 VGND.n2181 VGND.t46 191.915
R320 VGND.n6048 VGND.t27 191.915
R321 VGND.n6048 VGND.t85 191.915
R322 VGND.n2106 VGND.t128 191.915
R323 VGND.n2106 VGND.t189 191.915
R324 VGND.n6207 VGND.t64 191.915
R325 VGND.n3472 VGND.t29 191.915
R326 VGND.n3472 VGND.t25 191.915
R327 VGND.n128 VGND.t82 191.915
R328 VGND.n128 VGND.t33 191.915
R329 VGND.n3267 VGND.t84 191.915
R330 VGND.n3267 VGND.t136 191.915
R331 VGND.n7566 VGND.t102 191.915
R332 VGND.n7566 VGND.t172 191.915
R333 VGND.n7750 VGND.t208 191.915
R334 VGND.n4031 VGND.t20 191.915
R335 VGND.n4031 VGND.t80 191.915
R336 VGND.n4164 VGND.t238 191.915
R337 VGND.n4164 VGND.t62 191.915
R338 VGND.n2909 VGND.t133 191.915
R339 VGND.n2909 VGND.t198 191.915
R340 VGND.n4259 VGND.t125 191.915
R341 VGND.n4259 VGND.t200 191.915
R342 VGND.n5095 VGND.t8 191.915
R343 VGND.n5095 VGND.t81 191.915
R344 VGND.n2774 VGND.t252 191.915
R345 VGND.n2774 VGND.t58 191.915
R346 VGND.n1496 VGND.t118 191.915
R347 VGND.n1496 VGND.t162 191.915
R348 VGND.n5176 VGND.t145 191.915
R349 VGND.n5176 VGND.t95 191.915
R350 VGND.n5366 VGND.t224 191.915
R351 VGND.n5366 VGND.t28 191.915
R352 VGND.n1702 VGND.t146 191.915
R353 VGND.n1702 VGND.t217 191.915
R354 VGND.n1263 VGND.t160 191.915
R355 VGND.n1263 VGND.t221 191.915
R356 VGND.n1869 VGND.t15 191.915
R357 VGND.n1869 VGND.t73 191.915
R358 VGND.n7915 VGND.t167 191.915
R359 VGND.n7915 VGND.t228 191.915
R360 VGND.n3970 VGND.t32 191.047
R361 VGND.n3840 VGND.t14 190.984
R362 VGND.n6505 VGND.t108 189.316
R363 VGND.n7399 VGND.t87 189.316
R364 VGND.n3914 VGND.t38 189.316
R365 VGND.n4718 VGND.t116 189.316
R366 VGND.n3169 VGND.t196 189.308
R367 VGND.n7973 VGND.t44 189.298
R368 VGND.n7374 VGND.t10 189.298
R369 VGND.n1649 VGND.t215 189.298
R370 VGND.n1103 VGND.t43 188.97
R371 VGND.n514 VGND.t157 186.719
R372 VGND.n646 VGND.t30 186.719
R373 VGND.n664 VGND.t114 186.719
R374 VGND.n669 VGND.t21 186.719
R375 VGND.n346 VGND.t31 186.719
R376 VGND.n301 VGND.t253 186.719
R377 VGND.n326 VGND.t37 186.719
R378 VGND.n7982 VGND.t176 186.719
R379 VGND.n6672 VGND.t227 186.719
R380 VGND.n6693 VGND.t150 186.719
R381 VGND.n6693 VGND.t69 186.719
R382 VGND.n6640 VGND.t177 186.719
R383 VGND.n6633 VGND.t42 186.719
R384 VGND.n6593 VGND.t56 186.719
R385 VGND.n6571 VGND.t131 186.719
R386 VGND.n6532 VGND.t65 186.719
R387 VGND.n916 VGND.t240 186.719
R388 VGND.n7234 VGND.t230 186.719
R389 VGND.n7056 VGND.t207 186.719
R390 VGND.n6958 VGND.t101 186.719
R391 VGND.n6923 VGND.t83 186.719
R392 VGND.n6063 VGND.t226 186.719
R393 VGND.n6056 VGND.t90 186.719
R394 VGND.n6189 VGND.t206 186.719
R395 VGND.n2051 VGND.t72 186.719
R396 VGND.n1223 VGND.t229 186.719
R397 VGND.n6263 VGND.t67 186.719
R398 VGND.n206 VGND.t4 186.719
R399 VGND.n228 VGND.t251 186.719
R400 VGND.n762 VGND.t190 186.719
R401 VGND.n778 VGND.t241 186.719
R402 VGND.n7379 VGND.t78 186.719
R403 VGND.n3205 VGND.t1 186.719
R404 VGND.n3229 VGND.t184 186.719
R405 VGND.n7661 VGND.t153 186.719
R406 VGND.n7683 VGND.t149 186.719
R407 VGND.n7811 VGND.t171 186.719
R408 VGND.n7630 VGND.t35 186.719
R409 VGND.n3143 VGND.t203 186.719
R410 VGND.n4445 VGND.t175 186.719
R411 VGND.n2983 VGND.t165 186.719
R412 VGND.n5085 VGND.t122 186.719
R413 VGND.n2762 VGND.t154 186.719
R414 VGND.n4981 VGND.t124 186.719
R415 VGND.n5028 VGND.t91 186.719
R416 VGND.n4736 VGND.t106 186.719
R417 VGND.n2628 VGND.t34 186.719
R418 VGND.n2485 VGND.t183 186.719
R419 VGND.n2667 VGND.t194 186.719
R420 VGND.n5375 VGND.t152 186.719
R421 VGND.n5399 VGND.t161 186.719
R422 VGND.n1798 VGND.t232 186.719
R423 VGND.n5762 VGND.t159 186.719
R424 VGND.n5916 VGND.t142 186.719
R425 VGND.n6349 VGND.t213 186.719
R426 VGND.n6367 VGND.t49 186.719
R427 VGND.n493 VGND.t168 183.082
R428 VGND.n436 VGND.t100 183.082
R429 VGND.n2183 VGND.t195 183.082
R430 VGND.n885 VGND.t0 183.082
R431 VGND.n7255 VGND.t2 183.082
R432 VGND.n7118 VGND.t163 183.082
R433 VGND.n1014 VGND.t88 183.082
R434 VGND.n6838 VGND.t111 183.082
R435 VGND.n1990 VGND.t110 183.082
R436 VGND.n1123 VGND.t26 183.082
R437 VGND.n3469 VGND.t245 183.082
R438 VGND.n126 VGND.t92 183.082
R439 VGND.n7564 VGND.t52 183.082
R440 VGND.n7658 VGND.t36 183.082
R441 VGND.n4160 VGND.t70 183.082
R442 VGND.n3632 VGND.t192 183.082
R443 VGND.n4269 VGND.t156 183.082
R444 VGND.n4568 VGND.t40 183.082
R445 VGND.n4478 VGND.t218 183.082
R446 VGND.n2975 VGND.t120 183.082
R447 VGND.n1484 VGND.t250 183.082
R448 VGND.n5173 VGND.t170 183.082
R449 VGND.n2511 VGND.t212 183.082
R450 VGND.n1456 VGND.t48 183.082
R451 VGND.n1401 VGND.t16 183.082
R452 VGND.n1398 VGND.t236 183.082
R453 VGND.n1373 VGND.t169 183.082
R454 VGND.n5841 VGND.t166 183.082
R455 VGND.n5926 VGND.t119 183.082
R456 VGND.n1179 VGND.t247 183.082
R457 VGND.n109 VGND.t86 163.852
R458 VGND.n1100 VGND.t139 150.213
R459 VGND.n4999 VGND.t233 148.862
R460 VGND.n6728 VGND.t75 148.846
R461 VGND.n4247 VGND.t144 148.843
R462 VGND.n5831 VGND.t129 148.843
R463 VGND.n6350 VGND.t219 147.3
R464 VGND.n4249 VGND.t231 147.28
R465 VGND.n7955 VGND.t54 147.28
R466 VGND.n7368 VGND 143.296
R467 VGND.n1829 VGND 143.296
R468 VGND.n577 VGND.t138 142.308
R469 VGND.n528 VGND.t94 142.308
R470 VGND.n408 VGND.t66 142.308
R471 VGND.n320 VGND.t182 142.308
R472 VGND.n2196 VGND.t220 142.308
R473 VGND.n968 VGND.t147 142.308
R474 VGND.n6845 VGND.t89 142.308
R475 VGND.n3344 VGND.t239 142.308
R476 VGND.n3413 VGND.t222 142.308
R477 VGND.n3373 VGND.t214 142.308
R478 VGND.n3197 VGND.t132 142.308
R479 VGND.n4035 VGND.t210 142.308
R480 VGND.n4050 VGND.t39 142.308
R481 VGND.n3822 VGND.t178 142.308
R482 VGND.n3850 VGND.t45 142.308
R483 VGND.n4257 VGND.t104 142.308
R484 VGND.n4575 VGND.t7 142.308
R485 VGND.n3004 VGND.t6 142.308
R486 VGND.n4540 VGND.t50 142.308
R487 VGND.n2812 VGND.t211 142.308
R488 VGND.n4773 VGND.t117 142.308
R489 VGND.n2624 VGND.t223 142.308
R490 VGND.n5454 VGND.t185 142.308
R491 VGND.n1755 VGND.t235 142.308
R492 VGND.n1749 VGND.t47 142.308
R493 VGND.n1266 VGND.t180 142.308
R494 VGND.n1943 VGND.t109 142.308
R495 VGND.n1912 VGND.t151 142.308
R496 VGND.n5737 VGND.t158 142.308
R497 VGND.n5891 VGND.t148 142.308
R498 VGND.n1926 VGND.t121 142.308
R499 VGND.n3693 VGND.n3677 124.692
R500 VGND.n2783 VGND.n2782 124.692
R501 VGND.n3692 VGND.n3691 114.398
R502 VGND.n2769 VGND.n2766 114.398
R503 VGND.n7331 VGND 109.317
R504 VGND.n896 VGND.t17 84.847
R505 VGND.n3447 VGND.t248 84.847
R506 VGND.n3261 VGND.t71 84.847
R507 VGND.n2929 VGND.t134 84.847
R508 VGND.n1364 VGND.t225 84.847
R509 VGND.n7784 VGND.t127 84.847
R510 VGND.n3809 VGND.t76 84.847
R511 VGND.n1257 VGND.t135 84.847
R512 VGND.n2085 VGND.t140 82.587
R513 VGND.n6044 VGND.t237 82.1249
R514 VGND.n113 VGND.t41 79.2407
R515 VGND.n4715 VGND.t5 79.2407
R516 VGND.n9 VGND.t57 79.2004
R517 VGND.n172 VGND.t18 79.2004
R518 VGND.n6489 VGND.t115 78.7329
R519 VGND.n1063 VGND.t107 78.7329
R520 VGND.n6162 VGND.t97 78.7329
R521 VGND.n188 VGND.t98 78.7329
R522 VGND.n107 VGND.t53 78.7329
R523 VGND.n4833 VGND.t60 78.7329
R524 VGND.n1602 VGND.t74 78.7329
R525 VGND.n3392 VGND.t51 78.7329
R526 VGND.n3657 VGND.t202 78.7329
R527 VGND.n5093 VGND.t126 78.7329
R528 VGND.n5409 VGND.t61 78.7329
R529 VGND.n1762 VGND.t79 78.7329
R530 VGND.n1064 VGND.t55 76.1558
R531 VGND.n637 VGND.n636 76.0005
R532 VGND.n7212 VGND.n7211 76.0005
R533 VGND.n7178 VGND.n7177 76.0005
R534 VGND.n974 VGND.n973 76.0005
R535 VGND.n1983 VGND.n1982 76.0005
R536 VGND.n3507 VGND.n3506 76.0005
R537 VGND.n3347 VGND.n3346 76.0005
R538 VGND.n758 VGND.n757 76.0005
R539 VGND.n804 VGND.n803 76.0005
R540 VGND.n3297 VGND.n3296 76.0005
R541 VGND.n76 VGND.n75 76.0005
R542 VGND.n4071 VGND.n4070 76.0005
R543 VGND.n3624 VGND.n3623 76.0005
R544 VGND.n3694 VGND.n3693 76.0005
R545 VGND.n3976 VGND.n3975 76.0005
R546 VGND.n3933 VGND.n3932 76.0005
R547 VGND.n4421 VGND.n4420 76.0005
R548 VGND.n3016 VGND.n3015 76.0005
R549 VGND.n3053 VGND.n3052 76.0005
R550 VGND.n2784 VGND.n2783 76.0005
R551 VGND.n4899 VGND.n4898 76.0005
R552 VGND.n1527 VGND.n1526 76.0005
R553 VGND.n2618 VGND.n2617 76.0005
R554 VGND.n2689 VGND.n2688 76.0005
R555 VGND.n5931 VGND.n5930 76.0005
R556 VGND.n5938 VGND.n5937 76.0005
R557 VGND.n7949 VGND.n7948 76.0005
R558 VGND.n6042 VGND.t96 75.1361
R559 VGND.n3628 VGND.t59 75.1361
R560 VGND.n1255 VGND.t244 75.1361
R561 VGND.n1758 VGND.t246 74.3808
R562 VGND.n5000 VGND.t130 74.2621
R563 VGND.n6665 VGND.t113 73.7268
R564 VGND.n4242 VGND.t254 73.7268
R565 VGND.n1101 VGND.t242 68.7721
R566 VGND.n1105 VGND.t12 64.3579
R567 VGND.n7337 VGND 36.3206
R568 VGND.n2031 VGND.n1991 34.6358
R569 VGND.n3951 VGND.n3150 34.6358
R570 VGND.n4563 VGND.n4562 34.6358
R571 VGND.n2993 VGND.n2976 34.6358
R572 VGND.n5475 VGND.n5474 34.6358
R573 VGND.n5522 VGND.n1448 34.6358
R574 VGND.n5607 VGND.n5606 34.6358
R575 VGND.n539 VGND.n439 34.6358
R576 VGND.n541 VGND.n540 34.6358
R577 VGND.n540 VGND.n539 34.6358
R578 VGND.n541 VGND.n437 34.6358
R579 VGND.n614 VGND.n613 34.6358
R580 VGND.n6782 VGND.n6781 34.6358
R581 VGND.n6781 VGND.n1036 34.6358
R582 VGND.n6605 VGND.n1043 34.6358
R583 VGND.n6468 VGND.n6467 34.6358
R584 VGND.n6945 VGND.n1011 34.6358
R585 VGND.n6173 VGND.n6172 34.6358
R586 VGND.n6173 VGND.n1233 34.6358
R587 VGND.n2119 VGND.n2118 34.6358
R588 VGND.n2027 VGND.n2026 34.6358
R589 VGND.n3492 VGND.n3491 34.6358
R590 VGND.n796 VGND.n179 34.6358
R591 VGND.n3280 VGND.n3279 34.6358
R592 VGND.n7776 VGND.n72 34.6358
R593 VGND.n4157 VGND.n3139 34.6358
R594 VGND.n3943 VGND.n3942 34.6358
R595 VGND.n2913 VGND.n2912 34.6358
R596 VGND.n2914 VGND.n2913 34.6358
R597 VGND.n2936 VGND.n2935 34.6358
R598 VGND.n2945 VGND.n2944 34.6358
R599 VGND.n4274 VGND.n4254 34.6358
R600 VGND.n4606 VGND.n4605 34.6358
R601 VGND.n4586 VGND.n4585 34.6358
R602 VGND.n4585 VGND.n2959 34.6358
R603 VGND.n4562 VGND.n4561 34.6358
R604 VGND.n4555 VGND.n2966 34.6358
R605 VGND.n3037 VGND.n3036 34.6358
R606 VGND.n4878 VGND.n2736 34.6358
R607 VGND.n4754 VGND.n4713 34.6358
R608 VGND.n1505 VGND.n1504 34.6358
R609 VGND.n1510 VGND.n1489 34.6358
R610 VGND.n1511 VGND.n1510 34.6358
R611 VGND.n1634 VGND.n1633 34.6358
R612 VGND.n5301 VGND.n5300 34.6358
R613 VGND.n2576 VGND.n2575 34.6358
R614 VGND.n2570 VGND.n2569 34.6358
R615 VGND.n5464 VGND.n5463 34.6358
R616 VGND.n5463 VGND.n1458 34.6358
R617 VGND.n5474 VGND.n1457 34.6358
R618 VGND.n5511 VGND.n5510 34.6358
R619 VGND.n5503 VGND.n5502 34.6358
R620 VGND.n5516 VGND.n5515 34.6358
R621 VGND.n5518 VGND.n1448 34.6358
R622 VGND.n5574 VGND.n1410 34.6358
R623 VGND.n5575 VGND.n5574 34.6358
R624 VGND.n5629 VGND.n5628 34.6358
R625 VGND.n1844 VGND.n1843 34.6358
R626 VGND.n1716 VGND.n1715 34.6358
R627 VGND.n5751 VGND.n5750 34.6358
R628 VGND.n5795 VGND.n1366 34.6358
R629 VGND.n5799 VGND.n1366 34.6358
R630 VGND.n5800 VGND.n5799 34.6358
R631 VGND.n5970 VGND.n5969 34.6358
R632 VGND.n1296 VGND.n1295 34.6358
R633 VGND.n6383 VGND.n6382 34.6358
R634 VGND.n7934 VGND.n7907 34.6358
R635 VGND.n7930 VGND.n7907 34.6358
R636 VGND.n7947 VGND.t105 34.2973
R637 VGND.n635 VGND.t99 34.2973
R638 VGND.n972 VGND.t188 34.2973
R639 VGND.n7176 VGND.t187 34.2973
R640 VGND.n7210 VGND.t234 34.2973
R641 VGND.n1981 VGND.t24 34.2973
R642 VGND.n3505 VGND.t249 34.2973
R643 VGND.n3345 VGND.t199 34.2973
R644 VGND.n802 VGND.t186 34.2973
R645 VGND.n756 VGND.t11 34.2973
R646 VGND.n3295 VGND.t197 34.2973
R647 VGND.n74 VGND.t143 34.2973
R648 VGND.n3622 VGND.t193 34.2973
R649 VGND.n4069 VGND.t22 34.2973
R650 VGND.n3692 VGND.t209 34.2973
R651 VGND.n3931 VGND.t179 34.2973
R652 VGND.n3974 VGND.t216 34.2973
R653 VGND.n3051 VGND.t112 34.2973
R654 VGND.n3014 VGND.t68 34.2973
R655 VGND.n4419 VGND.t103 34.2973
R656 VGND.n2769 VGND.t23 34.2973
R657 VGND.n4897 VGND.t77 34.2973
R658 VGND.n2687 VGND.t204 34.2973
R659 VGND.n1525 VGND.t19 34.2973
R660 VGND.n2616 VGND.t3 34.2973
R661 VGND.n5936 VGND.t13 34.2973
R662 VGND.n5929 VGND.t173 34.2973
R663 VGND.n3179 VGND.n3174 33.5064
R664 VGND.n5523 VGND.n5522 33.5064
R665 VGND.n3704 VGND.n3703 32.377
R666 VGND.n4275 VGND.n4274 32.0005
R667 VGND.n1627 VGND.n1578 31.624
R668 VGND.n1133 VGND.n1132 30.4946
R669 VGND.n2590 VGND.n2589 29.7417
R670 VGND.n1839 VGND.n1751 29.7417
R671 VGND.n4822 VGND.n2872 28.9887
R672 VGND.n6463 VGND.n1107 28.9887
R673 VGND.n6855 VGND 28.9887
R674 VGND.n3425 VGND 28.9887
R675 VGND.n2569 VGND.n2427 28.9887
R676 VGND.n1740 VGND 28.9887
R677 VGND.n7647 VGND.n109 28.9689
R678 VGND.n3720 VGND.n3675 28.6616
R679 VGND.n6618 VGND.n1064 28.4695
R680 VGND.n7076 VGND 28.2358
R681 VGND VGND.n1011 28.2358
R682 VGND.n2914 VGND 28.2358
R683 VGND.n7924 VGND.n7909 28.2358
R684 VGND VGND.n5568 28.2358
R685 VGND.n4561 VGND 27.8593
R686 VGND VGND.n2966 27.8593
R687 VGND.n5623 VGND.n5622 27.4829
R688 VGND.n3062 VGND 27.4829
R689 VGND.n7442 VGND.n7441 26.7299
R690 VGND.n6970 VGND.n1003 26.7299
R691 VGND.n7578 VGND.n7562 26.7299
R692 VGND.n1641 VGND.n1576 26.7299
R693 VGND.n5589 VGND.n5588 26.7299
R694 VGND.n7043 VGND.n7041 26.6009
R695 VGND.n6946 VGND.n6945 26.6009
R696 VGND.n4157 VGND.n4156 26.6009
R697 VGND.n5012 VGND.n5011 26.6009
R698 VGND.n908 VGND.n907 26.314
R699 VGND.n6183 VGND.n6182 26.314
R700 VGND.n2042 VGND.n2041 26.314
R701 VGND.n2989 VGND.n2976 26.314
R702 VGND.n4744 VGND.n4743 26.314
R703 VGND.n5757 VGND.n5756 26.314
R704 VGND.n6379 VGND.n6378 26.314
R705 VGND.n3487 VGND.n3467 25.977
R706 VGND.n1616 VGND.n1579 25.977
R707 VGND.n5575 VGND.n1409 25.977
R708 VGND.n5583 VGND.n1404 25.977
R709 VGND.n2188 VGND.n2178 25.7355
R710 VGND.n4569 VGND.n2898 25.7355
R711 VGND.n4563 VGND.n2962 25.7355
R712 VGND.n5607 VGND.n1399 25.7355
R713 VGND.n6768 VGND.n6767 25.7355
R714 VGND.n7112 VGND.n7111 25.7355
R715 VGND.n2037 VGND.n2036 25.7355
R716 VGND.n2032 VGND.n2031 25.7355
R717 VGND.n2999 VGND.n2997 25.7355
R718 VGND.n5182 VGND.n5181 25.7355
R719 VGND.n2507 VGND.n2506 25.7355
R720 VGND.n5481 VGND.n5480 25.7355
R721 VGND.n5598 VGND.n5597 25.7355
R722 VGND.n5603 VGND.n5602 25.7355
R723 VGND.n4573 VGND.n2898 25.6926
R724 VGND.n5787 VGND.n1371 25.6926
R725 VGND.n7077 VGND.n7076 25.6926
R726 VGND.n6850 VGND.n6835 25.6926
R727 VGND.n2092 VGND.n2091 25.6926
R728 VGND.n3426 VGND.n3425 25.6926
R729 VGND.n3418 VGND.n3417 25.6926
R730 VGND.n846 VGND.n800 25.6926
R731 VGND.n4041 VGND.n4040 25.6926
R732 VGND.n4056 VGND.n4055 25.6926
R733 VGND.n3820 VGND.n3663 25.6926
R734 VGND.n2935 VGND.n2901 25.6926
R735 VGND.n4580 VGND.n2960 25.6926
R736 VGND.n2795 VGND.n2794 25.6926
R737 VGND.n4886 VGND.n4885 25.6926
R738 VGND.n4826 VGND.n2872 25.6926
R739 VGND.n4755 VGND.n4754 25.6926
R740 VGND.n2662 VGND.n2423 25.6926
R741 VGND.n2605 VGND.n2604 25.6926
R742 VGND.n5459 VGND.n1458 25.6926
R743 VGND.n1941 VGND.n1940 25.6926
R744 VGND.n1948 VGND.n1922 25.6926
R745 VGND.n1883 VGND.n1882 25.6926
R746 VGND.n5969 VGND.n5927 25.6926
R747 VGND.n1932 VGND.n1931 25.6926
R748 VGND.n903 VGND.n902 25.6005
R749 VGND.n6177 VGND.n1233 25.6005
R750 VGND.n3180 VGND.n3179 25.6005
R751 VGND.n1511 VGND.n1488 25.6005
R752 VGND.n7936 VGND.n7935 25.6005
R753 VGND.n7929 VGND.n7928 25.6005
R754 VGND.n7920 VGND.n7919 25.6005
R755 VGND.n4551 VGND.n4550 25.4884
R756 VGND.n4968 VGND.n4966 25.4715
R757 VGND.n613 VGND.n411 25.4203
R758 VGND.n3067 VGND.n3065 25.4203
R759 VGND.n5861 VGND.n5859 25.4203
R760 VGND.n7442 VGND.n7427 25.224
R761 VGND.n502 VGND.n449 25.224
R762 VGND.n6794 VGND.n6793 25.224
R763 VGND.n6966 VGND.n6965 25.224
R764 VGND.n6966 VGND.n1003 25.224
R765 VGND.n3491 VGND.n3467 25.224
R766 VGND.n3828 VGND.n3827 25.224
R767 VGND.n3829 VGND.n3828 25.224
R768 VGND.n4845 VGND.n4844 25.224
R769 VGND.n5188 VGND.n5187 25.224
R770 VGND.n1641 VGND.n1640 25.224
R771 VGND.n5588 VGND.n1403 25.224
R772 VGND.n6387 VGND.n6386 25.224
R773 VGND.n7766 VGND.n7765 24.9894
R774 VGND.n3942 VGND.n3633 24.9894
R775 VGND.n3061 VGND.n2973 24.9894
R776 VGND.n1520 VGND.n1519 24.9894
R777 VGND.n2662 VGND.n2422 24.9894
R778 VGND.n6178 VGND.n1232 24.8476
R779 VGND.n4882 VGND.n4881 24.8476
R780 VGND.n5569 VGND.n1411 24.8476
R781 VGND.n6602 VGND.n1043 24.6184
R782 VGND.n1127 VGND.n1121 24.4711
R783 VGND.n3814 VGND.n3665 24.4711
R784 VGND.n2919 VGND.n2906 24.4711
R785 VGND.n2919 VGND.n2918 24.4711
R786 VGND.n1505 VGND.n1490 24.4711
R787 VGND.n1504 VGND.n1492 24.4711
R788 VGND.n1634 VGND.n1577 24.4711
R789 VGND.n1706 VGND.n1701 24.4711
R790 VGND.n5836 VGND.n1362 24.4711
R791 VGND.n5859 VGND.n1359 24.4711
R792 VGND.n7930 VGND.n7929 24.4711
R793 VGND.n1106 VGND.n1105 24.2743
R794 VGND.n7446 VGND.n7427 24.0946
R795 VGND.n6856 VGND.n6855 24.0946
R796 VGND.n6178 VGND.n6177 24.0946
R797 VGND.n3816 VGND.n3663 24.0946
R798 VGND.n2918 VGND.n2907 24.0946
R799 VGND.n4620 VGND.n4619 24.0946
R800 VGND.n1707 VGND.n1706 24.0946
R801 VGND.n7935 VGND.n7934 24.0946
R802 VGND.n2912 VGND.n2909 23.7181
R803 VGND.n4875 VGND.n2736 23.7181
R804 VGND.n534 VGND.n16 23.7181
R805 VGND.n439 VGND.n16 23.7181
R806 VGND.n895 VGND.n894 23.7181
R807 VGND.n7198 VGND.n7197 23.7181
R808 VGND.n7038 VGND.n7037 23.7181
R809 VGND.n6203 VGND.n1224 23.7181
R810 VGND.n2071 VGND.n1985 23.7181
R811 VGND.n847 VGND.n179 23.7181
R812 VGND.n847 VGND.n846 23.7181
R813 VGND.n7794 VGND.n70 23.7181
R814 VGND.n3666 VGND.n3665 23.7181
R815 VGND.n4403 VGND.n4246 23.7181
R816 VGND.n4391 VGND.n4390 23.7181
R817 VGND.n4386 VGND.n4385 23.7181
R818 VGND.n4407 VGND.n4246 23.7181
R819 VGND.n3037 VGND.n2897 23.7181
R820 VGND.n5095 VGND.n5094 23.7181
R821 VGND.n4993 VGND.n2737 23.7181
R822 VGND.n5002 VGND.n5001 23.7181
R823 VGND.n5305 VGND.n1575 23.7181
R824 VGND.n5305 VGND.n5304 23.7181
R825 VGND.n5502 VGND.n1450 23.7181
R826 VGND.n5582 VGND.n1405 23.7181
R827 VGND.n5583 VGND.n5582 23.7181
R828 VGND.n1404 VGND.n1403 23.7181
R829 VGND.n5629 VGND.n1396 23.7181
R830 VGND.n1702 VGND.n1701 23.7181
R831 VGND.n1259 VGND.n1258 23.7181
R832 VGND.n1869 VGND.n1868 23.7181
R833 VGND.n5839 VGND.n1362 23.7181
R834 VGND.n534 VGND.n533 23.4101
R835 VGND.n4181 VGND.n4180 23.1002
R836 VGND.n4556 VGND.n4555 22.9652
R837 VGND.n7447 VGND.n7446 22.9652
R838 VGND.n6772 VGND.n6771 22.9652
R839 VGND.n2994 VGND.n2993 22.9652
R840 VGND.n2580 VGND 22.9652
R841 VGND.n556 VGND.n555 22.5887
R842 VGND.n4875 VGND.n4874 22.5887
R843 VGND.n551 VGND.n434 22.2123
R844 VGND.n555 VGND.n434 22.2123
R845 VGND.n2189 VGND.n2188 22.2123
R846 VGND.n2190 VGND.n2189 22.2123
R847 VGND.n6464 VGND.n6463 22.2123
R848 VGND.n894 VGND.n883 22.2123
R849 VGND.n890 VGND.n883 22.2123
R850 VGND.n6851 VGND.n6850 22.2123
R851 VGND.n6852 VGND.n6851 22.2123
R852 VGND.n2092 VGND.n1976 22.2123
R853 VGND.n2026 VGND.n1992 22.2123
R854 VGND.n3725 VGND.n3724 22.2123
R855 VGND.n2924 VGND.n2903 22.2123
R856 VGND.n5099 VGND.n5094 22.2123
R857 VGND.n5100 VGND.n5099 22.2123
R858 VGND.n2795 VGND.n2763 22.2123
R859 VGND.n5186 VGND.n5172 22.2123
R860 VGND.n5182 VGND.n5172 22.2123
R861 VGND.n1260 VGND.n1259 22.2123
R862 VGND.n1873 VGND.n1868 22.2123
R863 VGND.n1874 VGND.n1873 22.2123
R864 VGND.n1295 VGND.n1253 22.2123
R865 VGND.n4837 VGND.n4836 21.5514
R866 VGND.n4995 VGND.n4993 21.5038
R867 VGND.n6478 VGND.n6477 21.4593
R868 VGND.n6182 VGND.n1232 21.4593
R869 VGND.n3700 VGND.n3699 21.4593
R870 VGND.n5491 VGND.n5490 21.4593
R871 VGND.n5511 VGND.n1449 21.4593
R872 VGND.n5824 VGND.n5822 20.7985
R873 VGND.n6619 VGND.n6618 20.5833
R874 VGND.n3684 VGND.n3146 20.422
R875 VGND.n5008 VGND.n5007 20.3299
R876 VGND.n2067 VGND.n2066 20.1888
R877 VGND.n6491 VGND.n1106 20.103
R878 VGND VGND.n550 20.0885
R879 VGND VGND.n889 20.0885
R880 VGND.n2193 VGND 20.0456
R881 VGND.n5103 VGND 20.0456
R882 VGND.n545 VGND.n437 19.9534
R883 VGND.n3816 VGND.n3815 19.9534
R884 VGND.n7928 VGND.n7909 19.9534
R885 VGND.n7919 VGND.n7914 19.9534
R886 VGND.n6965 VGND.n6964 19.914
R887 VGND.n501 VGND.n450 19.577
R888 VGND.n903 VGND.n879 19.577
R889 VGND.n3475 VGND.n3470 19.577
R890 VGND.n1581 VGND.n1580 19.577
R891 VGND.n1411 VGND.n1410 19.577
R892 VGND VGND.n1867 19.577
R893 VGND.n7936 VGND.n7905 19.577
R894 VGND.n7923 VGND.n7922 19.577
R895 VGND.n6353 VGND.n6350 19.3766
R896 VGND.n546 VGND.n545 19.3355
R897 VGND.n7253 VGND 19.3355
R898 VGND.n6902 VGND 19.3355
R899 VGND.n7572 VGND.n7571 19.3355
R900 VGND.n625 VGND.n624 19.2926
R901 VGND.n7100 VGND.n7099 19.2926
R902 VGND VGND.n6171 19.2926
R903 VGND.n3518 VGND.n3465 19.2926
R904 VGND.n3829 VGND.n3659 19.2926
R905 VGND.n6203 VGND.n6202 18.824
R906 VGND.n3439 VGND.n3438 18.824
R907 VGND.n3379 VGND.n3378 18.824
R908 VGND.n3181 VGND.n3180 18.824
R909 VGND.n4557 VGND.n4556 18.824
R910 VGND.n7186 VGND.n7185 18.5894
R911 VGND.n3403 VGND.n3402 18.5894
R912 VGND.n831 VGND.n830 18.5894
R913 VGND.n5846 VGND.n1360 18.5826
R914 VGND VGND.n501 18.4476
R915 VGND.n879 VGND 18.4476
R916 VGND.n6971 VGND 18.4476
R917 VGND.n3264 VGND 18.4476
R918 VGND.n2771 VGND 18.4476
R919 VGND.n7905 VGND 18.4476
R920 VGND.n3724 VGND.n3675 18.3426
R921 VGND.n313 VGND.n308 18.2791
R922 VGND.n3224 VGND.n3223 18.2791
R923 VGND.n3247 VGND.n3246 18.2791
R924 VGND.n5079 VGND.n2731 18.2791
R925 VGND.n5391 VGND.n5390 18.2791
R926 VGND.n4869 VGND.n4868 18.0711
R927 VGND.n5187 VGND 18.0711
R928 VGND.n1628 VGND.n1627 18.0711
R929 VGND.n6223 VGND.n6222 18.0105
R930 VGND.n7649 VGND.n7647 17.9905
R931 VGND.n110 VGND.n109 17.9122
R932 VGND.n3827 VGND.n3661 17.7867
R933 VGND.n4409 VGND.n4407 17.7459
R934 VGND.n6910 VGND.n6908 17.7007
R935 VGND.n134 VGND.n133 17.7007
R936 VGND.n2655 VGND.n2654 17.6577
R937 VGND.n1817 VGND.n1816 17.6577
R938 VGND.n6353 VGND.n6352 17.6081
R939 VGND.n6202 VGND.n6201 17.5656
R940 VGND.n5900 VGND.n1320 17.4535
R941 VGND.n7430 VGND.n7429 17.3181
R942 VGND.n2107 VGND.n2106 17.3181
R943 VGND.n4164 VGND.n4163 17.3181
R944 VGND.n1496 VGND.n1495 17.3181
R945 VGND.n5192 VGND.n5191 17.3181
R946 VGND.n7915 VGND.n7914 17.3181
R947 VGND.n6685 VGND.n6684 17.1563
R948 VGND.n5113 VGND.n5112 17.0312
R949 VGND.n2682 VGND.n2681 16.9545
R950 VGND.n7221 VGND.n7219 16.9545
R951 VGND.n4452 VGND.n4451 16.9331
R952 VGND.n6843 VGND.n6837 16.7924
R953 VGND.n3959 VGND.n3958 16.7924
R954 VGND.n4267 VGND.n4258 16.7924
R955 VGND.n1538 VGND.n1537 16.7924
R956 VGND.n3378 VGND.n3377 16.6573
R957 VGND.n6085 VGND.n6084 16.6081
R958 VGND.n1291 VGND.n1290 16.6081
R959 VGND.n4385 VGND.n4250 16.5652
R960 VGND.n1831 VGND.n1827 16.5652
R961 VGND.n4048 VGND.n4047 16.2808
R962 VGND.n1856 VGND.n1855 16.2808
R963 VGND.n4430 VGND.n4428 16.1971
R964 VGND.n508 VGND.n507 16.1492
R965 VGND.n2493 VGND.n2492 16.1492
R966 VGND.n5484 VGND.n1454 15.9473
R967 VGND.n1822 VGND.n1753 15.9044
R968 VGND.n5952 VGND.n5951 15.9044
R969 VGND.n3007 VGND.n3003 15.9033
R970 VGND.n6077 VGND.n6076 15.8505
R971 VGND.n3991 VGND.n3990 15.8505
R972 VGND.n1283 VGND.n1282 15.8505
R973 VGND.n7245 VGND.n7244 15.7728
R974 VGND.n7067 VGND.n7066 15.7728
R975 VGND.n681 VGND.n14 15.6833
R976 VGND.n3292 VGND.n3291 15.5776
R977 VGND.n3484 VGND.n3468 15.5708
R978 VGND.n3433 VGND.n3432 15.5279
R979 VGND.n2906 VGND.n2905 15.4358
R980 VGND.n1451 VGND.n1450 15.4358
R981 VGND.n6934 VGND.n6933 15.3963
R982 VGND.n6049 VGND.n6048 15.3963
R983 VGND.n4136 VGND.n3145 15.3963
R984 VGND.n4989 VGND.n2737 15.3963
R985 VGND.n5367 VGND.n5366 15.3963
R986 VGND.n5612 VGND.n1397 15.1944
R987 VGND.n902 VGND.n901 15.1514
R988 VGND.n1271 VGND.n1261 15.1514
R989 VGND.n5743 VGND.n1376 15.1514
R990 VGND.n2604 VGND.n2426 15.0593
R991 VGND.n4581 VGND 15.0593
R992 VGND.n2763 VGND 15.0593
R993 VGND.n1878 VGND.n1867 15.0593
R994 VGND.n3500 VGND.n3499 14.8247
R995 VGND.n4064 VGND.n4063 14.8247
R996 VGND.n2182 VGND.n2181 14.8179
R997 VGND.n1173 VGND.n1172 14.8179
R998 VGND.n6285 VGND.n1124 14.8179
R999 VGND.n129 VGND.n128 14.8179
R1000 VGND.n7567 VGND.n7566 14.8179
R1001 VGND.n5177 VGND.n5176 14.8179
R1002 VGND.n5984 VGND.n5983 14.8179
R1003 VGND.n6285 VGND.n6284 14.8179
R1004 VGND.n630 VGND.n15 14.775
R1005 VGND.n7200 VGND.n7198 14.775
R1006 VGND.n7093 VGND.n7092 14.775
R1007 VGND.n7752 VGND.n7750 14.775
R1008 VGND.n4034 VGND.n4031 14.775
R1009 VGND.n3983 VGND.n3982 14.775
R1010 VGND.n4261 VGND.n4259 14.775
R1011 VGND.n3041 VGND.n2897 14.775
R1012 VGND.n1264 VGND.n1263 14.775
R1013 VGND.n6288 VGND.n1121 14.6829
R1014 VGND.n1840 VGND.n1839 14.6829
R1015 VGND.n1940 VGND.n1923 14.6829
R1016 VGND.n7924 VGND.n7923 14.6829
R1017 VGND.n1793 VGND.n1792 14.6434
R1018 VGND.n5037 VGND.n5036 14.6237
R1019 VGND.n3440 VGND.n3439 14.3662
R1020 VGND.n5491 VGND.n1453 14.3064
R1021 VGND.n3185 VGND.n3172 14.1532
R1022 VGND.n406 VGND.n15 14.0717
R1023 VGND.n7092 VGND.n7091 14.0717
R1024 VGND.n2072 VGND.n2071 14.0717
R1025 VGND.n3480 VGND.n3479 14.065
R1026 VGND.n6663 VGND.n6662 14.0503
R1027 VGND.n1275 VGND.n1261 13.9299
R1028 VGND.n2903 VGND.n2902 13.5534
R1029 VGND.n4002 VGND.n4001 13.3188
R1030 VGND.n3699 VGND.n3698 13.3188
R1031 VGND.n6935 VGND.n6934 13.177
R1032 VGND.n3472 VGND.n3471 13.177
R1033 VGND.n3385 VGND.n3384 13.177
R1034 VGND.n3267 VGND.n3266 13.177
R1035 VGND.n2774 VGND.n2773 13.177
R1036 VGND.n5291 VGND.n5290 13.1375
R1037 VGND.n5847 VGND.n5846 13.0724
R1038 VGND.n5980 VGND.n5979 12.8663
R1039 VGND.n3840 VGND.n3839 12.8336
R1040 VGND.n449 VGND.n448 12.8005
R1041 VGND.n507 VGND.n448 12.8005
R1042 VGND.n6207 VGND.n1224 12.8005
R1043 VGND.n1976 VGND.n1975 12.8005
R1044 VGND.n4029 VGND.n4028 12.8005
R1045 VGND.n4176 VGND.n4162 12.5591
R1046 VGND.n3805 VGND.n3804 12.5161
R1047 VGND.n3266 VGND.n3265 12.424
R1048 VGND.n4558 VGND.n4557 12.424
R1049 VGND.n2773 VGND.n2772 12.424
R1050 VGND.n1879 VGND.n1878 12.424
R1051 VGND.n7922 VGND.n7921 12.424
R1052 VGND.n3804 VGND.n3148 12.0476
R1053 VGND.n1409 VGND.n1408 12.0476
R1054 VGND.n3025 VGND.n3024 11.8129
R1055 VGND.n3388 VGND.n3385 11.7989
R1056 VGND.n1788 VGND.n1787 11.7989
R1057 VGND.n1610 VGND.n1581 11.7632
R1058 VGND.n3410 VGND.n3408 11.7567
R1059 VGND.n3479 VGND.n3470 11.6711
R1060 VGND.n5984 VGND.n1318 11.5582
R1061 VGND.n4270 VGND.n4254 11.4282
R1062 VGND.n1788 VGND.n1757 11.2946
R1063 VGND.n5953 VGND.n5952 11.2946
R1064 VGND.n7921 VGND.n7920 11.2946
R1065 VGND.n5781 VGND.n5780 11.2885
R1066 VGND.n527 VGND.n526 11.2456
R1067 VGND.n6494 VGND.n1106 11.0824
R1068 VGND.n2085 VGND.n2084 11.0085
R1069 VGND.n4169 VGND.n4168 10.9181
R1070 VGND.n1276 VGND.n1275 10.9181
R1071 VGND.n742 VGND.n181 10.9091
R1072 VGND.n2084 VGND.n1979 10.8605
R1073 VGND.n4390 VGND.n4247 10.7135
R1074 VGND.n4386 VGND.n4249 10.7135
R1075 VGND.n5832 VGND.n5831 10.7135
R1076 VGND.n788 VGND.n787 10.5417
R1077 VGND.n5855 VGND.n1359 10.5417
R1078 VGND.n787 VGND.n180 10.4353
R1079 VGND.n659 VGND.n401 10.3645
R1080 VGND.n6584 VGND.n6582 10.3645
R1081 VGND.n3841 VGND.n3149 10.3645
R1082 VGND.n191 VGND.n177 10.333
R1083 VGND.n5954 VGND.n5953 10.307
R1084 VGND.n6495 VGND.n6494 10.2786
R1085 VGND.n6729 VGND.n6727 10.2477
R1086 VGND.n1715 VGND.n1700 10.1652
R1087 VGND.n192 VGND.n191 10.1609
R1088 VGND.n7669 VGND.n7668 10.1609
R1089 VGND.n3815 VGND.n3814 9.78874
R1090 VGND.n1169 VGND.n1168 9.41227
R1091 VGND.n4168 VGND.n4163 9.41227
R1092 VGND.n5836 VGND.n5835 9.41227
R1093 VGND.n2801 VGND.n2800 9.37278
R1094 VGND.n244 VGND.n243 9.3005
R1095 VGND.n254 VGND.n253 9.3005
R1096 VGND.n246 VGND.n245 9.3005
R1097 VGND.n811 VGND.n810 9.3005
R1098 VGND.n3372 VGND.n3371 9.3005
R1099 VGND.n809 VGND.n808 9.3005
R1100 VGND.n3370 VGND.n3369 9.3005
R1101 VGND.n147 VGND.n146 9.3005
R1102 VGND.n145 VGND.n144 9.3005
R1103 VGND.n7699 VGND.n7698 9.3005
R1104 VGND.n7701 VGND.n7700 9.3005
R1105 VGND.n7709 VGND.n7708 9.3005
R1106 VGND.n7835 VGND.n7834 9.3005
R1107 VGND.n3177 VGND.n3174 9.3005
R1108 VGND.n7837 VGND.n7836 9.3005
R1109 VGND.n3176 VGND.n3175 9.3005
R1110 VGND.n3599 VGND.n3598 9.3005
R1111 VGND.n3601 VGND.n3600 9.3005
R1112 VGND.n7830 VGND.n7829 9.3005
R1113 VGND.n7828 VGND.n7827 9.3005
R1114 VGND.n3766 VGND.n3765 9.3005
R1115 VGND.n3880 VGND.n3879 9.3005
R1116 VGND.n3882 VGND.n3881 9.3005
R1117 VGND.n4104 VGND.n4103 9.3005
R1118 VGND.n4102 VGND.n4101 9.3005
R1119 VGND.n3875 VGND.n3874 9.3005
R1120 VGND.n3873 VGND.n3872 9.3005
R1121 VGND.n3768 VGND.n3767 9.3005
R1122 VGND.n4205 VGND.n4204 9.3005
R1123 VGND.n4207 VGND.n4206 9.3005
R1124 VGND.n4184 VGND.n4183 9.3005
R1125 VGND.n4182 VGND.n4181 9.3005
R1126 VGND.n2979 VGND.n2977 9.3005
R1127 VGND.n4480 VGND.n4479 9.3005
R1128 VGND.n4531 VGND.n4530 9.3005
R1129 VGND.n4548 VGND.n4547 9.3005
R1130 VGND.n4529 VGND.n4528 9.3005
R1131 VGND.n2971 VGND.n2970 9.3005
R1132 VGND.n4550 VGND.n4549 9.3005
R1133 VGND.n4278 VGND.n4277 9.3005
R1134 VGND.n4276 VGND.n4275 9.3005
R1135 VGND.n4966 VGND.n4965 9.3005
R1136 VGND.n5146 VGND.n5145 9.3005
R1137 VGND.n4909 VGND.n4908 9.3005
R1138 VGND.n2853 VGND.n2852 9.3005
R1139 VGND.n2851 VGND.n2850 9.3005
R1140 VGND.n4964 VGND.n4963 9.3005
R1141 VGND.n5148 VGND.n5147 9.3005
R1142 VGND.n4948 VGND.n4947 9.3005
R1143 VGND.n5116 VGND.n5115 9.3005
R1144 VGND.n5114 VGND.n5113 9.3005
R1145 VGND.n4823 VGND.n4822 9.3005
R1146 VGND.n4820 VGND.n2735 9.3005
R1147 VGND.n4770 VGND.n4769 9.3005
R1148 VGND.n4772 VGND.n4771 9.3005
R1149 VGND.n4781 VGND.n4780 9.3005
R1150 VGND.n2565 VGND.n2421 9.3005
R1151 VGND.n2630 VGND.n2629 9.3005
R1152 VGND.n1591 VGND.n1590 9.3005
R1153 VGND.n1589 VGND.n1588 9.3005
R1154 VGND.n5261 VGND.n5260 9.3005
R1155 VGND.n2567 VGND.n2427 9.3005
R1156 VGND.n2543 VGND.n2542 9.3005
R1157 VGND.n2541 VGND.n2540 9.3005
R1158 VGND.n5195 VGND.n5194 9.3005
R1159 VGND.n5193 VGND.n5192 9.3005
R1160 VGND.n2707 VGND.n2706 9.3005
R1161 VGND.n2705 VGND.n2704 9.3005
R1162 VGND.n5448 VGND.n5447 9.3005
R1163 VGND.n5450 VGND.n5449 9.3005
R1164 VGND.n5524 VGND.n5523 9.3005
R1165 VGND.n5526 VGND.n5525 9.3005
R1166 VGND.n5532 VGND.n5531 9.3005
R1167 VGND.n5534 VGND.n5533 9.3005
R1168 VGND.n5561 VGND.n5560 9.3005
R1169 VGND.n5559 VGND.n5558 9.3005
R1170 VGND.n1766 VGND.n1765 9.3005
R1171 VGND.n2354 VGND.n2353 9.3005
R1172 VGND.n2352 VGND.n2351 9.3005
R1173 VGND.n1723 VGND.n1722 9.3005
R1174 VGND.n1721 VGND.n1720 9.3005
R1175 VGND.n5901 VGND.n5900 9.3005
R1176 VGND.n5720 VGND.n5679 9.3005
R1177 VGND.n5882 VGND.n5881 9.3005
R1178 VGND.n5880 VGND.n5879 9.3005
R1179 VGND.n1357 VGND.n1356 9.3005
R1180 VGND.n5899 VGND.n5898 9.3005
R1181 VGND.n5711 VGND.n5710 9.3005
R1182 VGND.n5713 VGND.n5712 9.3005
R1183 VGND.n5678 VGND.n5677 9.3005
R1184 VGND.n2310 VGND.n2309 9.3005
R1185 VGND.n2308 VGND.n2307 9.3005
R1186 VGND.n1890 VGND.n1889 9.3005
R1187 VGND.n1888 VGND.n1887 9.3005
R1188 VGND.n6229 VGND.n6228 9.3005
R1189 VGND.n6231 VGND.n6230 9.3005
R1190 VGND.n6236 VGND.n6235 9.3005
R1191 VGND.n6088 VGND.n6087 9.3005
R1192 VGND.n6090 VGND.n6089 9.3005
R1193 VGND.n6224 VGND.n6223 9.3005
R1194 VGND.n6226 VGND.n6225 9.3005
R1195 VGND.n6238 VGND.n6237 9.3005
R1196 VGND.n2278 VGND.n2277 9.3005
R1197 VGND.n2276 VGND.n2275 9.3005
R1198 VGND.n2128 VGND.n2127 9.3005
R1199 VGND.n2126 VGND.n2125 9.3005
R1200 VGND.n7002 VGND.n7001 9.3005
R1201 VGND.n7120 VGND.n7119 9.3005
R1202 VGND.n7273 VGND.n7272 9.3005
R1203 VGND.n7275 VGND.n7274 9.3005
R1204 VGND.n7168 VGND.n7167 9.3005
R1205 VGND.n7166 VGND.n7165 9.3005
R1206 VGND.n7117 VGND.n7116 9.3005
R1207 VGND.n7125 VGND.n7124 9.3005
R1208 VGND.n7000 VGND.n6999 9.3005
R1209 VGND.n7012 VGND.n7011 9.3005
R1210 VGND.n7010 VGND.n7009 9.3005
R1211 VGND.n6878 VGND.n6877 9.3005
R1212 VGND.n1018 VGND.n1017 9.3005
R1213 VGND.n6861 VGND.n6860 9.3005
R1214 VGND.n6859 VGND.n6858 9.3005
R1215 VGND.n6459 VGND.n1041 9.3005
R1216 VGND.n6560 VGND.n6559 9.3005
R1217 VGND.n6580 VGND.n1067 9.3005
R1218 VGND.n6537 VGND.n6536 9.3005
R1219 VGND.n6461 VGND.n1107 9.3005
R1220 VGND.n6418 VGND.n6417 9.3005
R1221 VGND.n6416 VGND.n6415 9.3005
R1222 VGND.n6408 VGND.n6407 9.3005
R1223 VGND.n6406 VGND.n6405 9.3005
R1224 VGND.n2234 VGND.n2233 9.3005
R1225 VGND.n2232 VGND.n2231 9.3005
R1226 VGND.n2202 VGND.n2201 9.3005
R1227 VGND.n2200 VGND.n2199 9.3005
R1228 VGND.n558 VGND.n557 9.3005
R1229 VGND.n370 VGND.n369 9.3005
R1230 VGND.n380 VGND.n379 9.3005
R1231 VGND.n372 VGND.n371 9.3005
R1232 VGND.n566 VGND.n565 9.3005
R1233 VGND.n561 VGND.n560 9.3005
R1234 VGND.n482 VGND.n481 9.3005
R1235 VGND.n480 VGND.n479 9.3005
R1236 VGND.n568 VGND.n567 9.3005
R1237 VGND.n414 VGND.n413 9.3005
R1238 VGND.n7450 VGND.n7449 9.3005
R1239 VGND.n7448 VGND.n7447 9.3005
R1240 VGND.n6522 VGND.n6521 9.28042
R1241 VGND.n7795 VGND.n7794 9.27112
R1242 VGND.n660 VGND.n659 9.24531
R1243 VGND.n5840 VGND.n5839 9.10662
R1244 VGND.n6582 VGND.n1067 9.09293
R1245 VGND.n3703 VGND 9.03579
R1246 VGND.n1792 VGND.n1757 9.03579
R1247 VGND.n1753 VGND.n1752 9.03579
R1248 VGND.n4084 VGND.n4083 9.02922
R1249 VGND.n2820 VGND.n2819 9.02922
R1250 VGND.n5416 VGND.n5415 9.02922
R1251 VGND.n6710 VGND.n6709 9.02922
R1252 VGND.n248 VGND.n247 9.0005
R1253 VGND.n242 VGND.n241 9.0005
R1254 VGND.n739 VGND.n738 9.0005
R1255 VGND.n45 VGND.n44 9.0005
R1256 VGND.n3368 VGND.n3367 9.0005
R1257 VGND.n3544 VGND.n3543 9.0005
R1258 VGND.n3534 VGND.n3533 9.0005
R1259 VGND.n816 VGND.n815 9.0005
R1260 VGND.n150 VGND.n149 9.0005
R1261 VGND.n7826 VGND.n7825 9.0005
R1262 VGND.n7697 VGND.n7696 9.0005
R1263 VGND.n7703 VGND.n7702 9.0005
R1264 VGND.n7716 VGND.n7715 9.0005
R1265 VGND.n7839 VGND.n7838 9.0005
R1266 VGND.n69 VGND.n68 9.0005
R1267 VGND.n3603 VGND.n3602 9.0005
R1268 VGND.n3597 VGND.n3596 9.0005
R1269 VGND.n3871 VGND.n3870 9.0005
R1270 VGND.n4187 VGND.n4186 9.0005
R1271 VGND.n4202 VGND.n4201 9.0005
R1272 VGND.n4209 VGND.n4208 9.0005
R1273 VGND.n3884 VGND.n3883 9.0005
R1274 VGND.n4100 VGND.n4099 9.0005
R1275 VGND.n4106 VGND.n4105 9.0005
R1276 VGND.n3770 VGND.n3769 9.0005
R1277 VGND.n3764 VGND.n3763 9.0005
R1278 VGND.n3068 VGND.n3067 9.0005
R1279 VGND.n4688 VGND.n4687 9.0005
R1280 VGND.n4280 VGND.n4279 9.0005
R1281 VGND.n4473 VGND.n4472 9.0005
R1282 VGND.n4488 VGND.n4487 9.0005
R1283 VGND.n4533 VGND.n4532 9.0005
R1284 VGND.n4546 VGND.n4545 9.0005
R1285 VGND.n5038 VGND.n5037 9.0005
R1286 VGND.n4962 VGND.n4961 9.0005
R1287 VGND.n4914 VGND.n4913 9.0005
R1288 VGND.n2849 VGND.n2848 9.0005
R1289 VGND.n5143 VGND.n5142 9.0005
R1290 VGND.n5150 VGND.n5149 9.0005
R1291 VGND.n4950 VGND.n4949 9.0005
R1292 VGND.n4819 VGND.n4818 9.0005
R1293 VGND.n4768 VGND.n4767 9.0005
R1294 VGND.n4775 VGND.n4774 9.0005
R1295 VGND.n4789 VGND.n4788 9.0005
R1296 VGND.n2528 VGND.n2527 9.0005
R1297 VGND.n2546 VGND.n2545 9.0005
R1298 VGND.n1593 VGND.n1592 9.0005
R1299 VGND.n2634 VGND.n2633 9.0005
R1300 VGND.n1587 VGND.n1586 9.0005
R1301 VGND.n2564 VGND.n2563 9.0005
R1302 VGND.n5198 VGND.n5197 9.0005
R1303 VGND.n2710 VGND.n2709 9.0005
R1304 VGND.n2703 VGND.n2702 9.0005
R1305 VGND.n1739 VGND.n1738 9.0005
R1306 VGND.n2357 VGND.n2356 9.0005
R1307 VGND.n2350 VGND.n2349 9.0005
R1308 VGND.n5563 VGND.n5562 9.0005
R1309 VGND.n5452 VGND.n5451 9.0005
R1310 VGND.n5446 VGND.n5445 9.0005
R1311 VGND.n5528 VGND.n5527 9.0005
R1312 VGND.n5536 VGND.n5535 9.0005
R1313 VGND.n5653 VGND.n5652 9.0005
R1314 VGND.n5897 VGND.n5896 9.0005
R1315 VGND.n5862 VGND.n5861 9.0005
R1316 VGND.n5734 VGND.n5733 9.0005
R1317 VGND.n1893 VGND.n1892 9.0005
R1318 VGND.n1921 VGND.n1909 9.0005
R1319 VGND.n2313 VGND.n2312 9.0005
R1320 VGND.n2306 VGND.n2305 9.0005
R1321 VGND.n5709 VGND.n5708 9.0005
R1322 VGND.n5884 VGND.n5883 9.0005
R1323 VGND.n1307 VGND.n1306 9.0005
R1324 VGND.n6006 VGND.n6005 9.0005
R1325 VGND.n5676 VGND.n5675 9.0005
R1326 VGND.n5722 VGND 9.0005
R1327 VGND VGND.n5721 9.0005
R1328 VGND.n1181 VGND.n1180 9.0005
R1329 VGND.n2131 VGND.n2130 9.0005
R1330 VGND.n2160 VGND.n2146 9.0005
R1331 VGND.n2281 VGND.n2280 9.0005
R1332 VGND.n2274 VGND.n2273 9.0005
R1333 VGND.n6227 VGND.n1219 9.0005
R1334 VGND.n6240 VGND.n6239 9.0005
R1335 VGND.n1236 VGND.n1235 9.0005
R1336 VGND.n6122 VGND.n6121 9.0005
R1337 VGND.n6092 VGND.n6091 9.0005
R1338 VGND.n6864 VGND.n6863 9.0005
R1339 VGND.n6881 VGND.n6880 9.0005
R1340 VGND.n6901 VGND.n6900 9.0005
R1341 VGND.n7129 VGND.n7128 9.0005
R1342 VGND.n7164 VGND.n7163 9.0005
R1343 VGND.n7271 VGND.n7270 9.0005
R1344 VGND.n7277 VGND.n7276 9.0005
R1345 VGND.n7115 VGND.n7114 9.0005
R1346 VGND.n6998 VGND.n6997 9.0005
R1347 VGND.n7004 VGND.n7003 9.0005
R1348 VGND.n7017 VGND.n7013 9.0005
R1349 VGND.n2204 VGND.n2203 9.0005
R1350 VGND.n2237 VGND.n2236 9.0005
R1351 VGND.n2230 VGND.n2229 9.0005
R1352 VGND.n6425 VGND.n6424 9.0005
R1353 VGND.n6541 VGND.n6540 9.0005
R1354 VGND.n6458 VGND.n6457 9.0005
R1355 VGND.n6404 VGND.n6403 9.0005
R1356 VGND.n6410 VGND.n6409 9.0005
R1357 VGND.n484 VGND.n483 9.0005
R1358 VGND.n562 VGND.n433 9.0005
R1359 VGND.n416 VGND.n411 9.0005
R1360 VGND.n7453 VGND.n7452 9.0005
R1361 VGND.n374 VGND.n373 9.0005
R1362 VGND.n368 VGND.n367 9.0005
R1363 VGND.n391 VGND.n390 9.0005
R1364 VGND.n570 VGND.n569 9.0005
R1365 VGND.n478 VGND.n477 9.0005
R1366 VGND.n784 VGND 8.99034
R1367 VGND.n7668 VGND 8.99034
R1368 VGND.n2905 VGND.n2904 8.65932
R1369 VGND.n6208 VGND.n6207 8.54875
R1370 VGND.n3994 VGND.n3627 8.36259
R1371 VGND.n7956 VGND.n7954 8.36259
R1372 VGND.n8 VGND 8.34833
R1373 VGND.n526 VGND.n442 8.23546
R1374 VGND.n522 VGND.n442 8.23546
R1375 VGND.n522 VGND.n521 8.23546
R1376 VGND.n521 VGND.n520 8.23546
R1377 VGND.n520 VGND.n444 8.23546
R1378 VGND.n516 VGND.n444 8.23546
R1379 VGND.n516 VGND.n515 8.23546
R1380 VGND.n513 VGND.n446 8.23546
R1381 VGND.n509 VGND.n446 8.23546
R1382 VGND.n509 VGND.n508 8.23546
R1383 VGND.n652 VGND.n402 8.23546
R1384 VGND.n652 VGND.n651 8.23546
R1385 VGND.n681 VGND.n680 8.23546
R1386 VGND.n7972 VGND.n13 8.23546
R1387 VGND.n13 VGND.n12 8.23546
R1388 VGND.n6684 VGND.n6657 8.23546
R1389 VGND.n6658 VGND.n6657 8.23546
R1390 VGND.n6679 VGND.n6658 8.23546
R1391 VGND.n6727 VGND.n1059 8.23546
R1392 VGND.n6584 VGND.n6583 8.23546
R1393 VGND.n6500 VGND.n6499 8.23546
R1394 VGND.n6504 VGND.n1103 8.23546
R1395 VGND.n6495 VGND.n1104 8.23546
R1396 VGND.n6499 VGND.n1104 8.23546
R1397 VGND.n7221 VGND.n7220 8.23546
R1398 VGND.n7043 VGND.n7042 8.23546
R1399 VGND.n6947 VGND.n6946 8.23546
R1400 VGND.n6947 VGND.n1009 8.23546
R1401 VGND.n6951 VGND.n1009 8.23546
R1402 VGND.n6952 VGND.n6951 8.23546
R1403 VGND.n6953 VGND.n6952 8.23546
R1404 VGND.n6953 VGND.n1007 8.23546
R1405 VGND.n6957 VGND.n1007 8.23546
R1406 VGND.n6960 VGND.n6959 8.23546
R1407 VGND.n6960 VGND.n1005 8.23546
R1408 VGND.n6964 VGND.n1005 8.23546
R1409 VGND.n6910 VGND.n6909 8.23546
R1410 VGND.n6053 VGND.n6046 8.23546
R1411 VGND.n6201 VGND.n1226 8.23546
R1412 VGND.n6197 VGND.n1226 8.23546
R1413 VGND.n6197 VGND.n6196 8.23546
R1414 VGND.n6196 VGND.n6195 8.23546
R1415 VGND.n6195 VGND.n1228 8.23546
R1416 VGND.n6191 VGND.n1228 8.23546
R1417 VGND.n6191 VGND.n6190 8.23546
R1418 VGND.n6188 VGND.n1230 8.23546
R1419 VGND.n6184 VGND.n1230 8.23546
R1420 VGND.n6184 VGND.n6183 8.23546
R1421 VGND.n2066 VGND.n1988 8.23546
R1422 VGND.n6219 VGND.n6218 8.23546
R1423 VGND.n6218 VGND.n6217 8.23546
R1424 VGND.n6217 VGND.n1221 8.23546
R1425 VGND.n6213 VGND.n1221 8.23546
R1426 VGND.n6213 VGND.n6212 8.23546
R1427 VGND.n6212 VGND.n6211 8.23546
R1428 VGND.n138 VGND.n124 8.23546
R1429 VGND.n139 VGND.n138 8.23546
R1430 VGND.n139 VGND.n123 8.23546
R1431 VGND.n143 VGND.n123 8.23546
R1432 VGND.n7373 VGND.n177 8.23546
R1433 VGND.n3240 VGND.n3201 8.23546
R1434 VGND.n3240 VGND.n3239 8.23546
R1435 VGND.n3224 VGND.n3202 8.23546
R1436 VGND.n3252 VGND.n3170 8.23546
R1437 VGND.n3200 VGND.n3170 8.23546
R1438 VGND.n3247 VGND.n3200 8.23546
R1439 VGND.n3186 VGND.n3185 8.23546
R1440 VGND.n3190 VGND.n3171 8.23546
R1441 VGND.n7649 VGND.n7648 8.23546
R1442 VGND.n4156 VGND.n3140 8.23546
R1443 VGND.n4151 VGND.n3141 8.23546
R1444 VGND.n4147 VGND.n3141 8.23546
R1445 VGND.n4147 VGND.n4146 8.23546
R1446 VGND.n4146 VGND.n4145 8.23546
R1447 VGND.n4142 VGND.n4141 8.23546
R1448 VGND.n4141 VGND.n4140 8.23546
R1449 VGND.n4140 VGND.n3145 8.23546
R1450 VGND.n3844 VGND.n3149 8.23546
R1451 VGND.n4430 VGND.n4429 8.23546
R1452 VGND.n4456 VGND.n4240 8.23546
R1453 VGND.n2986 VGND.n2984 8.23546
R1454 VGND.n2986 VGND.n2985 8.23546
R1455 VGND.n5084 VGND.n2729 8.23546
R1456 VGND.n5080 VGND.n5079 8.23546
R1457 VGND.n4968 VGND.n4967 8.23546
R1458 VGND.n4978 VGND.n2855 8.23546
R1459 VGND.n4979 VGND.n4978 8.23546
R1460 VGND.n4982 VGND.n4979 8.23546
R1461 VGND.n4730 VGND.n4729 8.23546
R1462 VGND.n4743 VGND.n4714 8.23546
R1463 VGND.n2731 VGND.n2730 8.23546
R1464 VGND.n5068 VGND.n5067 8.23546
R1465 VGND.n5067 VGND.n2733 8.23546
R1466 VGND.n5286 VGND.n5285 8.23546
R1467 VGND.n5286 VGND.n1648 8.23546
R1468 VGND.n5290 VGND.n1648 8.23546
R1469 VGND.n2650 VGND.n2625 8.23546
R1470 VGND.n2650 VGND.n2649 8.23546
R1471 VGND.n2492 VGND.n2463 8.23546
R1472 VGND.n2681 VGND.n2417 8.23546
R1473 VGND.n2417 VGND.n2416 8.23546
R1474 VGND.n2666 VGND.n2419 8.23546
R1475 VGND.n2466 VGND.n2419 8.23546
R1476 VGND.n2467 VGND.n2466 8.23546
R1477 VGND.n5390 VGND.n5364 8.23546
R1478 VGND.n5406 VGND.n5363 8.23546
R1479 VGND.n1793 VGND.n1756 8.23546
R1480 VGND.n5757 VGND.n1374 8.23546
R1481 VGND.n5904 VGND.n1320 8.23546
R1482 VGND.n5906 VGND.n5904 8.23546
R1483 VGND.n5906 VGND.n5905 8.23546
R1484 VGND.n5914 VGND.n1319 8.23546
R1485 VGND.n5915 VGND.n5914 8.23546
R1486 VGND.n5918 VGND.n5917 8.23546
R1487 VGND.n5921 VGND.n1318 8.23546
R1488 VGND.n6378 VGND.n6346 8.23546
R1489 VGND.n5036 VGND.n5035 8.23409
R1490 VGND.n7942 VGND.n7941 8.0482
R1491 VGND.n3265 VGND.n3264 7.90638
R1492 VGND.n4162 VGND.n4161 7.90638
R1493 VGND.n2772 VGND.n2771 7.90638
R1494 VGND.n4729 VGND.n4716 7.77299
R1495 VGND.n496 VGND.n451 7.65637
R1496 VGND.n144 VGND.n143 7.60889
R1497 VGND.n6077 VGND.n6042 7.56414
R1498 VGND.n3990 VGND.n3628 7.56414
R1499 VGND.n1283 VGND.n1255 7.56414
R1500 VGND.n5791 VGND.n5790 7.52991
R1501 VGND.n6357 VGND.n6356 7.47675
R1502 VGND.n6072 VGND.n6045 7.42364
R1503 VGND.n5134 VGND.n5133 7.34036
R1504 VGND.n2086 VGND.n2085 7.23528
R1505 VGND VGND.n4580 7.15344
R1506 VGND VGND.n3061 7.15344
R1507 VGND.n2799 VGND 7.15344
R1508 VGND.n680 VGND.n679 7.15139
R1509 VGND.n2649 VGND.n2626 7.15139
R1510 VGND.n343 VGND.n299 7.11268
R1511 VGND.n6641 VGND.n6639 7.11268
R1512 VGND.n6054 VGND.n6053 7.11268
R1513 VGND.n779 VGND.n776 7.11268
R1514 VGND.n3860 VGND.n3652 7.11268
R1515 VGND.n6374 VGND.n6373 7.11268
R1516 VGND.n7656 VGND.n108 6.90655
R1517 VGND.n7662 VGND.n7659 6.90655
R1518 VGND.n4460 VGND.n4456 6.90655
R1519 VGND VGND.n4151 6.89281
R1520 VGND.n2982 VGND.n2977 6.89281
R1521 VGND.n651 VGND.n403 6.88949
R1522 VGND.n314 VGND.n307 6.88949
R1523 VGND.n6679 VGND.n6678 6.88949
R1524 VGND.n3191 VGND.n3190 6.88949
R1525 VGND.n3844 VGND.n3656 6.88949
R1526 VGND.n4437 VGND.n4436 6.88949
R1527 VGND.n2810 VGND.n2809 6.88949
R1528 VGND.n5407 VGND.n5406 6.88949
R1529 VGND.n6045 VGND.n6044 6.85195
R1530 VGND.n6043 VGND.n6042 6.82364
R1531 VGND.n3628 VGND.n3627 6.82364
R1532 VGND.n1256 VGND.n1255 6.82364
R1533 VGND.n4558 VGND 6.77697
R1534 VGND.n4551 VGND 6.77697
R1535 VGND.n1617 VGND.n1616 6.77697
R1536 VGND.n655 VGND 6.71379
R1537 VGND.n344 VGND 6.71379
R1538 VGND.n314 VGND 6.71379
R1539 VGND.n4436 VGND 6.71379
R1540 VGND.n7989 VGND.n10 6.65013
R1541 VGND.n7388 VGND.n173 6.65013
R1542 VGND.n6219 VGND 6.62428
R1543 VGND.n6521 VGND.n1100 6.61527
R1544 VGND.n6729 VGND.n6728 6.57117
R1545 VGND.n6518 VGND.n1100 6.57117
R1546 VGND.n6518 VGND.n6517 6.57117
R1547 VGND.n3861 VGND 6.53477
R1548 VGND.n3841 VGND.n3840 6.44345
R1549 VGND.n502 VGND 6.4005
R1550 VGND.n550 VGND.n435 6.4005
R1551 VGND.n2184 VGND.n2182 6.4005
R1552 VGND.n889 VGND.n884 6.4005
R1553 VGND.n907 VGND 6.4005
R1554 VGND VGND.n7252 6.4005
R1555 VGND.n7073 VGND 6.4005
R1556 VGND VGND.n6970 6.4005
R1557 VGND.n6941 VGND 6.4005
R1558 VGND.n6839 VGND.n6837 6.4005
R1559 VGND.n6172 VGND 6.4005
R1560 VGND.n784 VGND.n180 6.4005
R1561 VGND.n4177 VGND.n4176 6.4005
R1562 VGND.n3700 VGND 6.4005
R1563 VGND.n3971 VGND.n3970 6.4005
R1564 VGND VGND.n2907 6.4005
R1565 VGND.n4268 VGND.n4267 6.4005
R1566 VGND.n5178 VGND.n5177 6.4005
R1567 VGND.n5569 VGND 6.4005
R1568 VGND.n5602 VGND.n1400 6.4005
R1569 VGND.n5612 VGND.n5611 6.4005
R1570 VGND.n5983 VGND.n5925 6.4005
R1571 VGND.n6767 VGND.n1039 6.4005
R1572 VGND.n7940 VGND 6.4005
R1573 VGND.n3484 VGND.n3483 6.4005
R1574 VGND.n4567 VGND.n2962 6.4005
R1575 VGND.n2999 VGND.n2998 6.4005
R1576 VGND.n5842 VGND.n5840 6.39431
R1577 VGND.n1257 VGND.n1256 6.38812
R1578 VGND.n6838 VGND 6.27264
R1579 VGND.n533 VGND.n440 6.26433
R1580 VGND.n2194 VGND.n2193 6.26433
R1581 VGND.n901 VGND.n881 6.26433
R1582 VGND.n7200 VGND.n7199 6.26433
R1583 VGND.n6844 VGND.n6843 6.26433
R1584 VGND.n6084 VGND.n6041 6.26433
R1585 VGND.n2091 VGND.n1977 6.26433
R1586 VGND.n3518 VGND.n3517 6.26433
R1587 VGND.n3410 VGND.n3409 6.26433
R1588 VGND.n3260 VGND.n3259 6.26433
R1589 VGND.n7752 VGND.n7751 6.26433
R1590 VGND.n4055 VGND.n4026 6.26433
R1591 VGND.n3685 VGND.n3684 6.26433
R1592 VGND.n3686 VGND.n3685 6.26433
R1593 VGND.n3821 VGND.n3820 6.26433
R1594 VGND.n3823 VGND.n3821 6.26433
R1595 VGND.n3833 VGND.n3659 6.26433
R1596 VGND.n3835 VGND.n3657 6.26433
R1597 VGND.n3839 VGND.n3657 6.26433
R1598 VGND.n2931 VGND.n2901 6.26433
R1599 VGND.n4262 VGND.n4261 6.26433
R1600 VGND.n4574 VGND.n4573 6.26433
R1601 VGND.n4409 VGND.n4408 6.26433
R1602 VGND.n3041 VGND.n3040 6.26433
R1603 VGND.n5104 VGND.n5103 6.26433
R1604 VGND.n5112 VGND.n5093 6.26433
R1605 VGND.n2794 VGND.n2764 6.26433
R1606 VGND.n2790 VGND.n2764 6.26433
R1607 VGND.n4995 VGND.n4994 6.26433
R1608 VGND.n4828 VGND.n4826 6.26433
R1609 VGND.n1537 VGND.n1485 6.26433
R1610 VGND.n1948 VGND.n1947 6.26433
R1611 VGND.n5824 VGND.n5823 6.26433
R1612 VGND.n1290 VGND.n1254 6.26433
R1613 VGND.n1931 VGND.n1924 6.26433
R1614 VGND.n529 VGND.n440 6.26433
R1615 VGND.n897 VGND.n881 6.26433
R1616 VGND.n6846 VGND.n6844 6.26433
R1617 VGND.n2080 VGND.n1979 6.26433
R1618 VGND.n3517 VGND.n3466 6.26433
R1619 VGND.n4037 VGND.n4036 6.26433
R1620 VGND.n3989 VGND.n3629 6.26433
R1621 VGND.n3686 VGND.n3680 6.26433
R1622 VGND.n3810 VGND.n3808 6.26433
R1623 VGND.n3834 VGND.n3833 6.26433
R1624 VGND.n3835 VGND.n3834 6.26433
R1625 VGND.n2931 VGND.n2930 6.26433
R1626 VGND.n4576 VGND.n4574 6.26433
R1627 VGND.n2790 VGND.n2789 6.26433
R1628 VGND.n4828 VGND.n4827 6.26433
R1629 VGND.n1533 VGND.n1532 6.26433
R1630 VGND.n2696 VGND.n2695 6.26433
R1631 VGND.n2695 VGND.n2405 6.26433
R1632 VGND.n1271 VGND.n1270 6.26433
R1633 VGND.n886 VGND.n885 6.2505
R1634 VGND.n220 VGND.n219 6.02861
R1635 VGND.n7626 VGND.n7623 6.02861
R1636 VGND.n333 VGND.n332 6.0286
R1637 VGND.n4047 VGND.n4027 6.02403
R1638 VGND.n2936 VGND.n2900 6.02403
R1639 VGND.n1580 VGND.n1579 6.02403
R1640 VGND VGND.n2579 6.02403
R1641 VGND.n321 VGND.n305 5.80542
R1642 VGND.n6627 VGND.n6626 5.80542
R1643 VGND.n198 VGND.n197 5.80542
R1644 VGND.n7675 VGND.n7674 5.80542
R1645 VGND.n2800 VGND 5.72682
R1646 VGND.n7941 VGND 5.72682
R1647 VGND.n2080 VGND.n2079 5.65809
R1648 VGND.n3302 VGND.n3301 5.65809
R1649 VGND.n7760 VGND.n7758 5.65809
R1650 VGND.n3996 VGND.n3994 5.65809
R1651 VGND.n3690 VGND.n3680 5.65809
R1652 VGND.n2789 VGND.n2788 5.65809
R1653 VGND.n2405 VGND.n2404 5.65809
R1654 VGND.n551 VGND 5.64756
R1655 VGND.n2190 VGND 5.64756
R1656 VGND.n890 VGND 5.64756
R1657 VGND.n6852 VGND 5.64756
R1658 VGND.n3422 VGND 5.64756
R1659 VGND.n5100 VGND 5.64756
R1660 VGND VGND.n5186 5.64756
R1661 VGND.n1874 VGND 5.64756
R1662 VGND.n2613 VGND.n2425 5.64169
R1663 VGND.n1532 VGND.n1487 5.62903
R1664 VGND.n7954 VGND.n20 5.62903
R1665 VGND.n7643 VGND.n7642 5.5878
R1666 VGND.n6512 VGND.n1042 5.53969
R1667 VGND.n765 VGND.n761 5.48128
R1668 VGND.n5001 VGND.n5000 5.35702
R1669 VGND.n2499 VGND.n2498 5.27109
R1670 VGND.n7758 VGND 5.24305
R1671 VGND.n1102 VGND.n1101 5.13241
R1672 VGND.n6616 VGND.n1066 5.12314
R1673 VGND.n4037 VGND 5.10688
R1674 VGND.n3808 VGND 5.10688
R1675 VGND.n5965 VGND 5.0388
R1676 VGND.n2781 VGND.n2770 5.03644
R1677 VGND.n3936 VGND.n3928 4.93346
R1678 VGND.n4136 VGND.n3146 4.89462
R1679 VGND.n7948 VGND.n7947 4.85762
R1680 VGND.n636 VGND.n635 4.85762
R1681 VGND.n973 VGND.n972 4.85762
R1682 VGND.n7177 VGND.n7176 4.85762
R1683 VGND.n7211 VGND.n7210 4.85762
R1684 VGND.n1982 VGND.n1981 4.85762
R1685 VGND.n3506 VGND.n3505 4.85762
R1686 VGND.n3346 VGND.n3345 4.85762
R1687 VGND.n803 VGND.n802 4.85762
R1688 VGND.n757 VGND.n756 4.85762
R1689 VGND.n3296 VGND.n3295 4.85762
R1690 VGND.n75 VGND.n74 4.85762
R1691 VGND.n3623 VGND.n3622 4.85762
R1692 VGND.n4070 VGND.n4069 4.85762
R1693 VGND.n3693 VGND.n3692 4.85762
R1694 VGND.n3932 VGND.n3931 4.85762
R1695 VGND.n3975 VGND.n3974 4.85762
R1696 VGND.n3052 VGND.n3051 4.85762
R1697 VGND.n3015 VGND.n3014 4.85762
R1698 VGND.n4420 VGND.n4419 4.85762
R1699 VGND.n2783 VGND.n2769 4.85762
R1700 VGND.n4898 VGND.n4897 4.85762
R1701 VGND.n2688 VGND.n2687 4.85762
R1702 VGND.n1526 VGND.n1525 4.85762
R1703 VGND.n2617 VGND.n2616 4.85762
R1704 VGND.n5937 VGND.n5936 4.85762
R1705 VGND.n5930 VGND.n5929 4.85762
R1706 VGND.n494 VGND.n493 4.8005
R1707 VGND.n436 VGND.n435 4.8005
R1708 VGND.n2184 VGND.n2183 4.8005
R1709 VGND.n885 VGND.n884 4.8005
R1710 VGND.n7256 VGND.n7255 4.8005
R1711 VGND.n6839 VGND.n6838 4.8005
R1712 VGND.n1990 VGND.n1989 4.8005
R1713 VGND.n1123 VGND.n1122 4.8005
R1714 VGND.n126 VGND.n125 4.8005
R1715 VGND.n7564 VGND.n7563 4.8005
R1716 VGND.n4177 VGND.n4160 4.8005
R1717 VGND.n3632 VGND.n3631 4.8005
R1718 VGND.n4269 VGND.n4268 4.8005
R1719 VGND.n4568 VGND.n4567 4.8005
R1720 VGND.n2998 VGND.n2975 4.8005
R1721 VGND.n5178 VGND.n5173 4.8005
R1722 VGND.n1456 VGND.n1455 4.8005
R1723 VGND.n5611 VGND.n1398 4.8005
R1724 VGND.n1373 VGND.n1372 4.8005
R1725 VGND.n5842 VGND.n5841 4.8005
R1726 VGND.n5926 VGND.n5925 4.8005
R1727 VGND.n1179 VGND.n1178 4.8005
R1728 VGND.n3019 VGND.n3012 4.76901
R1729 VGND.n4402 VGND.n4401 4.72253
R1730 VGND.n400 VGND.n399 4.67352
R1731 VGND.n338 VGND.n337 4.67352
R1732 VGND.n339 VGND.n338 4.67352
R1733 VGND.n328 VGND.n327 4.67352
R1734 VGND.n328 VGND.n303 4.67352
R1735 VGND.n7988 VGND.n7987 4.67352
R1736 VGND.n1061 VGND.n1060 4.67352
R1737 VGND.n6071 VGND.n6070 4.67352
R1738 VGND.n186 VGND.n185 4.67352
R1739 VGND.n184 VGND.n183 4.67352
R1740 VGND.n764 VGND.n763 4.67352
R1741 VGND.n175 VGND.n174 4.67352
R1742 VGND.n7617 VGND.n7616 4.67352
R1743 VGND.n7625 VGND.n7624 4.67352
R1744 VGND.n3856 VGND.n3855 4.67352
R1745 VGND.n6348 VGND.n6347 4.67352
R1746 VGND.n679 VGND.n400 4.67352
R1747 VGND.n334 VGND.n333 4.67352
R1748 VGND.n339 VGND.n299 4.67352
R1749 VGND.n325 VGND.n305 4.67352
R1750 VGND.n332 VGND.n303 4.67352
R1751 VGND.n7989 VGND.n7988 4.67352
R1752 VGND.n6639 VGND.n1061 4.67352
R1753 VGND.n6072 VGND.n6071 4.67352
R1754 VGND.n212 VGND.n186 4.67352
R1755 VGND.n219 VGND.n184 4.67352
R1756 VGND.n765 VGND.n764 4.67352
R1757 VGND.n7375 VGND.n175 4.67352
R1758 VGND.n7618 VGND.n7617 4.67352
R1759 VGND.n7626 VGND.n7625 4.67352
R1760 VGND.n3855 VGND.n3854 4.67352
R1761 VGND.n3856 VGND.n3652 4.67352
R1762 VGND.n643 VGND.n642 4.65776
R1763 VGND.n5036 VGND.n5034 4.65281
R1764 VGND.n3441 VGND.n3440 4.65209
R1765 VGND.n2613 VGND.n2612 4.65207
R1766 VGND.n4428 VGND.n4427 4.65146
R1767 VGND.n787 VGND.n786 4.6505
R1768 VGND.n789 VGND.n788 4.6505
R1769 VGND.n847 VGND.n799 4.6505
R1770 VGND.n830 VGND.n829 4.6505
R1771 VGND.n828 VGND.n807 4.6505
R1772 VGND.n193 VGND.n192 4.6505
R1773 VGND.n197 VGND.n196 4.6505
R1774 VGND.n199 VGND.n198 4.6505
R1775 VGND.n201 VGND.n200 4.6505
R1776 VGND.n203 VGND.n202 4.6505
R1777 VGND.n205 VGND.n204 4.6505
R1778 VGND.n208 VGND.n207 4.6505
R1779 VGND.n212 VGND.n211 4.6505
R1780 VGND.n215 VGND.n214 4.6505
R1781 VGND.n219 VGND.n218 4.6505
R1782 VGND.n221 VGND.n220 4.6505
R1783 VGND.n223 VGND.n222 4.6505
R1784 VGND.n225 VGND.n224 4.6505
R1785 VGND.n227 VGND.n226 4.6505
R1786 VGND.n230 VGND.n229 4.6505
R1787 VGND.n745 VGND.n744 4.6505
R1788 VGND.n753 VGND.n752 4.6505
R1789 VGND.n766 VGND.n765 4.6505
R1790 VGND.n770 VGND.n769 4.6505
R1791 VGND.n772 VGND.n771 4.6505
R1792 VGND.n774 VGND.n773 4.6505
R1793 VGND.n776 VGND.n775 4.6505
R1794 VGND.n780 VGND.n779 4.6505
R1795 VGND.n783 VGND.n782 4.6505
R1796 VGND.n3378 VGND.n3349 4.6505
R1797 VGND.n3384 VGND.n3383 4.6505
R1798 VGND.n3385 VGND.n3348 4.6505
R1799 VGND.n3404 VGND.n3403 4.6505
R1800 VGND.n3408 VGND.n3407 4.6505
R1801 VGND.n3434 VGND.n3433 4.6505
R1802 VGND.n3436 VGND.n3435 4.6505
R1803 VGND.n3439 VGND.n3342 4.6505
R1804 VGND.n3520 VGND.n3465 4.6505
R1805 VGND.n3499 VGND.n3498 4.6505
R1806 VGND.n3489 VGND.n3467 4.6505
R1807 VGND.n3486 VGND.n3468 4.6505
R1808 VGND.n3479 VGND.n3478 4.6505
R1809 VGND.n3477 VGND.n3470 4.6505
R1810 VGND.n3474 VGND.n3471 4.6505
R1811 VGND.n3519 VGND.n3518 4.6505
R1812 VGND.n3517 VGND.n3516 4.6505
R1813 VGND.n3514 VGND.n3513 4.6505
R1814 VGND.n3512 VGND.n3511 4.6505
R1815 VGND.n3509 VGND.n3508 4.6505
R1816 VGND.n3504 VGND.n3503 4.6505
R1817 VGND.n3501 VGND.n3500 4.6505
R1818 VGND.n3497 VGND.n3496 4.6505
R1819 VGND.n3495 VGND.n3494 4.6505
R1820 VGND.n3493 VGND.n3492 4.6505
R1821 VGND.n3491 VGND.n3490 4.6505
R1822 VGND.n3488 VGND.n3487 4.6505
R1823 VGND.n3485 VGND.n3484 4.6505
R1824 VGND.n3481 VGND.n3480 4.6505
R1825 VGND.n3476 VGND.n3475 4.6505
R1826 VGND.n3537 VGND.n3536 4.6505
R1827 VGND.n3375 VGND.n3374 4.6505
R1828 VGND.n3377 VGND.n3376 4.6505
R1829 VGND.n3380 VGND.n3379 4.6505
R1830 VGND.n3382 VGND.n3381 4.6505
R1831 VGND.n3389 VGND.n3388 4.6505
R1832 VGND.n3393 VGND.n3392 4.6505
R1833 VGND.n3396 VGND.n3395 4.6505
R1834 VGND.n3397 VGND.n848 4.6505
R1835 VGND.n3400 VGND.n3399 4.6505
R1836 VGND.n3406 VGND.n3405 4.6505
R1837 VGND.n3411 VGND.n3410 4.6505
R1838 VGND.n3415 VGND.n3414 4.6505
R1839 VGND.n3417 VGND.n3416 4.6505
R1840 VGND.n3419 VGND.n3418 4.6505
R1841 VGND.n3421 VGND.n3420 4.6505
R1842 VGND.n3423 VGND.n3422 4.6505
R1843 VGND.n3425 VGND.n3424 4.6505
R1844 VGND.n3427 VGND.n3426 4.6505
R1845 VGND.n3429 VGND.n3428 4.6505
R1846 VGND.n3432 VGND.n3431 4.6505
R1847 VGND.n3438 VGND.n3437 4.6505
R1848 VGND.n3443 VGND.n3442 4.6505
R1849 VGND.n3445 VGND.n3444 4.6505
R1850 VGND.n832 VGND.n831 4.6505
R1851 VGND.n837 VGND.n836 4.6505
R1852 VGND.n839 VGND.n838 4.6505
R1853 VGND.n841 VGND.n840 4.6505
R1854 VGND.n843 VGND.n842 4.6505
R1855 VGND.n844 VGND.n800 4.6505
R1856 VGND.n846 VGND.n845 4.6505
R1857 VGND.n798 VGND.n179 4.6505
R1858 VGND.n797 VGND.n796 4.6505
R1859 VGND.n795 VGND.n794 4.6505
R1860 VGND.n793 VGND.n792 4.6505
R1861 VGND.n791 VGND.n790 4.6505
R1862 VGND.n130 VGND.n129 4.6505
R1863 VGND.n133 VGND.n132 4.6505
R1864 VGND.n135 VGND.n134 4.6505
R1865 VGND.n138 VGND.n137 4.6505
R1866 VGND.n140 VGND.n139 4.6505
R1867 VGND.n143 VGND.n142 4.6505
R1868 VGND.n7394 VGND.n7393 4.6505
R1869 VGND.n7392 VGND.n7391 4.6505
R1870 VGND.n7389 VGND.n7388 4.6505
R1871 VGND.n7387 VGND.n7386 4.6505
R1872 VGND.n7385 VGND.n7384 4.6505
R1873 VGND.n7383 VGND.n7382 4.6505
R1874 VGND.n7381 VGND.n7380 4.6505
R1875 VGND.n7376 VGND.n7375 4.6505
R1876 VGND.n7373 VGND.n176 4.6505
R1877 VGND.n189 VGND.n177 4.6505
R1878 VGND.n7787 VGND.n7786 4.6505
R1879 VGND.n7789 VGND.n7788 4.6505
R1880 VGND.n7791 VGND.n7790 4.6505
R1881 VGND.n7794 VGND.n7793 4.6505
R1882 VGND.n7573 VGND.n7572 4.6505
R1883 VGND.n7575 VGND.n7574 4.6505
R1884 VGND.n7647 VGND.n7646 4.6505
R1885 VGND.n7650 VGND.n7649 4.6505
R1886 VGND.n7652 VGND.n108 4.6505
R1887 VGND.n7656 VGND.n7655 4.6505
R1888 VGND.n7663 VGND.n7662 4.6505
R1889 VGND.n7666 VGND.n7665 4.6505
R1890 VGND.n7670 VGND.n7669 4.6505
R1891 VGND.n7674 VGND.n7673 4.6505
R1892 VGND.n7676 VGND.n7675 4.6505
R1893 VGND.n7678 VGND.n7677 4.6505
R1894 VGND.n7680 VGND.n7679 4.6505
R1895 VGND.n7682 VGND.n7681 4.6505
R1896 VGND.n7685 VGND.n7684 4.6505
R1897 VGND.n7753 VGND.n7752 4.6505
R1898 VGND.n7756 VGND.n7755 4.6505
R1899 VGND.n7758 VGND.n7757 4.6505
R1900 VGND.n7761 VGND.n7760 4.6505
R1901 VGND.n7765 VGND.n7764 4.6505
R1902 VGND.n7778 VGND.n7777 4.6505
R1903 VGND.n7780 VGND.n7779 4.6505
R1904 VGND.n7782 VGND.n7781 4.6505
R1905 VGND.n3180 VGND.n3173 4.6505
R1906 VGND.n3183 VGND.n3172 4.6505
R1907 VGND.n3185 VGND.n3184 4.6505
R1908 VGND.n3291 VGND.n3290 4.6505
R1909 VGND.n3272 VGND.n3263 4.6505
R1910 VGND.n3271 VGND.n3264 4.6505
R1911 VGND.n3270 VGND.n3265 4.6505
R1912 VGND.n3269 VGND.n3266 4.6505
R1913 VGND.n3307 VGND.n3306 4.6505
R1914 VGND.n3305 VGND.n3304 4.6505
R1915 VGND.n3303 VGND.n3302 4.6505
R1916 VGND.n3301 VGND.n3300 4.6505
R1917 VGND.n3299 VGND.n3298 4.6505
R1918 VGND.n3289 VGND.n3288 4.6505
R1919 VGND.n3287 VGND.n3286 4.6505
R1920 VGND.n3285 VGND.n3284 4.6505
R1921 VGND.n3283 VGND.n3282 4.6505
R1922 VGND.n3281 VGND.n3280 4.6505
R1923 VGND.n3279 VGND.n3278 4.6505
R1924 VGND.n3277 VGND.n3260 4.6505
R1925 VGND.n3275 VGND.n3274 4.6505
R1926 VGND.n3324 VGND.n3323 4.6505
R1927 VGND.n3179 VGND.n3178 4.6505
R1928 VGND.n3182 VGND.n3181 4.6505
R1929 VGND.n3187 VGND.n3186 4.6505
R1930 VGND.n3190 VGND.n3189 4.6505
R1931 VGND.n3192 VGND.n3191 4.6505
R1932 VGND.n3199 VGND.n3198 4.6505
R1933 VGND.n3252 VGND.n3251 4.6505
R1934 VGND.n3250 VGND.n3170 4.6505
R1935 VGND.n3248 VGND.n3247 4.6505
R1936 VGND.n3246 VGND.n3245 4.6505
R1937 VGND.n3244 VGND.n3243 4.6505
R1938 VGND.n3241 VGND.n3240 4.6505
R1939 VGND.n3239 VGND.n3238 4.6505
R1940 VGND.n3237 VGND.n3236 4.6505
R1941 VGND.n3235 VGND.n3234 4.6505
R1942 VGND.n3233 VGND.n3232 4.6505
R1943 VGND.n3231 VGND.n3230 4.6505
R1944 VGND.n3228 VGND.n3227 4.6505
R1945 VGND.n3225 VGND.n3224 4.6505
R1946 VGND.n3223 VGND.n3222 4.6505
R1947 VGND.n3221 VGND.n3220 4.6505
R1948 VGND.n3219 VGND.n3218 4.6505
R1949 VGND.n3217 VGND.n3216 4.6505
R1950 VGND.n3215 VGND.n3214 4.6505
R1951 VGND.n3213 VGND.n3212 4.6505
R1952 VGND.n3211 VGND.n3210 4.6505
R1953 VGND.n3209 VGND.n3208 4.6505
R1954 VGND.n3207 VGND.n3206 4.6505
R1955 VGND.n3204 VGND.n3203 4.6505
R1956 VGND.n3162 VGND.n3161 4.6505
R1957 VGND.n7817 VGND.n7816 4.6505
R1958 VGND.n7815 VGND.n7814 4.6505
R1959 VGND.n7813 VGND.n7812 4.6505
R1960 VGND.n7810 VGND.n7809 4.6505
R1961 VGND.n7808 VGND.n7807 4.6505
R1962 VGND.n7806 VGND.n7805 4.6505
R1963 VGND.n7804 VGND.n7803 4.6505
R1964 VGND.n7802 VGND.n7801 4.6505
R1965 VGND.n7800 VGND.n7799 4.6505
R1966 VGND.n7798 VGND.n7797 4.6505
R1967 VGND.n7796 VGND.n7795 4.6505
R1968 VGND.n7792 VGND.n70 4.6505
R1969 VGND.n7776 VGND.n7775 4.6505
R1970 VGND.n7774 VGND.n72 4.6505
R1971 VGND.n7773 VGND.n7772 4.6505
R1972 VGND.n7771 VGND.n7770 4.6505
R1973 VGND.n7769 VGND.n7768 4.6505
R1974 VGND.n7767 VGND.n7766 4.6505
R1975 VGND.n7568 VGND.n7567 4.6505
R1976 VGND.n7571 VGND.n7570 4.6505
R1977 VGND.n7576 VGND.n7562 4.6505
R1978 VGND.n7578 VGND.n7577 4.6505
R1979 VGND.n7580 VGND.n7579 4.6505
R1980 VGND.n7583 VGND.n7582 4.6505
R1981 VGND.n7619 VGND.n7618 4.6505
R1982 VGND.n7623 VGND.n7622 4.6505
R1983 VGND.n7627 VGND.n7626 4.6505
R1984 VGND.n7632 VGND.n7631 4.6505
R1985 VGND.n7634 VGND.n7633 4.6505
R1986 VGND.n7636 VGND.n7635 4.6505
R1987 VGND.n7638 VGND.n7637 4.6505
R1988 VGND.n7640 VGND.n7639 4.6505
R1989 VGND.n7644 VGND.n7643 4.6505
R1990 VGND.n3804 VGND.n3803 4.6505
R1991 VGND.n3814 VGND.n3813 4.6505
R1992 VGND.n3817 VGND.n3816 4.6505
R1993 VGND.n3827 VGND.n3826 4.6505
R1994 VGND.n3830 VGND.n3829 4.6505
R1995 VGND.n4159 VGND.n3139 4.6505
R1996 VGND.n3682 VGND.n3146 4.6505
R1997 VGND.n3699 VGND.n3676 4.6505
R1998 VGND.n3703 VGND.n3702 4.6505
R1999 VGND.n3726 VGND.n3725 4.6505
R2000 VGND.n4166 VGND.n4163 4.6505
R2001 VGND.n4168 VGND.n4167 4.6505
R2002 VGND.n4170 VGND.n4169 4.6505
R2003 VGND.n4174 VGND.n4162 4.6505
R2004 VGND.n4143 VGND.n4142 4.6505
R2005 VGND.n3685 VGND.n3681 4.6505
R2006 VGND.n3696 VGND.n3695 4.6505
R2007 VGND.n3709 VGND.n3708 4.6505
R2008 VGND.n3719 VGND.n3718 4.6505
R2009 VGND.n3806 VGND.n3805 4.6505
R2010 VGND.n3808 VGND.n3807 4.6505
R2011 VGND.n3811 VGND.n3810 4.6505
R2012 VGND.n3820 VGND.n3819 4.6505
R2013 VGND.n3821 VGND.n3662 4.6505
R2014 VGND.n3824 VGND.n3823 4.6505
R2015 VGND.n3825 VGND.n3661 4.6505
R2016 VGND.n3831 VGND.n3659 4.6505
R2017 VGND.n3833 VGND.n3832 4.6505
R2018 VGND.n3834 VGND.n3658 4.6505
R2019 VGND.n3836 VGND.n3835 4.6505
R2020 VGND.n3837 VGND.n3657 4.6505
R2021 VGND.n3839 VGND.n3838 4.6505
R2022 VGND.n3843 VGND.n3149 4.6505
R2023 VGND.n3845 VGND.n3844 4.6505
R2024 VGND.n3846 VGND.n3656 4.6505
R2025 VGND.n3848 VGND.n3847 4.6505
R2026 VGND.n3849 VGND.n3655 4.6505
R2027 VGND.n3852 VGND.n3851 4.6505
R2028 VGND.n3854 VGND.n3853 4.6505
R2029 VGND.n3855 VGND.n3653 4.6505
R2030 VGND.n3857 VGND.n3856 4.6505
R2031 VGND.n3858 VGND.n3652 4.6505
R2032 VGND.n3862 VGND.n3861 4.6505
R2033 VGND.n3948 VGND.n3947 4.6505
R2034 VGND.n3984 VGND.n3983 4.6505
R2035 VGND.n4003 VGND.n4002 4.6505
R2036 VGND.n4063 VGND.n4062 4.6505
R2037 VGND.n4047 VGND.n4046 4.6505
R2038 VGND.n4045 VGND.n4027 4.6505
R2039 VGND.n4044 VGND.n4028 4.6505
R2040 VGND.n4043 VGND.n4029 4.6505
R2041 VGND.n4082 VGND.n4081 4.6505
R2042 VGND.n4080 VGND.n4079 4.6505
R2043 VGND.n4078 VGND.n4077 4.6505
R2044 VGND.n4076 VGND.n4075 4.6505
R2045 VGND.n4073 VGND.n4072 4.6505
R2046 VGND.n4068 VGND.n4067 4.6505
R2047 VGND.n4065 VGND.n4064 4.6505
R2048 VGND.n4061 VGND.n4060 4.6505
R2049 VGND.n4059 VGND.n4058 4.6505
R2050 VGND.n4057 VGND.n4056 4.6505
R2051 VGND.n4055 VGND.n4054 4.6505
R2052 VGND.n4052 VGND.n4051 4.6505
R2053 VGND.n4049 VGND.n4048 4.6505
R2054 VGND.n4042 VGND.n4041 4.6505
R2055 VGND.n4040 VGND.n4039 4.6505
R2056 VGND.n4038 VGND.n4037 4.6505
R2057 VGND.n4036 VGND.n4030 4.6505
R2058 VGND.n4034 VGND.n4033 4.6505
R2059 VGND.n4024 VGND.n4023 4.6505
R2060 VGND.n3926 VGND.n3925 4.6505
R2061 VGND.n3928 VGND.n3927 4.6505
R2062 VGND.n3937 VGND.n3936 4.6505
R2063 VGND.n3940 VGND.n3633 4.6505
R2064 VGND.n3942 VGND.n3941 4.6505
R2065 VGND.n3944 VGND.n3943 4.6505
R2066 VGND.n3946 VGND.n3945 4.6505
R2067 VGND.n3950 VGND.n3949 4.6505
R2068 VGND.n3952 VGND.n3951 4.6505
R2069 VGND.n3953 VGND.n3150 4.6505
R2070 VGND.n3955 VGND.n3954 4.6505
R2071 VGND.n3958 VGND.n3957 4.6505
R2072 VGND.n3960 VGND.n3959 4.6505
R2073 VGND.n3962 VGND.n3961 4.6505
R2074 VGND.n3964 VGND.n3963 4.6505
R2075 VGND.n3966 VGND.n3965 4.6505
R2076 VGND.n3978 VGND.n3977 4.6505
R2077 VGND.n3980 VGND.n3630 4.6505
R2078 VGND.n3982 VGND.n3981 4.6505
R2079 VGND.n3986 VGND.n3985 4.6505
R2080 VGND.n3989 VGND.n3988 4.6505
R2081 VGND.n3994 VGND.n3993 4.6505
R2082 VGND.n3997 VGND.n3996 4.6505
R2083 VGND.n4001 VGND.n4000 4.6505
R2084 VGND.n3860 VGND.n3859 4.6505
R2085 VGND.n3828 VGND.n3660 4.6505
R2086 VGND.n3818 VGND.n3663 4.6505
R2087 VGND.n3815 VGND.n3664 4.6505
R2088 VGND VGND.n3665 4.6505
R2089 VGND.n3724 VGND.n3723 4.6505
R2090 VGND.n3722 VGND.n3675 4.6505
R2091 VGND.n3721 VGND.n3720 4.6505
R2092 VGND.n3717 VGND.n3716 4.6505
R2093 VGND.n3715 VGND.n3714 4.6505
R2094 VGND.n3713 VGND.n3712 4.6505
R2095 VGND.n3711 VGND.n3710 4.6505
R2096 VGND.n3707 VGND.n3706 4.6505
R2097 VGND.n3705 VGND.n3704 4.6505
R2098 VGND.n3701 VGND.n3700 4.6505
R2099 VGND.n3698 VGND.n3697 4.6505
R2100 VGND.n3679 VGND.n3678 4.6505
R2101 VGND.n3690 VGND.n3689 4.6505
R2102 VGND.n3688 VGND.n3680 4.6505
R2103 VGND.n3687 VGND.n3686 4.6505
R2104 VGND.n3684 VGND.n3683 4.6505
R2105 VGND.n4138 VGND.n3145 4.6505
R2106 VGND.n4140 VGND.n4139 4.6505
R2107 VGND.n4141 VGND.n3144 4.6505
R2108 VGND.n4145 VGND.n4144 4.6505
R2109 VGND.n4146 VGND.n3142 4.6505
R2110 VGND.n4148 VGND.n4147 4.6505
R2111 VGND.n4149 VGND.n3141 4.6505
R2112 VGND.n4151 VGND.n4150 4.6505
R2113 VGND.n4153 VGND.n4152 4.6505
R2114 VGND.n4156 VGND.n4155 4.6505
R2115 VGND.n4158 VGND.n4157 4.6505
R2116 VGND.n4172 VGND.n4171 4.6505
R2117 VGND.n4176 VGND.n4175 4.6505
R2118 VGND.n4178 VGND.n4177 4.6505
R2119 VGND.n4180 VGND.n4179 4.6505
R2120 VGND.n4137 VGND.n4136 4.6505
R2121 VGND.n2995 VGND.n2994 4.6505
R2122 VGND.n3026 VGND.n3025 4.6505
R2123 VGND.n3039 VGND.n2897 4.6505
R2124 VGND.n4383 VGND.n4250 4.6505
R2125 VGND.n4387 VGND.n4386 4.6505
R2126 VGND.n4392 VGND.n4391 4.6505
R2127 VGND.n4400 VGND.n4399 4.6505
R2128 VGND.n4413 VGND.n4412 4.6505
R2129 VGND.n4438 VGND.n4437 4.6505
R2130 VGND.n4440 VGND.n4439 4.6505
R2131 VGND.n4442 VGND.n4441 4.6505
R2132 VGND.n4444 VGND.n4443 4.6505
R2133 VGND.n4447 VGND.n4446 4.6505
R2134 VGND.n4451 VGND.n4450 4.6505
R2135 VGND.n4456 VGND.n4455 4.6505
R2136 VGND.n2987 VGND.n2986 4.6505
R2137 VGND.n2991 VGND.n2976 4.6505
R2138 VGND.n3008 VGND.n3007 4.6505
R2139 VGND.n3012 VGND.n3011 4.6505
R2140 VGND.n3063 VGND.n3062 4.6505
R2141 VGND.n4556 VGND.n2965 4.6505
R2142 VGND.n4557 VGND.n2964 4.6505
R2143 VGND.n4582 VGND.n4581 4.6505
R2144 VGND.n4589 VGND.n4588 4.6505
R2145 VGND.n4593 VGND.n4592 4.6505
R2146 VGND.n4599 VGND.n4598 4.6505
R2147 VGND.n4607 VGND.n4606 4.6505
R2148 VGND.n4609 VGND.n4608 4.6505
R2149 VGND.n4611 VGND.n4610 4.6505
R2150 VGND.n4615 VGND.n4614 4.6505
R2151 VGND.n4619 VGND.n4618 4.6505
R2152 VGND.n2938 VGND.n2900 4.6505
R2153 VGND.n2926 VGND.n2903 4.6505
R2154 VGND.n2923 VGND.n2904 4.6505
R2155 VGND.n2922 VGND.n2905 4.6505
R2156 VGND.n2921 VGND.n2906 4.6505
R2157 VGND.n2918 VGND.n2917 4.6505
R2158 VGND.n2946 VGND.n2945 4.6505
R2159 VGND.n2944 VGND.n2943 4.6505
R2160 VGND.n2942 VGND.n2941 4.6505
R2161 VGND.n2940 VGND.n2939 4.6505
R2162 VGND.n2937 VGND.n2936 4.6505
R2163 VGND.n2935 VGND.n2934 4.6505
R2164 VGND.n2933 VGND.n2901 4.6505
R2165 VGND.n2932 VGND.n2931 4.6505
R2166 VGND.n2925 VGND.n2924 4.6505
R2167 VGND.n2920 VGND.n2919 4.6505
R2168 VGND.n2916 VGND.n2907 4.6505
R2169 VGND.n2915 VGND.n2914 4.6505
R2170 VGND.n2913 VGND.n2908 4.6505
R2171 VGND.n2912 VGND.n2911 4.6505
R2172 VGND.n4553 VGND.n2966 4.6505
R2173 VGND.n4555 VGND.n4554 4.6505
R2174 VGND.n4559 VGND.n4558 4.6505
R2175 VGND.n4561 VGND.n4560 4.6505
R2176 VGND.n4562 VGND.n2963 4.6505
R2177 VGND.n4564 VGND.n4563 4.6505
R2178 VGND.n4565 VGND.n2962 4.6505
R2179 VGND.n4567 VGND.n4566 4.6505
R2180 VGND.n4570 VGND.n4569 4.6505
R2181 VGND.n4571 VGND.n2898 4.6505
R2182 VGND.n4573 VGND.n4572 4.6505
R2183 VGND.n4574 VGND.n2961 4.6505
R2184 VGND.n4577 VGND.n4576 4.6505
R2185 VGND.n4578 VGND.n2960 4.6505
R2186 VGND.n4580 VGND.n4579 4.6505
R2187 VGND.n4583 VGND.n2959 4.6505
R2188 VGND.n4585 VGND.n4584 4.6505
R2189 VGND.n4587 VGND.n4586 4.6505
R2190 VGND.n4591 VGND.n4590 4.6505
R2191 VGND.n4595 VGND.n4594 4.6505
R2192 VGND.n4597 VGND.n4596 4.6505
R2193 VGND.n4601 VGND.n4600 4.6505
R2194 VGND.n4603 VGND.n4602 4.6505
R2195 VGND.n4605 VGND.n4604 4.6505
R2196 VGND.n4613 VGND.n4612 4.6505
R2197 VGND.n4617 VGND.n4616 4.6505
R2198 VGND.n4621 VGND.n4620 4.6505
R2199 VGND.n4552 VGND.n4551 4.6505
R2200 VGND.n3065 VGND.n3064 4.6505
R2201 VGND.n3061 VGND.n3060 4.6505
R2202 VGND.n3059 VGND.n2973 4.6505
R2203 VGND.n3058 VGND.n3057 4.6505
R2204 VGND.n3055 VGND.n3054 4.6505
R2205 VGND.n3050 VGND.n3049 4.6505
R2206 VGND.n3047 VGND.n3046 4.6505
R2207 VGND.n3045 VGND.n3044 4.6505
R2208 VGND.n3042 VGND.n3041 4.6505
R2209 VGND.n3038 VGND.n3037 4.6505
R2210 VGND.n3036 VGND.n3035 4.6505
R2211 VGND.n3034 VGND.n3033 4.6505
R2212 VGND.n3032 VGND.n3031 4.6505
R2213 VGND.n3030 VGND.n3029 4.6505
R2214 VGND.n3028 VGND.n3027 4.6505
R2215 VGND.n3024 VGND.n3023 4.6505
R2216 VGND.n3020 VGND.n3019 4.6505
R2217 VGND.n3003 VGND.n3002 4.6505
R2218 VGND.n3000 VGND.n2999 4.6505
R2219 VGND.n2997 VGND.n2996 4.6505
R2220 VGND.n2993 VGND.n2992 4.6505
R2221 VGND.n2990 VGND.n2989 4.6505
R2222 VGND.n2982 VGND.n2981 4.6505
R2223 VGND.n4453 VGND.n4452 4.6505
R2224 VGND.n4436 VGND.n4435 4.6505
R2225 VGND.n4434 VGND.n4433 4.6505
R2226 VGND.n4431 VGND.n4430 4.6505
R2227 VGND.n4426 VGND.n4425 4.6505
R2228 VGND.n4423 VGND.n4422 4.6505
R2229 VGND.n4418 VGND.n4417 4.6505
R2230 VGND.n4415 VGND.n4414 4.6505
R2231 VGND.n4410 VGND.n4409 4.6505
R2232 VGND.n4407 VGND.n4406 4.6505
R2233 VGND.n4404 VGND.n4403 4.6505
R2234 VGND.n4398 VGND.n4397 4.6505
R2235 VGND.n4396 VGND.n4395 4.6505
R2236 VGND.n4394 VGND.n4393 4.6505
R2237 VGND.n4390 VGND.n4389 4.6505
R2238 VGND.n4385 VGND.n4384 4.6505
R2239 VGND.n4261 VGND 4.6505
R2240 VGND.n4263 VGND.n4262 4.6505
R2241 VGND.n4265 VGND.n4258 4.6505
R2242 VGND.n4267 VGND.n4266 4.6505
R2243 VGND.n4271 VGND.n4270 4.6505
R2244 VGND.n4272 VGND.n4254 4.6505
R2245 VGND.n4274 VGND.n4273 4.6505
R2246 VGND.n4405 VGND.n4246 4.6505
R2247 VGND.n4991 VGND.n2737 4.6505
R2248 VGND.n5005 VGND.n5004 4.6505
R2249 VGND.n4846 VGND.n4845 4.6505
R2250 VGND.n4850 VGND.n4849 4.6505
R2251 VGND.n4854 VGND.n4853 4.6505
R2252 VGND.n4866 VGND.n4865 4.6505
R2253 VGND.n4868 VGND.n4867 4.6505
R2254 VGND.n4872 VGND.n4871 4.6505
R2255 VGND.n4876 VGND.n4875 4.6505
R2256 VGND.n4881 VGND.n4880 4.6505
R2257 VGND.n5092 VGND.n2728 4.6505
R2258 VGND.n5099 VGND.n5098 4.6505
R2259 VGND.n5091 VGND.n5090 4.6505
R2260 VGND.n5089 VGND.n5088 4.6505
R2261 VGND.n5087 VGND.n5086 4.6505
R2262 VGND.n5084 VGND.n5083 4.6505
R2263 VGND.n5081 VGND.n5080 4.6505
R2264 VGND.n5079 VGND.n5078 4.6505
R2265 VGND.n4842 VGND.n4841 4.6505
R2266 VGND.n4887 VGND.n4886 4.6505
R2267 VGND.n4889 VGND.n4888 4.6505
R2268 VGND.n4891 VGND.n4890 4.6505
R2269 VGND.n4893 VGND.n4892 4.6505
R2270 VGND.n4896 VGND.n4895 4.6505
R2271 VGND.n4901 VGND.n4900 4.6505
R2272 VGND.n4907 VGND.n4906 4.6505
R2273 VGND.n4969 VGND.n4968 4.6505
R2274 VGND.n4972 VGND.n4971 4.6505
R2275 VGND.n4974 VGND.n4973 4.6505
R2276 VGND.n4975 VGND.n2855 4.6505
R2277 VGND.n4978 VGND.n4977 4.6505
R2278 VGND.n4983 VGND.n4982 4.6505
R2279 VGND.n4986 VGND.n4985 4.6505
R2280 VGND.n4988 VGND.n4987 4.6505
R2281 VGND.n4990 VGND.n4989 4.6505
R2282 VGND.n4996 VGND.n4995 4.6505
R2283 VGND.n5013 VGND.n5012 4.6505
R2284 VGND.n5015 VGND.n5014 4.6505
R2285 VGND.n5017 VGND.n5016 4.6505
R2286 VGND.n5019 VGND.n5018 4.6505
R2287 VGND.n5021 VGND.n5020 4.6505
R2288 VGND.n5023 VGND.n5022 4.6505
R2289 VGND.n5025 VGND.n5024 4.6505
R2290 VGND.n5027 VGND.n5026 4.6505
R2291 VGND.n5030 VGND.n5029 4.6505
R2292 VGND.n5032 VGND.n5031 4.6505
R2293 VGND.n2797 VGND.n2763 4.6505
R2294 VGND.n2779 VGND.n2770 4.6505
R2295 VGND.n2778 VGND.n2771 4.6505
R2296 VGND.n2777 VGND.n2772 4.6505
R2297 VGND.n2776 VGND.n2773 4.6505
R2298 VGND.n2796 VGND.n2795 4.6505
R2299 VGND.n2794 VGND.n2793 4.6505
R2300 VGND.n2792 VGND.n2764 4.6505
R2301 VGND.n2791 VGND.n2790 4.6505
R2302 VGND.n2789 VGND.n2765 4.6505
R2303 VGND.n2788 VGND.n2787 4.6505
R2304 VGND.n2786 VGND.n2785 4.6505
R2305 VGND.n2768 VGND.n2767 4.6505
R2306 VGND.n2781 VGND.n2780 4.6505
R2307 VGND.n2759 VGND.n2758 4.6505
R2308 VGND.n2818 VGND.n2817 4.6505
R2309 VGND.n2816 VGND.n2815 4.6505
R2310 VGND.n2814 VGND.n2813 4.6505
R2311 VGND.n2811 VGND.n2810 4.6505
R2312 VGND.n2809 VGND.n2808 4.6505
R2313 VGND.n2806 VGND.n2805 4.6505
R2314 VGND.n2804 VGND.n2803 4.6505
R2315 VGND.n2802 VGND.n2801 4.6505
R2316 VGND.n2799 VGND.n2798 4.6505
R2317 VGND.n5011 VGND.n5010 4.6505
R2318 VGND.n5009 VGND.n5008 4.6505
R2319 VGND.n5007 VGND.n5006 4.6505
R2320 VGND.n5003 VGND.n5002 4.6505
R2321 VGND.n4993 VGND.n4992 4.6505
R2322 VGND.n4885 VGND.n4884 4.6505
R2323 VGND.n4883 VGND.n4882 4.6505
R2324 VGND.n4879 VGND.n4878 4.6505
R2325 VGND.n4877 VGND.n2736 4.6505
R2326 VGND.n4874 VGND.n4873 4.6505
R2327 VGND.n4870 VGND.n4869 4.6505
R2328 VGND.n4864 VGND.n4863 4.6505
R2329 VGND.n4862 VGND.n4861 4.6505
R2330 VGND.n4860 VGND.n4859 4.6505
R2331 VGND.n4858 VGND.n4857 4.6505
R2332 VGND.n4856 VGND.n4855 4.6505
R2333 VGND.n4852 VGND.n4851 4.6505
R2334 VGND.n4848 VGND.n4847 4.6505
R2335 VGND.n4844 VGND.n4843 4.6505
R2336 VGND.n4840 VGND.n4839 4.6505
R2337 VGND.n5097 VGND.n5094 4.6505
R2338 VGND.n5101 VGND.n5100 4.6505
R2339 VGND.n5103 VGND.n5102 4.6505
R2340 VGND.n5105 VGND.n5104 4.6505
R2341 VGND.n5107 VGND.n5106 4.6505
R2342 VGND.n5109 VGND.n5108 4.6505
R2343 VGND.n5112 VGND.n5111 4.6505
R2344 VGND.n4838 VGND.n4837 4.6505
R2345 VGND.n4832 VGND.n4831 4.6505
R2346 VGND.n4836 VGND.n4835 4.6505
R2347 VGND.n4834 VGND.n4833 4.6505
R2348 VGND.n4829 VGND.n4828 4.6505
R2349 VGND.n4826 VGND.n4825 4.6505
R2350 VGND.n4824 VGND.n2872 4.6505
R2351 VGND.n4756 VGND.n4755 4.6505
R2352 VGND.n4754 VGND.n4753 4.6505
R2353 VGND.n4752 VGND.n4713 4.6505
R2354 VGND.n4751 VGND.n4750 4.6505
R2355 VGND.n4749 VGND.n4748 4.6505
R2356 VGND.n4747 VGND.n4746 4.6505
R2357 VGND.n4745 VGND.n4744 4.6505
R2358 VGND.n4729 VGND.n4728 4.6505
R2359 VGND.n4731 VGND.n4730 4.6505
R2360 VGND.n4733 VGND.n4732 4.6505
R2361 VGND.n4735 VGND.n4734 4.6505
R2362 VGND.n4738 VGND.n4737 4.6505
R2363 VGND.n4740 VGND.n4739 4.6505
R2364 VGND.n4743 VGND.n4742 4.6505
R2365 VGND.n4722 VGND.n4721 4.6505
R2366 VGND.n4726 VGND.n4725 4.6505
R2367 VGND.n5077 VGND.n2731 4.6505
R2368 VGND.n5075 VGND.n5074 4.6505
R2369 VGND.n5073 VGND.n5072 4.6505
R2370 VGND.n5071 VGND.n5070 4.6505
R2371 VGND.n5069 VGND.n5068 4.6505
R2372 VGND.n5067 VGND.n2732 4.6505
R2373 VGND.n4717 VGND.n2733 4.6505
R2374 VGND.n2494 VGND.n2493 4.6505
R2375 VGND.n2498 VGND.n2497 4.6505
R2376 VGND.n2500 VGND.n2499 4.6505
R2377 VGND.n2502 VGND.n2501 4.6505
R2378 VGND.n2504 VGND.n2503 4.6505
R2379 VGND.n5184 VGND.n5172 4.6505
R2380 VGND.n5187 VGND.n5171 4.6505
R2381 VGND.n2470 VGND.n2469 4.6505
R2382 VGND.n2472 VGND.n2471 4.6505
R2383 VGND.n2474 VGND.n2473 4.6505
R2384 VGND.n2476 VGND.n2475 4.6505
R2385 VGND.n2478 VGND.n2477 4.6505
R2386 VGND.n2480 VGND.n2479 4.6505
R2387 VGND.n2482 VGND.n2481 4.6505
R2388 VGND.n2484 VGND.n2483 4.6505
R2389 VGND.n2487 VGND.n2486 4.6505
R2390 VGND.n2489 VGND.n2488 4.6505
R2391 VGND.n2492 VGND.n2491 4.6505
R2392 VGND.n5292 VGND.n5291 4.6505
R2393 VGND.n5298 VGND.n5297 4.6505
R2394 VGND.n5305 VGND.n1647 4.6505
R2395 VGND.n1643 VGND.n1576 4.6505
R2396 VGND.n1640 VGND.n1639 4.6505
R2397 VGND.n1636 VGND.n1577 4.6505
R2398 VGND.n1627 VGND.n1626 4.6505
R2399 VGND.n1616 VGND.n1615 4.6505
R2400 VGND.n1613 VGND.n1580 4.6505
R2401 VGND.n1612 VGND.n1581 4.6505
R2402 VGND.n5283 VGND.n5282 4.6505
R2403 VGND.n5285 VGND.n5284 4.6505
R2404 VGND.n5287 VGND.n5286 4.6505
R2405 VGND.n5290 VGND.n5289 4.6505
R2406 VGND.n1635 VGND.n1634 4.6505
R2407 VGND.n1631 VGND.n1630 4.6505
R2408 VGND.n1609 VGND.n1608 4.6505
R2409 VGND.n1556 VGND.n1555 4.6505
R2410 VGND.n1513 VGND.n1488 4.6505
R2411 VGND.n1502 VGND.n1492 4.6505
R2412 VGND.n1498 VGND.n1495 4.6505
R2413 VGND.n1499 VGND.n1494 4.6505
R2414 VGND.n1500 VGND.n1493 4.6505
R2415 VGND.n1504 VGND.n1503 4.6505
R2416 VGND.n1506 VGND.n1505 4.6505
R2417 VGND.n1507 VGND.n1490 4.6505
R2418 VGND.n1508 VGND.n1489 4.6505
R2419 VGND.n1510 VGND.n1509 4.6505
R2420 VGND.n1512 VGND.n1511 4.6505
R2421 VGND.n1515 VGND.n1514 4.6505
R2422 VGND.n1539 VGND.n1538 4.6505
R2423 VGND.n1537 VGND.n1536 4.6505
R2424 VGND.n1534 VGND.n1533 4.6505
R2425 VGND.n1532 VGND.n1531 4.6505
R2426 VGND.n1529 VGND.n1528 4.6505
R2427 VGND.n1524 VGND.n1523 4.6505
R2428 VGND.n1521 VGND.n1520 4.6505
R2429 VGND.n1519 VGND.n1518 4.6505
R2430 VGND.n1517 VGND.n1516 4.6505
R2431 VGND.n1603 VGND.n1602 4.6505
R2432 VGND.n1605 VGND.n1604 4.6505
R2433 VGND.n1607 VGND.n1606 4.6505
R2434 VGND.n1611 VGND.n1610 4.6505
R2435 VGND.n1618 VGND.n1617 4.6505
R2436 VGND.n1620 VGND.n1619 4.6505
R2437 VGND.n1622 VGND.n1621 4.6505
R2438 VGND.n1624 VGND.n1623 4.6505
R2439 VGND.n1625 VGND.n1578 4.6505
R2440 VGND.n1629 VGND.n1628 4.6505
R2441 VGND.n1633 VGND.n1632 4.6505
R2442 VGND.n1638 VGND.n1637 4.6505
R2443 VGND.n1642 VGND.n1641 4.6505
R2444 VGND.n1645 VGND.n1644 4.6505
R2445 VGND.n1646 VGND.n1575 4.6505
R2446 VGND.n5304 VGND.n5303 4.6505
R2447 VGND.n5302 VGND.n5301 4.6505
R2448 VGND.n5300 VGND.n5299 4.6505
R2449 VGND.n5296 VGND.n5295 4.6505
R2450 VGND.n5294 VGND.n5293 4.6505
R2451 VGND.n2573 VGND.n2572 4.6505
R2452 VGND.n2575 VGND.n2574 4.6505
R2453 VGND.n2577 VGND.n2576 4.6505
R2454 VGND.n2579 VGND.n2578 4.6505
R2455 VGND.n2581 VGND.n2580 4.6505
R2456 VGND.n2583 VGND.n2582 4.6505
R2457 VGND.n2585 VGND.n2584 4.6505
R2458 VGND.n2587 VGND.n2586 4.6505
R2459 VGND.n2589 VGND.n2588 4.6505
R2460 VGND.n2591 VGND.n2590 4.6505
R2461 VGND.n2593 VGND.n2592 4.6505
R2462 VGND.n2595 VGND.n2594 4.6505
R2463 VGND.n2597 VGND.n2596 4.6505
R2464 VGND.n2599 VGND.n2598 4.6505
R2465 VGND.n2601 VGND.n2600 4.6505
R2466 VGND.n2602 VGND.n2426 4.6505
R2467 VGND.n2604 VGND.n2603 4.6505
R2468 VGND.n2606 VGND.n2605 4.6505
R2469 VGND.n2608 VGND.n2607 4.6505
R2470 VGND.n2610 VGND.n2609 4.6505
R2471 VGND.n2621 VGND.n2620 4.6505
R2472 VGND.n2622 VGND.n2422 4.6505
R2473 VGND.n2662 VGND.n2661 4.6505
R2474 VGND.n2660 VGND.n2423 4.6505
R2475 VGND.n2659 VGND.n2658 4.6505
R2476 VGND.n2656 VGND.n2655 4.6505
R2477 VGND.n2654 VGND.n2653 4.6505
R2478 VGND.n2651 VGND.n2650 4.6505
R2479 VGND.n2649 VGND.n2648 4.6505
R2480 VGND.n2647 VGND.n2626 4.6505
R2481 VGND.n2646 VGND.n2645 4.6505
R2482 VGND.n2644 VGND.n2643 4.6505
R2483 VGND.n2569 VGND.n2568 4.6505
R2484 VGND.n2571 VGND.n2570 4.6505
R2485 VGND.n2510 VGND.n2509 4.6505
R2486 VGND.n2508 VGND.n2507 4.6505
R2487 VGND.n2506 VGND.n2505 4.6505
R2488 VGND.n2496 VGND.n2495 4.6505
R2489 VGND.n5177 VGND.n5174 4.6505
R2490 VGND.n5179 VGND.n5178 4.6505
R2491 VGND.n5181 VGND.n5180 4.6505
R2492 VGND.n5183 VGND.n5182 4.6505
R2493 VGND.n5186 VGND.n5185 4.6505
R2494 VGND.n5189 VGND.n5188 4.6505
R2495 VGND.n5191 VGND.n5190 4.6505
R2496 VGND.n2695 VGND.n2694 4.6505
R2497 VGND.n2693 VGND.n2405 4.6505
R2498 VGND.n2691 VGND.n2690 4.6505
R2499 VGND.n2686 VGND.n2685 4.6505
R2500 VGND.n2683 VGND.n2682 4.6505
R2501 VGND.n2681 VGND.n2680 4.6505
R2502 VGND.n2679 VGND.n2417 4.6505
R2503 VGND.n2677 VGND.n2676 4.6505
R2504 VGND.n2675 VGND.n2674 4.6505
R2505 VGND.n2673 VGND.n2672 4.6505
R2506 VGND.n2671 VGND.n2670 4.6505
R2507 VGND.n2669 VGND.n2668 4.6505
R2508 VGND.n2666 VGND.n2418 4.6505
R2509 VGND.n2464 VGND.n2419 4.6505
R2510 VGND.n2468 VGND.n2467 4.6505
R2511 VGND.n1858 VGND.n1750 4.6505
R2512 VGND.n1855 VGND.n1854 4.6505
R2513 VGND.n1839 VGND.n1838 4.6505
R2514 VGND.n1827 VGND.n1826 4.6505
R2515 VGND.n1824 VGND.n1753 4.6505
R2516 VGND.n1792 VGND.n1791 4.6505
R2517 VGND.n1790 VGND.n1757 4.6505
R2518 VGND.n1706 VGND.n1705 4.6505
R2519 VGND.n1710 VGND.n1709 4.6505
R2520 VGND.n1713 VGND.n1700 4.6505
R2521 VGND.n1857 VGND.n1856 4.6505
R2522 VGND.n1849 VGND.n1848 4.6505
R2523 VGND.n1789 VGND.n1788 4.6505
R2524 VGND.n1787 VGND.n1786 4.6505
R2525 VGND.n1785 VGND.n1784 4.6505
R2526 VGND.n5628 VGND.n5627 4.6505
R2527 VGND.n5622 VGND.n5621 4.6505
R2528 VGND.n5614 VGND.n1397 4.6505
R2529 VGND.n5591 VGND.n1402 4.6505
R2530 VGND.n5588 VGND.n5587 4.6505
R2531 VGND.n5585 VGND.n1404 4.6505
R2532 VGND.n5582 VGND.n5581 4.6505
R2533 VGND.n5579 VGND.n1407 4.6505
R2534 VGND.n5578 VGND.n1408 4.6505
R2535 VGND.n5577 VGND.n1409 4.6505
R2536 VGND.n5571 VGND.n1411 4.6505
R2537 VGND.n5513 VGND.n1449 4.6505
R2538 VGND.n5500 VGND.n1450 4.6505
R2539 VGND.n5499 VGND.n1451 4.6505
R2540 VGND.n5496 VGND.n1452 4.6505
R2541 VGND.n5493 VGND.n1453 4.6505
R2542 VGND.n5490 VGND.n5489 4.6505
R2543 VGND.n5486 VGND.n1454 4.6505
R2544 VGND.n5403 VGND.n5402 4.6505
R2545 VGND.n5401 VGND.n5400 4.6505
R2546 VGND.n5398 VGND.n5397 4.6505
R2547 VGND.n5396 VGND.n5395 4.6505
R2548 VGND.n5394 VGND.n5393 4.6505
R2549 VGND.n5392 VGND.n5391 4.6505
R2550 VGND.n5390 VGND.n5389 4.6505
R2551 VGND.n5387 VGND.n5386 4.6505
R2552 VGND.n5385 VGND.n5384 4.6505
R2553 VGND.n5383 VGND.n5382 4.6505
R2554 VGND.n5381 VGND.n5380 4.6505
R2555 VGND.n5379 VGND.n5378 4.6505
R2556 VGND.n5377 VGND.n5376 4.6505
R2557 VGND.n5374 VGND.n5373 4.6505
R2558 VGND.n5372 VGND.n5371 4.6505
R2559 VGND.n5370 VGND.n5369 4.6505
R2560 VGND.n5368 VGND.n5367 4.6505
R2561 VGND.n5424 VGND.n5423 4.6505
R2562 VGND.n5414 VGND.n5413 4.6505
R2563 VGND.n5412 VGND.n5411 4.6505
R2564 VGND.n5410 VGND.n5409 4.6505
R2565 VGND.n5408 VGND.n5407 4.6505
R2566 VGND.n5406 VGND.n5405 4.6505
R2567 VGND.n5522 VGND.n5521 4.6505
R2568 VGND.n5520 VGND.n1448 4.6505
R2569 VGND.n5519 VGND.n5518 4.6505
R2570 VGND.n5517 VGND.n5516 4.6505
R2571 VGND.n5515 VGND.n5514 4.6505
R2572 VGND.n5512 VGND.n5511 4.6505
R2573 VGND.n5510 VGND.n5509 4.6505
R2574 VGND.n5508 VGND.n5507 4.6505
R2575 VGND.n5506 VGND.n5505 4.6505
R2576 VGND.n5504 VGND.n5503 4.6505
R2577 VGND.n5502 VGND.n5501 4.6505
R2578 VGND.n5498 VGND.n5497 4.6505
R2579 VGND.n5495 VGND.n5494 4.6505
R2580 VGND.n5492 VGND.n5491 4.6505
R2581 VGND.n5488 VGND.n5487 4.6505
R2582 VGND.n5485 VGND.n5484 4.6505
R2583 VGND.n5482 VGND.n5481 4.6505
R2584 VGND.n5480 VGND.n5479 4.6505
R2585 VGND.n5478 VGND.n5477 4.6505
R2586 VGND.n5476 VGND.n5475 4.6505
R2587 VGND.n5474 VGND.n5473 4.6505
R2588 VGND.n5472 VGND.n1457 4.6505
R2589 VGND.n5471 VGND.n5470 4.6505
R2590 VGND.n5469 VGND.n5468 4.6505
R2591 VGND.n5467 VGND.n5466 4.6505
R2592 VGND.n5465 VGND.n5464 4.6505
R2593 VGND.n5463 VGND.n5462 4.6505
R2594 VGND.n5461 VGND.n1458 4.6505
R2595 VGND.n5460 VGND.n5459 4.6505
R2596 VGND.n5458 VGND.n5457 4.6505
R2597 VGND.n5456 VGND.n5455 4.6505
R2598 VGND.n5626 VGND.n5625 4.6505
R2599 VGND.n5624 VGND.n5623 4.6505
R2600 VGND.n5620 VGND.n5619 4.6505
R2601 VGND.n5618 VGND.n5617 4.6505
R2602 VGND.n5616 VGND.n5615 4.6505
R2603 VGND.n5613 VGND.n5612 4.6505
R2604 VGND.n5611 VGND.n5610 4.6505
R2605 VGND.n5608 VGND.n5607 4.6505
R2606 VGND.n5606 VGND.n5605 4.6505
R2607 VGND.n5604 VGND.n5603 4.6505
R2608 VGND.n5602 VGND.n5601 4.6505
R2609 VGND.n5599 VGND.n5598 4.6505
R2610 VGND.n5597 VGND.n5596 4.6505
R2611 VGND.n5595 VGND.n5594 4.6505
R2612 VGND.n5593 VGND.n5592 4.6505
R2613 VGND.n5590 VGND.n5589 4.6505
R2614 VGND.n5586 VGND.n1403 4.6505
R2615 VGND.n5584 VGND.n5583 4.6505
R2616 VGND.n5580 VGND.n1405 4.6505
R2617 VGND.n5576 VGND.n5575 4.6505
R2618 VGND.n5574 VGND.n5573 4.6505
R2619 VGND.n5572 VGND.n1410 4.6505
R2620 VGND.n5570 VGND.n5569 4.6505
R2621 VGND.n5568 VGND.n5567 4.6505
R2622 VGND.n5566 VGND.n5565 4.6505
R2623 VGND.n5630 VGND.n5629 4.6505
R2624 VGND.n1794 VGND.n1793 4.6505
R2625 VGND.n1797 VGND.n1796 4.6505
R2626 VGND.n1800 VGND.n1799 4.6505
R2627 VGND.n1802 VGND.n1801 4.6505
R2628 VGND.n1804 VGND.n1803 4.6505
R2629 VGND.n1806 VGND.n1805 4.6505
R2630 VGND.n1808 VGND.n1807 4.6505
R2631 VGND.n1810 VGND.n1809 4.6505
R2632 VGND.n1812 VGND.n1811 4.6505
R2633 VGND.n1814 VGND.n1813 4.6505
R2634 VGND.n1816 VGND.n1815 4.6505
R2635 VGND.n1818 VGND.n1817 4.6505
R2636 VGND.n1821 VGND.n1820 4.6505
R2637 VGND.n1823 VGND.n1822 4.6505
R2638 VGND.n1834 VGND.n1833 4.6505
R2639 VGND.n1836 VGND.n1835 4.6505
R2640 VGND.n1837 VGND.n1751 4.6505
R2641 VGND.n1841 VGND.n1840 4.6505
R2642 VGND.n1843 VGND.n1842 4.6505
R2643 VGND.n1845 VGND.n1844 4.6505
R2644 VGND.n1847 VGND.n1846 4.6505
R2645 VGND.n1851 VGND.n1850 4.6505
R2646 VGND.n1853 VGND.n1852 4.6505
R2647 VGND.n1704 VGND.n1701 4.6505
R2648 VGND.n1708 VGND.n1707 4.6505
R2649 VGND.n1712 VGND.n1711 4.6505
R2650 VGND.n1715 VGND.n1714 4.6505
R2651 VGND.n1717 VGND.n1716 4.6505
R2652 VGND.n1719 VGND.n1718 4.6505
R2653 VGND.n1832 VGND.n1831 4.6505
R2654 VGND.n5984 VGND.n5924 4.6505
R2655 VGND.n5953 VGND.n5934 4.6505
R2656 VGND.n5952 VGND.n5935 4.6505
R2657 VGND.n5794 VGND.n5793 4.6505
R2658 VGND.n5813 VGND.n5812 4.6505
R2659 VGND.n5817 VGND.n5816 4.6505
R2660 VGND.n5820 VGND.n1365 4.6505
R2661 VGND.n5822 VGND.n5821 4.6505
R2662 VGND.n5835 VGND.n5834 4.6505
R2663 VGND.n5837 VGND.n5836 4.6505
R2664 VGND.n5839 VGND.n5838 4.6505
R2665 VGND.n5846 VGND.n5845 4.6505
R2666 VGND.n5856 VGND.n5855 4.6505
R2667 VGND.n5857 VGND.n1359 4.6505
R2668 VGND.n1950 VGND.n1922 4.6505
R2669 VGND.n5748 VGND.n1375 4.6505
R2670 VGND.n5745 VGND.n1376 4.6505
R2671 VGND.n1873 VGND.n1872 4.6505
R2672 VGND.n1876 VGND.n1867 4.6505
R2673 VGND.n1878 VGND.n1877 4.6505
R2674 VGND.n1880 VGND.n1879 4.6505
R2675 VGND.n5754 VGND.n5753 4.6505
R2676 VGND.n5833 VGND.n5832 4.6505
R2677 VGND.n5902 VGND.n1320 4.6505
R2678 VGND.n5904 VGND.n5903 4.6505
R2679 VGND.n5907 VGND.n5906 4.6505
R2680 VGND.n5910 VGND.n5909 4.6505
R2681 VGND.n5911 VGND.n1319 4.6505
R2682 VGND.n5914 VGND.n5913 4.6505
R2683 VGND.n5919 VGND.n5918 4.6505
R2684 VGND.n5922 VGND.n5921 4.6505
R2685 VGND.n5923 VGND.n1318 4.6505
R2686 VGND.n5983 VGND.n5982 4.6505
R2687 VGND VGND.n5925 4.6505
R2688 VGND.n5981 VGND.n5980 4.6505
R2689 VGND.n5967 VGND.n5927 4.6505
R2690 VGND.n5966 VGND.n5965 4.6505
R2691 VGND.n5964 VGND.n5963 4.6505
R2692 VGND.n5962 VGND.n5961 4.6505
R2693 VGND.n5960 VGND.n5959 4.6505
R2694 VGND.n5955 VGND.n5954 4.6505
R2695 VGND.n1293 VGND.n1253 4.6505
R2696 VGND.n1279 VGND.n1259 4.6505
R2697 VGND.n1278 VGND.n1260 4.6505
R2698 VGND.n1275 VGND.n1274 4.6505
R2699 VGND.n1273 VGND.n1261 4.6505
R2700 VGND.n1310 VGND.n1309 4.6505
R2701 VGND.n1297 VGND.n1296 4.6505
R2702 VGND.n1295 VGND.n1294 4.6505
R2703 VGND.n1292 VGND.n1291 4.6505
R2704 VGND.n1290 VGND.n1289 4.6505
R2705 VGND.n1287 VGND.n1286 4.6505
R2706 VGND.n1285 VGND.n1284 4.6505
R2707 VGND.n1277 VGND.n1276 4.6505
R2708 VGND.n1272 VGND.n1271 4.6505
R2709 VGND.n1268 VGND.n1267 4.6505
R2710 VGND.n1265 VGND.n1264 4.6505
R2711 VGND.n1247 VGND.n1246 4.6505
R2712 VGND.n5940 VGND.n5939 4.6505
R2713 VGND.n5943 VGND.n5942 4.6505
R2714 VGND.n5945 VGND.n5944 4.6505
R2715 VGND.n5947 VGND.n5946 4.6505
R2716 VGND.n5949 VGND.n5948 4.6505
R2717 VGND.n5951 VGND.n5950 4.6505
R2718 VGND.n5969 VGND.n5968 4.6505
R2719 VGND.n5971 VGND.n5970 4.6505
R2720 VGND.n5973 VGND.n5972 4.6505
R2721 VGND.n5975 VGND.n5974 4.6505
R2722 VGND.n5977 VGND.n5976 4.6505
R2723 VGND.n5979 VGND.n5978 4.6505
R2724 VGND.n5859 VGND.n5858 4.6505
R2725 VGND.n5854 VGND.n5853 4.6505
R2726 VGND.n5852 VGND.n5851 4.6505
R2727 VGND.n5850 VGND.n5849 4.6505
R2728 VGND.n5848 VGND.n5847 4.6505
R2729 VGND.n5844 VGND.n1360 4.6505
R2730 VGND.n5843 VGND.n5842 4.6505
R2731 VGND VGND.n1362 4.6505
R2732 VGND.n5828 VGND.n5827 4.6505
R2733 VGND.n5825 VGND.n5824 4.6505
R2734 VGND.n5819 VGND.n5818 4.6505
R2735 VGND.n5815 VGND.n5814 4.6505
R2736 VGND.n5811 VGND.n5810 4.6505
R2737 VGND.n5809 VGND.n5808 4.6505
R2738 VGND.n5807 VGND.n5806 4.6505
R2739 VGND.n5805 VGND.n5804 4.6505
R2740 VGND.n5803 VGND.n5802 4.6505
R2741 VGND.n5801 VGND.n5800 4.6505
R2742 VGND.n5799 VGND.n5798 4.6505
R2743 VGND.n5797 VGND.n1366 4.6505
R2744 VGND.n5796 VGND.n5795 4.6505
R2745 VGND.n5792 VGND.n5791 4.6505
R2746 VGND.n5742 VGND.n5741 4.6505
R2747 VGND.n5744 VGND.n5743 4.6505
R2748 VGND.n5747 VGND.n5746 4.6505
R2749 VGND.n5750 VGND.n5749 4.6505
R2750 VGND.n5752 VGND.n5751 4.6505
R2751 VGND.n5756 VGND.n5755 4.6505
R2752 VGND.n5758 VGND.n5757 4.6505
R2753 VGND.n5761 VGND.n5760 4.6505
R2754 VGND.n5764 VGND.n5763 4.6505
R2755 VGND.n5766 VGND.n5765 4.6505
R2756 VGND.n5768 VGND.n5767 4.6505
R2757 VGND.n5770 VGND.n5769 4.6505
R2758 VGND.n5772 VGND.n5771 4.6505
R2759 VGND.n5774 VGND.n5773 4.6505
R2760 VGND.n5776 VGND.n5775 4.6505
R2761 VGND.n5778 VGND.n5777 4.6505
R2762 VGND.n5780 VGND.n5779 4.6505
R2763 VGND.n5782 VGND.n5781 4.6505
R2764 VGND.n5785 VGND.n5784 4.6505
R2765 VGND.n1940 VGND.n1939 4.6505
R2766 VGND.n1942 VGND.n1941 4.6505
R2767 VGND.n1945 VGND.n1944 4.6505
R2768 VGND.n1949 VGND.n1948 4.6505
R2769 VGND.n1871 VGND.n1868 4.6505
R2770 VGND.n1875 VGND.n1874 4.6505
R2771 VGND.n1882 VGND.n1881 4.6505
R2772 VGND.n1884 VGND.n1883 4.6505
R2773 VGND.n1886 VGND.n1885 4.6505
R2774 VGND.n1938 VGND.n1923 4.6505
R2775 VGND.n1937 VGND.n1936 4.6505
R2776 VGND.n1935 VGND.n1934 4.6505
R2777 VGND.n1933 VGND.n1932 4.6505
R2778 VGND.n1925 VGND.n1371 4.6505
R2779 VGND.n1928 VGND.n1927 4.6505
R2780 VGND.n1931 VGND.n1930 4.6505
R2781 VGND.n5787 VGND.n5786 4.6505
R2782 VGND.n1126 VGND.n1121 4.6505
R2783 VGND.n1134 VGND.n1133 4.6505
R2784 VGND.n1142 VGND.n1141 4.6505
R2785 VGND.n1150 VGND.n1149 4.6505
R2786 VGND.n1168 VGND.n1167 4.6505
R2787 VGND.n1170 VGND.n1169 4.6505
R2788 VGND.n1172 VGND.n1171 4.6505
R2789 VGND.n6285 VGND.n1177 4.6505
R2790 VGND.n2094 VGND.n1976 4.6505
R2791 VGND.n2108 VGND.n2107 4.6505
R2792 VGND.n2112 VGND.n2111 4.6505
R2793 VGND.n2116 VGND.n2115 4.6505
R2794 VGND.n2091 VGND.n2090 4.6505
R2795 VGND.n2088 VGND.n2087 4.6505
R2796 VGND.n2081 VGND.n2080 4.6505
R2797 VGND.n2040 VGND.n2039 4.6505
R2798 VGND.n2036 VGND.n2035 4.6505
R2799 VGND.n2033 VGND.n2032 4.6505
R2800 VGND.n2031 VGND.n2030 4.6505
R2801 VGND.n1130 VGND.n1129 4.6505
R2802 VGND.n1164 VGND.n1163 4.6505
R2803 VGND.n6201 VGND.n6200 4.6505
R2804 VGND.n6120 VGND.n6119 4.6505
R2805 VGND.n6086 VGND.n6085 4.6505
R2806 VGND.n6084 VGND.n6083 4.6505
R2807 VGND.n6081 VGND.n6080 4.6505
R2808 VGND.n6079 VGND.n6078 4.6505
R2809 VGND.n6073 VGND.n6072 4.6505
R2810 VGND.n6067 VGND.n6066 4.6505
R2811 VGND.n6065 VGND.n6064 4.6505
R2812 VGND.n6062 VGND.n6061 4.6505
R2813 VGND.n6060 VGND.n6059 4.6505
R2814 VGND.n6058 VGND.n6057 4.6505
R2815 VGND.n6055 VGND.n6054 4.6505
R2816 VGND.n6053 VGND.n6052 4.6505
R2817 VGND.n6050 VGND.n6049 4.6505
R2818 VGND.n6163 VGND.n6162 4.6505
R2819 VGND.n6165 VGND.n6164 4.6505
R2820 VGND.n6167 VGND.n6166 4.6505
R2821 VGND.n6169 VGND.n6168 4.6505
R2822 VGND.n6171 VGND.n6170 4.6505
R2823 VGND.n6172 VGND.n1234 4.6505
R2824 VGND.n6174 VGND.n6173 4.6505
R2825 VGND.n6175 VGND.n1233 4.6505
R2826 VGND.n6177 VGND.n6176 4.6505
R2827 VGND.n6179 VGND.n6178 4.6505
R2828 VGND.n6180 VGND.n1232 4.6505
R2829 VGND.n6199 VGND.n1226 4.6505
R2830 VGND.n6198 VGND.n6197 4.6505
R2831 VGND.n6196 VGND.n1227 4.6505
R2832 VGND.n6195 VGND.n6194 4.6505
R2833 VGND.n6193 VGND.n1228 4.6505
R2834 VGND.n6192 VGND.n6191 4.6505
R2835 VGND.n6190 VGND.n1229 4.6505
R2836 VGND.n6188 VGND.n6187 4.6505
R2837 VGND.n6186 VGND.n1230 4.6505
R2838 VGND.n6185 VGND.n6184 4.6505
R2839 VGND.n6183 VGND.n1231 4.6505
R2840 VGND.n6182 VGND.n6181 4.6505
R2841 VGND.n6202 VGND.n1225 4.6505
R2842 VGND.n6220 VGND.n6219 4.6505
R2843 VGND.n6218 VGND.n1220 4.6505
R2844 VGND.n6217 VGND.n6216 4.6505
R2845 VGND.n6215 VGND.n1221 4.6505
R2846 VGND.n6214 VGND.n6213 4.6505
R2847 VGND.n6212 VGND.n1222 4.6505
R2848 VGND.n6211 VGND.n6210 4.6505
R2849 VGND.n6209 VGND.n6208 4.6505
R2850 VGND.n6205 VGND.n1224 4.6505
R2851 VGND.n6204 VGND.n6203 4.6505
R2852 VGND.n6222 VGND.n6221 4.6505
R2853 VGND.n6265 VGND.n6264 4.6505
R2854 VGND.n6267 VGND.n6266 4.6505
R2855 VGND.n6269 VGND.n6268 4.6505
R2856 VGND.n6271 VGND.n6270 4.6505
R2857 VGND.n6273 VGND.n6272 4.6505
R2858 VGND.n6275 VGND.n6274 4.6505
R2859 VGND.n6277 VGND.n6276 4.6505
R2860 VGND.n6279 VGND.n6278 4.6505
R2861 VGND.n6281 VGND.n6280 4.6505
R2862 VGND.n6284 VGND.n6283 4.6505
R2863 VGND.n1176 VGND.n1124 4.6505
R2864 VGND.n1174 VGND.n1173 4.6505
R2865 VGND.n1166 VGND.n1165 4.6505
R2866 VGND.n1162 VGND.n1161 4.6505
R2867 VGND.n1160 VGND.n1159 4.6505
R2868 VGND.n1158 VGND.n1157 4.6505
R2869 VGND.n1156 VGND.n1155 4.6505
R2870 VGND.n1154 VGND.n1153 4.6505
R2871 VGND.n1152 VGND.n1151 4.6505
R2872 VGND.n1148 VGND.n1147 4.6505
R2873 VGND.n1146 VGND.n1145 4.6505
R2874 VGND.n1144 VGND.n1143 4.6505
R2875 VGND.n1140 VGND.n1139 4.6505
R2876 VGND.n1138 VGND.n1137 4.6505
R2877 VGND.n1136 VGND.n1135 4.6505
R2878 VGND.n1132 VGND.n1131 4.6505
R2879 VGND.n1128 VGND.n1127 4.6505
R2880 VGND.n2026 VGND.n2025 4.6505
R2881 VGND.n2028 VGND.n2027 4.6505
R2882 VGND.n2029 VGND.n1991 4.6505
R2883 VGND.n2038 VGND.n2037 4.6505
R2884 VGND.n2043 VGND.n2042 4.6505
R2885 VGND.n2046 VGND.n2045 4.6505
R2886 VGND.n2048 VGND.n2047 4.6505
R2887 VGND.n2050 VGND.n2049 4.6505
R2888 VGND.n2053 VGND.n2052 4.6505
R2889 VGND.n2055 VGND.n2054 4.6505
R2890 VGND.n2057 VGND.n2056 4.6505
R2891 VGND.n2059 VGND.n2058 4.6505
R2892 VGND.n2061 VGND.n2060 4.6505
R2893 VGND.n2063 VGND.n2062 4.6505
R2894 VGND.n2066 VGND.n2065 4.6505
R2895 VGND.n2068 VGND.n2067 4.6505
R2896 VGND.n2069 VGND.n1985 4.6505
R2897 VGND.n2071 VGND.n2070 4.6505
R2898 VGND.n2075 VGND.n2074 4.6505
R2899 VGND.n2077 VGND.n2076 4.6505
R2900 VGND.n2082 VGND.n1979 4.6505
R2901 VGND.n2093 VGND.n2092 4.6505
R2902 VGND.n2110 VGND.n2109 4.6505
R2903 VGND.n2114 VGND.n2113 4.6505
R2904 VGND.n2118 VGND.n2117 4.6505
R2905 VGND.n2120 VGND.n2119 4.6505
R2906 VGND.n2122 VGND.n2121 4.6505
R2907 VGND.n2124 VGND.n2123 4.6505
R2908 VGND.n6851 VGND.n6834 4.6505
R2909 VGND.n6857 VGND.n6856 4.6505
R2910 VGND.n6934 VGND.n1013 4.6505
R2911 VGND.n6936 VGND.n6935 4.6505
R2912 VGND.n6940 VGND.n6939 4.6505
R2913 VGND.n6965 VGND.n1004 4.6505
R2914 VGND.n6968 VGND.n1003 4.6505
R2915 VGND.n6972 VGND.n6971 4.6505
R2916 VGND.n7068 VGND.n7067 4.6505
R2917 VGND.n7072 VGND.n7071 4.6505
R2918 VGND.n7092 VGND.n970 4.6505
R2919 VGND.n7101 VGND.n7100 4.6505
R2920 VGND.n7105 VGND.n7104 4.6505
R2921 VGND.n7109 VGND.n7108 4.6505
R2922 VGND.n887 VGND.n884 4.6505
R2923 VGND.n889 VGND.n888 4.6505
R2924 VGND.n891 VGND.n890 4.6505
R2925 VGND.n892 VGND.n883 4.6505
R2926 VGND.n894 VGND.n893 4.6505
R2927 VGND.n898 VGND.n897 4.6505
R2928 VGND.n899 VGND.n881 4.6505
R2929 VGND.n901 VGND.n900 4.6505
R2930 VGND.n902 VGND.n880 4.6505
R2931 VGND.n904 VGND.n903 4.6505
R2932 VGND.n905 VGND.n879 4.6505
R2933 VGND.n907 VGND.n906 4.6505
R2934 VGND.n909 VGND.n908 4.6505
R2935 VGND.n911 VGND.n910 4.6505
R2936 VGND.n913 VGND.n912 4.6505
R2937 VGND.n915 VGND.n914 4.6505
R2938 VGND.n918 VGND.n917 4.6505
R2939 VGND.n920 VGND.n919 4.6505
R2940 VGND.n922 VGND.n921 4.6505
R2941 VGND.n924 VGND.n923 4.6505
R2942 VGND.n926 VGND.n925 4.6505
R2943 VGND.n928 VGND.n927 4.6505
R2944 VGND.n930 VGND.n929 4.6505
R2945 VGND.n7316 VGND.n7315 4.6505
R2946 VGND.n7257 VGND.n7256 4.6505
R2947 VGND.n7254 VGND.n7253 4.6505
R2948 VGND.n7252 VGND.n7251 4.6505
R2949 VGND.n7250 VGND.n7249 4.6505
R2950 VGND.n7248 VGND.n7247 4.6505
R2951 VGND.n7246 VGND.n7245 4.6505
R2952 VGND.n7244 VGND.n7243 4.6505
R2953 VGND.n7242 VGND.n7241 4.6505
R2954 VGND.n7240 VGND.n7239 4.6505
R2955 VGND.n7238 VGND.n7237 4.6505
R2956 VGND.n7236 VGND.n7235 4.6505
R2957 VGND.n7233 VGND.n7232 4.6505
R2958 VGND.n7231 VGND.n7230 4.6505
R2959 VGND.n7229 VGND.n7228 4.6505
R2960 VGND.n7227 VGND.n7226 4.6505
R2961 VGND.n7225 VGND.n7224 4.6505
R2962 VGND.n7222 VGND.n7221 4.6505
R2963 VGND.n7219 VGND.n7218 4.6505
R2964 VGND.n7217 VGND.n7216 4.6505
R2965 VGND.n7214 VGND.n7213 4.6505
R2966 VGND.n7209 VGND.n7208 4.6505
R2967 VGND.n7206 VGND.n7205 4.6505
R2968 VGND.n7204 VGND.n7203 4.6505
R2969 VGND.n7201 VGND.n7200 4.6505
R2970 VGND.n7198 VGND.n942 4.6505
R2971 VGND.n7197 VGND.n7196 4.6505
R2972 VGND.n7195 VGND.n7194 4.6505
R2973 VGND.n7193 VGND.n7192 4.6505
R2974 VGND.n7191 VGND.n7190 4.6505
R2975 VGND.n7189 VGND.n7188 4.6505
R2976 VGND.n7187 VGND.n7186 4.6505
R2977 VGND.n7185 VGND.n7184 4.6505
R2978 VGND.n7183 VGND.n7182 4.6505
R2979 VGND.n7180 VGND.n7179 4.6505
R2980 VGND.n7175 VGND.n7174 4.6505
R2981 VGND.n7172 VGND.n7171 4.6505
R2982 VGND.n7170 VGND.n7169 4.6505
R2983 VGND.n7039 VGND.n7038 4.6505
R2984 VGND.n7041 VGND.n7040 4.6505
R2985 VGND.n7044 VGND.n7043 4.6505
R2986 VGND.n7047 VGND.n7046 4.6505
R2987 VGND.n7049 VGND.n7048 4.6505
R2988 VGND.n7051 VGND.n7050 4.6505
R2989 VGND.n7053 VGND.n7052 4.6505
R2990 VGND.n7055 VGND.n7054 4.6505
R2991 VGND.n7058 VGND.n7057 4.6505
R2992 VGND.n7060 VGND.n7059 4.6505
R2993 VGND.n7062 VGND.n7061 4.6505
R2994 VGND.n7064 VGND.n7063 4.6505
R2995 VGND.n7066 VGND.n7065 4.6505
R2996 VGND.n7070 VGND.n7069 4.6505
R2997 VGND.n7074 VGND.n7073 4.6505
R2998 VGND.n7076 VGND.n7075 4.6505
R2999 VGND.n7078 VGND.n7077 4.6505
R3000 VGND.n7080 VGND.n7079 4.6505
R3001 VGND.n7082 VGND.n7081 4.6505
R3002 VGND.n7084 VGND.n7083 4.6505
R3003 VGND.n7087 VGND.n7086 4.6505
R3004 VGND.n7091 VGND.n7090 4.6505
R3005 VGND.n7094 VGND.n7093 4.6505
R3006 VGND.n7096 VGND.n7095 4.6505
R3007 VGND.n7099 VGND.n7098 4.6505
R3008 VGND.n7103 VGND.n7102 4.6505
R3009 VGND.n7107 VGND.n7106 4.6505
R3010 VGND.n7111 VGND.n7110 4.6505
R3011 VGND.n7113 VGND.n7112 4.6505
R3012 VGND.n6906 VGND.n6905 4.6505
R3013 VGND.n6908 VGND.n6907 4.6505
R3014 VGND.n6911 VGND.n6910 4.6505
R3015 VGND.n6914 VGND.n6913 4.6505
R3016 VGND.n6916 VGND.n6915 4.6505
R3017 VGND.n6918 VGND.n6917 4.6505
R3018 VGND.n6920 VGND.n6919 4.6505
R3019 VGND.n6922 VGND.n6921 4.6505
R3020 VGND.n6925 VGND.n6924 4.6505
R3021 VGND.n6927 VGND.n6926 4.6505
R3022 VGND.n6929 VGND.n6928 4.6505
R3023 VGND.n6931 VGND.n6930 4.6505
R3024 VGND.n6933 VGND.n6932 4.6505
R3025 VGND.n6938 VGND.n6937 4.6505
R3026 VGND.n6942 VGND.n6941 4.6505
R3027 VGND.n6943 VGND.n1011 4.6505
R3028 VGND.n6945 VGND.n6944 4.6505
R3029 VGND.n6946 VGND.n1010 4.6505
R3030 VGND.n6948 VGND.n6947 4.6505
R3031 VGND.n6949 VGND.n1009 4.6505
R3032 VGND.n6951 VGND.n6950 4.6505
R3033 VGND.n6952 VGND.n1008 4.6505
R3034 VGND.n6954 VGND.n6953 4.6505
R3035 VGND.n6955 VGND.n1007 4.6505
R3036 VGND.n6957 VGND.n6956 4.6505
R3037 VGND.n6959 VGND.n1006 4.6505
R3038 VGND.n6961 VGND.n6960 4.6505
R3039 VGND.n6962 VGND.n1005 4.6505
R3040 VGND.n6964 VGND.n6963 4.6505
R3041 VGND.n6967 VGND.n6966 4.6505
R3042 VGND.n6970 VGND.n6969 4.6505
R3043 VGND.n6974 VGND.n6973 4.6505
R3044 VGND.n6840 VGND.n6839 4.6505
R3045 VGND.n6841 VGND.n6837 4.6505
R3046 VGND.n6843 VGND.n6842 4.6505
R3047 VGND.n6844 VGND.n6836 4.6505
R3048 VGND.n6847 VGND.n6846 4.6505
R3049 VGND.n6848 VGND.n6835 4.6505
R3050 VGND.n6850 VGND.n6849 4.6505
R3051 VGND.n6853 VGND.n6852 4.6505
R3052 VGND.n6855 VGND.n6854 4.6505
R3053 VGND.n6793 VGND.n6792 4.6505
R3054 VGND.n6774 VGND.n1037 4.6505
R3055 VGND.n6771 VGND.n6770 4.6505
R3056 VGND.n2189 VGND.n2177 4.6505
R3057 VGND.n6465 VGND.n6464 4.6505
R3058 VGND.n6477 VGND.n6476 4.6505
R3059 VGND.n6708 VGND.n6656 4.6505
R3060 VGND.n6680 VGND.n6679 4.6505
R3061 VGND.n6678 VGND.n6677 4.6505
R3062 VGND.n6674 VGND.n6673 4.6505
R3063 VGND.n6671 VGND.n6670 4.6505
R3064 VGND.n6669 VGND.n6668 4.6505
R3065 VGND.n6667 VGND.n6666 4.6505
R3066 VGND.n6664 VGND.n6663 4.6505
R3067 VGND.n6707 VGND.n6706 4.6505
R3068 VGND.n6705 VGND.n6704 4.6505
R3069 VGND.n6703 VGND.n6702 4.6505
R3070 VGND.n6701 VGND.n6700 4.6505
R3071 VGND.n6699 VGND.n6698 4.6505
R3072 VGND.n6697 VGND.n6696 4.6505
R3073 VGND.n6695 VGND.n6694 4.6505
R3074 VGND.n6692 VGND.n6691 4.6505
R3075 VGND.n6690 VGND.n6689 4.6505
R3076 VGND.n6688 VGND.n6687 4.6505
R3077 VGND.n6686 VGND.n6685 4.6505
R3078 VGND.n6684 VGND.n6683 4.6505
R3079 VGND.n6682 VGND.n6657 4.6505
R3080 VGND.n6608 VGND.n6607 4.6505
R3081 VGND.n6610 VGND.n6609 4.6505
R3082 VGND.n6612 VGND.n6611 4.6505
R3083 VGND.n6614 VGND.n6613 4.6505
R3084 VGND.n6618 VGND.n6617 4.6505
R3085 VGND.n6620 VGND.n6619 4.6505
R3086 VGND.n6622 VGND.n6621 4.6505
R3087 VGND.n6626 VGND.n6625 4.6505
R3088 VGND.n6628 VGND.n6627 4.6505
R3089 VGND.n6630 VGND.n6629 4.6505
R3090 VGND.n6632 VGND.n6631 4.6505
R3091 VGND.n6635 VGND.n6634 4.6505
R3092 VGND.n6639 VGND.n6638 4.6505
R3093 VGND.n6642 VGND.n6641 4.6505
R3094 VGND.n6727 VGND.n6726 4.6505
R3095 VGND.n6585 VGND.n6584 4.6505
R3096 VGND.n6588 VGND.n6587 4.6505
R3097 VGND.n6590 VGND.n6589 4.6505
R3098 VGND.n6592 VGND.n6591 4.6505
R3099 VGND.n6595 VGND.n6594 4.6505
R3100 VGND.n6597 VGND.n6596 4.6505
R3101 VGND.n6599 VGND.n6598 4.6505
R3102 VGND.n6601 VGND.n6600 4.6505
R3103 VGND.n6603 VGND.n6602 4.6505
R3104 VGND.n6604 VGND.n1043 4.6505
R3105 VGND.n6606 VGND.n6605 4.6505
R3106 VGND.n6467 VGND.n6466 4.6505
R3107 VGND.n6469 VGND.n6468 4.6505
R3108 VGND.n6471 VGND.n6470 4.6505
R3109 VGND.n6473 VGND.n6472 4.6505
R3110 VGND.n6475 VGND.n6474 4.6505
R3111 VGND.n6479 VGND.n6478 4.6505
R3112 VGND.n6481 VGND.n6480 4.6505
R3113 VGND.n6483 VGND.n6482 4.6505
R3114 VGND.n6485 VGND.n6484 4.6505
R3115 VGND.n6492 VGND.n6491 4.6505
R3116 VGND.n6496 VGND.n6495 4.6505
R3117 VGND.n6499 VGND.n6498 4.6505
R3118 VGND.n6501 VGND.n6500 4.6505
R3119 VGND.n6504 VGND.n6503 4.6505
R3120 VGND.n6507 VGND.n6506 4.6505
R3121 VGND.n6513 VGND.n6512 4.6505
R3122 VGND.n6514 VGND.n1042 4.6505
R3123 VGND.n6516 VGND.n6515 4.6505
R3124 VGND.n6523 VGND.n6522 4.6505
R3125 VGND.n6525 VGND.n6524 4.6505
R3126 VGND.n6527 VGND.n6526 4.6505
R3127 VGND.n6529 VGND.n6528 4.6505
R3128 VGND.n6531 VGND.n6530 4.6505
R3129 VGND.n6534 VGND.n6533 4.6505
R3130 VGND.n6463 VGND.n6462 4.6505
R3131 VGND.n6392 VGND.n6391 4.6505
R3132 VGND.n6390 VGND.n6389 4.6505
R3133 VGND.n6769 VGND.n6768 4.6505
R3134 VGND.n6773 VGND.n6772 4.6505
R3135 VGND.n6776 VGND.n6775 4.6505
R3136 VGND.n6778 VGND.n6777 4.6505
R3137 VGND.n6779 VGND.n1036 4.6505
R3138 VGND.n6781 VGND.n6780 4.6505
R3139 VGND.n6783 VGND.n6782 4.6505
R3140 VGND.n6785 VGND.n6784 4.6505
R3141 VGND.n6787 VGND.n6786 4.6505
R3142 VGND.n6789 VGND.n6788 4.6505
R3143 VGND.n6791 VGND.n6790 4.6505
R3144 VGND.n2182 VGND.n2179 4.6505
R3145 VGND.n2185 VGND.n2184 4.6505
R3146 VGND.n2186 VGND.n2178 4.6505
R3147 VGND.n2188 VGND.n2187 4.6505
R3148 VGND.n2191 VGND.n2190 4.6505
R3149 VGND.n2193 VGND.n2192 4.6505
R3150 VGND.n2195 VGND.n2194 4.6505
R3151 VGND.n2198 VGND.n2197 4.6505
R3152 VGND.n6388 VGND.n6387 4.6505
R3153 VGND.n6386 VGND.n6385 4.6505
R3154 VGND.n6384 VGND.n6383 4.6505
R3155 VGND.n6382 VGND.n6381 4.6505
R3156 VGND.n6380 VGND.n6379 4.6505
R3157 VGND.n6378 VGND.n6377 4.6505
R3158 VGND.n6375 VGND.n6374 4.6505
R3159 VGND.n6358 VGND.n6357 4.6505
R3160 VGND.n6360 VGND.n6359 4.6505
R3161 VGND.n6362 VGND.n6361 4.6505
R3162 VGND.n6364 VGND.n6363 4.6505
R3163 VGND.n6366 VGND.n6365 4.6505
R3164 VGND.n6369 VGND.n6368 4.6505
R3165 VGND.n6373 VGND.n6372 4.6505
R3166 VGND.n6354 VGND.n6353 4.6505
R3167 VGND.n6767 VGND.n1038 4.6505
R3168 VGND.n6351 VGND.n1039 4.6505
R3169 VGND.n553 VGND.n434 4.6505
R3170 VGND.n545 VGND.n544 4.6505
R3171 VGND.n536 VGND.n16 4.6505
R3172 VGND.n507 VGND.n506 4.6505
R3173 VGND.n505 VGND.n448 4.6505
R3174 VGND.n504 VGND.n449 4.6505
R3175 VGND.n501 VGND.n500 4.6505
R3176 VGND.n498 VGND.n451 4.6505
R3177 VGND.n632 VGND.n15 4.6505
R3178 VGND.n624 VGND.n623 4.6505
R3179 VGND.n616 VGND.n409 4.6505
R3180 VGND.n7972 VGND.n11 4.6505
R3181 VGND.n7431 VGND.n7430 4.6505
R3182 VGND.n7435 VGND.n7434 4.6505
R3183 VGND.n7439 VGND.n7438 4.6505
R3184 VGND.n7443 VGND.n7442 4.6505
R3185 VGND.n7446 VGND.n7445 4.6505
R3186 VGND.n7990 VGND.n7989 4.6505
R3187 VGND.n7984 VGND.n7983 4.6505
R3188 VGND.n7981 VGND.n7980 4.6505
R3189 VGND.n7979 VGND.n7978 4.6505
R3190 VGND.n7977 VGND.n7976 4.6505
R3191 VGND.n7975 VGND.n7974 4.6505
R3192 VGND.n309 VGND.n13 4.6505
R3193 VGND.n311 VGND.n308 4.6505
R3194 VGND.n313 VGND.n312 4.6505
R3195 VGND.n315 VGND.n314 4.6505
R3196 VGND.n316 VGND.n307 4.6505
R3197 VGND.n318 VGND.n317 4.6505
R3198 VGND.n319 VGND.n306 4.6505
R3199 VGND.n322 VGND.n321 4.6505
R3200 VGND.n323 VGND.n305 4.6505
R3201 VGND.n325 VGND.n324 4.6505
R3202 VGND.n327 VGND.n304 4.6505
R3203 VGND.n329 VGND.n328 4.6505
R3204 VGND.n330 VGND.n303 4.6505
R3205 VGND.n332 VGND.n331 4.6505
R3206 VGND.n333 VGND.n302 4.6505
R3207 VGND.n335 VGND.n334 4.6505
R3208 VGND.n337 VGND.n336 4.6505
R3209 VGND.n338 VGND.n300 4.6505
R3210 VGND.n340 VGND.n339 4.6505
R3211 VGND.n341 VGND.n299 4.6505
R3212 VGND.n343 VGND.n342 4.6505
R3213 VGND.n345 VGND.n344 4.6505
R3214 VGND.n348 VGND.n347 4.6505
R3215 VGND.n682 VGND.n681 4.6505
R3216 VGND.n679 VGND.n678 4.6505
R3217 VGND.n675 VGND.n674 4.6505
R3218 VGND.n673 VGND.n672 4.6505
R3219 VGND.n671 VGND.n670 4.6505
R3220 VGND.n668 VGND.n667 4.6505
R3221 VGND.n666 VGND.n665 4.6505
R3222 VGND.n663 VGND.n662 4.6505
R3223 VGND.n661 VGND.n660 4.6505
R3224 VGND.n657 VGND.n401 4.6505
R3225 VGND.n656 VGND.n655 4.6505
R3226 VGND.n653 VGND.n652 4.6505
R3227 VGND.n651 VGND.n650 4.6505
R3228 VGND.n649 VGND.n403 4.6505
R3229 VGND.n648 VGND.n647 4.6505
R3230 VGND.n634 VGND.n633 4.6505
R3231 VGND.n550 VGND.n549 4.6505
R3232 VGND.n533 VGND.n532 4.6505
R3233 VGND.n495 VGND.n494 4.6505
R3234 VGND.n497 VGND.n496 4.6505
R3235 VGND.n499 VGND.n450 4.6505
R3236 VGND.n503 VGND.n502 4.6505
R3237 VGND.n508 VGND.n447 4.6505
R3238 VGND.n510 VGND.n509 4.6505
R3239 VGND.n511 VGND.n446 4.6505
R3240 VGND.n513 VGND.n512 4.6505
R3241 VGND.n515 VGND.n445 4.6505
R3242 VGND.n517 VGND.n516 4.6505
R3243 VGND.n518 VGND.n444 4.6505
R3244 VGND.n520 VGND.n519 4.6505
R3245 VGND.n521 VGND.n443 4.6505
R3246 VGND.n523 VGND.n522 4.6505
R3247 VGND.n524 VGND.n442 4.6505
R3248 VGND.n526 VGND.n525 4.6505
R3249 VGND.n527 VGND.n441 4.6505
R3250 VGND.n530 VGND.n529 4.6505
R3251 VGND.n531 VGND.n440 4.6505
R3252 VGND.n535 VGND.n534 4.6505
R3253 VGND.n537 VGND.n439 4.6505
R3254 VGND.n539 VGND.n538 4.6505
R3255 VGND.n540 VGND.n438 4.6505
R3256 VGND.n542 VGND.n541 4.6505
R3257 VGND.n543 VGND.n437 4.6505
R3258 VGND.n547 VGND.n546 4.6505
R3259 VGND.n548 VGND.n435 4.6505
R3260 VGND.n552 VGND.n551 4.6505
R3261 VGND.n555 VGND.n554 4.6505
R3262 VGND.n613 VGND.n612 4.6505
R3263 VGND.n615 VGND.n614 4.6505
R3264 VGND.n618 VGND.n617 4.6505
R3265 VGND.n620 VGND.n619 4.6505
R3266 VGND.n622 VGND.n621 4.6505
R3267 VGND.n626 VGND.n625 4.6505
R3268 VGND.n629 VGND.n628 4.6505
R3269 VGND.n631 VGND.n630 4.6505
R3270 VGND VGND.n406 4.6505
R3271 VGND.n7433 VGND.n7432 4.6505
R3272 VGND.n7437 VGND.n7436 4.6505
R3273 VGND.n7441 VGND.n7440 4.6505
R3274 VGND.n7444 VGND.n7427 4.6505
R3275 VGND.n7954 VGND.n7953 4.6505
R3276 VGND.n7951 VGND.n7950 4.6505
R3277 VGND.n7946 VGND.n7945 4.6505
R3278 VGND.n7943 VGND.n7942 4.6505
R3279 VGND.n7940 VGND.n7939 4.6505
R3280 VGND.n7938 VGND.n7905 4.6505
R3281 VGND.n7937 VGND.n7936 4.6505
R3282 VGND.n7935 VGND.n7906 4.6505
R3283 VGND.n7934 VGND.n7933 4.6505
R3284 VGND.n7932 VGND.n7907 4.6505
R3285 VGND.n7931 VGND.n7930 4.6505
R3286 VGND.n7929 VGND.n7908 4.6505
R3287 VGND.n7928 VGND.n7927 4.6505
R3288 VGND.n7926 VGND.n7909 4.6505
R3289 VGND.n7925 VGND.n7924 4.6505
R3290 VGND.n7923 VGND.n7910 4.6505
R3291 VGND.n7922 VGND.n7911 4.6505
R3292 VGND.n7921 VGND.n7912 4.6505
R3293 VGND.n7920 VGND.n7913 4.6505
R3294 VGND.n7919 VGND.n7918 4.6505
R3295 VGND.n7917 VGND.n7914 4.6505
R3296 VGND.n233 VGND.n232 4.57427
R3297 VGND.n3463 VGND.n849 4.57427
R3298 VGND.n3364 VGND.n3363 4.57427
R3299 VGND.n7401 VGND.n7400 4.57427
R3300 VGND.n7512 VGND.n7511 4.57427
R3301 VGND.n7688 VGND.n7687 4.57427
R3302 VGND.n3332 VGND.n3255 4.57427
R3303 VGND.n7847 VGND.n7846 4.57427
R3304 VGND.n7596 VGND.n7595 4.57427
R3305 VGND.n4215 VGND.n4214 4.57427
R3306 VGND.n4130 VGND.n4129 4.57427
R3307 VGND.n3918 VGND.n3917 4.57427
R3308 VGND.n3779 VGND.n3778 4.57427
R3309 VGND.n4194 VGND.n4193 4.57427
R3310 VGND.n4461 VGND.n4460 4.57427
R3311 VGND.n4681 VGND.n4680 4.57427
R3312 VGND.n4542 VGND.n4541 4.57427
R3313 VGND.n4381 VGND.n4380 4.57427
R3314 VGND.n4365 VGND.n4364 4.57427
R3315 VGND.n5156 VGND.n5155 4.57427
R3316 VGND.n5061 VGND.n5060 4.57427
R3317 VGND.n4958 VGND.n4957 4.57427
R3318 VGND.n5135 VGND.n5134 4.57427
R3319 VGND.n4759 VGND.n4758 4.57427
R3320 VGND.n2515 VGND.n2512 4.57427
R3321 VGND.n5275 VGND.n5274 4.57427
R3322 VGND.n5309 VGND.n5308 4.57427
R3323 VGND.n2393 VGND.n2392 4.57427
R3324 VGND.n2697 VGND.n2696 4.57427
R3325 VGND.n1782 VGND.n1764 4.57427
R3326 VGND.n2344 VGND.n2343 4.57427
R3327 VGND.n5338 VGND.n5337 4.57427
R3328 VGND.n5544 VGND.n5543 4.57427
R3329 VGND.n1741 VGND.n1740 4.57427
R3330 VGND.n5739 VGND.n5738 4.57427
R3331 VGND.n5893 VGND.n5892 4.57427
R3332 VGND.n5988 VGND.n5987 4.57427
R3333 VGND.n2300 VGND.n2299 4.57427
R3334 VGND.n1914 VGND.n1913 4.57427
R3335 VGND.n2023 VGND.n1992 4.57427
R3336 VGND.n1975 VGND.n1974 4.57427
R3337 VGND.n6248 VGND.n6247 4.57427
R3338 VGND.n2151 VGND.n2150 4.57427
R3339 VGND.n6110 VGND.n6109 4.57427
R3340 VGND.n7325 VGND.n7324 4.57427
R3341 VGND.n7160 VGND.n7159 4.57427
R3342 VGND.n6989 VGND.n6988 4.57427
R3343 VGND.n6903 VGND.n6902 4.57427
R3344 VGND.n6871 VGND.n6870 4.57427
R3345 VGND.n6395 VGND.n6394 4.57427
R3346 VGND.n6575 VGND.n6574 4.57427
R3347 VGND.n6795 VGND.n6794 4.57427
R3348 VGND.n2220 VGND.n2219 4.57427
R3349 VGND.n359 VGND.n358 4.57427
R3350 VGND.n7966 VGND.n7965 4.57427
R3351 VGND.n579 VGND.n578 4.57427
R3352 VGND.n7460 VGND.n7459 4.57427
R3353 VGND.n3800 VGND.n3148 4.57412
R3354 VGND.n5790 VGND.n1369 4.57412
R3355 VGND.n7037 VGND.n7036 4.57412
R3356 VGND.n685 VGND.n14 4.57412
R3357 VGND.n710 VGND.n178 4.57412
R3358 VGND.n7746 VGND.n80 4.57412
R3359 VGND.n5633 VGND.n1396 4.57412
R3360 VGND.n6289 VGND.n6288 4.57412
R3361 VGND.n1066 VGND.n1065 4.5622
R3362 VGND.n6078 VGND.n6077 4.5622
R3363 VGND.n3990 VGND.n3989 4.5622
R3364 VGND.n1284 VGND.n1283 4.5622
R3365 VGND.n2206 VGND.n2205 4.53348
R3366 VGND.n4282 VGND.n4281 4.53348
R3367 VGND.n5126 VGND.n5125 4.53348
R3368 VGND.n1737 VGND.n1736 4.53348
R3369 VGND.n6799 VGND.n6798 4.5303
R3370 VGND.n2095 VGND.n1973 4.5303
R3371 VGND.n2415 VGND.n2414 4.5303
R3372 VGND.n5282 VGND.n5281 4.52113
R3373 VGND.n5822 VGND.n1365 4.51815
R3374 VGND.n3730 VGND.n3729 4.5005
R3375 VGND.n4484 VGND.n4483 4.5005
R3376 VGND.n4785 VGND.n4784 4.5005
R3377 VGND.n2550 VGND.n2549 4.5005
R3378 VGND.n5648 VGND.n5647 4.5005
R3379 VGND.n5696 VGND.n5695 4.5005
R3380 VGND.n7015 VGND.n7014 4.5005
R3381 VGND.n6422 VGND.n6421 4.5005
R3382 VGND.n396 VGND.n395 4.5005
R3383 VGND.n6280 VGND.n6279 4.49598
R3384 VGND.n1102 VGND.n1042 4.42603
R3385 VGND.n5274 VGND.n5271 4.41955
R3386 VGND.n6517 VGND.n6516 4.28986
R3387 VGND.n897 VGND.n896 4.28986
R3388 VGND.n2087 VGND.n2086 4.28986
R3389 VGND.n3810 VGND.n3809 4.28986
R3390 VGND.n2930 VGND.n2929 4.28986
R3391 VGND.n5827 VGND.n1364 4.28986
R3392 VGND.n1759 VGND.n1758 4.18553
R3393 VGND.n6119 VGND.n6118 4.14168
R3394 VGND.n3536 VGND.n3535 4.14168
R3395 VGND.n1492 VGND.n1491 4.14168
R3396 VGND.n1309 VGND.n1308 4.14168
R3397 VGND.n515 VGND.n514 4.11798
R3398 VGND.n514 VGND.n513 4.11798
R3399 VGND.n347 VGND.n346 4.11798
R3400 VGND.n6641 VGND.n6640 4.11798
R3401 VGND.n6640 VGND.n1059 4.11798
R3402 VGND.n6594 VGND.n6593 4.11798
R3403 VGND.n917 VGND.n916 4.11798
R3404 VGND.n7235 VGND.n7234 4.11798
R3405 VGND.n7057 VGND.n7056 4.11798
R3406 VGND.n6958 VGND.n6957 4.11798
R3407 VGND.n6959 VGND.n6958 4.11798
R3408 VGND.n6924 VGND.n6923 4.11798
R3409 VGND.n6190 VGND.n6189 4.11798
R3410 VGND.n6189 VGND.n6188 4.11798
R3411 VGND.n2052 VGND.n2051 4.11798
R3412 VGND.n6211 VGND.n1223 4.11798
R3413 VGND.n6208 VGND.n1223 4.11798
R3414 VGND.n779 VGND.n778 4.11798
R3415 VGND.n778 VGND.n777 4.11798
R3416 VGND.n3206 VGND.n3205 4.11798
R3417 VGND.n3230 VGND.n3229 4.11798
R3418 VGND.n7662 VGND.n7661 4.11798
R3419 VGND.n7661 VGND.n7660 4.11798
R3420 VGND.n7812 VGND.n7811 4.11798
R3421 VGND.n4145 VGND.n3143 4.11798
R3422 VGND.n4142 VGND.n3143 4.11798
R3423 VGND.n2983 VGND.n2982 4.11798
R3424 VGND.n2984 VGND.n2983 4.11798
R3425 VGND.n5086 VGND.n5085 4.11798
R3426 VGND.n5085 VGND.n5084 4.11798
R3427 VGND.n2809 VGND.n2762 4.11798
R3428 VGND.n2762 VGND.n2761 4.11798
R3429 VGND.n4982 VGND.n4981 4.11798
R3430 VGND.n4981 VGND.n4980 4.11798
R3431 VGND.n5029 VGND.n5028 4.11798
R3432 VGND.n4737 VGND.n4736 4.11798
R3433 VGND.n2486 VGND.n2485 4.11798
R3434 VGND.n2668 VGND.n2667 4.11798
R3435 VGND.n2667 VGND.n2666 4.11798
R3436 VGND.n5376 VGND.n5375 4.11798
R3437 VGND.n5400 VGND.n5399 4.11798
R3438 VGND.n1799 VGND.n1798 4.11798
R3439 VGND.n5763 VGND.n5762 4.11798
R3440 VGND.n5916 VGND.n5915 4.11798
R3441 VGND.n5918 VGND.n5916 4.11798
R3442 VGND.n6264 VGND.n6263 4.11798
R3443 VGND.n6356 VGND.n6350 4.09013
R3444 VGND.n8 VGND.n3 4.07323
R3445 VGND.n896 VGND.n895 4.07323
R3446 VGND.n3448 VGND.n3447 4.07323
R3447 VGND.n3262 VGND.n3261 4.07323
R3448 VGND.n7785 VGND.n7784 4.07323
R3449 VGND.n3809 VGND.n3666 4.07323
R3450 VGND.n4248 VGND.n4247 4.07323
R3451 VGND.n4249 VGND.n4248 4.07323
R3452 VGND.n5830 VGND.n1364 4.07323
R3453 VGND.n5831 VGND.n5830 4.07323
R3454 VGND.n1258 VGND.n1257 4.07323
R3455 VGND.n7956 VGND.n7955 4.07323
R3456 VGND.n6505 VGND.n6504 4.03876
R3457 VGND.n7400 VGND.n7399 4.03876
R3458 VGND.n4718 VGND.n2733 4.03876
R3459 VGND.n7657 VGND.n7656 4.01961
R3460 VGND.n7973 VGND.n7972 3.97459
R3461 VGND.n7374 VGND.n7373 3.97459
R3462 VGND.n5285 VGND.n1649 3.97459
R3463 VGND.n641 VGND.n640 3.96548
R3464 VGND.n318 VGND.n307 3.96548
R3465 VGND.n319 VGND.n318 3.96548
R3466 VGND.n6678 VGND.n6660 3.96548
R3467 VGND.n6660 VGND.n6659 3.96548
R3468 VGND.n1063 VGND.n1062 3.96548
R3469 VGND.n6626 VGND.n1063 3.96548
R3470 VGND.n6511 VGND.n6510 3.96548
R3471 VGND.n6512 VGND.n6511 3.96548
R3472 VGND.n188 VGND.n187 3.96548
R3473 VGND.n197 VGND.n188 3.96548
R3474 VGND.n744 VGND.n743 3.96548
R3475 VGND.n743 VGND.n742 3.96548
R3476 VGND.n3196 VGND.n3195 3.96548
R3477 VGND.n107 VGND.n106 3.96548
R3478 VGND.n7674 VGND.n107 3.96548
R3479 VGND.n3848 VGND.n3656 3.96548
R3480 VGND.n3849 VGND.n3848 3.96548
R3481 VGND.n4451 VGND.n4243 3.96548
R3482 VGND.n4721 VGND.n4720 3.96548
R3483 VGND.n4720 VGND.n4719 3.96548
R3484 VGND.n6574 VGND.n6573 3.9624
R3485 VGND.n5274 VGND.n5273 3.9624
R3486 VGND.n3252 VGND.n3169 3.96015
R3487 VGND.n642 VGND.n641 3.89322
R3488 VGND.n3279 VGND.n3260 3.85748
R3489 VGND.n7777 VGND.n7776 3.85748
R3490 VGND.n3925 VGND.n3924 3.83619
R3491 VGND.n3263 VGND.n3262 3.76521
R3492 VGND.n7786 VGND.n7785 3.76521
R3493 VGND.n4460 VGND.n4459 3.7575
R3494 VGND.n7582 VGND.n7581 3.6638
R3495 VGND.n1232 VGND 3.56771
R3496 VGND.n1878 VGND 3.56771
R3497 VGND.n7595 VGND.n7594 3.53451
R3498 VGND.n639 VGND.n638 3.50735
R3499 VGND.n2078 VGND.n2077 3.50735
R3500 VGND.n3298 VGND.n3256 3.50735
R3501 VGND.n3691 VGND.n3679 3.50735
R3502 VGND.n3977 VGND.n3969 3.50735
R3503 VGND.n3935 VGND.n3934 3.50735
R3504 VGND.n3018 VGND.n3017 3.50735
R3505 VGND.n2785 VGND.n2766 3.50735
R3506 VGND.n2615 VGND.n2614 3.50735
R3507 VGND.n6489 VGND.n6488 3.44377
R3508 VGND.n3388 VGND.n3387 3.44377
R3509 VGND.n3387 VGND.n3386 3.44377
R3510 VGND.n3007 VGND.n3006 3.44377
R3511 VGND.n3006 VGND.n3005 3.44377
R3512 VGND.n155 VGND.n154 3.4105
R3513 VGND VGND.n7495 3.4105
R3514 VGND.n7879 VGND.n7878 3.4105
R3515 VGND.n3559 VGND.n3558 3.4105
R3516 VGND.n3361 VGND.n3360 3.4105
R3517 VGND.n7405 VGND.n7404 3.4105
R3518 VGND.n714 VGND.n713 3.4105
R3519 VGND.n3592 VGND.n3591 3.4105
R3520 VGND.n7743 VGND.n7742 3.4105
R3521 VGND.n3910 VGND.n3909 3.4105
R3522 VGND.n4088 VGND.n4087 3.4105
R3523 VGND.n4126 VGND.n4125 3.4105
R3524 VGND.n3797 VGND.n3796 3.4105
R3525 VGND.n4360 VGND.n4359 3.4105
R3526 VGND.n4649 VGND.n4648 3.4105
R3527 VGND.n4691 VGND.n4690 3.4105
R3528 VGND.n2844 VGND.n2843 3.4105
R3529 VGND.n5057 VGND.n5056 3.4105
R3530 VGND.n2824 VGND.n2823 3.4105
R3531 VGND.n4910 VGND.n2857 3.4105
R3532 VGND.n4948 VGND.n4946 3.4105
R3533 VGND.n4816 VGND.n4815 3.4105
R3534 VGND.n5202 VGND.n5201 3.4105
R3535 VGND.n2714 VGND 3.4105
R3536 VGND.n1572 VGND.n1571 3.4105
R3537 VGND.n1582 VGND.n1481 3.4105
R3538 VGND.n2561 VGND.n2560 3.4105
R3539 VGND.n2400 VGND.n2399 3.4105
R3540 VGND.n1735 VGND.n1734 3.4105
R3541 VGND.n2360 VGND 3.4105
R3542 VGND.n5419 VGND.n5418 3.4105
R3543 VGND.n5430 VGND.n5429 3.4105
R3544 VGND.n5441 VGND.n5440 3.4105
R3545 VGND.n5645 VGND.n5644 3.4105
R3546 VGND.n1747 VGND.n1746 3.4105
R3547 VGND.n6001 VGND.n6000 3.4105
R3548 VGND.n1898 VGND.n1897 3.4105
R3549 VGND.n2317 VGND 3.4105
R3550 VGND.n5674 VGND.n5673 3.4105
R3551 VGND.n1920 VGND.n1919 3.4105
R3552 VGND.n5686 VGND.n5685 3.4105
R3553 VGND.n2135 VGND.n2134 3.4105
R3554 VGND.n2285 VGND 3.4105
R3555 VGND.n2272 VGND.n2271 3.4105
R3556 VGND.n2159 VGND.n2158 3.4105
R3557 VGND.n2098 VGND.n2097 3.4105
R3558 VGND.n6302 VGND.n6301 3.4105
R3559 VGND.n6102 VGND.n6101 3.4105
R3560 VGND.n6899 VGND.n6898 3.4105
R3561 VGND.n7281 VGND.n940 3.4105
R3562 VGND.n7031 VGND.n7030 3.4105
R3563 VGND.n2215 VGND.n2214 3.4105
R3564 VGND.n6714 VGND.n6713 3.4105
R3565 VGND.n6755 VGND.n6754 3.4105
R3566 VGND.n6455 VGND.n6454 3.4105
R3567 VGND.n8005 VGND.n8004 3.4105
R3568 VGND.n473 VGND.n472 3.4105
R3569 VGND.n7464 VGND.n7463 3.4105
R3570 VGND.n689 VGND.n688 3.4105
R3571 VGND.n7511 VGND.n7510 3.36212
R3572 VGND.n3917 VGND.n3916 3.36212
R3573 VGND.n3479 VGND 3.29747
R3574 VGND.n3263 VGND 3.29747
R3575 VGND.n2770 VGND 3.29747
R3576 VGND.n1402 VGND 3.29747
R3577 VGND.n1764 VGND.n1763 3.21921
R3578 VGND.n637 VGND.n634 3.2005
R3579 VGND.n975 VGND.n974 3.2005
R3580 VGND.n2074 VGND.n1983 3.2005
R3581 VGND.n3400 VGND.n3347 3.2005
R3582 VGND.n805 VGND.n804 3.2005
R3583 VGND.n3297 VGND.n3294 3.2005
R3584 VGND.n77 VGND.n76 3.2005
R3585 VGND.n3625 VGND.n3624 3.2005
R3586 VGND.n3695 VGND.n3694 3.2005
R3587 VGND.n3976 VGND.n3973 3.2005
R3588 VGND.n3933 VGND.n3930 3.2005
R3589 VGND.n3016 VGND.n3013 3.2005
R3590 VGND.n2784 VGND.n2768 3.2005
R3591 VGND.n2620 VGND.n2618 3.2005
R3592 VGND.n5932 VGND.n5931 3.2005
R3593 VGND.n528 VGND.n527 3.13242
R3594 VGND.n625 VGND.n408 3.13242
R3595 VGND.n7099 VGND.n968 3.13242
R3596 VGND.n6845 VGND.n6835 3.13242
R3597 VGND.n3432 VGND.n3344 3.13242
R3598 VGND.n4035 VGND.n4034 3.13242
R3599 VGND.n3822 VGND.n3661 3.13242
R3600 VGND.n4258 VGND.n4257 3.13242
R3601 VGND.n4575 VGND.n2960 3.13242
R3602 VGND.n2655 VGND.n2624 3.13242
R3603 VGND.n1817 VGND.n1755 3.13242
R3604 VGND.n1913 VGND.n1912 3.13242
R3605 VGND.n1926 VGND.n1371 3.13242
R3606 VGND.n529 VGND.n528 3.13241
R3607 VGND.n578 VGND.n577 3.13241
R3608 VGND.n408 VGND.n407 3.13241
R3609 VGND.n2197 VGND.n2196 3.13241
R3610 VGND.n968 VGND.n967 3.13241
R3611 VGND.n6846 VGND.n6845 3.13241
R3612 VGND.n3344 VGND.n3343 3.13241
R3613 VGND.n3414 VGND.n3413 3.13241
R3614 VGND.n3374 VGND.n3373 3.13241
R3615 VGND.n4036 VGND.n4035 3.13241
R3616 VGND.n4051 VGND.n4050 3.13241
R3617 VGND.n3823 VGND.n3822 3.13241
R3618 VGND.n4257 VGND.n4256 3.13241
R3619 VGND.n4576 VGND.n4575 3.13241
R3620 VGND.n4541 VGND.n4540 3.13241
R3621 VGND.n5000 VGND 3.13241
R3622 VGND.n2624 VGND.n2623 3.13241
R3623 VGND.n5455 VGND.n5454 3.13241
R3624 VGND.n1755 VGND.n1754 3.13241
R3625 VGND.n1750 VGND.n1749 3.13241
R3626 VGND.n1267 VGND.n1266 3.13241
R3627 VGND.n1944 VGND.n1943 3.13241
R3628 VGND.n5738 VGND.n5737 3.13241
R3629 VGND.n5892 VGND.n5891 3.13241
R3630 VGND.n1927 VGND.n1926 3.13241
R3631 VGND.n7 VGND.n6 3.06298
R3632 VGND.n4374 VGND.n4252 3.06297
R3633 VGND.n6322 VGND.n6306 3.06215
R3634 VGND.n3758 VGND.n3727 3.06214
R3635 VGND.n818 VGND.n817 3.06214
R3636 VGND.n7974 VGND.n7973 3.05276
R3637 VGND.n7375 VGND.n7374 3.05276
R3638 VGND.n5282 VGND.n1649 3.05276
R3639 VGND.n2024 VGND.n2019 3.01896
R3640 VGND.n3781 VGND.n3780 3.01896
R3641 VGND.n2517 VGND.n2516 3.01896
R3642 VGND.n5740 VGND.n1377 3.01896
R3643 VGND.n6987 VGND.n6986 3.01896
R3644 VGND.n357 VGND.n356 3.01896
R3645 VGND.n7658 VGND.n7657 3.01483
R3646 VGND.n7882 VGND.n7881 3.0005
R3647 VGND.n3886 VGND.n3885 3.0005
R3648 VGND.n2712 VGND.n2711 3.0005
R3649 VGND.n5718 VGND.n5717 3.0005
R3650 VGND.n2315 VGND.n2314 3.0005
R3651 VGND.n6319 VGND.n6318 3.0005
R3652 VGND.n2283 VGND.n2282 3.0005
R3653 VGND.n7153 VGND.n7152 3.0005
R3654 VGND.n6883 VGND.n6882 3.0005
R3655 VGND.n2239 VGND.n2238 3.0005
R3656 VGND.n8020 VGND.n8019 3.0005
R3657 VGND.n5000 VGND.n4999 2.9514
R3658 VGND.n7642 VGND.n110 2.90959
R3659 VGND.n557 VGND.n556 2.90012
R3660 VGND.n406 VGND.n404 2.89365
R3661 VGND.n7091 VGND.n976 2.89365
R3662 VGND.n2073 VGND.n2072 2.89365
R3663 VGND.n3402 VGND.n3401 2.89365
R3664 VGND.n831 VGND.n806 2.89365
R3665 VGND.n3293 VGND.n3292 2.89365
R3666 VGND.n7765 VGND.n78 2.89365
R3667 VGND.n4001 VGND.n3626 2.89365
R3668 VGND.n3698 VGND.n3677 2.89365
R3669 VGND.n3024 VGND.n2974 2.89365
R3670 VGND.n2782 VGND.n2781 2.89365
R3671 VGND.n2619 VGND.n2422 2.89365
R3672 VGND.n5954 VGND.n5933 2.89365
R3673 VGND.n7750 VGND.n79 2.8567
R3674 VGND.n3198 VGND.n3169 2.84782
R3675 VGND.n6506 VGND.n6505 2.77203
R3676 VGND.n3917 VGND.n3914 2.77203
R3677 VGND.n4721 VGND.n4718 2.77203
R3678 VGND.n3394 VGND.n848 2.76214
R3679 VGND.n4905 VGND.n4904 2.71831
R3680 VGND.n2800 VGND.n2799 2.63579
R3681 VGND.n7941 VGND.n7940 2.63579
R3682 VGND.n755 VGND.n754 2.55412
R3683 VGND.n738 VGND.n737 2.47351
R3684 VGND.n3461 VGND.n3460 2.47351
R3685 VGND.n7717 VGND.n7716 2.47351
R3686 VGND.n3335 VGND.n3334 2.47351
R3687 VGND.n3757 VGND.n3756 2.47351
R3688 VGND.n4112 VGND.n4111 2.47351
R3689 VGND.n4489 VGND.n4488 2.47351
R3690 VGND.n4629 VGND.n4628 2.47351
R3691 VGND.n2834 VGND.n2833 2.47351
R3692 VGND.n4790 VGND.n4789 2.47351
R3693 VGND.n2547 VGND.n2546 2.47351
R3694 VGND.n5312 VGND.n5311 2.47351
R3695 VGND.n5333 VGND.n5332 2.47351
R3696 VGND.n5654 VGND.n5653 2.47351
R3697 VGND.n5709 VGND.n5707 2.47351
R3698 VGND.n5991 VGND.n5990 2.47351
R3699 VGND.n6324 VGND.n6323 2.47351
R3700 VGND.n6105 VGND.n6104 2.47351
R3701 VGND.n7283 VGND.n7282 2.47351
R3702 VGND.n7018 VGND.n7017 2.47351
R3703 VGND.n6426 VGND.n6425 2.47351
R3704 VGND.n6741 VGND.n6740 2.47351
R3705 VGND.n391 VGND.n388 2.47351
R3706 VGND.n459 VGND.n458 2.47351
R3707 VGND.n1066 VGND.n1064 2.44756
R3708 VGND VGND.n7 2.36572
R3709 VGND.n670 VGND.n669 2.33701
R3710 VGND.n665 VGND.n664 2.33701
R3711 VGND.n334 VGND.n301 2.33701
R3712 VGND.n337 VGND.n301 2.33701
R3713 VGND.n326 VGND.n325 2.33701
R3714 VGND.n327 VGND.n326 2.33701
R3715 VGND.n7983 VGND.n7982 2.33701
R3716 VGND.n6694 VGND.n6693 2.33701
R3717 VGND.n6634 VGND.n6633 2.33701
R3718 VGND.n6533 VGND.n6532 2.33701
R3719 VGND.n6574 VGND.n6571 2.33701
R3720 VGND.n6064 VGND.n6063 2.33701
R3721 VGND.n6057 VGND.n6056 2.33701
R3722 VGND.n207 VGND.n206 2.33701
R3723 VGND.n229 VGND.n228 2.33701
R3724 VGND.n763 VGND.n762 2.33701
R3725 VGND.n7380 VGND.n7379 2.33701
R3726 VGND.n7684 VGND.n7683 2.33701
R3727 VGND.n7631 VGND.n7630 2.33701
R3728 VGND.n6368 VGND.n6367 2.33701
R3729 VGND.n6349 VGND.n6348 2.33701
R3730 VGND.n6373 VGND.n6349 2.33701
R3731 VGND.n759 VGND.n758 2.33067
R3732 VGND.n191 VGND.n190 2.29662
R3733 VGND.n785 VGND.n784 2.29662
R3734 VGND.n7668 VGND.n7667 2.29662
R3735 VGND.n7614 VGND.n7613 2.29662
R3736 VGND.n3842 VGND.n3841 2.29662
R3737 VGND.n2084 VGND.n2083 2.29662
R3738 VGND.n6582 VGND.n6581 2.29662
R3739 VGND.n6494 VGND.n6493 2.29662
R3740 VGND.n6519 VGND.n6518 2.29662
R3741 VGND.n6521 VGND.n6520 2.29662
R3742 VGND.n7992 VGND.n3 2.29662
R3743 VGND.n659 VGND.n658 2.29662
R3744 VGND.n5001 VGND.n2854 2.29643
R3745 VGND.n6761 VGND.n6760 2.2824
R3746 VGND.n4672 VGND.n4671 2.2824
R3747 VGND.n7957 VGND.n7956 2.28222
R3748 VGND.n4655 VGND.n4654 2.28171
R3749 VGND.n3564 VGND.n3448 2.28159
R3750 VGND.n6730 VGND.n6729 2.28159
R3751 VGND.n2534 VGND.n2462 2.28155
R3752 VGND.n6313 VGND.n6307 2.28144
R3753 VGND.n7615 VGND.n7614 2.26126
R3754 VGND.n1245 VGND.n1244 2.23612
R3755 VGND.n761 VGND.n760 2.10723
R3756 VGND.n6571 VGND.n6570 2.08304
R3757 VGND.n4242 VGND.n4241 2.06919
R3758 VGND.n3971 VGND.n3630 2.01694
R3759 VGND.n647 VGND.n646 1.98299
R3760 VGND.n320 VGND.n319 1.98299
R3761 VGND.n321 VGND.n320 1.98299
R3762 VGND.n6673 VGND.n6672 1.98299
R3763 VGND.n3197 VGND.n3196 1.98299
R3764 VGND.n3198 VGND.n3197 1.98299
R3765 VGND.n3850 VGND.n3849 1.98299
R3766 VGND.n3851 VGND.n3850 1.98299
R3767 VGND.n4446 VGND.n4445 1.98299
R3768 VGND.n2813 VGND.n2812 1.98299
R3769 VGND.n4774 VGND.n4773 1.97497
R3770 VGND.n6666 VGND.n6665 1.8968
R3771 VGND.n4243 VGND.n4242 1.8968
R3772 VGND VGND.n1739 1.88285
R3773 VGND.n6516 VGND.n1102 1.8388
R3774 VGND.n6490 VGND.n6489 1.79699
R3775 VGND.n3005 VGND.n3004 1.72214
R3776 VGND VGND.n3860 1.7012
R3777 VGND.n2629 VGND.n2628 1.67669
R3778 VGND.n6491 VGND.n6490 1.64728
R3779 VGND.n6222 VGND 1.61169
R3780 VGND.n546 VGND.n436 1.6005
R3781 VGND.n2183 VGND.n2178 1.6005
R3782 VGND.n6908 VGND.n1014 1.6005
R3783 VGND.n2032 VGND.n1990 1.6005
R3784 VGND.n1124 VGND.n1123 1.6005
R3785 VGND.n3480 VGND.n3469 1.6005
R3786 VGND.n133 VGND.n126 1.6005
R3787 VGND.n7571 VGND.n7564 1.6005
R3788 VGND.n4180 VGND.n4160 1.6005
R3789 VGND.n3958 VGND.n3632 1.6005
R3790 VGND.n4270 VGND.n4269 1.6005
R3791 VGND.n4569 VGND.n4568 1.6005
R3792 VGND.n3003 VGND.n2975 1.6005
R3793 VGND.n1538 VGND.n1484 1.6005
R3794 VGND.n5181 VGND.n5173 1.6005
R3795 VGND.n2512 VGND.n2511 1.6005
R3796 VGND.n5481 VGND.n1456 1.6005
R3797 VGND.n5598 VGND.n1401 1.6005
R3798 VGND.n1399 VGND.n1398 1.6005
R3799 VGND.n5781 VGND.n1373 1.6005
R3800 VGND.n5841 VGND.n1360 1.6005
R3801 VGND.n5980 VGND.n5926 1.6005
R3802 VGND.n6280 VGND.n1179 1.6005
R3803 VGND VGND.n401 1.52218
R3804 VGND VGND.n343 1.52218
R3805 VGND.n4433 VGND 1.52218
R3806 VGND VGND.n313 1.52218
R3807 VGND.n128 VGND.n127 1.50673
R3808 VGND.n7566 VGND.n7565 1.50646
R3809 VGND.n4165 VGND.n4164 1.50646
R3810 VGND.n4260 VGND.n4259 1.50646
R3811 VGND.n5096 VGND.n5095 1.50646
R3812 VGND.n5176 VGND.n5175 1.50646
R3813 VGND.n1703 VGND.n1702 1.50646
R3814 VGND.n1870 VGND.n1869 1.50646
R3815 VGND.n2106 VGND.n2105 1.50646
R3816 VGND.n2181 VGND.n2180 1.50646
R3817 VGND.n7429 VGND.n7428 1.50646
R3818 VGND VGND.n3263 1.50638
R3819 VGND VGND.n2770 1.50638
R3820 VGND.n7645 VGND.n110 1.49961
R3821 VGND.n3273 VGND.n3262 1.49961
R3822 VGND.n3992 VGND.n3627 1.49961
R3823 VGND.n4388 VGND.n4248 1.49961
R3824 VGND.n2927 VGND.n2902 1.49961
R3825 VGND.n5830 VGND.n5829 1.49961
R3826 VGND.n1281 VGND.n1256 1.49961
R3827 VGND.n1280 VGND.n1258 1.49961
R3828 VGND.n6075 VGND.n6043 1.49961
R3829 VGND.n6074 VGND.n6045 1.49961
R3830 VGND.n6207 VGND.n6206 1.49961
R3831 VGND.n6356 VGND.n6355 1.49961
R3832 VGND.n895 VGND.n882 1.49933
R3833 VGND.n3473 VGND.n3472 1.49932
R3834 VGND.n7750 VGND.n7749 1.49932
R3835 VGND.n7785 VGND.n7783 1.49932
R3836 VGND.n3268 VGND.n3267 1.49932
R3837 VGND.n3812 VGND.n3666 1.49932
R3838 VGND.n4032 VGND.n4031 1.49932
R3839 VGND.n2910 VGND.n2909 1.49932
R3840 VGND.n2775 VGND.n2774 1.49932
R3841 VGND.n1497 VGND.n1496 1.49932
R3842 VGND.n5366 VGND.n5365 1.49932
R3843 VGND.n1263 VGND.n1262 1.49932
R3844 VGND.n6048 VGND.n6047 1.49932
R3845 VGND.n6662 VGND.n6661 1.49932
R3846 VGND.n7916 VGND.n7915 1.49932
R3847 VGND.n213 VGND.n212 1.46398
R3848 VGND.n214 VGND.n213 1.42915
R3849 VGND.n3854 VGND.n3654 1.40924
R3850 VGND.n6904 VGND.n1015 1.35467
R3851 VGND.n7514 VGND.n7513 1.35465
R3852 VGND.n7612 VGND.n7561 1.35465
R3853 VGND.n4217 VGND.n4216 1.35465
R3854 VGND.n4382 VGND.n4251 1.35465
R3855 VGND.n5158 VGND.n5157 1.35465
R3856 VGND.n2342 VGND.n2341 1.35465
R3857 VGND.n2298 VGND.n2297 1.35465
R3858 VGND.n7999 VGND.n7998 1.35465
R3859 VGND.n5564 VGND.n5556 1.35464
R3860 VGND.n7131 VGND.n7130 1.35464
R3861 VGND.n6543 VGND.n6542 1.35464
R3862 VGND.n827 VGND.n826 1.35464
R3863 VGND.n7824 VGND.n7823 1.35464
R3864 VGND.n3869 VGND.n3868 1.35464
R3865 VGND.n3070 VGND.n3069 1.35464
R3866 VGND.n4919 VGND.n4918 1.35464
R3867 VGND.n2642 VGND.n2641 1.35464
R3868 VGND.n5864 VGND.n5863 1.35464
R3869 VGND.n6262 VGND.n6261 1.35464
R3870 VGND.n611 VGND.n610 1.35464
R3871 VGND.n1551 VGND.n1550 1.35459
R3872 VGND.n7311 VGND.n7310 1.35459
R3873 VGND.n7903 VGND.n7902 1.35459
R3874 VGND.n6124 VGND.n6123 1.35457
R3875 VGND.n3532 VGND.n3531 1.35457
R3876 VGND.n3319 VGND.n3318 1.35457
R3877 VGND.n4669 VGND.n4668 1.35457
R3878 VGND.n1305 VGND.n1304 1.35457
R3879 VGND.n5040 VGND.n5039 1.35455
R3880 VGND.n1601 VGND.n1600 1.35455
R3881 VGND.n6011 VGND.n6010 1.35455
R3882 VGND.n6161 VGND.n6160 1.35455
R3883 VGND.n7269 VGND.n7268 1.35455
R3884 VGND.n492 VGND.n491 1.35455
R3885 VGND.n3567 VGND.n3566 1.35455
R3886 VGND.n3605 VGND.n3604 1.35455
R3887 VGND.n4098 VGND.n4097 1.35455
R3888 VGND.n4658 VGND.n4657 1.35455
R3889 VGND.n5453 VGND.n1459 1.35455
R3890 VGND.n6724 VGND.n6723 1.35455
R3891 VGND.n7641 VGND.n7640 1.3469
R3892 VGND VGND.n783 1.34316
R3893 VGND.n7665 VGND 1.34316
R3894 VGND.n4152 VGND 1.34316
R3895 VGND.n7618 VGND.n7615 1.29559
R3896 VGND.n3982 VGND.n3630 1.27173
R3897 VGND.n3851 VGND.n3654 1.26145
R3898 VGND.n744 VGND.n741 1.25033
R3899 VGND VGND.n5927 1.22603
R3900 VGND.n740 VGND.n739 1.1942
R3901 VGND.n7715 VGND.n7714 1.1942
R3902 VGND.n3366 VGND.n3355 1.17646
R3903 VGND.n7850 VGND.n7849 1.17646
R3904 VGND.n3920 VGND.n3634 1.17646
R3905 VGND.n4544 VGND.n4525 1.17646
R3906 VGND.n5547 VGND.n5546 1.17646
R3907 VGND.n6251 VGND.n6250 1.17646
R3908 VGND.n7162 VGND.n943 1.17646
R3909 VGND.n6577 VGND.n6556 1.17646
R3910 VGND.n4960 VGND.n2856 1.17642
R3911 VGND.n5277 VGND.n5257 1.17642
R3912 VGND.n5895 VGND.n5876 1.17642
R3913 VGND.n582 VGND.n581 1.17642
R3914 VGND.n4040 VGND 1.15795
R3915 VGND.n3805 VGND 1.15795
R3916 VGND.n4994 VGND 1.15795
R3917 VGND.n634 VGND.n404 1.14023
R3918 VGND.n7216 VGND.n7215 1.14023
R3919 VGND.n7182 VGND.n7181 1.14023
R3920 VGND.n976 VGND.n975 1.14023
R3921 VGND.n2074 VGND.n2073 1.14023
R3922 VGND.n3503 VGND.n3502 1.14023
R3923 VGND.n3401 VGND.n3400 1.14023
R3924 VGND.n806 VGND.n805 1.14023
R3925 VGND.n3294 VGND.n3293 1.14023
R3926 VGND.n78 VGND.n77 1.14023
R3927 VGND.n4067 VGND.n4066 1.14023
R3928 VGND.n3626 VGND.n3625 1.14023
R3929 VGND.n3695 VGND.n3677 1.14023
R3930 VGND.n3973 VGND.n3972 1.14023
R3931 VGND.n3930 VGND.n3929 1.14023
R3932 VGND.n4425 VGND.n4424 1.14023
R3933 VGND.n3013 VGND.n2974 1.14023
R3934 VGND.n3057 VGND.n3056 1.14023
R3935 VGND.n2782 VGND.n2768 1.14023
R3936 VGND.n4906 VGND.n4905 1.14023
R3937 VGND.n1523 VGND.n1522 1.14023
R3938 VGND.n2620 VGND.n2619 1.14023
R3939 VGND.n2685 VGND.n2684 1.14023
R3940 VGND.n5933 VGND.n5932 1.14023
R3941 VGND.n1246 VGND.n1245 1.14023
R3942 VGND.n7945 VGND.n7944 1.14023
R3943 VGND.n3352 VGND.n40 1.13896
R3944 VGND.n7854 VGND.n7853 1.13896
R3945 VGND.n3901 VGND.n3900 1.13896
R3946 VGND.n4522 VGND.n4521 1.13896
R3947 VGND.n5047 VGND.n2827 1.13896
R3948 VGND.n5639 VGND.n1388 1.13896
R3949 VGND.n6018 VGND.n1241 1.13896
R3950 VGND.n5047 VGND.n5046 1.13896
R3951 VGND.n6018 VGND.n6017 1.13896
R3952 VGND.n4521 VGND.n3076 1.13896
R3953 VGND.n3901 VGND.n3644 1.13896
R3954 VGND.n7854 VGND.n50 1.13896
R3955 VGND.n822 VGND.n40 1.13896
R3956 VGND.n4926 VGND.n4925 1.13896
R3957 VGND.n5871 VGND.n5870 1.13896
R3958 VGND.n4354 VGND.n4353 1.13896
R3959 VGND.n3130 VGND.n3129 1.13896
R3960 VGND.n7556 VGND.n7555 1.13896
R3961 VGND.n163 VGND.n162 1.13896
R3962 VGND.n5119 VGND.n2719 1.13896
R3963 VGND.n1726 VGND.n1693 1.13896
R3964 VGND.n1906 VGND.n1905 1.13896
R3965 VGND.n7025 VGND.n7024 1.13896
R3966 VGND.n2887 VGND.n2886 1.13896
R3967 VGND.n3789 VGND.n3788 1.13896
R3968 VGND.n7735 VGND.n7734 1.13896
R3969 VGND.n726 VGND.n725 1.13896
R3970 VGND.n4808 VGND.n4807 1.13896
R3971 VGND.n1388 VGND.n1387 1.13896
R3972 VGND.n5728 VGND.n5727 1.13896
R3973 VGND.n3528 VGND.n3339 1.13885
R3974 VGND.n3315 VGND.n3158 1.13885
R3975 VGND.n4092 VGND.n4091 1.13885
R3976 VGND.n4665 VGND.n4664 1.13885
R3977 VGND.n5359 VGND.n5358 1.13885
R3978 VGND.n5551 VGND.n5550 1.13885
R3979 VGND.n6718 VGND.n6717 1.13885
R3980 VGND.n7307 VGND.n7306 1.13885
R3981 VGND.n487 VGND.n36 1.13885
R3982 VGND.n7143 VGND.n7142 1.13885
R3983 VGND.n606 VGND.n605 1.13885
R3984 VGND.n2209 VGND.n1026 1.13885
R3985 VGND.n6827 VGND.n6826 1.13885
R3986 VGND.n351 VGND.n293 1.13885
R3987 VGND.n6449 VGND.n6448 1.13885
R3988 VGND.n6802 VGND.n6801 1.13717
R3989 VGND.n6549 VGND.n6548 1.13717
R3990 VGND.n2100 VGND.n2099 1.13717
R3991 VGND.n6298 VGND.n6297 1.13717
R3992 VGND.n3571 VGND.n3570 1.13717
R3993 VGND.n7516 VGND.n7515 1.13717
R3994 VGND.n716 VGND.n715 1.13717
R3995 VGND.n3609 VGND.n3608 1.13717
R3996 VGND.n7560 VGND.n7559 1.13717
R3997 VGND.n7739 VGND.n7738 1.13717
R3998 VGND.n4096 VGND.n4095 1.13717
R3999 VGND.n4219 VGND.n4218 1.13717
R4000 VGND.n3793 VGND.n3792 1.13717
R4001 VGND.n4662 VGND.n4661 1.13717
R4002 VGND.n4351 VGND.n4350 1.13717
R4003 VGND.n4693 VGND.n4692 1.13717
R4004 VGND.n5160 VGND.n5159 1.13717
R4005 VGND.n4812 VGND.n4811 1.13717
R4006 VGND.n2870 VGND.n2869 1.13717
R4007 VGND.n5256 VGND.n5255 1.13717
R4008 VGND.n2412 VGND.n2411 1.13717
R4009 VGND.n5356 VGND.n5355 1.13717
R4010 VGND.n5555 VGND.n5554 1.13717
R4011 VGND.n2340 VGND.n2339 1.13717
R4012 VGND.n2296 VGND.n2295 1.13717
R4013 VGND.n5692 VGND.n5691 1.13717
R4014 VGND.n5875 VGND.n5874 1.13717
R4015 VGND.n6722 VGND.n6721 1.13717
R4016 VGND.n7267 VGND.n7266 1.13717
R4017 VGND.n7901 VGND.n7900 1.13717
R4018 VGND.n32 VGND.n31 1.13717
R4019 VGND.n471 VGND.n470 1.13717
R4020 VGND.n6153 VGND.n1239 1.13717
R4021 VGND.n6146 VGND.n6143 1.13717
R4022 VGND.n6126 VGND.n6125 1.13717
R4023 VGND.n6159 VGND.n6158 1.13717
R4024 VGND.n5045 VGND.n5043 1.13717
R4025 VGND.n4647 VGND.n4646 1.13717
R4026 VGND.n4640 VGND.n4639 1.13717
R4027 VGND.n4667 VGND.n4666 1.13717
R4028 VGND.n4115 VGND.n4114 1.13717
R4029 VGND.n4122 VGND.n4121 1.13717
R4030 VGND.n4090 VGND.n4089 1.13717
R4031 VGND.n3590 VGND.n3589 1.13717
R4032 VGND.n3583 VGND.n3582 1.13717
R4033 VGND.n3317 VGND.n3316 1.13717
R4034 VGND.n3557 VGND.n3556 1.13717
R4035 VGND.n3550 VGND.n3549 1.13717
R4036 VGND.n3530 VGND.n3529 1.13717
R4037 VGND.n5052 VGND.n5051 1.13717
R4038 VGND.n2826 VGND.n2825 1.13717
R4039 VGND.n2842 VGND.n2841 1.13717
R4040 VGND.n1549 VGND.n1548 1.13717
R4041 VGND.n1567 VGND.n1566 1.13717
R4042 VGND.n5319 VGND.n5314 1.13717
R4043 VGND.n1599 VGND.n1598 1.13717
R4044 VGND.n6016 VGND.n6014 1.13717
R4045 VGND.n5439 VGND.n5438 1.13717
R4046 VGND.n5432 VGND.n5431 1.13717
R4047 VGND.n5361 VGND.n5360 1.13717
R4048 VGND.n6744 VGND.n6743 1.13717
R4049 VGND.n6751 VGND.n6750 1.13717
R4050 VGND.n6716 VGND.n6715 1.13717
R4051 VGND.n1303 VGND.n1302 1.13717
R4052 VGND.n6032 VGND.n6031 1.13717
R4053 VGND.n5999 VGND.n5998 1.13717
R4054 VGND.n7309 VGND.n7308 1.13717
R4055 VGND.n7304 VGND.n7301 1.13717
R4056 VGND.n7286 VGND.n7285 1.13717
R4057 VGND.n490 VGND.n489 1.13717
R4058 VGND.n7136 VGND.n7135 1.13717
R4059 VGND.n584 VGND.n583 1.13717
R4060 VGND.n424 VGND.n423 1.13717
R4061 VGND.n603 VGND.n602 1.13717
R4062 VGND.n7141 VGND.n7140 1.13717
R4063 VGND.n7148 VGND.n7147 1.13717
R4064 VGND.n6260 VGND.n6259 1.13717
R4065 VGND.n5251 VGND.n5249 1.13717
R4066 VGND.n4524 VGND.n4523 1.13717
R4067 VGND.n3091 VGND.n3088 1.13717
R4068 VGND.n4519 VGND.n4515 1.13717
R4069 VGND.n3075 VGND.n3073 1.13717
R4070 VGND.n3899 VGND.n3898 1.13717
R4071 VGND.n3907 VGND.n3906 1.13717
R4072 VGND.n3894 VGND.n3890 1.13717
R4073 VGND.n3867 VGND.n3866 1.13717
R4074 VGND.n7852 VGND.n7851 1.13717
R4075 VGND.n64 VGND.n61 1.13717
R4076 VGND.n7868 VGND.n7864 1.13717
R4077 VGND.n7822 VGND.n7821 1.13717
R4078 VGND.n3354 VGND.n3353 1.13717
R4079 VGND.n7876 VGND.n7875 1.13717
R4080 VGND.n7890 VGND.n7886 1.13717
R4081 VGND.n825 VGND.n824 1.13717
R4082 VGND.n4934 VGND.n4933 1.13717
R4083 VGND.n4941 VGND.n4940 1.13717
R4084 VGND.n4924 VGND.n4922 1.13717
R4085 VGND.n2640 VGND.n2639 1.13717
R4086 VGND.n5232 VGND.n5231 1.13717
R4087 VGND.n1347 VGND.n1346 1.13717
R4088 VGND.n1353 VGND.n1340 1.13717
R4089 VGND.n1440 VGND.n1439 1.13717
R4090 VGND.n1425 VGND.n1424 1.13717
R4091 VGND.n5549 VGND.n5548 1.13717
R4092 VGND.n1096 VGND.n1093 1.13717
R4093 VGND.n1082 VGND.n1081 1.13717
R4094 VGND.n6555 VGND.n6554 1.13717
R4095 VGND.n5869 VGND.n5867 1.13717
R4096 VGND.n6253 VGND.n6252 1.13717
R4097 VGND.n1215 VGND.n1214 1.13717
R4098 VGND.n1198 VGND.n1197 1.13717
R4099 VGND.n955 VGND.n954 1.13717
R4100 VGND.n609 VGND.n608 1.13717
R4101 VGND.n2266 VGND.n2265 1.13717
R4102 VGND.n2288 VGND.n2287 1.13717
R4103 VGND.n1692 VGND.n1690 1.13717
R4104 VGND.n2717 VGND.n2716 1.13717
R4105 VGND.n4305 VGND.n4304 1.13717
R4106 VGND.n4311 VGND.n4297 1.13717
R4107 VGND.n4357 VGND.n4356 1.13717
R4108 VGND.n3113 VGND.n3112 1.13717
R4109 VGND.n3119 VGND.n3105 1.13717
R4110 VGND.n3128 VGND.n3126 1.13717
R4111 VGND.n7539 VGND.n7538 1.13717
R4112 VGND.n7545 VGND.n7531 1.13717
R4113 VGND.n7554 VGND.n7552 1.13717
R4114 VGND.n7484 VGND.n7483 1.13717
R4115 VGND.n7491 VGND.n7490 1.13717
R4116 VGND.n161 VGND.n159 1.13717
R4117 VGND.n4332 VGND.n4331 1.13717
R4118 VGND.n4338 VGND.n4324 1.13717
R4119 VGND.n5122 VGND.n5121 1.13717
R4120 VGND.n2370 VGND.n2369 1.13717
R4121 VGND.n2376 VGND.n2362 1.13717
R4122 VGND.n1729 VGND.n1728 1.13717
R4123 VGND.n2251 VGND.n2250 1.13717
R4124 VGND.n2257 VGND.n2243 1.13717
R4125 VGND.n2212 VGND.n2211 1.13717
R4126 VGND.n2327 VGND.n2326 1.13717
R4127 VGND.n2333 VGND.n2319 1.13717
R4128 VGND.n1904 VGND.n1902 1.13717
R4129 VGND.n5206 VGND.n5205 1.13717
R4130 VGND.n2138 VGND.n2137 1.13717
R4131 VGND.n8015 VGND.n8014 1.13717
R4132 VGND.n7469 VGND.n7468 1.13717
R4133 VGND.n6815 VGND.n6812 1.13717
R4134 VGND.n6825 VGND.n6824 1.13717
R4135 VGND.n6895 VGND.n6894 1.13717
R4136 VGND.n6888 VGND.n6887 1.13717
R4137 VGND.n6984 VGND.n6983 1.13717
R4138 VGND.n691 VGND.n690 1.13717
R4139 VGND.n387 VGND.n386 1.13717
R4140 VGND.n291 VGND.n290 1.13717
R4141 VGND.n7027 VGND.n7026 1.13717
R4142 VGND.n7022 VGND.n7019 1.13717
R4143 VGND.n6328 VGND.n6325 1.13717
R4144 VGND.n2011 VGND.n2010 1.13717
R4145 VGND.n2525 VGND.n2524 1.13717
R4146 VGND.n4491 VGND.n4490 1.13717
R4147 VGND.n4497 VGND.n4235 1.13717
R4148 VGND.n2885 VGND.n2883 1.13717
R4149 VGND.n3754 VGND.n3753 1.13717
R4150 VGND.n3747 VGND.n3746 1.13717
R4151 VGND.n3787 VGND.n3785 1.13717
R4152 VGND.n7719 VGND.n7718 1.13717
R4153 VGND.n7725 VGND.n102 1.13717
R4154 VGND.n7733 VGND.n7731 1.13717
R4155 VGND.n735 VGND.n734 1.13717
R4156 VGND.n728 VGND.n271 1.13717
R4157 VGND.n724 VGND.n722 1.13717
R4158 VGND.n4792 VGND.n4791 1.13717
R4159 VGND.n4798 VGND.n4709 1.13717
R4160 VGND.n4806 VGND.n4804 1.13717
R4161 VGND.n5641 VGND.n5640 1.13717
R4162 VGND.n5658 VGND.n5655 1.13717
R4163 VGND.n2451 VGND.n2447 1.13717
R4164 VGND.n1386 VGND.n1384 1.13717
R4165 VGND.n5705 VGND.n5704 1.13717
R4166 VGND.n5725 VGND.n5724 1.13717
R4167 VGND.n5731 VGND.n5730 1.13717
R4168 VGND.n2557 VGND.n2556 1.13717
R4169 VGND.n2461 VGND.n2460 1.13717
R4170 VGND.n1676 VGND.n1675 1.13717
R4171 VGND.n2017 VGND.n2016 1.13717
R4172 VGND.n992 VGND.n991 1.13717
R4173 VGND.n354 VGND.n353 1.13717
R4174 VGND.n6341 VGND.n6338 1.13717
R4175 VGND.n6451 VGND.n6450 1.13717
R4176 VGND.n6428 VGND.n6427 1.13717
R4177 VGND.n6445 VGND.n6444 1.13717
R4178 VGND.n7305 VGND.n7304 1.1368
R4179 VGND.n470 VGND.n464 1.1368
R4180 VGND.n7147 VGND.n7144 1.1368
R4181 VGND.n4520 VGND.n4519 1.1368
R4182 VGND.n3895 VGND.n3894 1.1368
R4183 VGND.n7869 VGND.n7868 1.1368
R4184 VGND.n7891 VGND.n7890 1.1368
R4185 VGND.n4940 VGND.n4927 1.1368
R4186 VGND.n1354 VGND.n1353 1.1368
R4187 VGND.n604 VGND.n603 1.1368
R4188 VGND.n4312 VGND.n4311 1.1368
R4189 VGND.n3120 VGND.n3119 1.1368
R4190 VGND.n7546 VGND.n7545 1.1368
R4191 VGND.n7490 VGND.n7476 1.1368
R4192 VGND.n4339 VGND.n4338 1.1368
R4193 VGND.n2377 VGND.n2376 1.1368
R4194 VGND.n2258 VGND.n2257 1.1368
R4195 VGND.n2334 VGND.n2333 1.1368
R4196 VGND.n7470 VGND.n7469 1.1368
R4197 VGND.n7023 VGND.n7022 1.1368
R4198 VGND.n4498 VGND.n4497 1.1368
R4199 VGND.n3747 VGND.n3674 1.1368
R4200 VGND.n7726 VGND.n7725 1.1368
R4201 VGND.n728 VGND.n727 1.1368
R4202 VGND.n4799 VGND.n4798 1.1368
R4203 VGND.n2452 VGND.n2451 1.1368
R4204 VGND.n5726 VGND.n5725 1.1368
R4205 VGND.n292 VGND.n291 1.1368
R4206 VGND.n4663 VGND.n4662 1.13669
R4207 VGND.n4646 VGND.n2954 1.13669
R4208 VGND.n4095 VGND.n4093 1.13669
R4209 VGND.n4115 VGND.n3613 1.13669
R4210 VGND.n3610 VGND.n3609 1.13669
R4211 VGND.n3589 VGND.n3575 1.13669
R4212 VGND.n3572 VGND.n3571 1.13669
R4213 VGND.n3556 VGND.n3456 1.13669
R4214 VGND.n5051 VGND.n5048 1.13669
R4215 VGND.n2841 VGND.n2747 1.13669
R4216 VGND.n5357 VGND.n5356 1.13669
R4217 VGND.n5438 VGND.n5324 1.13669
R4218 VGND.n6721 VGND.n6719 1.13669
R4219 VGND.n6744 VGND.n1050 1.13669
R4220 VGND.n6033 VGND.n6032 1.13669
R4221 VGND.n5998 VGND.n1240 1.13669
R4222 VGND.n7266 VGND.n936 1.13669
R4223 VGND.n7900 VGND.n7898 1.13669
R4224 VGND.n3092 VGND.n3091 1.13669
R4225 VGND.n3906 VGND.n3903 1.13669
R4226 VGND.n65 VGND.n64 1.13669
R4227 VGND.n7875 VGND.n7872 1.13669
R4228 VGND.n2871 VGND.n2870 1.13669
R4229 VGND.n5874 VGND.n5872 1.13669
R4230 VGND.n5554 VGND.n5552 1.13669
R4231 VGND.n1441 VGND.n1440 1.13669
R4232 VGND.n6554 VGND.n6552 1.13669
R4233 VGND.n6550 VGND.n6549 1.13669
R4234 VGND.n7137 VGND.n7136 1.13669
R4235 VGND.n585 VGND.n584 1.13669
R4236 VGND.n4352 VGND.n4351 1.13669
R4237 VGND.n4220 VGND.n4219 1.13669
R4238 VGND.n7559 VGND.n7557 1.13669
R4239 VGND.n7517 VGND.n7516 1.13669
R4240 VGND.n5161 VGND.n5160 1.13669
R4241 VGND.n2339 VGND.n2337 1.13669
R4242 VGND.n6803 VGND.n6802 1.13669
R4243 VGND.n2295 VGND.n2293 1.13669
R4244 VGND.n6816 VGND.n6815 1.13669
R4245 VGND.n6888 VGND.n6828 1.13669
R4246 VGND.n4694 VGND.n4693 1.13669
R4247 VGND.n3792 VGND.n3790 1.13669
R4248 VGND.n7738 VGND.n7736 1.13669
R4249 VGND.n717 VGND.n716 1.13669
R4250 VGND.n4811 VGND.n4809 1.13669
R4251 VGND.n5659 VGND.n5658 1.13669
R4252 VGND.n5691 VGND.n1379 1.13669
R4253 VGND.n6983 VGND.n983 1.13669
R4254 VGND.n692 VGND.n691 1.13669
R4255 VGND.n6342 VGND.n6341 1.13669
R4256 VGND.n6447 VGND.n6445 1.13669
R4257 VGND VGND.n6901 1.12991
R4258 VGND.n7390 VGND.n173 1.09272
R4259 VGND.n4999 VGND.n4998 1.09272
R4260 VGND.n4727 VGND.n4716 1.09272
R4261 VGND.n7991 VGND.n10 1.09272
R4262 VGND.n1760 VGND.n1759 1.08588
R4263 VGND.n7315 VGND.n7314 1.07463
R4264 VGND.n2758 VGND.n2757 1.07463
R4265 VGND.n7755 VGND 1.02178
R4266 VGND.n3395 VGND.n3394 1.00931
R4267 VGND.n7659 VGND.n7658 1.00528
R4268 VGND.n7315 VGND.n7313 0.985115
R4269 VGND.n2758 VGND.n2756 0.985115
R4270 VGND.n5652 VGND.n5651 0.973599
R4271 VGND.n10 VGND.n9 0.892621
R4272 VGND.n173 VGND.n172 0.892621
R4273 VGND.n3972 VGND.n3971 0.877212
R4274 VGND.n7614 VGND.n113 0.853833
R4275 VGND.n4716 VGND.n4715 0.853833
R4276 VGND.n1555 VGND.n1554 0.835283
R4277 VGND.n638 VGND.n637 0.833377
R4278 VGND.n7213 VGND.n7212 0.833377
R4279 VGND.n7179 VGND.n7178 0.833377
R4280 VGND.n974 VGND.n971 0.833377
R4281 VGND.n2077 VGND.n1983 0.833377
R4282 VGND.n3508 VGND.n3507 0.833377
R4283 VGND.n3347 VGND.n848 0.833377
R4284 VGND.n804 VGND.n801 0.833377
R4285 VGND.n3298 VGND.n3297 0.833377
R4286 VGND.n76 VGND.n73 0.833377
R4287 VGND.n4072 VGND.n4071 0.833377
R4288 VGND.n3624 VGND.n3621 0.833377
R4289 VGND.n3694 VGND.n3679 0.833377
R4290 VGND.n3977 VGND.n3976 0.833377
R4291 VGND.n3934 VGND.n3933 0.833377
R4292 VGND.n4422 VGND.n4421 0.833377
R4293 VGND.n3017 VGND.n3016 0.833377
R4294 VGND.n3054 VGND.n3053 0.833377
R4295 VGND.n2785 VGND.n2784 0.833377
R4296 VGND.n4900 VGND.n4899 0.833377
R4297 VGND.n1528 VGND.n1527 0.833377
R4298 VGND.n2618 VGND.n2615 0.833377
R4299 VGND.n2690 VGND.n2689 0.833377
R4300 VGND.n5931 VGND.n5928 0.833377
R4301 VGND.n5939 VGND.n5938 0.833377
R4302 VGND.n7950 VGND.n7949 0.833377
R4303 VGND.n760 VGND.n759 0.830425
R4304 VGND.n3323 VGND.n3322 0.817521
R4305 VGND.n4023 VGND.n4022 0.817521
R4306 VGND.n5423 VGND.n5422 0.817521
R4307 VGND.n753 VGND.n181 0.798505
R4308 VGND.n7119 VGND.n7118 0.765717
R4309 VGND.n1555 VGND.n1553 0.765717
R4310 VGND.n3323 VGND.n3321 0.749436
R4311 VGND.n5423 VGND.n5421 0.749436
R4312 VGND.n4023 VGND.n4021 0.732971
R4313 VGND.n6573 VGND.n6572 0.711611
R4314 VGND.n5273 VGND.n5272 0.711611
R4315 VGND.n758 VGND.n755 0.606984
R4316 VGND.n3916 VGND.n3915 0.603867
R4317 VGND.n4903 VGND.n4902 0.570363
R4318 VGND.n4501 VGND.n4222 0.546928
R4319 VGND.n7474 VGND.n38 0.546928
R4320 VGND.n7208 VGND.n7207 0.526527
R4321 VGND.n7174 VGND.n7173 0.526527
R4322 VGND.n7086 VGND.n7085 0.526527
R4323 VGND.n2079 VGND.n2078 0.526527
R4324 VGND.n3511 VGND.n3510 0.526527
R4325 VGND.n836 VGND.n835 0.526527
R4326 VGND.n3301 VGND.n3256 0.526527
R4327 VGND.n7760 VGND.n7759 0.526527
R4328 VGND.n4075 VGND.n4074 0.526527
R4329 VGND.n3996 VGND.n3995 0.526527
R4330 VGND.n3691 VGND.n3690 0.526527
R4331 VGND.n3936 VGND.n3935 0.526527
R4332 VGND.n4417 VGND.n4416 0.526527
R4333 VGND.n3019 VGND.n3018 0.526527
R4334 VGND.n3049 VGND.n3048 0.526527
R4335 VGND.n2788 VGND.n2766 0.526527
R4336 VGND.n4895 VGND.n4894 0.526527
R4337 VGND.n2404 VGND.n2403 0.526527
R4338 VGND.n5959 VGND.n5958 0.526527
R4339 VGND.n5942 VGND.n5941 0.526527
R4340 VGND.n1487 VGND.n1486 0.526125
R4341 VGND.n20 VGND.n19 0.526125
R4342 VGND.n2614 VGND.n2613 0.525887
R4343 VGND.n3969 VGND.n3968 0.523356
R4344 VGND.n642 VGND.n639 0.519731
R4345 VGND.n5721 VGND.n5720 0.477096
R4346 VGND.n4458 VGND.n4457 0.43736
R4347 VGND.n7594 VGND.n7593 0.431476
R4348 VGND.n4479 VGND.n4478 0.393674
R4349 VGND.n7510 VGND.n7509 0.388379
R4350 VGND.n7508 VGND.n7507 0.388379
R4351 VGND.n754 VGND.n753 0.383542
R4352 VGND.n1545 VGND.n1473 0.3805
R4353 VGND.n1597 VGND.n1473 0.3805
R4354 VGND.n1566 VGND.n1473 0.3805
R4355 VGND.n5253 VGND.n5252 0.3805
R4356 VGND.n5252 VGND.n1653 0.3805
R4357 VGND.n5252 VGND.n5251 0.3805
R4358 VGND.n5208 VGND.n5207 0.3805
R4359 VGND.n5208 VGND.n1692 0.3805
R4360 VGND.n5208 VGND.n1680 0.3805
R4361 VGND.n2523 VGND.n1677 0.3805
R4362 VGND.n1677 VGND.n1676 0.3805
R4363 VGND.n2554 VGND.n1677 0.3805
R4364 VGND.n1762 VGND.n1761 0.374769
R4365 VGND.n4503 VGND.n4501 0.356928
R4366 VGND.n4503 VGND.n4502 0.356928
R4367 VGND.n7894 VGND.n38 0.356928
R4368 VGND.n7895 VGND.n7894 0.356928
R4369 VGND.n5210 VGND.n5209 0.352216
R4370 VGND.n1968 VGND.n1966 0.352216
R4371 VGND.n1243 VGND.n1242 0.351185
R4372 VGND.n5213 VGND.n5212 0.347759
R4373 VGND.n1964 VGND.n1963 0.347759
R4374 VGND.n1657 VGND.n1656 0.34771
R4375 VGND.n1961 VGND.n1960 0.34507
R4376 VGND.n5320 VGND.n5319 0.342516
R4377 VGND.n5233 VGND.n5232 0.342516
R4378 VGND.n2718 VGND.n2717 0.342516
R4379 VGND.n2460 VGND.n2456 0.342516
R4380 VGND.n6148 VGND.n6127 0.341811
R4381 VGND.n6258 VGND.n6256 0.341811
R4382 VGND.n6256 VGND.n6255 0.341811
R4383 VGND.n2102 VGND.n2101 0.341811
R4384 VGND.n6295 VGND.n1113 0.341811
R4385 VGND.n2289 VGND.n2288 0.31175
R4386 VGND.n2011 VGND.n1998 0.31175
R4387 VGND.n1216 VGND.n1215 0.311379
R4388 VGND.n1199 VGND.n1198 0.311379
R4389 VGND.n6147 VGND.n6146 0.311321
R4390 VGND.n6153 VGND.n6149 0.311321
R4391 VGND.n2265 VGND.n2262 0.311321
R4392 VGND.n6329 VGND.n6328 0.311321
R4393 VGND.n1244 VGND.n1243 0.307349
R4394 VGND.n7128 VGND.n7127 0.278761
R4395 VGND VGND.n7390 0.274365
R4396 VGND.n4727 VGND 0.274365
R4397 VGND.n411 VGND.n410 0.27284
R4398 VGND.n3067 VGND.n3066 0.27284
R4399 VGND.n5861 VGND.n5860 0.27284
R4400 VGND.n390 VGND.n389 0.269031
R4401 VGND.n4459 VGND.n4458 0.262616
R4402 VGND.n1761 VGND.n1760 0.262488
R4403 VGND.n6570 VGND.n6569 0.254468
R4404 VGND.n5271 VGND.n5270 0.254468
R4405 VGND.n4502 VGND 0.242831
R4406 VGND.n7895 VGND 0.242831
R4407 VGND.n3275 VGND.n3273 0.239569
R4408 VGND.n2928 VGND.n2927 0.239569
R4409 VGND.n6616 VGND.n6615 0.239569
R4410 VGND.n1958 VGND 0.239202
R4411 VGND.n898 VGND.n882 0.238116
R4412 VGND.n7783 VGND.n7782 0.237885
R4413 VGND.n3812 VGND.n3811 0.237885
R4414 VGND.n1654 VGND 0.237242
R4415 VGND.n4998 VGND 0.236604
R4416 VGND VGND.n7991 0.236604
R4417 VGND.n1763 VGND.n1762 0.225061
R4418 VGND.n7509 VGND.n7508 0.215988
R4419 VGND.n4788 VGND.n4787 0.204755
R4420 VGND.n6540 VGND.n6539 0.203675
R4421 VGND.n2633 VGND.n2632 0.203675
R4422 VGND.n7390 VGND 0.196835
R4423 VGND.n4998 VGND 0.196835
R4424 VGND VGND.n4727 0.196835
R4425 VGND.n7991 VGND 0.196835
R4426 VGND.n4504 VGND.n4503 0.1905
R4427 VGND.n7894 VGND.n7893 0.1905
R4428 VGND.n7896 VGND.n7895 0.1905
R4429 VGND.n4501 VGND.n4500 0.1905
R4430 VGND.n694 VGND.n38 0.1905
R4431 VGND.n3446 VGND.n3445 0.180551
R4432 VGND.n7645 VGND 0.179673
R4433 VGND.n3992 VGND 0.179673
R4434 VGND.n4388 VGND 0.179673
R4435 VGND.n5829 VGND 0.179673
R4436 VGND VGND.n1281 0.179673
R4437 VGND VGND.n1280 0.179673
R4438 VGND.n6206 VGND 0.179673
R4439 VGND VGND.n6075 0.179673
R4440 VGND VGND.n6074 0.179673
R4441 VGND.n6355 VGND 0.179673
R4442 VGND.n4687 VGND.n4686 0.179521
R4443 VGND VGND.n7916 0.178345
R4444 VGND VGND.n3473 0.177989
R4445 VGND.n7749 VGND 0.177989
R4446 VGND VGND.n3268 0.177989
R4447 VGND VGND.n4032 0.177989
R4448 VGND VGND.n2910 0.177989
R4449 VGND VGND.n2775 0.177989
R4450 VGND VGND.n1497 0.177989
R4451 VGND.n5365 VGND 0.177989
R4452 VGND.n1262 VGND 0.177989
R4453 VGND.n6047 VGND 0.177989
R4454 VGND.n6661 VGND 0.177989
R4455 VGND.n4904 VGND.n4903 0.175842
R4456 VGND.n127 VGND 0.171261
R4457 VGND.n7565 VGND 0.171212
R4458 VGND VGND.n4165 0.171212
R4459 VGND VGND.n4260 0.171212
R4460 VGND VGND.n5096 0.171212
R4461 VGND.n5175 VGND 0.171212
R4462 VGND VGND.n1703 0.171212
R4463 VGND VGND.n1870 0.171212
R4464 VGND.n2105 VGND 0.171212
R4465 VGND.n2180 VGND 0.171212
R4466 VGND.n7428 VGND 0.171212
R4467 VGND.n7613 VGND.n7612 0.165322
R4468 VGND.n7999 VGND.n7992 0.165322
R4469 VGND.n6581 VGND 0.158415
R4470 VGND.n658 VGND 0.158415
R4471 VGND.n739 VGND.n182 0.152881
R4472 VGND.n7715 VGND.n7713 0.152881
R4473 VGND.n3574 VGND.n3573 0.151488
R4474 VGND.n3612 VGND.n3611 0.151488
R4475 VGND.n2956 VGND.n2955 0.151488
R4476 VGND.n5350 VGND.n5349 0.151488
R4477 VGND.n6647 VGND.n937 0.151488
R4478 VGND.n7871 VGND.n7870 0.151488
R4479 VGND.n3646 VGND.n3645 0.151488
R4480 VGND.n3077 VGND.n2860 0.151488
R4481 VGND.n1416 VGND.n1415 0.151488
R4482 VGND.n1087 VGND.n961 0.151488
R4483 VGND.n7519 VGND.n7518 0.151488
R4484 VGND.n3093 VGND.n121 0.151488
R4485 VGND.n4341 VGND.n4340 0.151488
R4486 VGND.n2336 VGND.n2335 0.151488
R4487 VGND.n6805 VGND.n6804 0.151488
R4488 VGND.n696 VGND.n89 0.151488
R4489 VGND.n3673 VGND.n88 0.151488
R4490 VGND.n4696 VGND.n4695 0.151488
R4491 VGND.n5661 VGND.n5660 0.151488
R4492 VGND.n6446 VGND.n984 0.151488
R4493 VGND.n5163 VGND.n5162 0.151341
R4494 VGND.n6129 VGND.n6128 0.148403
R4495 VGND.n1200 VGND.n1086 0.148403
R4496 VGND.n2260 VGND.n2259 0.148403
R4497 VGND.n6332 VGND.n6331 0.148403
R4498 VGND.n6035 VGND.n6034 0.145562
R4499 VGND.n1329 VGND.n1328 0.145562
R4500 VGND.n2292 VGND.n2291 0.145562
R4501 VGND.n1996 VGND.n1995 0.145562
R4502 VGND VGND.n882 0.141328
R4503 VGND.n5323 VGND.n5322 0.141179
R4504 VGND.n5215 VGND.n5214 0.141179
R4505 VGND.n2379 VGND.n2378 0.141179
R4506 VGND.n2454 VGND.n2453 0.141179
R4507 VGND VGND.n7645 0.140863
R4508 VGND.n3273 VGND 0.140863
R4509 VGND VGND.n3992 0.140863
R4510 VGND VGND.n4388 0.140863
R4511 VGND.n2927 VGND 0.140863
R4512 VGND.n5829 VGND 0.140863
R4513 VGND.n1281 VGND 0.140863
R4514 VGND.n1280 VGND 0.140863
R4515 VGND.n6206 VGND 0.140863
R4516 VGND.n6075 VGND 0.140863
R4517 VGND.n6074 VGND 0.140863
R4518 VGND VGND.n6616 0.140863
R4519 VGND.n6355 VGND 0.140863
R4520 VGND.n3473 VGND 0.140584
R4521 VGND.n7749 VGND 0.140584
R4522 VGND.n7783 VGND 0.140584
R4523 VGND.n3268 VGND 0.140584
R4524 VGND VGND.n3812 0.140584
R4525 VGND.n4032 VGND 0.140584
R4526 VGND.n2910 VGND 0.140584
R4527 VGND.n2775 VGND 0.140584
R4528 VGND.n1497 VGND 0.140584
R4529 VGND.n5365 VGND 0.140584
R4530 VGND.n1262 VGND 0.140584
R4531 VGND.n6047 VGND 0.140584
R4532 VGND.n6661 VGND 0.140584
R4533 VGND.n7916 VGND 0.140228
R4534 VGND.n7904 VGND.n7903 0.136751
R4535 VGND.n4487 VGND.n4486 0.131558
R4536 VGND.n3566 VGND.n3446 0.127051
R4537 VGND.n741 VGND.n740 0.126617
R4538 VGND.n7714 VGND.n79 0.126617
R4539 VGND.n7642 VGND.n7641 0.126304
R4540 VGND.n4008 VGND.n4007 0.122994
R4541 VGND.n4505 VGND.n4504 0.122994
R4542 VGND.n4285 VGND.n4222 0.122994
R4543 VGND.n4500 VGND.n4499 0.122994
R4544 VGND.n190 VGND 0.120655
R4545 VGND.n785 VGND 0.120655
R4546 VGND.n7667 VGND 0.120655
R4547 VGND.n3842 VGND 0.120655
R4548 VGND.n2083 VGND 0.120655
R4549 VGND.n6493 VGND 0.120655
R4550 VGND.n6519 VGND 0.120655
R4551 VGND.n6520 VGND 0.120655
R4552 VGND.n131 VGND.n130 0.120292
R4553 VGND.n132 VGND.n131 0.120292
R4554 VGND.n136 VGND.n135 0.120292
R4555 VGND.n137 VGND.n136 0.120292
R4556 VGND.n142 VGND.n141 0.120292
R4557 VGND.n7394 VGND.n7392 0.120292
R4558 VGND.n7389 VGND.n7387 0.120292
R4559 VGND.n7387 VGND.n7385 0.120292
R4560 VGND.n7385 VGND.n7383 0.120292
R4561 VGND.n7383 VGND.n7381 0.120292
R4562 VGND.n7381 VGND.n7378 0.120292
R4563 VGND.n7378 VGND.n7377 0.120292
R4564 VGND.n7377 VGND.n7376 0.120292
R4565 VGND.n194 VGND.n193 0.120292
R4566 VGND.n195 VGND.n194 0.120292
R4567 VGND.n196 VGND.n195 0.120292
R4568 VGND.n201 VGND.n199 0.120292
R4569 VGND.n203 VGND.n201 0.120292
R4570 VGND.n205 VGND.n203 0.120292
R4571 VGND.n208 VGND.n205 0.120292
R4572 VGND.n209 VGND.n208 0.120292
R4573 VGND.n210 VGND.n209 0.120292
R4574 VGND.n211 VGND.n210 0.120292
R4575 VGND.n216 VGND.n215 0.120292
R4576 VGND.n217 VGND.n216 0.120292
R4577 VGND.n218 VGND.n217 0.120292
R4578 VGND.n223 VGND.n221 0.120292
R4579 VGND.n225 VGND.n223 0.120292
R4580 VGND.n227 VGND.n225 0.120292
R4581 VGND.n230 VGND.n227 0.120292
R4582 VGND.n746 VGND.n745 0.120292
R4583 VGND.n747 VGND.n746 0.120292
R4584 VGND.n752 VGND.n748 0.120292
R4585 VGND.n752 VGND.n751 0.120292
R4586 VGND.n751 VGND.n750 0.120292
R4587 VGND.n750 VGND.n749 0.120292
R4588 VGND.n767 VGND.n766 0.120292
R4589 VGND.n768 VGND.n767 0.120292
R4590 VGND.n770 VGND.n768 0.120292
R4591 VGND.n772 VGND.n770 0.120292
R4592 VGND.n774 VGND.n772 0.120292
R4593 VGND.n775 VGND.n774 0.120292
R4594 VGND.n781 VGND.n780 0.120292
R4595 VGND.n782 VGND.n781 0.120292
R4596 VGND.n791 VGND.n789 0.120292
R4597 VGND.n793 VGND.n791 0.120292
R4598 VGND.n795 VGND.n793 0.120292
R4599 VGND.n797 VGND.n795 0.120292
R4600 VGND.n844 VGND.n843 0.120292
R4601 VGND.n843 VGND.n841 0.120292
R4602 VGND.n841 VGND.n839 0.120292
R4603 VGND.n839 VGND.n837 0.120292
R4604 VGND.n837 VGND.n834 0.120292
R4605 VGND.n834 VGND.n833 0.120292
R4606 VGND.n833 VGND.n832 0.120292
R4607 VGND.n829 VGND.n828 0.120292
R4608 VGND.n3376 VGND.n3375 0.120292
R4609 VGND.n3382 VGND.n3380 0.120292
R4610 VGND.n3383 VGND.n3382 0.120292
R4611 VGND.n3390 VGND.n3389 0.120292
R4612 VGND.n3391 VGND.n3390 0.120292
R4613 VGND.n3393 VGND.n3391 0.120292
R4614 VGND.n3396 VGND.n3393 0.120292
R4615 VGND.n3399 VGND.n3398 0.120292
R4616 VGND.n3406 VGND.n3404 0.120292
R4617 VGND.n3407 VGND.n3406 0.120292
R4618 VGND.n3412 VGND.n3411 0.120292
R4619 VGND.n3415 VGND.n3412 0.120292
R4620 VGND.n3416 VGND.n3415 0.120292
R4621 VGND.n3421 VGND.n3419 0.120292
R4622 VGND.n3423 VGND.n3421 0.120292
R4623 VGND.n3429 VGND.n3427 0.120292
R4624 VGND.n3430 VGND.n3429 0.120292
R4625 VGND.n3431 VGND.n3430 0.120292
R4626 VGND.n3436 VGND.n3434 0.120292
R4627 VGND.n3437 VGND.n3436 0.120292
R4628 VGND.n3443 VGND.n3441 0.120292
R4629 VGND.n3445 VGND.n3443 0.120292
R4630 VGND.n3516 VGND.n3515 0.120292
R4631 VGND.n3515 VGND.n3514 0.120292
R4632 VGND.n3514 VGND.n3512 0.120292
R4633 VGND.n3512 VGND.n3509 0.120292
R4634 VGND.n3509 VGND.n3504 0.120292
R4635 VGND.n3504 VGND.n3501 0.120292
R4636 VGND.n3498 VGND.n3497 0.120292
R4637 VGND.n3497 VGND.n3495 0.120292
R4638 VGND.n3495 VGND.n3493 0.120292
R4639 VGND.n3488 VGND.n3486 0.120292
R4640 VGND.n3485 VGND.n3482 0.120292
R4641 VGND.n3482 VGND.n3481 0.120292
R4642 VGND.n3476 VGND.n3474 0.120292
R4643 VGND.n7569 VGND.n7568 0.120292
R4644 VGND.n7570 VGND.n7569 0.120292
R4645 VGND.n7575 VGND.n7573 0.120292
R4646 VGND.n7576 VGND.n7575 0.120292
R4647 VGND.n7583 VGND.n7580 0.120292
R4648 VGND.n7620 VGND.n7619 0.120292
R4649 VGND.n7621 VGND.n7620 0.120292
R4650 VGND.n7622 VGND.n7621 0.120292
R4651 VGND.n7628 VGND.n7627 0.120292
R4652 VGND.n7629 VGND.n7628 0.120292
R4653 VGND.n7632 VGND.n7629 0.120292
R4654 VGND.n7634 VGND.n7632 0.120292
R4655 VGND.n7636 VGND.n7634 0.120292
R4656 VGND.n7638 VGND.n7636 0.120292
R4657 VGND.n7639 VGND.n7638 0.120292
R4658 VGND.n7651 VGND.n7650 0.120292
R4659 VGND.n7652 VGND.n7651 0.120292
R4660 VGND.n7655 VGND.n7654 0.120292
R4661 VGND.n7654 VGND.n7653 0.120292
R4662 VGND.n7664 VGND.n7663 0.120292
R4663 VGND.n7666 VGND.n7664 0.120292
R4664 VGND.n7671 VGND.n7670 0.120292
R4665 VGND.n7672 VGND.n7671 0.120292
R4666 VGND.n7673 VGND.n7672 0.120292
R4667 VGND.n7678 VGND.n7676 0.120292
R4668 VGND.n7680 VGND.n7678 0.120292
R4669 VGND.n7682 VGND.n7680 0.120292
R4670 VGND.n7685 VGND.n7682 0.120292
R4671 VGND.n7754 VGND.n7753 0.120292
R4672 VGND.n7756 VGND.n7754 0.120292
R4673 VGND.n7762 VGND.n7761 0.120292
R4674 VGND.n7763 VGND.n7762 0.120292
R4675 VGND.n7764 VGND.n7763 0.120292
R4676 VGND.n7769 VGND.n7767 0.120292
R4677 VGND.n7771 VGND.n7769 0.120292
R4678 VGND.n7773 VGND.n7771 0.120292
R4679 VGND.n7774 VGND.n7773 0.120292
R4680 VGND.n7780 VGND.n7778 0.120292
R4681 VGND.n7782 VGND.n7780 0.120292
R4682 VGND.n7789 VGND.n7787 0.120292
R4683 VGND.n7791 VGND.n7789 0.120292
R4684 VGND.n7792 VGND.n7791 0.120292
R4685 VGND.n7798 VGND.n7796 0.120292
R4686 VGND.n7800 VGND.n7798 0.120292
R4687 VGND.n7802 VGND.n7800 0.120292
R4688 VGND.n7804 VGND.n7802 0.120292
R4689 VGND.n7806 VGND.n7804 0.120292
R4690 VGND.n7808 VGND.n7806 0.120292
R4691 VGND.n7810 VGND.n7808 0.120292
R4692 VGND.n7813 VGND.n7810 0.120292
R4693 VGND.n7815 VGND.n7813 0.120292
R4694 VGND.n7817 VGND.n7815 0.120292
R4695 VGND.n3183 VGND.n3182 0.120292
R4696 VGND.n3189 VGND.n3188 0.120292
R4697 VGND.n3193 VGND.n3192 0.120292
R4698 VGND.n3194 VGND.n3193 0.120292
R4699 VGND.n3199 VGND.n3194 0.120292
R4700 VGND.n3249 VGND.n3248 0.120292
R4701 VGND.n3245 VGND.n3244 0.120292
R4702 VGND.n3244 VGND.n3242 0.120292
R4703 VGND.n3242 VGND.n3241 0.120292
R4704 VGND.n3238 VGND.n3237 0.120292
R4705 VGND.n3237 VGND.n3235 0.120292
R4706 VGND.n3235 VGND.n3233 0.120292
R4707 VGND.n3233 VGND.n3231 0.120292
R4708 VGND.n3231 VGND.n3228 0.120292
R4709 VGND.n3228 VGND.n3226 0.120292
R4710 VGND.n3226 VGND.n3225 0.120292
R4711 VGND.n3222 VGND.n3221 0.120292
R4712 VGND.n3221 VGND.n3219 0.120292
R4713 VGND.n3219 VGND.n3217 0.120292
R4714 VGND.n3217 VGND.n3215 0.120292
R4715 VGND.n3215 VGND.n3213 0.120292
R4716 VGND.n3213 VGND.n3211 0.120292
R4717 VGND.n3211 VGND.n3209 0.120292
R4718 VGND.n3209 VGND.n3207 0.120292
R4719 VGND.n3207 VGND.n3204 0.120292
R4720 VGND.n3204 VGND.n3162 0.120292
R4721 VGND.n3307 VGND.n3305 0.120292
R4722 VGND.n3305 VGND.n3303 0.120292
R4723 VGND.n3299 VGND.n3257 0.120292
R4724 VGND.n3258 VGND.n3257 0.120292
R4725 VGND.n3290 VGND.n3289 0.120292
R4726 VGND.n3289 VGND.n3287 0.120292
R4727 VGND.n3287 VGND.n3285 0.120292
R4728 VGND.n3285 VGND.n3283 0.120292
R4729 VGND.n3283 VGND.n3281 0.120292
R4730 VGND.n3277 VGND.n3276 0.120292
R4731 VGND.n3276 VGND.n3275 0.120292
R4732 VGND.n3271 VGND.n3270 0.120292
R4733 VGND.n3270 VGND.n3269 0.120292
R4734 VGND.n4172 VGND.n4170 0.120292
R4735 VGND.n4173 VGND.n4172 0.120292
R4736 VGND.n4174 VGND.n4173 0.120292
R4737 VGND.n4155 VGND.n4154 0.120292
R4738 VGND.n4154 VGND.n4153 0.120292
R4739 VGND.n4150 VGND.n4149 0.120292
R4740 VGND.n4149 VGND.n4148 0.120292
R4741 VGND.n4148 VGND.n3142 0.120292
R4742 VGND.n4144 VGND.n3142 0.120292
R4743 VGND.n4144 VGND.n4143 0.120292
R4744 VGND.n4143 VGND.n3144 0.120292
R4745 VGND.n4139 VGND.n3144 0.120292
R4746 VGND.n4139 VGND.n4138 0.120292
R4747 VGND.n3683 VGND.n3681 0.120292
R4748 VGND.n3687 VGND.n3681 0.120292
R4749 VGND.n3688 VGND.n3687 0.120292
R4750 VGND.n3689 VGND.n3688 0.120292
R4751 VGND.n3689 VGND.n3678 0.120292
R4752 VGND.n3696 VGND.n3678 0.120292
R4753 VGND.n3697 VGND.n3696 0.120292
R4754 VGND.n3701 VGND.n3676 0.120292
R4755 VGND.n3707 VGND.n3705 0.120292
R4756 VGND.n3709 VGND.n3707 0.120292
R4757 VGND.n3711 VGND.n3709 0.120292
R4758 VGND.n3713 VGND.n3711 0.120292
R4759 VGND.n3715 VGND.n3713 0.120292
R4760 VGND.n3717 VGND.n3715 0.120292
R4761 VGND.n3719 VGND.n3717 0.120292
R4762 VGND.n3721 VGND.n3719 0.120292
R4763 VGND.n3813 VGND.n3664 0.120292
R4764 VGND.n3817 VGND.n3664 0.120292
R4765 VGND.n3819 VGND.n3662 0.120292
R4766 VGND.n3824 VGND.n3662 0.120292
R4767 VGND.n3825 VGND.n3824 0.120292
R4768 VGND.n3830 VGND.n3660 0.120292
R4769 VGND.n3832 VGND.n3831 0.120292
R4770 VGND.n3832 VGND.n3658 0.120292
R4771 VGND.n3836 VGND.n3658 0.120292
R4772 VGND.n3837 VGND.n3836 0.120292
R4773 VGND.n3847 VGND.n3846 0.120292
R4774 VGND.n3847 VGND.n3655 0.120292
R4775 VGND.n3852 VGND.n3655 0.120292
R4776 VGND.n3853 VGND.n3653 0.120292
R4777 VGND.n3857 VGND.n3653 0.120292
R4778 VGND.n3858 VGND.n3857 0.120292
R4779 VGND.n3927 VGND.n3926 0.120292
R4780 VGND.n3938 VGND.n3937 0.120292
R4781 VGND.n3939 VGND.n3938 0.120292
R4782 VGND.n3940 VGND.n3939 0.120292
R4783 VGND.n3946 VGND.n3944 0.120292
R4784 VGND.n3948 VGND.n3946 0.120292
R4785 VGND.n3950 VGND.n3948 0.120292
R4786 VGND.n3952 VGND.n3950 0.120292
R4787 VGND.n3956 VGND.n3955 0.120292
R4788 VGND.n3957 VGND.n3956 0.120292
R4789 VGND.n3962 VGND.n3960 0.120292
R4790 VGND.n3964 VGND.n3962 0.120292
R4791 VGND.n3966 VGND.n3964 0.120292
R4792 VGND.n3967 VGND.n3966 0.120292
R4793 VGND.n3978 VGND.n3967 0.120292
R4794 VGND.n3980 VGND.n3979 0.120292
R4795 VGND.n3986 VGND.n3984 0.120292
R4796 VGND.n3987 VGND.n3986 0.120292
R4797 VGND.n3988 VGND.n3987 0.120292
R4798 VGND.n3998 VGND.n3997 0.120292
R4799 VGND.n3999 VGND.n3998 0.120292
R4800 VGND.n4000 VGND.n3999 0.120292
R4801 VGND.n4082 VGND.n4080 0.120292
R4802 VGND.n4080 VGND.n4078 0.120292
R4803 VGND.n4078 VGND.n4076 0.120292
R4804 VGND.n4076 VGND.n4073 0.120292
R4805 VGND.n4073 VGND.n4068 0.120292
R4806 VGND.n4068 VGND.n4065 0.120292
R4807 VGND.n4062 VGND.n4061 0.120292
R4808 VGND.n4061 VGND.n4059 0.120292
R4809 VGND.n4059 VGND.n4057 0.120292
R4810 VGND.n4054 VGND.n4053 0.120292
R4811 VGND.n4053 VGND.n4052 0.120292
R4812 VGND.n4052 VGND.n4049 0.120292
R4813 VGND.n4045 VGND.n4044 0.120292
R4814 VGND.n4043 VGND.n4042 0.120292
R4815 VGND.n4038 VGND.n4030 0.120292
R4816 VGND.n4033 VGND.n4030 0.120292
R4817 VGND.n4264 VGND.n4263 0.120292
R4818 VGND.n4265 VGND.n4264 0.120292
R4819 VGND.n4271 VGND.n4255 0.120292
R4820 VGND.n4394 VGND.n4392 0.120292
R4821 VGND.n4396 VGND.n4394 0.120292
R4822 VGND.n4398 VGND.n4396 0.120292
R4823 VGND.n4400 VGND.n4398 0.120292
R4824 VGND.n4402 VGND.n4400 0.120292
R4825 VGND.n4404 VGND.n4402 0.120292
R4826 VGND.n4411 VGND.n4410 0.120292
R4827 VGND.n4413 VGND.n4411 0.120292
R4828 VGND.n4415 VGND.n4413 0.120292
R4829 VGND.n4418 VGND.n4415 0.120292
R4830 VGND.n4423 VGND.n4418 0.120292
R4831 VGND.n4426 VGND.n4423 0.120292
R4832 VGND.n4427 VGND.n4426 0.120292
R4833 VGND.n4432 VGND.n4431 0.120292
R4834 VGND.n4434 VGND.n4432 0.120292
R4835 VGND.n4440 VGND.n4438 0.120292
R4836 VGND.n4442 VGND.n4440 0.120292
R4837 VGND.n4444 VGND.n4442 0.120292
R4838 VGND.n4447 VGND.n4444 0.120292
R4839 VGND.n4448 VGND.n4447 0.120292
R4840 VGND.n4449 VGND.n4448 0.120292
R4841 VGND.n4450 VGND.n4449 0.120292
R4842 VGND.n4454 VGND.n4453 0.120292
R4843 VGND.n4455 VGND.n4454 0.120292
R4844 VGND.n2981 VGND.n2980 0.120292
R4845 VGND.n2988 VGND.n2987 0.120292
R4846 VGND.n2990 VGND.n2988 0.120292
R4847 VGND.n2996 VGND.n2995 0.120292
R4848 VGND.n3001 VGND.n3000 0.120292
R4849 VGND.n3009 VGND.n3008 0.120292
R4850 VGND.n3010 VGND.n3009 0.120292
R4851 VGND.n3011 VGND.n3010 0.120292
R4852 VGND.n3021 VGND.n3020 0.120292
R4853 VGND.n3022 VGND.n3021 0.120292
R4854 VGND.n3028 VGND.n3026 0.120292
R4855 VGND.n3030 VGND.n3028 0.120292
R4856 VGND.n3032 VGND.n3030 0.120292
R4857 VGND.n3034 VGND.n3032 0.120292
R4858 VGND.n3035 VGND.n3034 0.120292
R4859 VGND.n3043 VGND.n3042 0.120292
R4860 VGND.n3045 VGND.n3043 0.120292
R4861 VGND.n3047 VGND.n3045 0.120292
R4862 VGND.n3050 VGND.n3047 0.120292
R4863 VGND.n3055 VGND.n3050 0.120292
R4864 VGND.n3058 VGND.n3055 0.120292
R4865 VGND.n3059 VGND.n3058 0.120292
R4866 VGND.n3064 VGND.n3063 0.120292
R4867 VGND.n4554 VGND.n4553 0.120292
R4868 VGND.n4554 VGND.n2965 0.120292
R4869 VGND.n2965 VGND.n2964 0.120292
R4870 VGND.n4560 VGND.n2963 0.120292
R4871 VGND.n4564 VGND.n2963 0.120292
R4872 VGND.n4566 VGND.n4565 0.120292
R4873 VGND.n4572 VGND.n2961 0.120292
R4874 VGND.n4577 VGND.n2961 0.120292
R4875 VGND.n4578 VGND.n4577 0.120292
R4876 VGND.n4583 VGND.n4582 0.120292
R4877 VGND.n4589 VGND.n4587 0.120292
R4878 VGND.n4591 VGND.n4589 0.120292
R4879 VGND.n4593 VGND.n4591 0.120292
R4880 VGND.n4595 VGND.n4593 0.120292
R4881 VGND.n4597 VGND.n4595 0.120292
R4882 VGND.n4599 VGND.n4597 0.120292
R4883 VGND.n4601 VGND.n4599 0.120292
R4884 VGND.n4603 VGND.n4601 0.120292
R4885 VGND.n4604 VGND.n4603 0.120292
R4886 VGND.n4609 VGND.n4607 0.120292
R4887 VGND.n4611 VGND.n4609 0.120292
R4888 VGND.n4613 VGND.n4611 0.120292
R4889 VGND.n4615 VGND.n4613 0.120292
R4890 VGND.n4617 VGND.n4615 0.120292
R4891 VGND.n4618 VGND.n4617 0.120292
R4892 VGND.n2943 VGND.n2942 0.120292
R4893 VGND.n2942 VGND.n2940 0.120292
R4894 VGND.n2940 VGND.n2938 0.120292
R4895 VGND.n2932 VGND.n2928 0.120292
R4896 VGND.n2925 VGND.n2923 0.120292
R4897 VGND.n2915 VGND.n2908 0.120292
R4898 VGND.n2911 VGND.n2908 0.120292
R4899 VGND.n5107 VGND.n5105 0.120292
R4900 VGND.n5109 VGND.n5107 0.120292
R4901 VGND.n5110 VGND.n5109 0.120292
R4902 VGND.n5111 VGND.n5110 0.120292
R4903 VGND.n5092 VGND.n5091 0.120292
R4904 VGND.n5091 VGND.n5089 0.120292
R4905 VGND.n5089 VGND.n5087 0.120292
R4906 VGND.n5083 VGND.n5082 0.120292
R4907 VGND.n5082 VGND.n5081 0.120292
R4908 VGND.n5077 VGND.n5076 0.120292
R4909 VGND.n5076 VGND.n5075 0.120292
R4910 VGND.n5075 VGND.n5073 0.120292
R4911 VGND.n5073 VGND.n5071 0.120292
R4912 VGND.n5071 VGND.n5069 0.120292
R4913 VGND.n4723 VGND.n4722 0.120292
R4914 VGND.n4724 VGND.n4723 0.120292
R4915 VGND.n4726 VGND.n4724 0.120292
R4916 VGND.n4733 VGND.n4731 0.120292
R4917 VGND.n4735 VGND.n4733 0.120292
R4918 VGND.n4738 VGND.n4735 0.120292
R4919 VGND.n4740 VGND.n4738 0.120292
R4920 VGND.n4741 VGND.n4740 0.120292
R4921 VGND.n4742 VGND.n4741 0.120292
R4922 VGND.n4747 VGND.n4745 0.120292
R4923 VGND.n4749 VGND.n4747 0.120292
R4924 VGND.n4751 VGND.n4749 0.120292
R4925 VGND.n4752 VGND.n4751 0.120292
R4926 VGND.n4830 VGND.n4829 0.120292
R4927 VGND.n4832 VGND.n4830 0.120292
R4928 VGND.n4834 VGND.n4832 0.120292
R4929 VGND.n4835 VGND.n4834 0.120292
R4930 VGND.n4840 VGND.n4838 0.120292
R4931 VGND.n4842 VGND.n4840 0.120292
R4932 VGND.n4843 VGND.n4842 0.120292
R4933 VGND.n4848 VGND.n4846 0.120292
R4934 VGND.n4850 VGND.n4848 0.120292
R4935 VGND.n4852 VGND.n4850 0.120292
R4936 VGND.n4854 VGND.n4852 0.120292
R4937 VGND.n4856 VGND.n4854 0.120292
R4938 VGND.n4858 VGND.n4856 0.120292
R4939 VGND.n4860 VGND.n4858 0.120292
R4940 VGND.n4862 VGND.n4860 0.120292
R4941 VGND.n4864 VGND.n4862 0.120292
R4942 VGND.n4866 VGND.n4864 0.120292
R4943 VGND.n4867 VGND.n4866 0.120292
R4944 VGND.n4872 VGND.n4870 0.120292
R4945 VGND.n4880 VGND.n4879 0.120292
R4946 VGND.n4884 VGND.n4883 0.120292
R4947 VGND.n4889 VGND.n4887 0.120292
R4948 VGND.n4891 VGND.n4889 0.120292
R4949 VGND.n4893 VGND.n4891 0.120292
R4950 VGND.n4896 VGND.n4893 0.120292
R4951 VGND.n4901 VGND.n4896 0.120292
R4952 VGND.n4907 VGND.n4901 0.120292
R4953 VGND.n4970 VGND.n4969 0.120292
R4954 VGND.n4972 VGND.n4970 0.120292
R4955 VGND.n4974 VGND.n4972 0.120292
R4956 VGND.n4975 VGND.n4974 0.120292
R4957 VGND.n4977 VGND.n4976 0.120292
R4958 VGND.n4984 VGND.n4983 0.120292
R4959 VGND.n4986 VGND.n4984 0.120292
R4960 VGND.n4988 VGND.n4986 0.120292
R4961 VGND.n4990 VGND.n4988 0.120292
R4962 VGND.n4997 VGND.n4996 0.120292
R4963 VGND.n5005 VGND.n5003 0.120292
R4964 VGND.n5006 VGND.n5005 0.120292
R4965 VGND.n5010 VGND.n5009 0.120292
R4966 VGND.n5015 VGND.n5013 0.120292
R4967 VGND.n5017 VGND.n5015 0.120292
R4968 VGND.n5019 VGND.n5017 0.120292
R4969 VGND.n5021 VGND.n5019 0.120292
R4970 VGND.n5023 VGND.n5021 0.120292
R4971 VGND.n5025 VGND.n5023 0.120292
R4972 VGND.n5027 VGND.n5025 0.120292
R4973 VGND.n5030 VGND.n5027 0.120292
R4974 VGND.n5032 VGND.n5030 0.120292
R4975 VGND.n5033 VGND.n5032 0.120292
R4976 VGND.n5034 VGND.n5033 0.120292
R4977 VGND.n2818 VGND.n2816 0.120292
R4978 VGND.n2816 VGND.n2814 0.120292
R4979 VGND.n2814 VGND.n2811 0.120292
R4980 VGND.n2808 VGND.n2807 0.120292
R4981 VGND.n2807 VGND.n2806 0.120292
R4982 VGND.n2806 VGND.n2804 0.120292
R4983 VGND.n2804 VGND.n2802 0.120292
R4984 VGND.n2797 VGND.n2796 0.120292
R4985 VGND.n2793 VGND.n2792 0.120292
R4986 VGND.n2792 VGND.n2791 0.120292
R4987 VGND.n2791 VGND.n2765 0.120292
R4988 VGND.n2787 VGND.n2765 0.120292
R4989 VGND.n2787 VGND.n2786 0.120292
R4990 VGND.n2786 VGND.n2767 0.120292
R4991 VGND.n2780 VGND.n2767 0.120292
R4992 VGND.n2778 VGND.n2777 0.120292
R4993 VGND.n2777 VGND.n2776 0.120292
R4994 VGND.n5179 VGND.n5174 0.120292
R4995 VGND.n5180 VGND.n5179 0.120292
R4996 VGND.n5184 VGND.n5183 0.120292
R4997 VGND.n5185 VGND.n5184 0.120292
R4998 VGND.n5190 VGND.n5189 0.120292
R4999 VGND.n2693 VGND.n2692 0.120292
R5000 VGND.n2692 VGND.n2691 0.120292
R5001 VGND.n2691 VGND.n2686 0.120292
R5002 VGND.n2686 VGND.n2683 0.120292
R5003 VGND.n2679 VGND.n2678 0.120292
R5004 VGND.n2678 VGND.n2677 0.120292
R5005 VGND.n2677 VGND.n2675 0.120292
R5006 VGND.n2675 VGND.n2673 0.120292
R5007 VGND.n2673 VGND.n2671 0.120292
R5008 VGND.n2671 VGND.n2669 0.120292
R5009 VGND.n2465 VGND.n2464 0.120292
R5010 VGND.n2472 VGND.n2470 0.120292
R5011 VGND.n2474 VGND.n2472 0.120292
R5012 VGND.n2476 VGND.n2474 0.120292
R5013 VGND.n2478 VGND.n2476 0.120292
R5014 VGND.n2480 VGND.n2478 0.120292
R5015 VGND.n2482 VGND.n2480 0.120292
R5016 VGND.n2484 VGND.n2482 0.120292
R5017 VGND.n2487 VGND.n2484 0.120292
R5018 VGND.n2489 VGND.n2487 0.120292
R5019 VGND.n2490 VGND.n2489 0.120292
R5020 VGND.n2491 VGND.n2490 0.120292
R5021 VGND.n2496 VGND.n2494 0.120292
R5022 VGND.n2497 VGND.n2496 0.120292
R5023 VGND.n2502 VGND.n2500 0.120292
R5024 VGND.n2504 VGND.n2502 0.120292
R5025 VGND.n2505 VGND.n2504 0.120292
R5026 VGND.n2510 VGND.n2508 0.120292
R5027 VGND.n2573 VGND.n2571 0.120292
R5028 VGND.n2574 VGND.n2573 0.120292
R5029 VGND.n2578 VGND.n2577 0.120292
R5030 VGND.n2583 VGND.n2581 0.120292
R5031 VGND.n2585 VGND.n2583 0.120292
R5032 VGND.n2587 VGND.n2585 0.120292
R5033 VGND.n2588 VGND.n2587 0.120292
R5034 VGND.n2593 VGND.n2591 0.120292
R5035 VGND.n2595 VGND.n2593 0.120292
R5036 VGND.n2597 VGND.n2595 0.120292
R5037 VGND.n2599 VGND.n2597 0.120292
R5038 VGND.n2601 VGND.n2599 0.120292
R5039 VGND.n2602 VGND.n2601 0.120292
R5040 VGND.n2608 VGND.n2606 0.120292
R5041 VGND.n2610 VGND.n2608 0.120292
R5042 VGND.n2611 VGND.n2610 0.120292
R5043 VGND.n2612 VGND.n2611 0.120292
R5044 VGND.n2621 VGND.n2424 0.120292
R5045 VGND.n2660 VGND.n2659 0.120292
R5046 VGND.n2659 VGND.n2657 0.120292
R5047 VGND.n2657 VGND.n2656 0.120292
R5048 VGND.n2653 VGND.n2652 0.120292
R5049 VGND.n2652 VGND.n2651 0.120292
R5050 VGND.n2647 VGND.n2646 0.120292
R5051 VGND.n2646 VGND.n2644 0.120292
R5052 VGND.n5288 VGND.n5287 0.120292
R5053 VGND.n5294 VGND.n5292 0.120292
R5054 VGND.n5296 VGND.n5294 0.120292
R5055 VGND.n5298 VGND.n5296 0.120292
R5056 VGND.n5299 VGND.n5298 0.120292
R5057 VGND.n5303 VGND.n5302 0.120292
R5058 VGND.n1646 VGND.n1645 0.120292
R5059 VGND.n1645 VGND.n1643 0.120292
R5060 VGND.n1638 VGND.n1636 0.120292
R5061 VGND.n1632 VGND.n1631 0.120292
R5062 VGND.n1631 VGND.n1629 0.120292
R5063 VGND.n1625 VGND.n1624 0.120292
R5064 VGND.n1624 VGND.n1622 0.120292
R5065 VGND.n1622 VGND.n1620 0.120292
R5066 VGND.n1620 VGND.n1618 0.120292
R5067 VGND.n1614 VGND.n1613 0.120292
R5068 VGND.n1611 VGND.n1609 0.120292
R5069 VGND.n1609 VGND.n1607 0.120292
R5070 VGND.n1607 VGND.n1605 0.120292
R5071 VGND.n1605 VGND.n1603 0.120292
R5072 VGND.n1536 VGND.n1535 0.120292
R5073 VGND.n1535 VGND.n1534 0.120292
R5074 VGND.n1531 VGND.n1530 0.120292
R5075 VGND.n1530 VGND.n1529 0.120292
R5076 VGND.n1529 VGND.n1524 0.120292
R5077 VGND.n1524 VGND.n1521 0.120292
R5078 VGND.n1518 VGND.n1517 0.120292
R5079 VGND.n1517 VGND.n1515 0.120292
R5080 VGND.n1515 VGND.n1513 0.120292
R5081 VGND.n1508 VGND.n1507 0.120292
R5082 VGND.n1502 VGND.n1501 0.120292
R5083 VGND.n1501 VGND.n1500 0.120292
R5084 VGND.n1500 VGND.n1499 0.120292
R5085 VGND.n1499 VGND.n1498 0.120292
R5086 VGND.n1710 VGND.n1708 0.120292
R5087 VGND.n1712 VGND.n1710 0.120292
R5088 VGND.n1713 VGND.n1712 0.120292
R5089 VGND.n1719 VGND.n1717 0.120292
R5090 VGND.n1858 VGND.n1857 0.120292
R5091 VGND.n1854 VGND.n1853 0.120292
R5092 VGND.n1853 VGND.n1851 0.120292
R5093 VGND.n1851 VGND.n1849 0.120292
R5094 VGND.n1849 VGND.n1847 0.120292
R5095 VGND.n1847 VGND.n1845 0.120292
R5096 VGND.n1842 VGND.n1841 0.120292
R5097 VGND.n1837 VGND.n1836 0.120292
R5098 VGND.n1836 VGND.n1834 0.120292
R5099 VGND.n1826 VGND.n1825 0.120292
R5100 VGND.n1825 VGND.n1824 0.120292
R5101 VGND.n1823 VGND.n1821 0.120292
R5102 VGND.n1821 VGND.n1819 0.120292
R5103 VGND.n1819 VGND.n1818 0.120292
R5104 VGND.n1815 VGND.n1814 0.120292
R5105 VGND.n1814 VGND.n1812 0.120292
R5106 VGND.n1812 VGND.n1810 0.120292
R5107 VGND.n1810 VGND.n1808 0.120292
R5108 VGND.n1808 VGND.n1806 0.120292
R5109 VGND.n1806 VGND.n1804 0.120292
R5110 VGND.n1804 VGND.n1802 0.120292
R5111 VGND.n1802 VGND.n1800 0.120292
R5112 VGND.n1800 VGND.n1797 0.120292
R5113 VGND.n1797 VGND.n1795 0.120292
R5114 VGND.n1795 VGND.n1794 0.120292
R5115 VGND.n1786 VGND.n1785 0.120292
R5116 VGND.n5627 VGND.n5626 0.120292
R5117 VGND.n5626 VGND.n5624 0.120292
R5118 VGND.n5621 VGND.n5620 0.120292
R5119 VGND.n5620 VGND.n5618 0.120292
R5120 VGND.n5618 VGND.n5616 0.120292
R5121 VGND.n5616 VGND.n5614 0.120292
R5122 VGND.n5610 VGND.n5609 0.120292
R5123 VGND.n5605 VGND.n5604 0.120292
R5124 VGND.n5601 VGND.n5600 0.120292
R5125 VGND.n5600 VGND.n5599 0.120292
R5126 VGND.n5596 VGND.n5595 0.120292
R5127 VGND.n5595 VGND.n5593 0.120292
R5128 VGND.n5593 VGND.n5591 0.120292
R5129 VGND.n5591 VGND.n5590 0.120292
R5130 VGND.n5580 VGND.n5579 0.120292
R5131 VGND.n5579 VGND.n5578 0.120292
R5132 VGND.n5567 VGND.n5566 0.120292
R5133 VGND.n5519 VGND.n5517 0.120292
R5134 VGND.n5514 VGND.n5513 0.120292
R5135 VGND.n5509 VGND.n5508 0.120292
R5136 VGND.n5508 VGND.n5506 0.120292
R5137 VGND.n5506 VGND.n5504 0.120292
R5138 VGND.n5498 VGND.n5496 0.120292
R5139 VGND.n5496 VGND.n5495 0.120292
R5140 VGND.n5495 VGND.n5493 0.120292
R5141 VGND.n5489 VGND.n5488 0.120292
R5142 VGND.n5488 VGND.n5486 0.120292
R5143 VGND.n5485 VGND.n5483 0.120292
R5144 VGND.n5483 VGND.n5482 0.120292
R5145 VGND.n5479 VGND.n5478 0.120292
R5146 VGND.n5478 VGND.n5476 0.120292
R5147 VGND.n5472 VGND.n5471 0.120292
R5148 VGND.n5471 VGND.n5469 0.120292
R5149 VGND.n5469 VGND.n5467 0.120292
R5150 VGND.n5467 VGND.n5465 0.120292
R5151 VGND.n5460 VGND.n5458 0.120292
R5152 VGND.n5458 VGND.n5456 0.120292
R5153 VGND.n5414 VGND.n5412 0.120292
R5154 VGND.n5412 VGND.n5410 0.120292
R5155 VGND.n5410 VGND.n5408 0.120292
R5156 VGND.n5405 VGND.n5404 0.120292
R5157 VGND.n5404 VGND.n5403 0.120292
R5158 VGND.n5403 VGND.n5401 0.120292
R5159 VGND.n5401 VGND.n5398 0.120292
R5160 VGND.n5398 VGND.n5396 0.120292
R5161 VGND.n5396 VGND.n5394 0.120292
R5162 VGND.n5394 VGND.n5392 0.120292
R5163 VGND.n5389 VGND.n5388 0.120292
R5164 VGND.n5388 VGND.n5387 0.120292
R5165 VGND.n5387 VGND.n5385 0.120292
R5166 VGND.n5385 VGND.n5383 0.120292
R5167 VGND.n5383 VGND.n5381 0.120292
R5168 VGND.n5381 VGND.n5379 0.120292
R5169 VGND.n5379 VGND.n5377 0.120292
R5170 VGND.n5377 VGND.n5374 0.120292
R5171 VGND.n5374 VGND.n5372 0.120292
R5172 VGND.n5372 VGND.n5370 0.120292
R5173 VGND.n5370 VGND.n5368 0.120292
R5174 VGND.n1881 VGND.n1880 0.120292
R5175 VGND.n1886 VGND.n1884 0.120292
R5176 VGND.n1949 VGND.n1946 0.120292
R5177 VGND.n1946 VGND.n1945 0.120292
R5178 VGND.n1945 VGND.n1942 0.120292
R5179 VGND.n1938 VGND.n1937 0.120292
R5180 VGND.n1937 VGND.n1935 0.120292
R5181 VGND.n1935 VGND.n1933 0.120292
R5182 VGND.n1930 VGND.n1929 0.120292
R5183 VGND.n1929 VGND.n1928 0.120292
R5184 VGND.n5785 VGND.n5783 0.120292
R5185 VGND.n5783 VGND.n5782 0.120292
R5186 VGND.n5779 VGND.n5778 0.120292
R5187 VGND.n5778 VGND.n5776 0.120292
R5188 VGND.n5776 VGND.n5774 0.120292
R5189 VGND.n5774 VGND.n5772 0.120292
R5190 VGND.n5772 VGND.n5770 0.120292
R5191 VGND.n5770 VGND.n5768 0.120292
R5192 VGND.n5768 VGND.n5766 0.120292
R5193 VGND.n5766 VGND.n5764 0.120292
R5194 VGND.n5764 VGND.n5761 0.120292
R5195 VGND.n5761 VGND.n5759 0.120292
R5196 VGND.n5759 VGND.n5758 0.120292
R5197 VGND.n5755 VGND.n5754 0.120292
R5198 VGND.n5754 VGND.n5752 0.120292
R5199 VGND.n5749 VGND.n5748 0.120292
R5200 VGND.n5748 VGND.n5747 0.120292
R5201 VGND.n5747 VGND.n5745 0.120292
R5202 VGND.n5744 VGND.n5742 0.120292
R5203 VGND.n5794 VGND.n5792 0.120292
R5204 VGND.n5796 VGND.n5794 0.120292
R5205 VGND.n5803 VGND.n5801 0.120292
R5206 VGND.n5805 VGND.n5803 0.120292
R5207 VGND.n5807 VGND.n5805 0.120292
R5208 VGND.n5809 VGND.n5807 0.120292
R5209 VGND.n5811 VGND.n5809 0.120292
R5210 VGND.n5813 VGND.n5811 0.120292
R5211 VGND.n5815 VGND.n5813 0.120292
R5212 VGND.n5817 VGND.n5815 0.120292
R5213 VGND.n5819 VGND.n5817 0.120292
R5214 VGND.n5820 VGND.n5819 0.120292
R5215 VGND.n5826 VGND.n5825 0.120292
R5216 VGND.n5828 VGND.n5826 0.120292
R5217 VGND VGND.n5837 0.120292
R5218 VGND.n5843 VGND.n1361 0.120292
R5219 VGND.n5850 VGND.n5848 0.120292
R5220 VGND.n5852 VGND.n5850 0.120292
R5221 VGND.n5854 VGND.n5852 0.120292
R5222 VGND.n5856 VGND.n5854 0.120292
R5223 VGND.n5908 VGND.n5907 0.120292
R5224 VGND.n5910 VGND.n5908 0.120292
R5225 VGND.n5911 VGND.n5910 0.120292
R5226 VGND.n5913 VGND.n5912 0.120292
R5227 VGND.n5920 VGND.n5919 0.120292
R5228 VGND.n5922 VGND.n5920 0.120292
R5229 VGND.n5982 VGND 0.120292
R5230 VGND.n5978 VGND.n5977 0.120292
R5231 VGND.n5977 VGND.n5975 0.120292
R5232 VGND.n5975 VGND.n5973 0.120292
R5233 VGND.n5973 VGND.n5971 0.120292
R5234 VGND.n5966 VGND.n5964 0.120292
R5235 VGND.n5964 VGND.n5962 0.120292
R5236 VGND.n5962 VGND.n5960 0.120292
R5237 VGND.n5960 VGND.n5957 0.120292
R5238 VGND.n5957 VGND.n5956 0.120292
R5239 VGND.n5956 VGND.n5955 0.120292
R5240 VGND.n5950 VGND.n5949 0.120292
R5241 VGND.n5949 VGND.n5947 0.120292
R5242 VGND.n5947 VGND.n5945 0.120292
R5243 VGND.n5945 VGND.n5943 0.120292
R5244 VGND.n5943 VGND.n5940 0.120292
R5245 VGND.n5940 VGND.n1247 0.120292
R5246 VGND.n1293 VGND.n1292 0.120292
R5247 VGND.n1289 VGND.n1288 0.120292
R5248 VGND.n1288 VGND.n1287 0.120292
R5249 VGND.n1287 VGND.n1285 0.120292
R5250 VGND.n1278 VGND.n1277 0.120292
R5251 VGND.n1272 VGND.n1269 0.120292
R5252 VGND.n1269 VGND.n1268 0.120292
R5253 VGND.n1268 VGND.n1265 0.120292
R5254 VGND.n2110 VGND.n2108 0.120292
R5255 VGND.n2112 VGND.n2110 0.120292
R5256 VGND.n2114 VGND.n2112 0.120292
R5257 VGND.n2116 VGND.n2114 0.120292
R5258 VGND.n2117 VGND.n2116 0.120292
R5259 VGND.n2122 VGND.n2120 0.120292
R5260 VGND.n2124 VGND.n2122 0.120292
R5261 VGND.n2090 VGND.n2089 0.120292
R5262 VGND.n2089 VGND.n2088 0.120292
R5263 VGND.n2088 VGND.n1978 0.120292
R5264 VGND.n2081 VGND.n1980 0.120292
R5265 VGND.n2075 VGND.n1984 0.120292
R5266 VGND.n2069 VGND.n2068 0.120292
R5267 VGND.n2065 VGND.n2064 0.120292
R5268 VGND.n2064 VGND.n2063 0.120292
R5269 VGND.n2063 VGND.n2061 0.120292
R5270 VGND.n2061 VGND.n2059 0.120292
R5271 VGND.n2059 VGND.n2057 0.120292
R5272 VGND.n2057 VGND.n2055 0.120292
R5273 VGND.n2055 VGND.n2053 0.120292
R5274 VGND.n2053 VGND.n2050 0.120292
R5275 VGND.n2050 VGND.n2048 0.120292
R5276 VGND.n2048 VGND.n2046 0.120292
R5277 VGND.n2046 VGND.n2044 0.120292
R5278 VGND.n2043 VGND.n2040 0.120292
R5279 VGND.n2040 VGND.n2038 0.120292
R5280 VGND.n2035 VGND.n2034 0.120292
R5281 VGND.n2034 VGND.n2033 0.120292
R5282 VGND.n2029 VGND.n2028 0.120292
R5283 VGND.n1130 VGND.n1128 0.120292
R5284 VGND.n1131 VGND.n1130 0.120292
R5285 VGND.n1136 VGND.n1134 0.120292
R5286 VGND.n1138 VGND.n1136 0.120292
R5287 VGND.n1140 VGND.n1138 0.120292
R5288 VGND.n1142 VGND.n1140 0.120292
R5289 VGND.n1144 VGND.n1142 0.120292
R5290 VGND.n1146 VGND.n1144 0.120292
R5291 VGND.n1148 VGND.n1146 0.120292
R5292 VGND.n1150 VGND.n1148 0.120292
R5293 VGND.n1152 VGND.n1150 0.120292
R5294 VGND.n1154 VGND.n1152 0.120292
R5295 VGND.n1156 VGND.n1154 0.120292
R5296 VGND.n1158 VGND.n1156 0.120292
R5297 VGND.n1160 VGND.n1158 0.120292
R5298 VGND.n1162 VGND.n1160 0.120292
R5299 VGND.n1164 VGND.n1162 0.120292
R5300 VGND.n1166 VGND.n1164 0.120292
R5301 VGND.n1171 VGND.n1170 0.120292
R5302 VGND.n1175 VGND.n1174 0.120292
R5303 VGND.n1176 VGND.n1175 0.120292
R5304 VGND.n6283 VGND.n6282 0.120292
R5305 VGND.n6282 VGND.n6281 0.120292
R5306 VGND.n6278 VGND.n6277 0.120292
R5307 VGND.n6277 VGND.n6275 0.120292
R5308 VGND.n6275 VGND.n6273 0.120292
R5309 VGND.n6273 VGND.n6271 0.120292
R5310 VGND.n6271 VGND.n6269 0.120292
R5311 VGND.n6269 VGND.n6267 0.120292
R5312 VGND.n6267 VGND.n6265 0.120292
R5313 VGND.n6220 VGND.n1220 0.120292
R5314 VGND.n6216 VGND.n1220 0.120292
R5315 VGND.n6216 VGND.n6215 0.120292
R5316 VGND.n6215 VGND.n6214 0.120292
R5317 VGND.n6214 VGND.n1222 0.120292
R5318 VGND.n6210 VGND.n1222 0.120292
R5319 VGND.n6210 VGND.n6209 0.120292
R5320 VGND.n6204 VGND.n1225 0.120292
R5321 VGND.n6200 VGND.n6199 0.120292
R5322 VGND.n6199 VGND.n6198 0.120292
R5323 VGND.n6198 VGND.n1227 0.120292
R5324 VGND.n6194 VGND.n1227 0.120292
R5325 VGND.n6193 VGND.n6192 0.120292
R5326 VGND.n6192 VGND.n1229 0.120292
R5327 VGND.n6187 VGND.n1229 0.120292
R5328 VGND.n6187 VGND.n6186 0.120292
R5329 VGND.n6186 VGND.n6185 0.120292
R5330 VGND.n6185 VGND.n1231 0.120292
R5331 VGND.n6181 VGND.n6180 0.120292
R5332 VGND.n6176 VGND.n6175 0.120292
R5333 VGND.n6175 VGND.n6174 0.120292
R5334 VGND.n6174 VGND.n1234 0.120292
R5335 VGND.n6170 VGND.n6169 0.120292
R5336 VGND.n6169 VGND.n6167 0.120292
R5337 VGND.n6167 VGND.n6165 0.120292
R5338 VGND.n6165 VGND.n6163 0.120292
R5339 VGND.n6083 VGND.n6082 0.120292
R5340 VGND.n6082 VGND.n6081 0.120292
R5341 VGND.n6081 VGND.n6079 0.120292
R5342 VGND.n6073 VGND.n6069 0.120292
R5343 VGND.n6069 VGND.n6068 0.120292
R5344 VGND.n6068 VGND.n6067 0.120292
R5345 VGND.n6067 VGND.n6065 0.120292
R5346 VGND.n6065 VGND.n6062 0.120292
R5347 VGND.n6062 VGND.n6060 0.120292
R5348 VGND.n6060 VGND.n6058 0.120292
R5349 VGND.n6058 VGND.n6055 0.120292
R5350 VGND.n6052 VGND.n6051 0.120292
R5351 VGND.n6051 VGND.n6050 0.120292
R5352 VGND.n6841 VGND.n6840 0.120292
R5353 VGND.n6842 VGND.n6836 0.120292
R5354 VGND.n6847 VGND.n6836 0.120292
R5355 VGND.n6848 VGND.n6847 0.120292
R5356 VGND.n6849 VGND.n6834 0.120292
R5357 VGND.n6853 VGND.n6834 0.120292
R5358 VGND.n6907 VGND.n6906 0.120292
R5359 VGND.n6912 VGND.n6911 0.120292
R5360 VGND.n6914 VGND.n6912 0.120292
R5361 VGND.n6916 VGND.n6914 0.120292
R5362 VGND.n6918 VGND.n6916 0.120292
R5363 VGND.n6920 VGND.n6918 0.120292
R5364 VGND.n6922 VGND.n6920 0.120292
R5365 VGND.n6925 VGND.n6922 0.120292
R5366 VGND.n6927 VGND.n6925 0.120292
R5367 VGND.n6929 VGND.n6927 0.120292
R5368 VGND.n6931 VGND.n6929 0.120292
R5369 VGND.n6932 VGND.n6931 0.120292
R5370 VGND.n6938 VGND.n6936 0.120292
R5371 VGND.n6940 VGND.n6938 0.120292
R5372 VGND.n6942 VGND.n6940 0.120292
R5373 VGND.n6944 VGND.n6943 0.120292
R5374 VGND.n6948 VGND.n1010 0.120292
R5375 VGND.n6949 VGND.n6948 0.120292
R5376 VGND.n6950 VGND.n6949 0.120292
R5377 VGND.n6950 VGND.n1008 0.120292
R5378 VGND.n6954 VGND.n1008 0.120292
R5379 VGND.n6955 VGND.n6954 0.120292
R5380 VGND.n6956 VGND.n6955 0.120292
R5381 VGND.n6956 VGND.n1006 0.120292
R5382 VGND.n6961 VGND.n1006 0.120292
R5383 VGND.n6962 VGND.n6961 0.120292
R5384 VGND.n6963 VGND.n6962 0.120292
R5385 VGND.n6967 VGND.n1004 0.120292
R5386 VGND.n6968 VGND.n6967 0.120292
R5387 VGND.n6974 VGND.n6972 0.120292
R5388 VGND.n7040 VGND.n7039 0.120292
R5389 VGND.n7045 VGND.n7044 0.120292
R5390 VGND.n7047 VGND.n7045 0.120292
R5391 VGND.n7049 VGND.n7047 0.120292
R5392 VGND.n7051 VGND.n7049 0.120292
R5393 VGND.n7053 VGND.n7051 0.120292
R5394 VGND.n7055 VGND.n7053 0.120292
R5395 VGND.n7058 VGND.n7055 0.120292
R5396 VGND.n7060 VGND.n7058 0.120292
R5397 VGND.n7062 VGND.n7060 0.120292
R5398 VGND.n7064 VGND.n7062 0.120292
R5399 VGND.n7065 VGND.n7064 0.120292
R5400 VGND.n7070 VGND.n7068 0.120292
R5401 VGND.n7072 VGND.n7070 0.120292
R5402 VGND.n7074 VGND.n7072 0.120292
R5403 VGND.n7080 VGND.n7078 0.120292
R5404 VGND.n7082 VGND.n7080 0.120292
R5405 VGND.n7084 VGND.n7082 0.120292
R5406 VGND.n7087 VGND.n7084 0.120292
R5407 VGND.n7088 VGND.n7087 0.120292
R5408 VGND.n7089 VGND.n7088 0.120292
R5409 VGND.n7090 VGND.n7089 0.120292
R5410 VGND.n7096 VGND.n7094 0.120292
R5411 VGND.n7097 VGND.n7096 0.120292
R5412 VGND.n7098 VGND.n7097 0.120292
R5413 VGND.n7103 VGND.n7101 0.120292
R5414 VGND.n7105 VGND.n7103 0.120292
R5415 VGND.n7107 VGND.n7105 0.120292
R5416 VGND.n7109 VGND.n7107 0.120292
R5417 VGND.n7110 VGND.n7109 0.120292
R5418 VGND.n7172 VGND.n7170 0.120292
R5419 VGND.n7175 VGND.n7172 0.120292
R5420 VGND.n7180 VGND.n7175 0.120292
R5421 VGND.n7183 VGND.n7180 0.120292
R5422 VGND.n7184 VGND.n7183 0.120292
R5423 VGND.n7189 VGND.n7187 0.120292
R5424 VGND.n7191 VGND.n7189 0.120292
R5425 VGND.n7193 VGND.n7191 0.120292
R5426 VGND.n7195 VGND.n7193 0.120292
R5427 VGND.n7196 VGND.n7195 0.120292
R5428 VGND.n7202 VGND.n7201 0.120292
R5429 VGND.n7204 VGND.n7202 0.120292
R5430 VGND.n7206 VGND.n7204 0.120292
R5431 VGND.n7209 VGND.n7206 0.120292
R5432 VGND.n7214 VGND.n7209 0.120292
R5433 VGND.n7217 VGND.n7214 0.120292
R5434 VGND.n7218 VGND.n7217 0.120292
R5435 VGND.n7223 VGND.n7222 0.120292
R5436 VGND.n7225 VGND.n7223 0.120292
R5437 VGND.n7227 VGND.n7225 0.120292
R5438 VGND.n7229 VGND.n7227 0.120292
R5439 VGND.n7231 VGND.n7229 0.120292
R5440 VGND.n7233 VGND.n7231 0.120292
R5441 VGND.n7236 VGND.n7233 0.120292
R5442 VGND.n7238 VGND.n7236 0.120292
R5443 VGND.n7240 VGND.n7238 0.120292
R5444 VGND.n7242 VGND.n7240 0.120292
R5445 VGND.n7243 VGND.n7242 0.120292
R5446 VGND.n7248 VGND.n7246 0.120292
R5447 VGND.n7250 VGND.n7248 0.120292
R5448 VGND.n7251 VGND.n7250 0.120292
R5449 VGND.n7257 VGND.n7254 0.120292
R5450 VGND.n930 VGND.n928 0.120292
R5451 VGND.n928 VGND.n926 0.120292
R5452 VGND.n926 VGND.n924 0.120292
R5453 VGND.n924 VGND.n922 0.120292
R5454 VGND.n922 VGND.n920 0.120292
R5455 VGND.n920 VGND.n918 0.120292
R5456 VGND.n918 VGND.n915 0.120292
R5457 VGND.n915 VGND.n913 0.120292
R5458 VGND.n913 VGND.n911 0.120292
R5459 VGND.n911 VGND.n909 0.120292
R5460 VGND.n905 VGND.n904 0.120292
R5461 VGND.n904 VGND.n880 0.120292
R5462 VGND.n900 VGND.n899 0.120292
R5463 VGND.n899 VGND.n898 0.120292
R5464 VGND.n893 VGND.n892 0.120292
R5465 VGND.n892 VGND.n891 0.120292
R5466 VGND.n888 VGND.n887 0.120292
R5467 VGND.n887 VGND.n886 0.120292
R5468 VGND.n2185 VGND.n2179 0.120292
R5469 VGND.n2186 VGND.n2185 0.120292
R5470 VGND.n2187 VGND.n2177 0.120292
R5471 VGND.n2191 VGND.n2177 0.120292
R5472 VGND.n2198 VGND.n2195 0.120292
R5473 VGND.n6792 VGND.n6791 0.120292
R5474 VGND.n6791 VGND.n6789 0.120292
R5475 VGND.n6789 VGND.n6787 0.120292
R5476 VGND.n6787 VGND.n6785 0.120292
R5477 VGND.n6785 VGND.n6783 0.120292
R5478 VGND.n6779 VGND.n6778 0.120292
R5479 VGND.n6778 VGND.n6776 0.120292
R5480 VGND.n6776 VGND.n6774 0.120292
R5481 VGND.n6774 VGND.n6773 0.120292
R5482 VGND.n6770 VGND.n6769 0.120292
R5483 VGND.n6360 VGND.n6358 0.120292
R5484 VGND.n6362 VGND.n6360 0.120292
R5485 VGND.n6364 VGND.n6362 0.120292
R5486 VGND.n6366 VGND.n6364 0.120292
R5487 VGND.n6369 VGND.n6366 0.120292
R5488 VGND.n6370 VGND.n6369 0.120292
R5489 VGND.n6371 VGND.n6370 0.120292
R5490 VGND.n6372 VGND.n6371 0.120292
R5491 VGND.n6376 VGND.n6375 0.120292
R5492 VGND.n6377 VGND.n6376 0.120292
R5493 VGND.n6381 VGND.n6380 0.120292
R5494 VGND.n6385 VGND.n6384 0.120292
R5495 VGND.n6390 VGND.n6388 0.120292
R5496 VGND.n6392 VGND.n6390 0.120292
R5497 VGND.n6466 VGND.n6465 0.120292
R5498 VGND.n6471 VGND.n6469 0.120292
R5499 VGND.n6473 VGND.n6471 0.120292
R5500 VGND.n6475 VGND.n6473 0.120292
R5501 VGND.n6476 VGND.n6475 0.120292
R5502 VGND.n6483 VGND.n6481 0.120292
R5503 VGND.n6485 VGND.n6483 0.120292
R5504 VGND.n6486 VGND.n6485 0.120292
R5505 VGND.n6487 VGND.n6486 0.120292
R5506 VGND.n6492 VGND.n6487 0.120292
R5507 VGND.n6498 VGND.n6497 0.120292
R5508 VGND.n6502 VGND.n6501 0.120292
R5509 VGND.n6503 VGND.n6502 0.120292
R5510 VGND.n6508 VGND.n6507 0.120292
R5511 VGND.n6509 VGND.n6508 0.120292
R5512 VGND.n6513 VGND.n6509 0.120292
R5513 VGND.n6525 VGND.n6523 0.120292
R5514 VGND.n6527 VGND.n6525 0.120292
R5515 VGND.n6529 VGND.n6527 0.120292
R5516 VGND.n6531 VGND.n6529 0.120292
R5517 VGND.n6534 VGND.n6531 0.120292
R5518 VGND.n6586 VGND.n6585 0.120292
R5519 VGND.n6588 VGND.n6586 0.120292
R5520 VGND.n6590 VGND.n6588 0.120292
R5521 VGND.n6592 VGND.n6590 0.120292
R5522 VGND.n6595 VGND.n6592 0.120292
R5523 VGND.n6597 VGND.n6595 0.120292
R5524 VGND.n6599 VGND.n6597 0.120292
R5525 VGND.n6601 VGND.n6599 0.120292
R5526 VGND.n6603 VGND.n6601 0.120292
R5527 VGND.n6608 VGND.n6606 0.120292
R5528 VGND.n6612 VGND.n6610 0.120292
R5529 VGND.n6614 VGND.n6612 0.120292
R5530 VGND.n6615 VGND.n6614 0.120292
R5531 VGND.n6622 VGND.n6620 0.120292
R5532 VGND.n6623 VGND.n6622 0.120292
R5533 VGND.n6624 VGND.n6623 0.120292
R5534 VGND.n6625 VGND.n6624 0.120292
R5535 VGND.n6630 VGND.n6628 0.120292
R5536 VGND.n6632 VGND.n6630 0.120292
R5537 VGND.n6635 VGND.n6632 0.120292
R5538 VGND.n6636 VGND.n6635 0.120292
R5539 VGND.n6637 VGND.n6636 0.120292
R5540 VGND.n6638 VGND.n6637 0.120292
R5541 VGND.n6726 VGND.n6643 0.120292
R5542 VGND.n6708 VGND.n6707 0.120292
R5543 VGND.n6707 VGND.n6705 0.120292
R5544 VGND.n6705 VGND.n6703 0.120292
R5545 VGND.n6703 VGND.n6701 0.120292
R5546 VGND.n6701 VGND.n6699 0.120292
R5547 VGND.n6699 VGND.n6697 0.120292
R5548 VGND.n6697 VGND.n6695 0.120292
R5549 VGND.n6695 VGND.n6692 0.120292
R5550 VGND.n6692 VGND.n6690 0.120292
R5551 VGND.n6690 VGND.n6688 0.120292
R5552 VGND.n6688 VGND.n6686 0.120292
R5553 VGND.n6682 VGND.n6681 0.120292
R5554 VGND.n6677 VGND.n6676 0.120292
R5555 VGND.n6676 VGND.n6675 0.120292
R5556 VGND.n6675 VGND.n6674 0.120292
R5557 VGND.n6674 VGND.n6671 0.120292
R5558 VGND.n6671 VGND.n6669 0.120292
R5559 VGND.n6669 VGND.n6667 0.120292
R5560 VGND.n6667 VGND.n6664 0.120292
R5561 VGND.n7433 VGND.n7431 0.120292
R5562 VGND.n7435 VGND.n7433 0.120292
R5563 VGND.n7437 VGND.n7435 0.120292
R5564 VGND.n7439 VGND.n7437 0.120292
R5565 VGND.n7440 VGND.n7439 0.120292
R5566 VGND.n7990 VGND.n7986 0.120292
R5567 VGND.n7986 VGND.n7985 0.120292
R5568 VGND.n7985 VGND.n7984 0.120292
R5569 VGND.n7984 VGND.n7981 0.120292
R5570 VGND.n7981 VGND.n7979 0.120292
R5571 VGND.n7979 VGND.n7977 0.120292
R5572 VGND.n7977 VGND.n7975 0.120292
R5573 VGND.n310 VGND.n309 0.120292
R5574 VGND.n311 VGND.n310 0.120292
R5575 VGND.n317 VGND.n316 0.120292
R5576 VGND.n317 VGND.n306 0.120292
R5577 VGND.n322 VGND.n306 0.120292
R5578 VGND.n324 VGND.n323 0.120292
R5579 VGND.n324 VGND.n304 0.120292
R5580 VGND.n329 VGND.n304 0.120292
R5581 VGND.n330 VGND.n329 0.120292
R5582 VGND.n331 VGND.n330 0.120292
R5583 VGND.n335 VGND.n302 0.120292
R5584 VGND.n336 VGND.n335 0.120292
R5585 VGND.n336 VGND.n300 0.120292
R5586 VGND.n340 VGND.n300 0.120292
R5587 VGND.n341 VGND.n340 0.120292
R5588 VGND.n348 VGND.n345 0.120292
R5589 VGND.n682 VGND.n398 0.120292
R5590 VGND.n678 VGND.n677 0.120292
R5591 VGND.n677 VGND.n676 0.120292
R5592 VGND.n676 VGND.n675 0.120292
R5593 VGND.n675 VGND.n673 0.120292
R5594 VGND.n673 VGND.n671 0.120292
R5595 VGND.n671 VGND.n668 0.120292
R5596 VGND.n668 VGND.n666 0.120292
R5597 VGND.n666 VGND.n663 0.120292
R5598 VGND.n663 VGND.n661 0.120292
R5599 VGND.n656 VGND.n654 0.120292
R5600 VGND.n654 VGND.n653 0.120292
R5601 VGND.n649 VGND.n648 0.120292
R5602 VGND.n648 VGND.n645 0.120292
R5603 VGND.n645 VGND.n644 0.120292
R5604 VGND.n644 VGND.n643 0.120292
R5605 VGND.n633 VGND.n405 0.120292
R5606 VGND.n633 VGND 0.120292
R5607 VGND.n631 VGND.n629 0.120292
R5608 VGND.n629 VGND.n627 0.120292
R5609 VGND.n627 VGND.n626 0.120292
R5610 VGND.n623 VGND.n622 0.120292
R5611 VGND.n622 VGND.n620 0.120292
R5612 VGND.n620 VGND.n618 0.120292
R5613 VGND.n618 VGND.n616 0.120292
R5614 VGND.n616 VGND.n615 0.120292
R5615 VGND.n548 VGND.n547 0.120292
R5616 VGND.n544 VGND.n543 0.120292
R5617 VGND.n543 VGND.n542 0.120292
R5618 VGND.n542 VGND.n438 0.120292
R5619 VGND.n538 VGND.n438 0.120292
R5620 VGND.n532 VGND.n531 0.120292
R5621 VGND.n531 VGND.n530 0.120292
R5622 VGND.n530 VGND.n441 0.120292
R5623 VGND.n525 VGND.n524 0.120292
R5624 VGND.n524 VGND.n523 0.120292
R5625 VGND.n523 VGND.n443 0.120292
R5626 VGND.n519 VGND.n443 0.120292
R5627 VGND.n519 VGND.n518 0.120292
R5628 VGND.n518 VGND.n517 0.120292
R5629 VGND.n517 VGND.n445 0.120292
R5630 VGND.n512 VGND.n445 0.120292
R5631 VGND.n512 VGND.n511 0.120292
R5632 VGND.n511 VGND.n510 0.120292
R5633 VGND.n510 VGND.n447 0.120292
R5634 VGND.n506 VGND.n505 0.120292
R5635 VGND.n505 VGND.n504 0.120292
R5636 VGND.n499 VGND.n498 0.120292
R5637 VGND.n497 VGND.n495 0.120292
R5638 VGND.n7953 VGND.n7952 0.120292
R5639 VGND.n7952 VGND.n7951 0.120292
R5640 VGND.n7951 VGND.n7946 0.120292
R5641 VGND.n7946 VGND.n7943 0.120292
R5642 VGND.n7938 VGND.n7937 0.120292
R5643 VGND.n7937 VGND.n7906 0.120292
R5644 VGND.n7932 VGND.n7931 0.120292
R5645 VGND.n7931 VGND.n7908 0.120292
R5646 VGND.n7927 VGND.n7908 0.120292
R5647 VGND.n7927 VGND.n7926 0.120292
R5648 VGND.n7912 VGND.n7911 0.120292
R5649 VGND.n7913 VGND.n7912 0.120292
R5650 VGND.n7918 VGND.n7917 0.120292
R5651 VGND VGND.n2854 0.12003
R5652 VGND.n3375 VGND.n3372 0.116385
R5653 VGND.n3926 VGND.n3923 0.116385
R5654 VGND.n5283 VGND.n5280 0.116385
R5655 VGND.n7170 VGND.n7168 0.116385
R5656 VGND.n5652 VGND.n5650 0.112781
R5657 VGND.n7584 VGND.n7583 0.111177
R5658 VGND.n1721 VGND.n1719 0.111177
R5659 VGND.n1888 VGND.n1886 0.111177
R5660 VGND.n2126 VGND.n2124 0.111177
R5661 VGND.n6859 VGND.n6857 0.111177
R5662 VGND.n2200 VGND.n2198 0.111177
R5663 VGND.n6393 VGND.n6392 0.106288
R5664 VGND.n231 VGND.n230 0.106288
R5665 VGND.n7686 VGND.n7685 0.106288
R5666 VGND.n3780 VGND.n3726 0.106288
R5667 VGND.n4757 VGND.n4756 0.106288
R5668 VGND.n2516 VGND.n2510 0.106288
R5669 VGND.n1785 VGND.n1783 0.106288
R5670 VGND.n5742 VGND.n5740 0.106288
R5671 VGND.n6987 VGND.n6974 0.106288
R5672 VGND.n357 VGND.n348 0.106288
R5673 VGND.n127 VGND 0.105074
R5674 VGND.n7513 VGND.n7394 0.105063
R5675 VGND.n4216 VGND.n4159 0.105063
R5676 VGND.n4383 VGND.n4382 0.105063
R5677 VGND.n5157 VGND.n5092 0.105063
R5678 VGND.n2342 VGND.n1858 0.105063
R5679 VGND.n2298 VGND.n1950 0.105063
R5680 VGND.n6906 VGND.n6904 0.104289
R5681 VGND.n7565 VGND 0.104136
R5682 VGND.n4165 VGND 0.104136
R5683 VGND.n4260 VGND 0.104136
R5684 VGND.n5096 VGND 0.104136
R5685 VGND.n5175 VGND 0.104136
R5686 VGND.n1703 VGND 0.104136
R5687 VGND.n1870 VGND 0.104136
R5688 VGND.n2105 VGND 0.104136
R5689 VGND.n2180 VGND 0.104136
R5690 VGND.n7428 VGND 0.104136
R5691 VGND.n7896 VGND.n37 0.103019
R5692 VGND.n7893 VGND.n7892 0.103019
R5693 VGND.n7475 VGND.n7474 0.103019
R5694 VGND.n695 VGND.n694 0.103019
R5695 VGND.n5101 VGND 0.0994583
R5696 VGND.n5605 VGND 0.0994583
R5697 VGND VGND.n5498 0.0994583
R5698 VGND.n141 VGND 0.0981562
R5699 VGND.n176 VGND 0.0981562
R5700 VGND.n193 VGND 0.0981562
R5701 VGND.n215 VGND 0.0981562
R5702 VGND.n221 VGND 0.0981562
R5703 VGND.n748 VGND 0.0981562
R5704 VGND.n780 VGND 0.0981562
R5705 VGND.n786 VGND 0.0981562
R5706 VGND.n3380 VGND 0.0981562
R5707 VGND VGND.n3477 0.0981562
R5708 VGND.n7627 VGND 0.0981562
R5709 VGND.n7644 VGND 0.0981562
R5710 VGND.n7646 VGND 0.0981562
R5711 VGND.n7670 VGND 0.0981562
R5712 VGND.n3182 VGND 0.0981562
R5713 VGND VGND.n3249 0.0981562
R5714 VGND.n3245 VGND 0.0981562
R5715 VGND.n3222 VGND 0.0981562
R5716 VGND VGND.n3271 0.0981562
R5717 VGND.n4170 VGND 0.0981562
R5718 VGND.n4179 VGND 0.0981562
R5719 VGND VGND.n4137 0.0981562
R5720 VGND.n3726 VGND 0.0981562
R5721 VGND.n3813 VGND 0.0981562
R5722 VGND VGND.n3660 0.0981562
R5723 VGND.n3859 VGND 0.0981562
R5724 VGND.n3937 VGND 0.0981562
R5725 VGND.n3944 VGND 0.0981562
R5726 VGND.n3997 VGND 0.0981562
R5727 VGND VGND.n4038 0.0981562
R5728 VGND.n4263 VGND 0.0981562
R5729 VGND VGND.n4255 0.0981562
R5730 VGND.n4273 VGND 0.0981562
R5731 VGND.n2991 VGND 0.0981562
R5732 VGND.n2995 VGND 0.0981562
R5733 VGND.n4587 VGND 0.0981562
R5734 VGND VGND.n2932 0.0981562
R5735 VGND.n2917 VGND 0.0981562
R5736 VGND VGND.n2915 0.0981562
R5737 VGND VGND.n5077 0.0981562
R5738 VGND.n4731 VGND 0.0981562
R5739 VGND.n4745 VGND 0.0981562
R5740 VGND.n4876 VGND 0.0981562
R5741 VGND.n2798 VGND 0.0981562
R5742 VGND VGND.n2778 0.0981562
R5743 VGND.n5189 VGND 0.0981562
R5744 VGND VGND.n2693 0.0981562
R5745 VGND.n2470 VGND 0.0981562
R5746 VGND.n2494 VGND 0.0981562
R5747 VGND.n2571 VGND 0.0981562
R5748 VGND.n5284 VGND 0.0981562
R5749 VGND.n5292 VGND 0.0981562
R5750 VGND.n1632 VGND 0.0981562
R5751 VGND VGND.n1502 0.0981562
R5752 VGND.n1705 VGND 0.0981562
R5753 VGND VGND.n1837 0.0981562
R5754 VGND.n1791 VGND 0.0981562
R5755 VGND VGND.n1790 0.0981562
R5756 VGND VGND.n5586 0.0981562
R5757 VGND VGND.n5570 0.0981562
R5758 VGND.n5509 VGND 0.0981562
R5759 VGND VGND.n5472 0.0981562
R5760 VGND.n5389 VGND 0.0981562
R5761 VGND.n1875 VGND 0.0981562
R5762 VGND VGND.n1938 0.0981562
R5763 VGND.n5755 VGND 0.0981562
R5764 VGND.n5837 VGND 0.0981562
R5765 VGND.n5848 VGND 0.0981562
R5766 VGND.n5924 VGND 0.0981562
R5767 VGND VGND.n1293 0.0981562
R5768 VGND VGND.n1278 0.0981562
R5769 VGND VGND.n2081 0.0981562
R5770 VGND VGND.n2043 0.0981562
R5771 VGND.n1170 VGND 0.0981562
R5772 VGND.n6181 VGND 0.0981562
R5773 VGND.n6052 VGND 0.0981562
R5774 VGND.n6840 VGND 0.0981562
R5775 VGND VGND.n1013 0.0981562
R5776 VGND VGND.n1004 0.0981562
R5777 VGND.n6972 VGND 0.0981562
R5778 VGND.n7068 VGND 0.0981562
R5779 VGND.n7246 VGND 0.0981562
R5780 VGND.n906 VGND 0.0981562
R5781 VGND VGND.n905 0.0981562
R5782 VGND.n6375 VGND 0.0981562
R5783 VGND.n6380 VGND 0.0981562
R5784 VGND.n6465 VGND 0.0981562
R5785 VGND.n6497 VGND 0.0981562
R5786 VGND.n6514 VGND 0.0981562
R5787 VGND.n6585 VGND 0.0981562
R5788 VGND.n6604 VGND 0.0981562
R5789 VGND.n6642 VGND 0.0981562
R5790 VGND.n6643 VGND 0.0981562
R5791 VGND.n6683 VGND 0.0981562
R5792 VGND VGND.n6682 0.0981562
R5793 VGND.n7444 VGND 0.0981562
R5794 VGND.n11 VGND 0.0981562
R5795 VGND.n312 VGND 0.0981562
R5796 VGND VGND.n302 0.0981562
R5797 VGND.n342 VGND 0.0981562
R5798 VGND.n345 VGND 0.0981562
R5799 VGND VGND.n657 0.0981562
R5800 VGND VGND.n656 0.0981562
R5801 VGND.n405 VGND 0.0981562
R5802 VGND.n506 VGND 0.0981562
R5803 VGND.n500 VGND 0.0981562
R5804 VGND VGND.n7938 0.0981562
R5805 VGND VGND.n7932 0.0981562
R5806 VGND.n7911 VGND 0.0981562
R5807 VGND VGND.n3488 0.0968542
R5808 VGND.n3188 VGND 0.0968542
R5809 VGND VGND.n4045 0.0968542
R5810 VGND.n4553 VGND 0.0968542
R5811 VGND.n4560 VGND 0.0968542
R5812 VGND VGND.n2925 0.0968542
R5813 VGND.n5287 VGND 0.0968542
R5814 VGND VGND.n1638 0.0968542
R5815 VGND VGND.n1614 0.0968542
R5816 VGND VGND.n1508 0.0968542
R5817 VGND VGND.n5519 0.0968542
R5818 VGND.n5489 VGND 0.0968542
R5819 VGND.n5801 VGND 0.0968542
R5820 VGND.n5907 VGND 0.0968542
R5821 VGND VGND.n5966 0.0968542
R5822 VGND VGND.n6220 0.0968542
R5823 VGND VGND.n552 0.0968542
R5824 VGND.n3862 VGND 0.0955521
R5825 VGND.n3063 VGND 0.0955521
R5826 VGND.n4582 VGND 0.0955521
R5827 VGND VGND.n2797 0.0955521
R5828 VGND.n1880 VGND 0.0955521
R5829 VGND.n5566 VGND.n5564 0.0946561
R5830 VGND.n7130 VGND.n7113 0.0946561
R5831 VGND.n6542 VGND.n6534 0.0946561
R5832 VGND.n828 VGND.n827 0.0946561
R5833 VGND.n7824 VGND.n7817 0.0946561
R5834 VGND.n3869 VGND.n3862 0.0946561
R5835 VGND.n4918 VGND.n4907 0.0946561
R5836 VGND.n2644 VGND.n2642 0.0946561
R5837 VGND.n6265 VGND.n6262 0.0946561
R5838 VGND.n5252 VGND.n5213 0.0942472
R5839 VGND.n1966 VGND.n1113 0.0942472
R5840 VGND.n5210 VGND.n1677 0.0942472
R5841 VGND.n1656 VGND.n1473 0.0940635
R5842 VGND VGND.n2024 0.0841522
R5843 VGND VGND.n785 0.0826382
R5844 VGND.n190 VGND 0.0826382
R5845 VGND.n7667 VGND 0.0826382
R5846 VGND.n7613 VGND 0.0826382
R5847 VGND VGND.n3842 0.0826382
R5848 VGND.n2083 VGND 0.0826382
R5849 VGND.n6493 VGND 0.0826382
R5850 VGND VGND.n6519 0.0826382
R5851 VGND.n6520 VGND 0.0826382
R5852 VGND.n6581 VGND 0.0826382
R5853 VGND.n658 VGND 0.0826382
R5854 VGND.n7992 VGND 0.0826382
R5855 VGND VGND.n7904 0.0826382
R5856 VGND.n2854 VGND 0.0822696
R5857 VGND.n3532 VGND.n3520 0.0772651
R5858 VGND.n3319 VGND.n3307 0.0772651
R5859 VGND.n4669 VGND.n2946 0.0772651
R5860 VGND.n1305 VGND.n1297 0.0772651
R5861 VGND.n6123 VGND.n6086 0.0772651
R5862 VGND.n1551 VGND.n1539 0.0764916
R5863 VGND.n7311 VGND.n930 0.0764916
R5864 VGND.n4960 VGND.n4959 0.0711194
R5865 VGND.n5277 VGND.n5276 0.0711194
R5866 VGND.n5895 VGND.n5894 0.0711194
R5867 VGND.n581 VGND.n580 0.0711194
R5868 VGND.n7849 VGND.n7848 0.0709266
R5869 VGND.n3920 VGND.n3919 0.0709266
R5870 VGND.n4544 VGND.n4543 0.0709266
R5871 VGND.n5546 VGND.n5545 0.0709266
R5872 VGND.n6250 VGND.n6249 0.0709266
R5873 VGND.n7162 VGND.n7161 0.0709266
R5874 VGND.n6577 VGND.n6576 0.0709266
R5875 VGND.n560 VGND.n559 0.0685851
R5876 VGND.n3604 VGND.n3162 0.0670478
R5877 VGND.n4098 VGND.n4003 0.0670478
R5878 VGND.n4657 VGND.n4621 0.0670478
R5879 VGND.n1603 VGND.n1601 0.0670478
R5880 VGND.n5456 VGND.n5453 0.0670478
R5881 VGND.n6010 VGND.n1247 0.0670478
R5882 VGND.n6163 VGND.n6161 0.0670478
R5883 VGND.n7269 VGND.n7257 0.0670478
R5884 VGND.n6725 VGND.n6724 0.0670478
R5885 VGND.n495 VGND.n492 0.0670478
R5886 VGND.n130 VGND 0.0603958
R5887 VGND.n135 VGND 0.0603958
R5888 VGND.n140 VGND 0.0603958
R5889 VGND.n142 VGND 0.0603958
R5890 VGND VGND.n7389 0.0603958
R5891 VGND.n189 VGND 0.0603958
R5892 VGND.n199 VGND 0.0603958
R5893 VGND.n745 VGND 0.0603958
R5894 VGND.n766 VGND 0.0603958
R5895 VGND.n789 VGND 0.0603958
R5896 VGND.n798 VGND 0.0603958
R5897 VGND.n799 VGND 0.0603958
R5898 VGND.n845 VGND 0.0603958
R5899 VGND VGND.n844 0.0603958
R5900 VGND.n829 VGND 0.0603958
R5901 VGND VGND.n3349 0.0603958
R5902 VGND VGND.n3348 0.0603958
R5903 VGND.n3389 VGND 0.0603958
R5904 VGND.n3397 VGND 0.0603958
R5905 VGND.n3399 VGND 0.0603958
R5906 VGND.n3404 VGND 0.0603958
R5907 VGND.n3411 VGND 0.0603958
R5908 VGND.n3419 VGND 0.0603958
R5909 VGND.n3424 VGND 0.0603958
R5910 VGND.n3427 VGND 0.0603958
R5911 VGND.n3434 VGND 0.0603958
R5912 VGND VGND.n3342 0.0603958
R5913 VGND.n3441 VGND 0.0603958
R5914 VGND VGND.n3519 0.0603958
R5915 VGND.n3516 VGND 0.0603958
R5916 VGND.n3498 VGND 0.0603958
R5917 VGND.n3490 VGND 0.0603958
R5918 VGND VGND.n3489 0.0603958
R5919 VGND.n3486 VGND 0.0603958
R5920 VGND VGND.n3485 0.0603958
R5921 VGND.n3478 VGND 0.0603958
R5922 VGND VGND.n3476 0.0603958
R5923 VGND.n7568 VGND 0.0603958
R5924 VGND.n7573 VGND 0.0603958
R5925 VGND.n7577 VGND 0.0603958
R5926 VGND.n7580 VGND 0.0603958
R5927 VGND.n7619 VGND 0.0603958
R5928 VGND.n7650 VGND 0.0603958
R5929 VGND.n7655 VGND 0.0603958
R5930 VGND.n7663 VGND 0.0603958
R5931 VGND.n7676 VGND 0.0603958
R5932 VGND.n7753 VGND 0.0603958
R5933 VGND.n7757 VGND 0.0603958
R5934 VGND.n7761 VGND 0.0603958
R5935 VGND.n7767 VGND 0.0603958
R5936 VGND.n7775 VGND 0.0603958
R5937 VGND.n7778 VGND 0.0603958
R5938 VGND.n7787 VGND 0.0603958
R5939 VGND.n7793 VGND 0.0603958
R5940 VGND.n7796 VGND 0.0603958
R5941 VGND.n3178 VGND 0.0603958
R5942 VGND VGND.n3173 0.0603958
R5943 VGND.n3184 VGND 0.0603958
R5944 VGND.n3184 VGND 0.0603958
R5945 VGND.n3187 VGND 0.0603958
R5946 VGND.n3189 VGND 0.0603958
R5947 VGND.n3192 VGND 0.0603958
R5948 VGND.n3251 VGND 0.0603958
R5949 VGND VGND.n3250 0.0603958
R5950 VGND.n3241 VGND 0.0603958
R5951 VGND.n3238 VGND 0.0603958
R5952 VGND.n3300 VGND 0.0603958
R5953 VGND VGND.n3299 0.0603958
R5954 VGND.n3290 VGND 0.0603958
R5955 VGND.n3278 VGND 0.0603958
R5956 VGND VGND.n3277 0.0603958
R5957 VGND VGND.n3272 0.0603958
R5958 VGND.n4166 VGND 0.0603958
R5959 VGND.n4167 VGND 0.0603958
R5960 VGND.n4175 VGND 0.0603958
R5961 VGND.n4175 VGND 0.0603958
R5962 VGND.n4178 VGND 0.0603958
R5963 VGND.n4159 VGND 0.0603958
R5964 VGND VGND.n4158 0.0603958
R5965 VGND.n4155 VGND 0.0603958
R5966 VGND.n4150 VGND 0.0603958
R5967 VGND.n3682 VGND 0.0603958
R5968 VGND.n3683 VGND 0.0603958
R5969 VGND VGND.n3676 0.0603958
R5970 VGND.n3702 VGND 0.0603958
R5971 VGND.n3705 VGND 0.0603958
R5972 VGND.n3722 VGND 0.0603958
R5973 VGND.n3723 VGND 0.0603958
R5974 VGND.n3803 VGND 0.0603958
R5975 VGND.n3806 VGND 0.0603958
R5976 VGND.n3807 VGND 0.0603958
R5977 VGND.n3811 VGND 0.0603958
R5978 VGND VGND.n3817 0.0603958
R5979 VGND.n3818 VGND 0.0603958
R5980 VGND.n3819 VGND 0.0603958
R5981 VGND.n3826 VGND 0.0603958
R5982 VGND VGND.n3830 0.0603958
R5983 VGND.n3831 VGND 0.0603958
R5984 VGND.n3838 VGND 0.0603958
R5985 VGND.n3843 VGND 0.0603958
R5986 VGND.n3845 VGND 0.0603958
R5987 VGND.n3846 VGND 0.0603958
R5988 VGND.n3853 VGND 0.0603958
R5989 VGND.n3941 VGND 0.0603958
R5990 VGND VGND.n3952 0.0603958
R5991 VGND.n3953 VGND 0.0603958
R5992 VGND.n3955 VGND 0.0603958
R5993 VGND.n3960 VGND 0.0603958
R5994 VGND.n3979 VGND 0.0603958
R5995 VGND.n3981 VGND 0.0603958
R5996 VGND.n3984 VGND 0.0603958
R5997 VGND.n3991 VGND 0.0603958
R5998 VGND.n3993 VGND 0.0603958
R5999 VGND.n4003 VGND 0.0603958
R6000 VGND.n4062 VGND 0.0603958
R6001 VGND.n4054 VGND 0.0603958
R6002 VGND.n4046 VGND 0.0603958
R6003 VGND.n4044 VGND 0.0603958
R6004 VGND VGND.n4043 0.0603958
R6005 VGND.n4039 VGND 0.0603958
R6006 VGND.n4266 VGND 0.0603958
R6007 VGND.n4272 VGND 0.0603958
R6008 VGND.n4273 VGND 0.0603958
R6009 VGND VGND.n4383 0.0603958
R6010 VGND.n4384 VGND 0.0603958
R6011 VGND.n4387 VGND 0.0603958
R6012 VGND.n4389 VGND 0.0603958
R6013 VGND.n4392 VGND 0.0603958
R6014 VGND.n4405 VGND 0.0603958
R6015 VGND.n4406 VGND 0.0603958
R6016 VGND.n4410 VGND 0.0603958
R6017 VGND.n4431 VGND 0.0603958
R6018 VGND.n4435 VGND 0.0603958
R6019 VGND.n4438 VGND 0.0603958
R6020 VGND.n4453 VGND 0.0603958
R6021 VGND.n2981 VGND 0.0603958
R6022 VGND.n2987 VGND 0.0603958
R6023 VGND.n2992 VGND 0.0603958
R6024 VGND.n3000 VGND 0.0603958
R6025 VGND VGND.n3001 0.0603958
R6026 VGND.n3002 VGND 0.0603958
R6027 VGND.n3008 VGND 0.0603958
R6028 VGND.n3020 VGND 0.0603958
R6029 VGND.n3023 VGND 0.0603958
R6030 VGND.n3026 VGND 0.0603958
R6031 VGND.n3038 VGND 0.0603958
R6032 VGND.n3039 VGND 0.0603958
R6033 VGND.n3042 VGND 0.0603958
R6034 VGND.n3060 VGND 0.0603958
R6035 VGND.n4552 VGND 0.0603958
R6036 VGND.n4559 VGND 0.0603958
R6037 VGND VGND.n4564 0.0603958
R6038 VGND.n4565 VGND 0.0603958
R6039 VGND.n4566 VGND 0.0603958
R6040 VGND.n4570 VGND 0.0603958
R6041 VGND.n4571 VGND 0.0603958
R6042 VGND.n4572 VGND 0.0603958
R6043 VGND.n4579 VGND 0.0603958
R6044 VGND VGND.n4583 0.0603958
R6045 VGND.n4584 VGND 0.0603958
R6046 VGND.n4607 VGND 0.0603958
R6047 VGND.n4621 VGND 0.0603958
R6048 VGND.n2943 VGND 0.0603958
R6049 VGND VGND.n2937 0.0603958
R6050 VGND.n2934 VGND 0.0603958
R6051 VGND VGND.n2933 0.0603958
R6052 VGND VGND.n2926 0.0603958
R6053 VGND.n2923 VGND 0.0603958
R6054 VGND VGND.n2922 0.0603958
R6055 VGND VGND.n2921 0.0603958
R6056 VGND VGND.n2920 0.0603958
R6057 VGND VGND.n2916 0.0603958
R6058 VGND.n2911 VGND 0.0603958
R6059 VGND.n5097 VGND 0.0603958
R6060 VGND.n5098 VGND 0.0603958
R6061 VGND.n5102 VGND 0.0603958
R6062 VGND.n5102 VGND 0.0603958
R6063 VGND.n5105 VGND 0.0603958
R6064 VGND.n5087 VGND 0.0603958
R6065 VGND.n5083 VGND 0.0603958
R6066 VGND.n5078 VGND 0.0603958
R6067 VGND.n2732 VGND 0.0603958
R6068 VGND.n4717 VGND 0.0603958
R6069 VGND.n4722 VGND 0.0603958
R6070 VGND.n4728 VGND 0.0603958
R6071 VGND.n4753 VGND 0.0603958
R6072 VGND.n4756 VGND 0.0603958
R6073 VGND.n4824 VGND 0.0603958
R6074 VGND VGND.n4824 0.0603958
R6075 VGND.n4825 VGND 0.0603958
R6076 VGND.n4829 VGND 0.0603958
R6077 VGND.n4838 VGND 0.0603958
R6078 VGND.n4846 VGND 0.0603958
R6079 VGND.n4870 VGND 0.0603958
R6080 VGND.n4873 VGND 0.0603958
R6081 VGND.n4877 VGND 0.0603958
R6082 VGND.n4879 VGND 0.0603958
R6083 VGND.n4880 VGND 0.0603958
R6084 VGND.n4883 VGND 0.0603958
R6085 VGND.n4887 VGND 0.0603958
R6086 VGND.n4969 VGND 0.0603958
R6087 VGND.n4977 VGND 0.0603958
R6088 VGND.n4983 VGND 0.0603958
R6089 VGND.n4991 VGND 0.0603958
R6090 VGND.n4992 VGND 0.0603958
R6091 VGND.n4996 VGND 0.0603958
R6092 VGND.n5003 VGND 0.0603958
R6093 VGND.n5009 VGND 0.0603958
R6094 VGND.n5013 VGND 0.0603958
R6095 VGND.n2808 VGND 0.0603958
R6096 VGND.n2796 VGND 0.0603958
R6097 VGND.n2793 VGND 0.0603958
R6098 VGND VGND.n2779 0.0603958
R6099 VGND VGND.n5174 0.0603958
R6100 VGND.n5183 VGND 0.0603958
R6101 VGND VGND.n5171 0.0603958
R6102 VGND.n5190 VGND 0.0603958
R6103 VGND.n2694 VGND 0.0603958
R6104 VGND.n2680 VGND 0.0603958
R6105 VGND.n2680 VGND 0.0603958
R6106 VGND VGND.n2679 0.0603958
R6107 VGND.n2418 VGND 0.0603958
R6108 VGND.n2464 VGND 0.0603958
R6109 VGND.n2468 VGND 0.0603958
R6110 VGND.n2500 VGND 0.0603958
R6111 VGND.n2508 VGND 0.0603958
R6112 VGND.n2568 VGND 0.0603958
R6113 VGND.n2574 VGND 0.0603958
R6114 VGND.n2577 VGND 0.0603958
R6115 VGND.n2581 VGND 0.0603958
R6116 VGND.n2591 VGND 0.0603958
R6117 VGND.n2603 VGND 0.0603958
R6118 VGND.n2606 VGND 0.0603958
R6119 VGND VGND.n2424 0.0603958
R6120 VGND.n2622 VGND 0.0603958
R6121 VGND.n2661 VGND 0.0603958
R6122 VGND VGND.n2660 0.0603958
R6123 VGND.n2653 VGND 0.0603958
R6124 VGND.n2651 VGND 0.0603958
R6125 VGND.n2648 VGND 0.0603958
R6126 VGND VGND.n2647 0.0603958
R6127 VGND VGND.n5288 0.0603958
R6128 VGND.n5289 VGND 0.0603958
R6129 VGND.n5302 VGND 0.0603958
R6130 VGND VGND.n1647 0.0603958
R6131 VGND VGND.n1646 0.0603958
R6132 VGND VGND.n1642 0.0603958
R6133 VGND.n1639 VGND 0.0603958
R6134 VGND.n1636 VGND 0.0603958
R6135 VGND VGND.n1635 0.0603958
R6136 VGND.n1626 VGND 0.0603958
R6137 VGND VGND.n1625 0.0603958
R6138 VGND.n1615 VGND 0.0603958
R6139 VGND.n1613 VGND 0.0603958
R6140 VGND VGND.n1612 0.0603958
R6141 VGND VGND.n1611 0.0603958
R6142 VGND.n1536 VGND 0.0603958
R6143 VGND.n1534 VGND 0.0603958
R6144 VGND.n1531 VGND 0.0603958
R6145 VGND.n1518 VGND 0.0603958
R6146 VGND VGND.n1512 0.0603958
R6147 VGND.n1509 VGND 0.0603958
R6148 VGND.n1507 VGND 0.0603958
R6149 VGND VGND.n1506 0.0603958
R6150 VGND.n1503 VGND 0.0603958
R6151 VGND.n1704 VGND 0.0603958
R6152 VGND.n1708 VGND 0.0603958
R6153 VGND VGND.n1713 0.0603958
R6154 VGND.n1714 VGND 0.0603958
R6155 VGND.n1717 VGND 0.0603958
R6156 VGND.n1854 VGND 0.0603958
R6157 VGND.n1842 VGND 0.0603958
R6158 VGND.n1838 VGND 0.0603958
R6159 VGND VGND.n1832 0.0603958
R6160 VGND.n1826 VGND 0.0603958
R6161 VGND VGND.n1823 0.0603958
R6162 VGND.n1815 VGND 0.0603958
R6163 VGND VGND.n1789 0.0603958
R6164 VGND.n1789 VGND 0.0603958
R6165 VGND.n1786 VGND 0.0603958
R6166 VGND VGND.n5630 0.0603958
R6167 VGND.n5627 VGND 0.0603958
R6168 VGND.n5624 VGND 0.0603958
R6169 VGND.n5621 VGND 0.0603958
R6170 VGND VGND.n5613 0.0603958
R6171 VGND.n5610 VGND 0.0603958
R6172 VGND VGND.n5608 0.0603958
R6173 VGND.n5601 VGND 0.0603958
R6174 VGND.n5596 VGND 0.0603958
R6175 VGND.n5587 VGND 0.0603958
R6176 VGND VGND.n5585 0.0603958
R6177 VGND VGND.n5584 0.0603958
R6178 VGND.n5581 VGND 0.0603958
R6179 VGND VGND.n5580 0.0603958
R6180 VGND VGND.n5577 0.0603958
R6181 VGND VGND.n5576 0.0603958
R6182 VGND.n5573 VGND 0.0603958
R6183 VGND.n5573 VGND 0.0603958
R6184 VGND VGND.n5572 0.0603958
R6185 VGND VGND.n5571 0.0603958
R6186 VGND.n5567 VGND 0.0603958
R6187 VGND.n5521 VGND 0.0603958
R6188 VGND VGND.n5520 0.0603958
R6189 VGND.n5517 VGND 0.0603958
R6190 VGND.n5514 VGND 0.0603958
R6191 VGND VGND.n5512 0.0603958
R6192 VGND.n5501 VGND 0.0603958
R6193 VGND VGND.n5500 0.0603958
R6194 VGND VGND.n5499 0.0603958
R6195 VGND VGND.n5492 0.0603958
R6196 VGND.n5486 VGND 0.0603958
R6197 VGND VGND.n5485 0.0603958
R6198 VGND.n5479 VGND 0.0603958
R6199 VGND.n5476 VGND 0.0603958
R6200 VGND.n5473 VGND 0.0603958
R6201 VGND.n5462 VGND 0.0603958
R6202 VGND.n5462 VGND 0.0603958
R6203 VGND VGND.n5461 0.0603958
R6204 VGND VGND.n5460 0.0603958
R6205 VGND.n5405 VGND 0.0603958
R6206 VGND.n1871 VGND 0.0603958
R6207 VGND.n1872 VGND 0.0603958
R6208 VGND.n1876 VGND 0.0603958
R6209 VGND VGND.n1876 0.0603958
R6210 VGND.n1877 VGND 0.0603958
R6211 VGND.n1881 VGND 0.0603958
R6212 VGND.n1884 VGND 0.0603958
R6213 VGND.n1950 VGND 0.0603958
R6214 VGND VGND.n1949 0.0603958
R6215 VGND.n1939 VGND 0.0603958
R6216 VGND.n1930 VGND 0.0603958
R6217 VGND VGND.n1925 0.0603958
R6218 VGND.n5786 VGND 0.0603958
R6219 VGND VGND.n5785 0.0603958
R6220 VGND.n5779 VGND 0.0603958
R6221 VGND.n5749 VGND 0.0603958
R6222 VGND VGND.n5744 0.0603958
R6223 VGND.n5792 VGND 0.0603958
R6224 VGND.n5797 VGND 0.0603958
R6225 VGND.n5798 VGND 0.0603958
R6226 VGND VGND.n5820 0.0603958
R6227 VGND.n5821 VGND 0.0603958
R6228 VGND.n5825 VGND 0.0603958
R6229 VGND.n5833 VGND 0.0603958
R6230 VGND.n5834 VGND 0.0603958
R6231 VGND.n5838 VGND 0.0603958
R6232 VGND VGND.n1361 0.0603958
R6233 VGND VGND.n5843 0.0603958
R6234 VGND.n5844 VGND 0.0603958
R6235 VGND.n5845 VGND 0.0603958
R6236 VGND VGND.n5856 0.0603958
R6237 VGND.n5857 VGND 0.0603958
R6238 VGND VGND.n5857 0.0603958
R6239 VGND.n5858 VGND 0.0603958
R6240 VGND.n5902 VGND 0.0603958
R6241 VGND.n5903 VGND 0.0603958
R6242 VGND VGND.n5911 0.0603958
R6243 VGND.n5913 VGND 0.0603958
R6244 VGND.n5919 VGND 0.0603958
R6245 VGND.n5923 VGND 0.0603958
R6246 VGND.n5982 VGND 0.0603958
R6247 VGND VGND.n5981 0.0603958
R6248 VGND.n5978 VGND 0.0603958
R6249 VGND.n5968 VGND 0.0603958
R6250 VGND VGND.n5967 0.0603958
R6251 VGND.n5934 VGND 0.0603958
R6252 VGND VGND.n5934 0.0603958
R6253 VGND.n5935 VGND 0.0603958
R6254 VGND.n5950 VGND 0.0603958
R6255 VGND.n1294 VGND 0.0603958
R6256 VGND.n1292 VGND 0.0603958
R6257 VGND.n1289 VGND 0.0603958
R6258 VGND.n1282 VGND 0.0603958
R6259 VGND VGND.n1279 0.0603958
R6260 VGND.n1277 VGND 0.0603958
R6261 VGND.n1274 VGND 0.0603958
R6262 VGND VGND.n1273 0.0603958
R6263 VGND VGND.n1272 0.0603958
R6264 VGND.n2108 VGND 0.0603958
R6265 VGND.n2120 VGND 0.0603958
R6266 VGND VGND.n2094 0.0603958
R6267 VGND.n2094 VGND 0.0603958
R6268 VGND VGND.n2093 0.0603958
R6269 VGND.n2090 VGND 0.0603958
R6270 VGND VGND.n2082 0.0603958
R6271 VGND VGND.n1980 0.0603958
R6272 VGND.n2076 VGND 0.0603958
R6273 VGND VGND.n2075 0.0603958
R6274 VGND.n2070 VGND 0.0603958
R6275 VGND VGND.n2069 0.0603958
R6276 VGND.n2065 VGND 0.0603958
R6277 VGND.n2035 VGND 0.0603958
R6278 VGND.n2030 VGND 0.0603958
R6279 VGND VGND.n2029 0.0603958
R6280 VGND.n2025 VGND 0.0603958
R6281 VGND.n1126 VGND 0.0603958
R6282 VGND.n1128 VGND 0.0603958
R6283 VGND.n1134 VGND 0.0603958
R6284 VGND.n1167 VGND 0.0603958
R6285 VGND.n1174 VGND 0.0603958
R6286 VGND.n1177 VGND 0.0603958
R6287 VGND.n6283 VGND 0.0603958
R6288 VGND.n6278 VGND 0.0603958
R6289 VGND.n6221 VGND 0.0603958
R6290 VGND.n6209 VGND 0.0603958
R6291 VGND VGND.n6205 0.0603958
R6292 VGND VGND.n6204 0.0603958
R6293 VGND.n6200 VGND 0.0603958
R6294 VGND VGND.n6193 0.0603958
R6295 VGND VGND.n6179 0.0603958
R6296 VGND.n6176 VGND 0.0603958
R6297 VGND.n6170 VGND 0.0603958
R6298 VGND.n6083 VGND 0.0603958
R6299 VGND.n6076 VGND 0.0603958
R6300 VGND VGND.n6073 0.0603958
R6301 VGND VGND.n6841 0.0603958
R6302 VGND.n6842 VGND 0.0603958
R6303 VGND.n6849 VGND 0.0603958
R6304 VGND.n6854 VGND 0.0603958
R6305 VGND.n6857 VGND 0.0603958
R6306 VGND.n6911 VGND 0.0603958
R6307 VGND.n6936 VGND 0.0603958
R6308 VGND.n6943 VGND 0.0603958
R6309 VGND VGND.n1010 0.0603958
R6310 VGND.n6969 VGND 0.0603958
R6311 VGND.n7039 VGND 0.0603958
R6312 VGND.n7044 VGND 0.0603958
R6313 VGND.n7075 VGND 0.0603958
R6314 VGND.n7078 VGND 0.0603958
R6315 VGND VGND.n970 0.0603958
R6316 VGND.n7094 VGND 0.0603958
R6317 VGND.n7101 VGND 0.0603958
R6318 VGND.n7113 VGND 0.0603958
R6319 VGND.n7187 VGND 0.0603958
R6320 VGND VGND.n942 0.0603958
R6321 VGND.n7201 VGND 0.0603958
R6322 VGND.n7222 VGND 0.0603958
R6323 VGND.n7254 VGND 0.0603958
R6324 VGND VGND.n880 0.0603958
R6325 VGND.n900 VGND 0.0603958
R6326 VGND.n893 VGND 0.0603958
R6327 VGND.n888 VGND 0.0603958
R6328 VGND VGND.n2179 0.0603958
R6329 VGND.n2187 VGND 0.0603958
R6330 VGND.n2192 VGND 0.0603958
R6331 VGND.n2195 VGND 0.0603958
R6332 VGND.n6792 VGND 0.0603958
R6333 VGND.n6780 VGND 0.0603958
R6334 VGND VGND.n6779 0.0603958
R6335 VGND.n6770 VGND 0.0603958
R6336 VGND.n1038 VGND 0.0603958
R6337 VGND.n6351 VGND 0.0603958
R6338 VGND.n6354 VGND 0.0603958
R6339 VGND.n6358 VGND 0.0603958
R6340 VGND.n6384 VGND 0.0603958
R6341 VGND.n6388 VGND 0.0603958
R6342 VGND.n6462 VGND 0.0603958
R6343 VGND.n6466 VGND 0.0603958
R6344 VGND.n6469 VGND 0.0603958
R6345 VGND.n6479 VGND 0.0603958
R6346 VGND.n6481 VGND 0.0603958
R6347 VGND.n6496 VGND 0.0603958
R6348 VGND.n6498 VGND 0.0603958
R6349 VGND.n6501 VGND 0.0603958
R6350 VGND.n6507 VGND 0.0603958
R6351 VGND.n6515 VGND 0.0603958
R6352 VGND.n6523 VGND 0.0603958
R6353 VGND.n6606 VGND 0.0603958
R6354 VGND.n6610 VGND 0.0603958
R6355 VGND.n6617 VGND 0.0603958
R6356 VGND.n6620 VGND 0.0603958
R6357 VGND.n6628 VGND 0.0603958
R6358 VGND.n6726 VGND 0.0603958
R6359 VGND VGND.n6725 0.0603958
R6360 VGND.n6681 VGND 0.0603958
R6361 VGND VGND.n6680 0.0603958
R6362 VGND.n6677 VGND 0.0603958
R6363 VGND.n7431 VGND 0.0603958
R6364 VGND.n7443 VGND 0.0603958
R6365 VGND.n7445 VGND 0.0603958
R6366 VGND.n7445 VGND 0.0603958
R6367 VGND VGND.n7990 0.0603958
R6368 VGND.n309 VGND 0.0603958
R6369 VGND.n315 VGND 0.0603958
R6370 VGND.n316 VGND 0.0603958
R6371 VGND.n323 VGND 0.0603958
R6372 VGND VGND.n682 0.0603958
R6373 VGND.n678 VGND 0.0603958
R6374 VGND.n653 VGND 0.0603958
R6375 VGND.n650 VGND 0.0603958
R6376 VGND VGND.n649 0.0603958
R6377 VGND VGND.n632 0.0603958
R6378 VGND VGND.n631 0.0603958
R6379 VGND.n623 VGND 0.0603958
R6380 VGND.n612 VGND 0.0603958
R6381 VGND.n554 VGND 0.0603958
R6382 VGND VGND.n553 0.0603958
R6383 VGND.n549 VGND 0.0603958
R6384 VGND.n549 VGND 0.0603958
R6385 VGND VGND.n548 0.0603958
R6386 VGND.n544 VGND 0.0603958
R6387 VGND VGND.n537 0.0603958
R6388 VGND VGND.n536 0.0603958
R6389 VGND VGND.n535 0.0603958
R6390 VGND.n532 VGND 0.0603958
R6391 VGND.n525 VGND 0.0603958
R6392 VGND VGND.n503 0.0603958
R6393 VGND VGND.n499 0.0603958
R6394 VGND.n498 VGND 0.0603958
R6395 VGND VGND.n497 0.0603958
R6396 VGND.n7953 VGND 0.0603958
R6397 VGND.n7939 VGND 0.0603958
R6398 VGND VGND.n7906 0.0603958
R6399 VGND.n7933 VGND 0.0603958
R6400 VGND.n7926 VGND 0.0603958
R6401 VGND VGND.n7925 0.0603958
R6402 VGND.n7910 VGND 0.0603958
R6403 VGND.n7918 VGND 0.0603958
R6404 VGND.n4965 VGND 0.0564896
R6405 VGND.n5209 VGND.n5208 0.0548679
R6406 VGND.n2102 VGND.n1968 0.0548679
R6407 VGND.n7512 VGND.n7506 0.0525833
R6408 VGND.n7611 VGND.n7610 0.0525833
R6409 VGND.n4215 VGND.n4213 0.0525833
R6410 VGND.n4381 VGND.n4379 0.0525833
R6411 VGND.n5156 VGND.n5154 0.0525833
R6412 VGND.n2698 VGND.n2697 0.0525833
R6413 VGND.n2345 VGND.n2344 0.0525833
R6414 VGND.n2301 VGND.n2300 0.0525833
R6415 VGND.n6903 VGND.n1016 0.0525833
R6416 VGND.n6795 VGND.n1035 0.0525833
R6417 VGND.n8001 VGND.n8000 0.0525833
R6418 VGND.n145 VGND 0.0512812
R6419 VGND.n4182 VGND 0.0512812
R6420 VGND.n4276 VGND 0.0512812
R6421 VGND.n5114 VGND 0.0512812
R6422 VGND.n5193 VGND 0.0512812
R6423 VGND.n7448 VGND 0.0512812
R6424 VGND.n7897 VGND.n7896 0.0489687
R6425 VGND.n7893 VGND.n39 0.0489687
R6426 VGND.n7474 VGND.n7473 0.0489687
R6427 VGND.n694 VGND.n693 0.0489687
R6428 VGND.n4084 VGND.n4082 0.0486771
R6429 VGND.n2820 VGND.n2818 0.0486771
R6430 VGND.n5415 VGND.n5414 0.0486771
R6431 VGND.n6710 VGND.n6708 0.0486771
R6432 VGND VGND.n4239 0.0463917
R6433 VGND.n153 VGND.n152 0.0460729
R6434 VGND.n707 VGND.n706 0.0460729
R6435 VGND.n7591 VGND.n7590 0.0460729
R6436 VGND.n7711 VGND.n81 0.0460729
R6437 VGND.n4191 VGND.n4190 0.0460729
R6438 VGND.n5131 VGND.n5130 0.0460729
R6439 VGND.n1896 VGND.n1895 0.0460729
R6440 VGND.n6868 VGND.n6867 0.0460729
R6441 VGND.n7457 VGND.n7456 0.0460729
R6442 VGND.n5039 VGND 0.0449123
R6443 VGND.n6740 VGND.n6735 0.0447708
R6444 VGND.n237 VGND.n236 0.0395625
R6445 VGND.n7692 VGND.n7691 0.0395625
R6446 VGND.n4465 VGND.n4464 0.0395625
R6447 VGND.n4763 VGND.n4762 0.0395625
R6448 VGND.n1779 VGND.n1778 0.0395625
R6449 VGND.n6399 VGND.n6398 0.0395625
R6450 VGND.n6812 VGND.n6811 0.0393514
R6451 VGND.n2212 VGND.n2208 0.0393514
R6452 VGND.n6555 VGND.n1071 0.0393514
R6453 VGND.n159 VGND.n158 0.0393514
R6454 VGND.n3354 VGND.n3350 0.0393514
R6455 VGND.n7552 VGND.n7551 0.0393514
R6456 VGND.n7851 VGND.n67 0.0393514
R6457 VGND.n3126 VGND.n3125 0.0393514
R6458 VGND.n3898 VGND.n3897 0.0393514
R6459 VGND.n4357 VGND.n4284 0.0393514
R6460 VGND.n4524 VGND.n2967 0.0393514
R6461 VGND.n5122 VGND.n5118 0.0393514
R6462 VGND.n2869 VGND.n2868 0.0393514
R6463 VGND.n5256 VGND.n1650 0.0393514
R6464 VGND.n5205 VGND.n5204 0.0393514
R6465 VGND.n5548 VGND.n1447 0.0393514
R6466 VGND.n1729 VGND.n1725 0.0393514
R6467 VGND.n1902 VGND.n1901 0.0393514
R6468 VGND.n5875 VGND.n1323 0.0393514
R6469 VGND.n6252 VGND.n1218 0.0393514
R6470 VGND.n7140 VGND.n7139 0.0393514
R6471 VGND.n583 VGND.n432 0.0393514
R6472 VGND.n7422 VGND.n7421 0.0393514
R6473 VGND.n6823 VGND.n6822 0.0376622
R6474 VGND.n1034 VGND.n1033 0.0376622
R6475 VGND.n1972 VGND.n1971 0.0376622
R6476 VGND.n171 VGND.n170 0.0376622
R6477 VGND.n117 VGND.n116 0.0376622
R6478 VGND.n3138 VGND.n3137 0.0376622
R6479 VGND.n4349 VGND.n4348 0.0376622
R6480 VGND.n2727 VGND.n2726 0.0376622
R6481 VGND.n2408 VGND.n2407 0.0376622
R6482 VGND.n1862 VGND.n1861 0.0376622
R6483 VGND.n1954 VGND.n1953 0.0376622
R6484 VGND.n7996 VGND.n7995 0.0376622
R6485 VGND.n3759 VGND.n3758 0.0373368
R6486 VGND.n3566 VGND.n3565 0.0371114
R6487 VGND.n3604 VGND.n3603 0.0371114
R6488 VGND.n4100 VGND.n4098 0.0371114
R6489 VGND.n4657 VGND.n4656 0.0371114
R6490 VGND.n5039 VGND.n5038 0.0371114
R6491 VGND.n1601 VGND.n1593 0.0371114
R6492 VGND.n5453 VGND.n5452 0.0371114
R6493 VGND.n6010 VGND.n6009 0.0371114
R6494 VGND.n6161 VGND.n1236 0.0371114
R6495 VGND.n7271 VGND.n7269 0.0371114
R6496 VGND.n6724 VGND.n1058 0.0371114
R6497 VGND.n492 VGND.n484 0.0371114
R6498 VGND.n6322 VGND.n6321 0.0370003
R6499 VGND.n7843 VGND.n7842 0.0369583
R6500 VGND.n4537 VGND.n4536 0.0369583
R6501 VGND.n4954 VGND.n4953 0.0369583
R6502 VGND.n5267 VGND.n5266 0.0369583
R6503 VGND.n5540 VGND.n5539 0.0369583
R6504 VGND.n5888 VGND.n5887 0.0369583
R6505 VGND.n6566 VGND.n6565 0.0369583
R6506 VGND.n574 VGND.n573 0.0369583
R6507 VGND.n3069 VGND 0.0347603
R6508 VGND.n5863 VGND 0.0347603
R6509 VGND VGND.n611 0.0347603
R6510 VGND.n3520 VGND 0.0343542
R6511 VGND.n3474 VGND 0.0343542
R6512 VGND.n2980 VGND 0.0343542
R6513 VGND.n2946 VGND 0.0343542
R6514 VGND.n2921 VGND 0.0343542
R6515 VGND.n4825 VGND 0.0343542
R6516 VGND VGND.n4872 0.0343542
R6517 VGND.n4884 VGND 0.0343542
R6518 VGND.n4976 VGND 0.0343542
R6519 VGND.n5010 VGND 0.0343542
R6520 VGND VGND.n2465 0.0343542
R6521 VGND VGND.n2621 0.0343542
R6522 VGND.n5303 VGND 0.0343542
R6523 VGND.n1705 VGND 0.0343542
R6524 VGND.n1841 VGND 0.0343542
R6525 VGND.n5586 VGND 0.0343542
R6526 VGND.n5513 VGND 0.0343542
R6527 VGND.n5912 VGND 0.0343542
R6528 VGND.n1297 VGND 0.0343542
R6529 VGND.n2068 VGND 0.0343542
R6530 VGND.n2028 VGND 0.0343542
R6531 VGND VGND.n1225 0.0343542
R6532 VGND.n6086 VGND 0.0343542
R6533 VGND.n6944 VGND 0.0343542
R6534 VGND.n7040 VGND 0.0343542
R6535 VGND.n6385 VGND 0.0343542
R6536 VGND VGND.n6608 0.0343542
R6537 VGND VGND.n7444 0.0343542
R6538 VGND VGND.n398 0.0343542
R6539 VGND.n500 VGND 0.0343542
R6540 VGND.n7917 VGND 0.0343542
R6541 VGND VGND.n176 0.0330521
R6542 VGND VGND.n799 0.0330521
R6543 VGND VGND.n3397 0.0330521
R6544 VGND VGND.n7644 0.0330521
R6545 VGND.n7793 VGND 0.0330521
R6546 VGND.n3251 VGND 0.0330521
R6547 VGND.n4137 VGND 0.0330521
R6548 VGND VGND.n3843 0.0330521
R6549 VGND VGND.n3953 0.0330521
R6550 VGND.n4362 VGND 0.0330521
R6551 VGND VGND.n4405 0.0330521
R6552 VGND VGND.n3039 0.0330521
R6553 VGND VGND.n4571 0.0330521
R6554 VGND VGND.n2732 0.0330521
R6555 VGND VGND.n4877 0.0330521
R6556 VGND VGND.n4991 0.0330521
R6557 VGND VGND.n2418 0.0330521
R6558 VGND.n2661 VGND 0.0330521
R6559 VGND.n1647 VGND 0.0330521
R6560 VGND VGND.n1732 0.0330521
R6561 VGND.n1832 VGND 0.0330521
R6562 VGND.n5581 VGND 0.0330521
R6563 VGND.n5500 VGND 0.0330521
R6564 VGND.n5786 VGND 0.0330521
R6565 VGND.n5838 VGND 0.0330521
R6566 VGND VGND.n5924 0.0330521
R6567 VGND.n2070 VGND 0.0330521
R6568 VGND VGND.n1177 0.0330521
R6569 VGND.n6205 VGND 0.0330521
R6570 VGND.n1013 VGND 0.0330521
R6571 VGND.n970 VGND 0.0330521
R6572 VGND.n942 VGND 0.0330521
R6573 VGND.n2217 VGND 0.0330521
R6574 VGND VGND.n1038 0.0330521
R6575 VGND VGND.n6514 0.0330521
R6576 VGND VGND.n6604 0.0330521
R6577 VGND VGND.n11 0.0330521
R6578 VGND.n632 VGND 0.0330521
R6579 VGND.n536 VGND 0.0330521
R6580 VGND.n6441 VGND.n6440 0.0325946
R6581 VGND.n3460 VGND.n3459 0.0325946
R6582 VGND.n268 VGND.n267 0.0325946
R6583 VGND.n3335 VGND.n3168 0.0325946
R6584 VGND.n99 VGND.n98 0.0325946
R6585 VGND.n4112 VGND.n3620 0.0325946
R6586 VGND.n3743 VGND.n3742 0.0325946
R6587 VGND.n4629 VGND.n4627 0.0325946
R6588 VGND.n4232 VGND.n4231 0.0325946
R6589 VGND.n4706 VGND.n4705 0.0325946
R6590 VGND.n2834 VGND.n2832 0.0325946
R6591 VGND.n5312 VGND.n1483 0.0325946
R6592 VGND.n5332 VGND.n5331 0.0325946
R6593 VGND.n2444 VGND.n2443 0.0325946
R6594 VGND.n5717 VGND.n5666 0.0325946
R6595 VGND.n5991 VGND.n1252 0.0325946
R6596 VGND.n6741 VGND.n1057 0.0325946
R6597 VGND.n459 VGND.n457 0.0325946
R6598 VGND.n287 VGND.n286 0.0325946
R6599 VGND.n6123 VGND.n6122 0.0317953
R6600 VGND.n3534 VGND.n3532 0.0317953
R6601 VGND.n3320 VGND.n3319 0.0317953
R6602 VGND.n4670 VGND.n4669 0.0317953
R6603 VGND.n1307 VGND.n1305 0.0317953
R6604 VGND VGND.n189 0.03175
R6605 VGND VGND.n798 0.03175
R6606 VGND.n845 VGND 0.03175
R6607 VGND.n3348 VGND 0.03175
R6608 VGND.n3424 VGND 0.03175
R6609 VGND.n3519 VGND 0.03175
R6610 VGND.n3490 VGND 0.03175
R6611 VGND.n7577 VGND 0.03175
R6612 VGND.n7600 VGND.n7599 0.03175
R6613 VGND.n7757 VGND 0.03175
R6614 VGND.n7775 VGND 0.03175
R6615 VGND.n3178 VGND 0.03175
R6616 VGND.n3300 VGND 0.03175
R6617 VGND.n3278 VGND 0.03175
R6618 VGND VGND.n4166 0.03175
R6619 VGND.n4198 VGND.n4197 0.03175
R6620 VGND VGND.n3682 0.03175
R6621 VGND.n3702 VGND 0.03175
R6622 VGND VGND.n3722 0.03175
R6623 VGND.n3803 VGND 0.03175
R6624 VGND.n3807 VGND 0.03175
R6625 VGND VGND.n3818 0.03175
R6626 VGND VGND.n3845 0.03175
R6627 VGND VGND.n3991 0.03175
R6628 VGND.n4369 VGND.n4368 0.03175
R6629 VGND VGND.n4387 0.03175
R6630 VGND.n4406 VGND 0.03175
R6631 VGND.n4435 VGND 0.03175
R6632 VGND VGND.n3038 0.03175
R6633 VGND.n2934 VGND 0.03175
R6634 VGND VGND.n5097 0.03175
R6635 VGND.n5139 VGND.n5138 0.03175
R6636 VGND VGND.n4717 0.03175
R6637 VGND.n4753 VGND 0.03175
R6638 VGND.n4992 VGND 0.03175
R6639 VGND.n2603 VGND 0.03175
R6640 VGND.n2648 VGND 0.03175
R6641 VGND.n1642 VGND 0.03175
R6642 VGND.n1626 VGND 0.03175
R6643 VGND.n1612 VGND 0.03175
R6644 VGND.n1512 VGND 0.03175
R6645 VGND.n1506 VGND 0.03175
R6646 VGND.n5584 VGND 0.03175
R6647 VGND.n5576 VGND 0.03175
R6648 VGND.n5572 VGND 0.03175
R6649 VGND.n5521 VGND 0.03175
R6650 VGND.n5501 VGND 0.03175
R6651 VGND.n5461 VGND 0.03175
R6652 VGND VGND.n1871 0.03175
R6653 VGND VGND.n1921 0.03175
R6654 VGND VGND.n5797 0.03175
R6655 VGND.n5821 VGND 0.03175
R6656 VGND.n5858 VGND 0.03175
R6657 VGND VGND.n5902 0.03175
R6658 VGND.n5968 VGND 0.03175
R6659 VGND VGND.n5935 0.03175
R6660 VGND.n1282 VGND 0.03175
R6661 VGND.n1273 VGND 0.03175
R6662 VGND VGND.n2160 0.03175
R6663 VGND.n2093 VGND 0.03175
R6664 VGND.n2076 VGND 0.03175
R6665 VGND VGND.n1126 0.03175
R6666 VGND.n6179 VGND 0.03175
R6667 VGND.n6076 VGND 0.03175
R6668 VGND.n6854 VGND 0.03175
R6669 VGND.n6875 VGND.n6874 0.03175
R6670 VGND.n7075 VGND 0.03175
R6671 VGND.n2192 VGND 0.03175
R6672 VGND.n2224 VGND.n2223 0.03175
R6673 VGND.n6780 VGND 0.03175
R6674 VGND VGND.n6351 0.03175
R6675 VGND.n6515 VGND 0.03175
R6676 VGND.n6680 VGND 0.03175
R6677 VGND VGND.n315 0.03175
R6678 VGND.n650 VGND 0.03175
R6679 VGND.n612 VGND 0.03175
R6680 VGND.n535 VGND 0.03175
R6681 VGND.n7925 VGND 0.03175
R6682 VGND.n7312 VGND.n7311 0.0315717
R6683 VGND.n7903 VGND.n18 0.0315717
R6684 VGND.n6421 VGND.n6420 0.0309054
R6685 VGND.n6822 VGND.n6821 0.0309054
R6686 VGND.n1033 VGND.n1032 0.0309054
R6687 VGND.n6547 VGND.n6546 0.0309054
R6688 VGND.n6546 VGND.n6545 0.0309054
R6689 VGND.n1071 VGND.n1070 0.0309054
R6690 VGND.n2002 VGND.n2001 0.0309054
R6691 VGND.n6317 VGND.n6316 0.0309054
R6692 VGND.n170 VGND.n169 0.0309054
R6693 VGND.n702 VGND.n701 0.0309054
R6694 VGND.n821 VGND.n820 0.0309054
R6695 VGND.n116 VGND.n115 0.0309054
R6696 VGND.n83 VGND.n82 0.0309054
R6697 VGND.n7819 VGND.n7818 0.0309054
R6698 VGND.n3137 VGND.n3136 0.0309054
R6699 VGND.n3729 VGND.n3728 0.0309054
R6700 VGND.n3864 VGND.n3863 0.0309054
R6701 VGND.n4348 VGND.n4347 0.0309054
R6702 VGND.n4483 VGND.n4482 0.0309054
R6703 VGND.n3072 VGND.n3071 0.0309054
R6704 VGND.n2726 VGND.n2725 0.0309054
R6705 VGND.n4784 VGND.n4783 0.0309054
R6706 VGND.n4921 VGND.n4920 0.0309054
R6707 VGND.n2868 VGND.n2867 0.0309054
R6708 VGND.n2636 VGND.n2635 0.0309054
R6709 VGND.n2430 VGND.n2429 0.0309054
R6710 VGND.n1413 VGND.n1412 0.0309054
R6711 VGND.n1447 VGND.n1446 0.0309054
R6712 VGND.n1861 VGND.n1860 0.0309054
R6713 VGND.n1392 VGND.n1391 0.0309054
R6714 VGND.n1953 VGND.n1952 0.0309054
R6715 VGND.n5695 VGND.n5694 0.0309054
R6716 VGND.n5866 VGND.n5865 0.0309054
R6717 VGND.n1323 VGND.n1322 0.0309054
R6718 VGND.n1183 VGND.n1182 0.0309054
R6719 VGND.n7134 VGND.n7133 0.0309054
R6720 VGND.n7133 VGND.n7132 0.0309054
R6721 VGND.n418 VGND.n417 0.0309054
R6722 VGND.n432 VGND.n431 0.0309054
R6723 VGND.n8019 VGND.n8018 0.0309054
R6724 VGND.n7995 VGND.n7994 0.0309054
R6725 VGND.n6977 VGND.n6976 0.0309054
R6726 VGND.n1000 VGND.n999 0.0309054
R6727 VGND.n395 VGND.n394 0.0309054
R6728 VGND.n3461 VGND 0.0304479
R6729 VGND.n3334 VGND 0.0304479
R6730 VGND.n4111 VGND 0.0304479
R6731 VGND.n4628 VGND 0.0304479
R6732 VGND.n2833 VGND 0.0304479
R6733 VGND.n5311 VGND 0.0304479
R6734 VGND.n5333 VGND 0.0304479
R6735 VGND.n5990 VGND 0.0304479
R6736 VGND.n6105 VGND 0.0304479
R6737 VGND.n7282 VGND 0.0304479
R6738 VGND.n458 VGND 0.0304479
R6739 VGND.n6420 VGND.n1109 0.0292162
R6740 VGND.n6293 VGND.n6292 0.0292162
R6741 VGND.n3570 VGND.n3569 0.0292162
R6742 VGND.n703 VGND.n702 0.0292162
R6743 VGND.n3608 VGND.n3607 0.0292162
R6744 VGND.n84 VGND.n83 0.0292162
R6745 VGND.n4096 VGND.n4005 0.0292162
R6746 VGND.n3728 VGND.n3668 0.0292162
R6747 VGND.n4661 VGND.n4660 0.0292162
R6748 VGND.n4482 VGND.n2892 0.0292162
R6749 VGND.n4783 VGND.n2874 0.0292162
R6750 VGND.n5043 VGND.n5042 0.0292162
R6751 VGND.n1599 VGND.n1595 0.0292162
R6752 VGND.n2553 VGND.n2552 0.0292162
R6753 VGND.n5355 VGND.n5354 0.0292162
R6754 VGND.n5637 VGND.n5636 0.0292162
R6755 VGND.n5694 VGND.n5693 0.0292162
R6756 VGND.n6014 VGND.n6013 0.0292162
R6757 VGND.n6159 VGND.n1237 0.0292162
R6758 VGND.n6097 VGND.n6096 0.0292162
R6759 VGND.n6722 VGND.n6645 0.0292162
R6760 VGND.n7267 VGND.n7261 0.0292162
R6761 VGND.n7260 VGND.n7259 0.0292162
R6762 VGND.n490 VGND.n486 0.0292162
R6763 VGND.n980 VGND.n979 0.0292162
R6764 VGND.n394 VGND.n296 0.0292162
R6765 VGND.n812 VGND.n811 0.0291458
R6766 VGND.n7835 VGND.n7833 0.0291458
R6767 VGND.n3880 VGND.n3878 0.0291458
R6768 VGND.n4529 VGND.n4527 0.0291458
R6769 VGND.n4910 VGND.n4909 0.0291458
R6770 VGND.n5261 VGND.n5259 0.0291458
R6771 VGND.n5532 VGND.n5530 0.0291458
R6772 VGND.n5880 VGND.n5878 0.0291458
R6773 VGND.n6236 VGND.n6234 0.0291458
R6774 VGND.n7121 VGND.n7120 0.0291458
R6775 VGND.n6560 VGND.n6558 0.0291458
R6776 VGND.n566 VGND.n564 0.0291458
R6777 VGND.n4009 VGND.n4008 0.0289937
R6778 VGND.n4222 VGND.n4221 0.0289937
R6779 VGND.n3775 VGND 0.0278438
R6780 VGND VGND.n2528 0.0278438
R6781 VGND.n5734 VGND 0.0278438
R6782 VGND VGND.n6992 0.0278438
R6783 VGND VGND.n362 0.0278438
R6784 VGND.n3356 VGND 0.0265417
R6785 VGND VGND.n3365 0.0265417
R6786 VGND.n3911 VGND 0.0265417
R6787 VGND.n6244 VGND 0.0265417
R6788 VGND.n7156 VGND 0.0265417
R6789 VGND.n4962 VGND.n4960 0.0264488
R6790 VGND.n5278 VGND.n5277 0.0264488
R6791 VGND.n5897 VGND.n5895 0.0264488
R6792 VGND.n581 VGND.n562 0.0264488
R6793 VGND.n6421 VGND.n6419 0.0258378
R6794 VGND.n6545 VGND.n6544 0.0258378
R6795 VGND.n1119 VGND.n1118 0.0258378
R6796 VGND.n3451 VGND.n3450 0.0258378
R6797 VGND.n815 VGND.n814 0.0258378
R6798 VGND.n3165 VGND.n3164 0.0258378
R6799 VGND.n7858 VGND.n7857 0.0258378
R6800 VGND.n3616 VGND.n3615 0.0258378
R6801 VGND.n3650 VGND.n3649 0.0258378
R6802 VGND.n4624 VGND.n4623 0.0258378
R6803 VGND.n4509 VGND.n4508 0.0258378
R6804 VGND.n4913 VGND.n4912 0.0258378
R6805 VGND.n2830 VGND.n2829 0.0258378
R6806 VGND.n2741 VGND.n2740 0.0258378
R6807 VGND.n5054 VGND.n5053 0.0258378
R6808 VGND.n5225 VGND.n5224 0.0258378
R6809 VGND.n1479 VGND.n1478 0.0258378
R6810 VGND.n1569 VGND.n1568 0.0258378
R6811 VGND.n2549 VGND.n2548 0.0258378
R6812 VGND.n1462 VGND.n1461 0.0258378
R6813 VGND.n1432 VGND.n1431 0.0258378
R6814 VGND.n5647 VGND.n1394 0.0258378
R6815 VGND.n1333 VGND.n1332 0.0258378
R6816 VGND.n1250 VGND.n1249 0.0258378
R6817 VGND.n6024 VGND.n6023 0.0258378
R6818 VGND.n6028 VGND.n6027 0.0258378
R6819 VGND.n1191 VGND.n1190 0.0258378
R6820 VGND.n6099 VGND.n6098 0.0258378
R6821 VGND.n6135 VGND.n6134 0.0258378
R6822 VGND.n6140 VGND.n6139 0.0258378
R6823 VGND.n1053 VGND.n1052 0.0258378
R6824 VGND.n7294 VGND.n7293 0.0258378
R6825 VGND.n7298 VGND.n7297 0.0258378
R6826 VGND.n454 VGND.n453 0.0258378
R6827 VGND.n22 VGND.n21 0.0258378
R6828 VGND.n595 VGND.n594 0.0258378
R6829 VGND.n7014 VGND.n1002 0.0258378
R6830 VGND.n395 VGND.n393 0.0258378
R6831 VGND.n3368 VGND.n3366 0.0256464
R6832 VGND.n7849 VGND.n69 0.0256464
R6833 VGND.n3921 VGND.n3920 0.0256464
R6834 VGND.n4546 VGND.n4544 0.0256464
R6835 VGND.n5546 VGND.n5528 0.0256464
R6836 VGND.n6250 VGND.n6227 0.0256464
R6837 VGND.n7164 VGND.n7162 0.0256464
R6838 VGND.n6578 VGND.n6577 0.0256464
R6839 VGND.n151 VGND.n150 0.0252396
R6840 VGND.n250 VGND.n249 0.0252396
R6841 VGND.n3462 VGND.n3461 0.0252396
R6842 VGND.n7588 VGND.n7587 0.0252396
R6843 VGND.n7705 VGND.n7704 0.0252396
R6844 VGND.n3334 VGND.n3333 0.0252396
R6845 VGND.n4188 VGND.n4187 0.0252396
R6846 VGND.n3762 VGND.n3761 0.0252396
R6847 VGND.n3859 VGND 0.0252396
R6848 VGND.n3876 VGND.n3875 0.0252396
R6849 VGND.n4111 VGND.n3151 0.0252396
R6850 VGND.n4475 VGND.n4474 0.0252396
R6851 VGND.n3060 VGND 0.0252396
R6852 VGND.n2971 VGND.n2969 0.0252396
R6853 VGND.n4579 VGND 0.0252396
R6854 VGND.n4628 VGND.n2899 0.0252396
R6855 VGND.n4777 VGND.n4776 0.0252396
R6856 VGND.n2833 VGND.n2738 0.0252396
R6857 VGND.n2798 VGND 0.0252396
R6858 VGND.n5199 VGND.n5198 0.0252396
R6859 VGND.n2537 VGND.n2536 0.0252396
R6860 VGND.n2630 VGND.n2627 0.0252396
R6861 VGND.n5311 VGND.n5310 0.0252396
R6862 VGND.n1770 VGND.n1769 0.0252396
R6863 VGND.n5559 VGND.n5557 0.0252396
R6864 VGND.n5334 VGND.n5333 0.0252396
R6865 VGND.n1877 VGND 0.0252396
R6866 VGND.n1894 VGND.n1893 0.0252396
R6867 VGND.n5719 VGND.n5718 0.0252396
R6868 VGND.n1357 VGND.n1355 0.0252396
R6869 VGND.n5990 VGND.n5989 0.0252396
R6870 VGND.n2132 VGND.n2131 0.0252396
R6871 VGND.n6319 VGND.n6315 0.0252396
R6872 VGND.n6232 VGND.n6231 0.0252396
R6873 VGND.n6106 VGND.n6105 0.0252396
R6874 VGND.n6865 VGND.n6864 0.0252396
R6875 VGND.n7006 VGND.n7005 0.0252396
R6876 VGND.n7125 VGND.n7123 0.0252396
R6877 VGND.n7282 VGND.n878 0.0252396
R6878 VGND.n6412 VGND.n6411 0.0252396
R6879 VGND.n6537 VGND.n6535 0.0252396
R6880 VGND.n6740 VGND.n6739 0.0252396
R6881 VGND.n7454 VGND.n7453 0.0252396
R6882 VGND.n376 VGND.n375 0.0252396
R6883 VGND.n414 VGND.n412 0.0252396
R6884 VGND.n458 VGND.n17 0.0252396
R6885 VGND VGND.n1551 0.0250613
R6886 VGND.n6830 VGND.n6829 0.0241486
R6887 VGND.n2172 VGND.n2171 0.0241486
R6888 VGND.n2156 VGND.n2155 0.0241486
R6889 VGND.n7396 VGND.n7395 0.0241486
R6890 VGND.n7883 VGND.n7882 0.0241486
R6891 VGND.n7523 VGND.n7522 0.0241486
R6892 VGND.n7861 VGND.n7860 0.0241486
R6893 VGND.n3097 VGND.n3096 0.0241486
R6894 VGND.n3887 VGND.n3886 0.0241486
R6895 VGND.n4289 VGND.n4288 0.0241486
R6896 VGND.n4512 VGND.n4511 0.0241486
R6897 VGND.n4316 VGND.n4315 0.0241486
R6898 VGND.n4945 VGND.n4944 0.0241486
R6899 VGND.n5228 VGND.n5227 0.0241486
R6900 VGND.n2397 VGND.n2396 0.0241486
R6901 VGND.n1436 VGND.n1435 0.0241486
R6902 VGND.n1744 VGND.n1743 0.0241486
R6903 VGND.n1917 VGND.n1916 0.0241486
R6904 VGND.n1337 VGND.n1336 0.0241486
R6905 VGND.n1194 VGND.n1193 0.0241486
R6906 VGND.n7152 VGND.n944 0.0241486
R6907 VGND.n599 VGND.n598 0.0241486
R6908 VGND.n7425 VGND.n7424 0.0241486
R6909 VGND.n7498 VGND.n7497 0.0239375
R6910 VGND.n252 VGND.n251 0.0239375
R6911 VGND.n3489 VGND 0.0239375
R6912 VGND.n7603 VGND.n7602 0.0239375
R6913 VGND.n7707 VGND.n7706 0.0239375
R6914 VGND VGND.n3187 0.0239375
R6915 VGND.n4202 VGND.n4200 0.0239375
R6916 VGND.n3760 VGND.n3759 0.0239375
R6917 VGND VGND.n3667 0.0239375
R6918 VGND.n4046 VGND 0.0239375
R6919 VGND.n4372 VGND.n4371 0.0239375
R6920 VGND.n4455 VGND 0.0239375
R6921 VGND.n4477 VGND.n4476 0.0239375
R6922 VGND VGND.n2895 0.0239375
R6923 VGND VGND.n3022 0.0239375
R6924 VGND VGND.n4552 0.0239375
R6925 VGND VGND.n4559 0.0239375
R6926 VGND.n2926 VGND 0.0239375
R6927 VGND.n5143 VGND.n5141 0.0239375
R6928 VGND.n5081 VGND 0.0239375
R6929 VGND.n4779 VGND.n4778 0.0239375
R6930 VGND VGND.n2873 0.0239375
R6931 VGND.n2712 VGND.n2710 0.0239375
R6932 VGND.n2539 VGND.n2538 0.0239375
R6933 VGND.n2551 VGND 0.0239375
R6934 VGND.n5284 VGND 0.0239375
R6935 VGND.n1639 VGND 0.0239375
R6936 VGND.n1615 VGND 0.0239375
R6937 VGND.n1509 VGND 0.0239375
R6938 VGND.n2358 VGND.n2357 0.0239375
R6939 VGND.n1768 VGND.n1767 0.0239375
R6940 VGND VGND.n5646 0.0239375
R6941 VGND.n5630 VGND 0.0239375
R6942 VGND.n5585 VGND 0.0239375
R6943 VGND.n5577 VGND 0.0239375
R6944 VGND.n5520 VGND 0.0239375
R6945 VGND.n5492 VGND 0.0239375
R6946 VGND.n2315 VGND.n2313 0.0239375
R6947 VGND.n5682 VGND 0.0239375
R6948 VGND.n5798 VGND 0.0239375
R6949 VGND.n5903 VGND 0.0239375
R6950 VGND.n5967 VGND 0.0239375
R6951 VGND.n2283 VGND.n2281 0.0239375
R6952 VGND VGND.n6303 0.0239375
R6953 VGND.n6221 VGND 0.0239375
R6954 VGND.n6882 VGND.n6881 0.0239375
R6955 VGND.n7008 VGND.n7007 0.0239375
R6956 VGND VGND.n978 0.0239375
R6957 VGND.n2238 VGND.n2237 0.0239375
R6958 VGND.n6414 VGND.n6413 0.0239375
R6959 VGND VGND.n1108 0.0239375
R6960 VGND.n8020 VGND.n0 0.0239375
R6961 VGND.n378 VGND.n377 0.0239375
R6962 VGND.n397 VGND 0.0239375
R6963 VGND.n553 VGND 0.0239375
R6964 VGND.n5564 VGND.n5563 0.0238078
R6965 VGND.n7130 VGND.n7129 0.0238078
R6966 VGND.n6542 VGND.n6541 0.0238078
R6967 VGND.n827 VGND.n819 0.0238078
R6968 VGND.n7826 VGND.n7824 0.0238078
R6969 VGND.n3871 VGND.n3869 0.0238078
R6970 VGND.n3069 VGND.n3068 0.0238078
R6971 VGND.n4918 VGND.n4917 0.0238078
R6972 VGND.n2642 VGND.n2634 0.0238078
R6973 VGND.n5863 VGND.n5862 0.0238078
R6974 VGND.n6262 VGND.n1181 0.0238078
R6975 VGND.n611 VGND.n416 0.0238078
R6976 VGND VGND.n2415 0.0231359
R6977 VGND.n2095 VGND 0.0231359
R6978 VGND.n6798 VGND 0.0231359
R6979 VGND.n132 VGND 0.0226354
R6980 VGND.n137 VGND 0.0226354
R6981 VGND VGND.n140 0.0226354
R6982 VGND.n7392 VGND 0.0226354
R6983 VGND.n7376 VGND 0.0226354
R6984 VGND.n196 VGND 0.0226354
R6985 VGND.n211 VGND 0.0226354
R6986 VGND.n218 VGND 0.0226354
R6987 VGND.n254 VGND.n252 0.0226354
R6988 VGND VGND.n747 0.0226354
R6989 VGND.n749 VGND 0.0226354
R6990 VGND.n775 VGND 0.0226354
R6991 VGND.n786 VGND 0.0226354
R6992 VGND VGND.n797 0.0226354
R6993 VGND.n832 VGND 0.0226354
R6994 VGND.n3376 VGND 0.0226354
R6995 VGND.n3349 VGND 0.0226354
R6996 VGND.n3383 VGND 0.0226354
R6997 VGND VGND.n3396 0.0226354
R6998 VGND.n3398 VGND 0.0226354
R6999 VGND.n3407 VGND 0.0226354
R7000 VGND.n3416 VGND 0.0226354
R7001 VGND.n3431 VGND 0.0226354
R7002 VGND.n3437 VGND 0.0226354
R7003 VGND.n3342 VGND 0.0226354
R7004 VGND.n3501 VGND 0.0226354
R7005 VGND.n3493 VGND 0.0226354
R7006 VGND.n3481 VGND 0.0226354
R7007 VGND.n3478 VGND 0.0226354
R7008 VGND.n3477 VGND 0.0226354
R7009 VGND.n7570 VGND 0.0226354
R7010 VGND VGND.n7576 0.0226354
R7011 VGND.n7622 VGND 0.0226354
R7012 VGND.n7639 VGND 0.0226354
R7013 VGND.n7646 VGND 0.0226354
R7014 VGND VGND.n7652 0.0226354
R7015 VGND.n7653 VGND 0.0226354
R7016 VGND.n7673 VGND 0.0226354
R7017 VGND.n7709 VGND.n7707 0.0226354
R7018 VGND.n7764 VGND 0.0226354
R7019 VGND VGND.n7774 0.0226354
R7020 VGND VGND.n7792 0.0226354
R7021 VGND.n3173 VGND 0.0226354
R7022 VGND VGND.n3183 0.0226354
R7023 VGND VGND.n3199 0.0226354
R7024 VGND.n3250 VGND 0.0226354
R7025 VGND.n3248 VGND 0.0226354
R7026 VGND.n3225 VGND 0.0226354
R7027 VGND.n3303 VGND 0.0226354
R7028 VGND VGND.n3258 0.0226354
R7029 VGND.n3281 VGND 0.0226354
R7030 VGND.n3272 VGND 0.0226354
R7031 VGND.n3269 VGND 0.0226354
R7032 VGND.n4167 VGND 0.0226354
R7033 VGND VGND.n4174 0.0226354
R7034 VGND VGND.n4178 0.0226354
R7035 VGND.n4179 VGND 0.0226354
R7036 VGND.n4158 VGND 0.0226354
R7037 VGND.n4138 VGND 0.0226354
R7038 VGND.n3697 VGND 0.0226354
R7039 VGND VGND.n3701 0.0226354
R7040 VGND.n3723 VGND 0.0226354
R7041 VGND.n3730 VGND 0.0226354
R7042 VGND VGND.n3806 0.0226354
R7043 VGND VGND.n3825 0.0226354
R7044 VGND.n3826 VGND 0.0226354
R7045 VGND VGND.n3837 0.0226354
R7046 VGND.n3838 VGND 0.0226354
R7047 VGND VGND.n3852 0.0226354
R7048 VGND VGND.n3858 0.0226354
R7049 VGND.n3927 VGND 0.0226354
R7050 VGND VGND.n3940 0.0226354
R7051 VGND.n3941 VGND 0.0226354
R7052 VGND.n3957 VGND 0.0226354
R7053 VGND VGND.n3978 0.0226354
R7054 VGND VGND.n3980 0.0226354
R7055 VGND.n3981 VGND 0.0226354
R7056 VGND.n3988 VGND 0.0226354
R7057 VGND.n3993 VGND 0.0226354
R7058 VGND.n4000 VGND 0.0226354
R7059 VGND.n4065 VGND 0.0226354
R7060 VGND.n4057 VGND 0.0226354
R7061 VGND.n4049 VGND 0.0226354
R7062 VGND.n4042 VGND 0.0226354
R7063 VGND.n4039 VGND 0.0226354
R7064 VGND.n4033 VGND 0.0226354
R7065 VGND VGND.n4265 0.0226354
R7066 VGND.n4266 VGND 0.0226354
R7067 VGND VGND.n4271 0.0226354
R7068 VGND VGND.n4272 0.0226354
R7069 VGND.n4384 VGND 0.0226354
R7070 VGND.n4389 VGND 0.0226354
R7071 VGND VGND.n4404 0.0226354
R7072 VGND.n4427 VGND 0.0226354
R7073 VGND VGND.n4434 0.0226354
R7074 VGND.n4450 VGND 0.0226354
R7075 VGND.n4480 VGND.n4477 0.0226354
R7076 VGND.n4484 VGND 0.0226354
R7077 VGND VGND.n2990 0.0226354
R7078 VGND VGND.n2991 0.0226354
R7079 VGND.n2992 VGND 0.0226354
R7080 VGND.n3002 VGND 0.0226354
R7081 VGND.n3011 VGND 0.0226354
R7082 VGND.n3023 VGND 0.0226354
R7083 VGND.n3035 VGND 0.0226354
R7084 VGND VGND.n3059 0.0226354
R7085 VGND.n3064 VGND 0.0226354
R7086 VGND VGND.n4570 0.0226354
R7087 VGND VGND.n4578 0.0226354
R7088 VGND.n4584 VGND 0.0226354
R7089 VGND.n4604 VGND 0.0226354
R7090 VGND.n4618 VGND 0.0226354
R7091 VGND.n2938 VGND 0.0226354
R7092 VGND.n2937 VGND 0.0226354
R7093 VGND.n2933 VGND 0.0226354
R7094 VGND.n2922 VGND 0.0226354
R7095 VGND.n2920 VGND 0.0226354
R7096 VGND.n2916 VGND 0.0226354
R7097 VGND.n5111 VGND 0.0226354
R7098 VGND.n5078 VGND 0.0226354
R7099 VGND.n5069 VGND 0.0226354
R7100 VGND VGND.n4726 0.0226354
R7101 VGND.n4728 VGND 0.0226354
R7102 VGND.n4742 VGND 0.0226354
R7103 VGND VGND.n4752 0.0226354
R7104 VGND.n4781 VGND.n4779 0.0226354
R7105 VGND.n4785 VGND 0.0226354
R7106 VGND.n4835 VGND 0.0226354
R7107 VGND.n4873 VGND 0.0226354
R7108 VGND VGND.n4876 0.0226354
R7109 VGND VGND.n4975 0.0226354
R7110 VGND VGND.n4997 0.0226354
R7111 VGND.n5006 VGND 0.0226354
R7112 VGND.n5034 VGND 0.0226354
R7113 VGND.n2811 VGND 0.0226354
R7114 VGND.n2802 VGND 0.0226354
R7115 VGND.n2780 VGND 0.0226354
R7116 VGND.n2779 VGND 0.0226354
R7117 VGND.n2776 VGND 0.0226354
R7118 VGND.n5180 VGND 0.0226354
R7119 VGND.n5171 VGND 0.0226354
R7120 VGND.n2694 VGND 0.0226354
R7121 VGND.n2683 VGND 0.0226354
R7122 VGND.n2669 VGND 0.0226354
R7123 VGND VGND.n2468 0.0226354
R7124 VGND.n2491 VGND 0.0226354
R7125 VGND.n2505 VGND 0.0226354
R7126 VGND.n2541 VGND.n2539 0.0226354
R7127 VGND VGND.n2550 0.0226354
R7128 VGND.n2568 VGND 0.0226354
R7129 VGND.n2588 VGND 0.0226354
R7130 VGND.n2612 VGND 0.0226354
R7131 VGND VGND.n2622 0.0226354
R7132 VGND.n2656 VGND 0.0226354
R7133 VGND VGND.n5283 0.0226354
R7134 VGND.n5289 VGND 0.0226354
R7135 VGND.n1643 VGND 0.0226354
R7136 VGND.n1635 VGND 0.0226354
R7137 VGND.n1629 VGND 0.0226354
R7138 VGND.n1618 VGND 0.0226354
R7139 VGND.n1539 VGND 0.0226354
R7140 VGND.n1521 VGND 0.0226354
R7141 VGND.n1513 VGND 0.0226354
R7142 VGND.n1503 VGND 0.0226354
R7143 VGND.n1498 VGND 0.0226354
R7144 VGND VGND.n1704 0.0226354
R7145 VGND.n1714 VGND 0.0226354
R7146 VGND.n1857 VGND 0.0226354
R7147 VGND.n1845 VGND 0.0226354
R7148 VGND.n1838 VGND 0.0226354
R7149 VGND.n1834 VGND 0.0226354
R7150 VGND.n1824 VGND 0.0226354
R7151 VGND.n1818 VGND 0.0226354
R7152 VGND.n1794 VGND 0.0226354
R7153 VGND.n1791 VGND 0.0226354
R7154 VGND.n1790 VGND 0.0226354
R7155 VGND.n1767 VGND.n1766 0.0226354
R7156 VGND.n5648 VGND 0.0226354
R7157 VGND.n5609 VGND 0.0226354
R7158 VGND.n5604 VGND 0.0226354
R7159 VGND.n5599 VGND 0.0226354
R7160 VGND.n5587 VGND 0.0226354
R7161 VGND.n5578 VGND 0.0226354
R7162 VGND.n5571 VGND 0.0226354
R7163 VGND.n5570 VGND 0.0226354
R7164 VGND.n5512 VGND 0.0226354
R7165 VGND.n5504 VGND 0.0226354
R7166 VGND.n5493 VGND 0.0226354
R7167 VGND.n5482 VGND 0.0226354
R7168 VGND.n5473 VGND 0.0226354
R7169 VGND.n5408 VGND 0.0226354
R7170 VGND.n5392 VGND 0.0226354
R7171 VGND.n5368 VGND 0.0226354
R7172 VGND.n1872 VGND 0.0226354
R7173 VGND.n1942 VGND 0.0226354
R7174 VGND.n1939 VGND 0.0226354
R7175 VGND.n1933 VGND 0.0226354
R7176 VGND.n1928 VGND 0.0226354
R7177 VGND.n1925 VGND 0.0226354
R7178 VGND.n5782 VGND 0.0226354
R7179 VGND.n5758 VGND 0.0226354
R7180 VGND.n5752 VGND 0.0226354
R7181 VGND.n5745 VGND 0.0226354
R7182 VGND.n5714 VGND.n5713 0.0226354
R7183 VGND.n5696 VGND 0.0226354
R7184 VGND VGND.n5796 0.0226354
R7185 VGND VGND.n5828 0.0226354
R7186 VGND VGND.n5833 0.0226354
R7187 VGND.n5834 VGND 0.0226354
R7188 VGND VGND.n5844 0.0226354
R7189 VGND.n5845 VGND 0.0226354
R7190 VGND VGND.n5923 0.0226354
R7191 VGND.n5981 VGND 0.0226354
R7192 VGND.n5971 VGND 0.0226354
R7193 VGND.n5955 VGND 0.0226354
R7194 VGND.n1294 VGND 0.0226354
R7195 VGND.n1285 VGND 0.0226354
R7196 VGND.n1279 VGND 0.0226354
R7197 VGND.n1274 VGND 0.0226354
R7198 VGND.n1265 VGND 0.0226354
R7199 VGND.n2117 VGND 0.0226354
R7200 VGND.n2096 VGND 0.0226354
R7201 VGND VGND.n1978 0.0226354
R7202 VGND.n2082 VGND 0.0226354
R7203 VGND VGND.n1984 0.0226354
R7204 VGND.n2044 VGND 0.0226354
R7205 VGND.n2038 VGND 0.0226354
R7206 VGND.n2033 VGND 0.0226354
R7207 VGND.n2030 VGND 0.0226354
R7208 VGND.n2025 VGND 0.0226354
R7209 VGND.n6304 VGND 0.0226354
R7210 VGND.n1131 VGND 0.0226354
R7211 VGND VGND.n1166 0.0226354
R7212 VGND.n1167 VGND 0.0226354
R7213 VGND.n1171 VGND 0.0226354
R7214 VGND VGND.n1176 0.0226354
R7215 VGND.n6281 VGND 0.0226354
R7216 VGND.n6194 VGND 0.0226354
R7217 VGND VGND.n1231 0.0226354
R7218 VGND VGND.n1234 0.0226354
R7219 VGND.n6079 VGND 0.0226354
R7220 VGND.n6055 VGND 0.0226354
R7221 VGND.n6050 VGND 0.0226354
R7222 VGND VGND.n6848 0.0226354
R7223 VGND.n6907 VGND 0.0226354
R7224 VGND.n6932 VGND 0.0226354
R7225 VGND VGND.n6942 0.0226354
R7226 VGND.n6963 VGND 0.0226354
R7227 VGND VGND.n6968 0.0226354
R7228 VGND.n6969 VGND 0.0226354
R7229 VGND.n7010 VGND.n7008 0.0226354
R7230 VGND.n7015 VGND 0.0226354
R7231 VGND.n7065 VGND 0.0226354
R7232 VGND VGND.n7074 0.0226354
R7233 VGND.n7090 VGND 0.0226354
R7234 VGND.n7098 VGND 0.0226354
R7235 VGND.n7110 VGND 0.0226354
R7236 VGND.n7184 VGND 0.0226354
R7237 VGND.n7196 VGND 0.0226354
R7238 VGND.n7218 VGND 0.0226354
R7239 VGND.n7243 VGND 0.0226354
R7240 VGND.n7251 VGND 0.0226354
R7241 VGND.n909 VGND 0.0226354
R7242 VGND.n906 VGND 0.0226354
R7243 VGND.n886 VGND 0.0226354
R7244 VGND VGND.n2186 0.0226354
R7245 VGND.n6783 VGND 0.0226354
R7246 VGND.n6773 VGND 0.0226354
R7247 VGND.n6769 VGND 0.0226354
R7248 VGND VGND.n6354 0.0226354
R7249 VGND.n6372 VGND 0.0226354
R7250 VGND.n6377 VGND 0.0226354
R7251 VGND.n6381 VGND 0.0226354
R7252 VGND.n6416 VGND.n6414 0.0226354
R7253 VGND.n6422 VGND 0.0226354
R7254 VGND.n6462 VGND 0.0226354
R7255 VGND.n6476 VGND 0.0226354
R7256 VGND VGND.n6479 0.0226354
R7257 VGND VGND.n6492 0.0226354
R7258 VGND VGND.n6496 0.0226354
R7259 VGND.n6503 VGND 0.0226354
R7260 VGND VGND.n6513 0.0226354
R7261 VGND VGND.n6603 0.0226354
R7262 VGND.n6617 VGND 0.0226354
R7263 VGND.n6625 VGND 0.0226354
R7264 VGND.n6638 VGND 0.0226354
R7265 VGND VGND.n6642 0.0226354
R7266 VGND.n6686 VGND 0.0226354
R7267 VGND.n6683 VGND 0.0226354
R7268 VGND.n6664 VGND 0.0226354
R7269 VGND.n7440 VGND 0.0226354
R7270 VGND VGND.n7443 0.0226354
R7271 VGND.n7975 VGND 0.0226354
R7272 VGND VGND.n311 0.0226354
R7273 VGND.n312 VGND 0.0226354
R7274 VGND VGND.n322 0.0226354
R7275 VGND.n331 VGND 0.0226354
R7276 VGND VGND.n341 0.0226354
R7277 VGND.n342 VGND 0.0226354
R7278 VGND.n380 VGND.n378 0.0226354
R7279 VGND VGND.n396 0.0226354
R7280 VGND.n661 VGND 0.0226354
R7281 VGND.n657 VGND 0.0226354
R7282 VGND.n643 VGND 0.0226354
R7283 VGND.n626 VGND 0.0226354
R7284 VGND.n615 VGND 0.0226354
R7285 VGND.n554 VGND 0.0226354
R7286 VGND.n547 VGND 0.0226354
R7287 VGND.n538 VGND 0.0226354
R7288 VGND.n537 VGND 0.0226354
R7289 VGND VGND.n441 0.0226354
R7290 VGND VGND.n447 0.0226354
R7291 VGND.n503 VGND 0.0226354
R7292 VGND.n7943 VGND 0.0226354
R7293 VGND.n7939 VGND 0.0226354
R7294 VGND.n7933 VGND 0.0226354
R7295 VGND VGND.n7910 0.0226354
R7296 VGND VGND.n7913 0.0226354
R7297 VGND.n6345 VGND.n6344 0.0224595
R7298 VGND.n6427 VGND.n6426 0.0224595
R7299 VGND.n6886 VGND.n6885 0.0224595
R7300 VGND.n1023 VGND.n1022 0.0224595
R7301 VGND.n2242 VGND.n2241 0.0224595
R7302 VGND.n2246 VGND.n2245 0.0224595
R7303 VGND.n1093 VGND.n1089 0.0224595
R7304 VGND.n1092 VGND.n1091 0.0224595
R7305 VGND.n1078 VGND.n1077 0.0224595
R7306 VGND.n2286 VGND.n2285 0.0224595
R7307 VGND.n2166 VGND.n2165 0.0224595
R7308 VGND.n6316 VGND.n1117 0.0224595
R7309 VGND.n6325 VGND.n6324 0.0224595
R7310 VGND.n3558 VGND.n3557 0.0224595
R7311 VGND.n3460 VGND.n3453 0.0224595
R7312 VGND.n3549 VGND.n3548 0.0224595
R7313 VGND.n7495 VGND.n7492 0.0224595
R7314 VGND.n7479 VGND.n7478 0.0224595
R7315 VGND.n258 VGND.n257 0.0224595
R7316 VGND.n737 VGND.n735 0.0224595
R7317 VGND.n7886 VGND.n43 0.0224595
R7318 VGND.n7885 VGND.n7884 0.0224595
R7319 VGND.n7878 VGND.n7877 0.0224595
R7320 VGND.n3591 VGND.n3590 0.0224595
R7321 VGND.n3336 VGND.n3335 0.0224595
R7322 VGND.n3582 VGND.n3581 0.0224595
R7323 VGND.n7530 VGND.n7529 0.0224595
R7324 VGND.n7534 VGND.n7533 0.0224595
R7325 VGND.n104 VGND.n103 0.0224595
R7326 VGND.n7718 VGND.n7717 0.0224595
R7327 VGND.n7864 VGND.n7859 0.0224595
R7328 VGND.n7863 VGND.n7862 0.0224595
R7329 VGND.n55 VGND.n54 0.0224595
R7330 VGND.n4114 VGND.n3618 0.0224595
R7331 VGND.n4113 VGND.n4112 0.0224595
R7332 VGND.n4125 VGND.n4122 0.0224595
R7333 VGND.n3104 VGND.n3103 0.0224595
R7334 VGND.n3108 VGND.n3107 0.0224595
R7335 VGND.n3733 VGND.n3732 0.0224595
R7336 VGND.n3756 VGND.n3754 0.0224595
R7337 VGND.n3890 VGND.n3651 0.0224595
R7338 VGND.n3889 VGND.n3888 0.0224595
R7339 VGND.n3909 VGND.n3908 0.0224595
R7340 VGND.n4648 VGND.n4647 0.0224595
R7341 VGND.n4630 VGND.n4629 0.0224595
R7342 VGND.n4639 VGND.n4638 0.0224595
R7343 VGND.n4296 VGND.n4295 0.0224595
R7344 VGND.n4300 VGND.n4299 0.0224595
R7345 VGND.n4237 VGND.n4236 0.0224595
R7346 VGND.n4490 VGND.n4489 0.0224595
R7347 VGND.n4515 VGND.n4510 0.0224595
R7348 VGND.n4514 VGND.n4513 0.0224595
R7349 VGND.n3082 VGND.n3081 0.0224595
R7350 VGND.n4323 VGND.n4322 0.0224595
R7351 VGND.n4327 VGND.n4326 0.0224595
R7352 VGND.n4711 VGND.n4710 0.0224595
R7353 VGND.n4791 VGND.n4790 0.0224595
R7354 VGND.n4941 VGND.n2857 0.0224595
R7355 VGND.n4946 VGND.n4942 0.0224595
R7356 VGND.n4929 VGND.n4928 0.0224595
R7357 VGND.n2843 VGND.n2842 0.0224595
R7358 VGND.n2835 VGND.n2834 0.0224595
R7359 VGND.n5056 VGND.n5052 0.0224595
R7360 VGND.n5231 VGND.n5226 0.0224595
R7361 VGND.n5230 VGND.n5229 0.0224595
R7362 VGND.n5243 VGND.n5242 0.0224595
R7363 VGND.n5314 VGND.n1481 0.0224595
R7364 VGND.n5313 VGND.n5312 0.0224595
R7365 VGND.n1571 VGND.n1567 0.0224595
R7366 VGND.n2715 VGND.n2714 0.0224595
R7367 VGND.n1684 VGND.n1683 0.0224595
R7368 VGND.n2431 VGND.n2430 0.0224595
R7369 VGND.n2547 VGND.n2461 0.0224595
R7370 VGND.n5440 VGND.n5439 0.0224595
R7371 VGND.n5332 VGND.n1464 0.0224595
R7372 VGND.n5431 VGND.n5430 0.0224595
R7373 VGND.n1439 VGND.n1433 0.0224595
R7374 VGND.n1438 VGND.n1437 0.0224595
R7375 VGND.n1420 VGND.n1419 0.0224595
R7376 VGND.n2361 VGND.n2360 0.0224595
R7377 VGND.n2365 VGND.n2364 0.0224595
R7378 VGND.n1393 VGND.n1392 0.0224595
R7379 VGND.n5655 VGND.n5654 0.0224595
R7380 VGND.n2318 VGND.n2317 0.0224595
R7381 VGND.n2322 VGND.n2321 0.0224595
R7382 VGND.n5699 VGND.n5698 0.0224595
R7383 VGND.n5707 VGND.n5705 0.0224595
R7384 VGND.n1340 VGND.n1334 0.0224595
R7385 VGND.n1339 VGND.n1338 0.0224595
R7386 VGND.n1342 VGND.n1341 0.0224595
R7387 VGND.n6000 VGND.n5999 0.0224595
R7388 VGND.n5992 VGND.n5991 0.0224595
R7389 VGND.n6031 VGND.n6030 0.0224595
R7390 VGND.n1197 VGND.n1192 0.0224595
R7391 VGND.n1196 VGND.n1195 0.0224595
R7392 VGND.n1208 VGND.n1207 0.0224595
R7393 VGND.n6101 VGND.n1239 0.0224595
R7394 VGND.n6104 VGND.n6103 0.0224595
R7395 VGND.n6143 VGND.n6142 0.0224595
R7396 VGND.n6743 VGND.n1055 0.0224595
R7397 VGND.n6742 VGND.n6741 0.0224595
R7398 VGND.n6754 VGND.n6751 0.0224595
R7399 VGND.n7285 VGND.n940 0.0224595
R7400 VGND.n7284 VGND.n7283 0.0224595
R7401 VGND.n7301 VGND.n7300 0.0224595
R7402 VGND.n472 VGND.n471 0.0224595
R7403 VGND.n460 VGND.n459 0.0224595
R7404 VGND.n31 VGND.n30 0.0224595
R7405 VGND.n954 VGND.n951 0.0224595
R7406 VGND.n953 VGND.n952 0.0224595
R7407 VGND.n7150 VGND.n7149 0.0224595
R7408 VGND.n602 VGND.n596 0.0224595
R7409 VGND.n601 VGND.n600 0.0224595
R7410 VGND.n420 VGND.n419 0.0224595
R7411 VGND.n7467 VGND.n7466 0.0224595
R7412 VGND.n8017 VGND.n8016 0.0224595
R7413 VGND.n1001 VGND.n1000 0.0224595
R7414 VGND.n7019 VGND.n7018 0.0224595
R7415 VGND.n383 VGND.n382 0.0224595
R7416 VGND.n388 VGND.n387 0.0224595
R7417 VGND.n236 VGND.n235 0.0213333
R7418 VGND.n7691 VGND.n7690 0.0213333
R7419 VGND VGND.n3721 0.0213333
R7420 VGND.n3776 VGND.n3775 0.0213333
R7421 VGND.n4464 VGND.n4463 0.0213333
R7422 VGND.n2996 VGND 0.0213333
R7423 VGND.n2964 VGND 0.0213333
R7424 VGND.n2917 VGND 0.0213333
R7425 VGND.n5098 VGND 0.0213333
R7426 VGND.n4762 VGND.n4761 0.0213333
R7427 VGND.n4843 VGND 0.0213333
R7428 VGND.n4867 VGND 0.0213333
R7429 VGND VGND.n4990 0.0213333
R7430 VGND.n2497 VGND 0.0213333
R7431 VGND.n2578 VGND 0.0213333
R7432 VGND VGND.n2602 0.0213333
R7433 VGND.n5299 VGND 0.0213333
R7434 VGND.n1780 VGND.n1779 0.0213333
R7435 VGND.n5614 VGND 0.0213333
R7436 VGND.n5613 VGND 0.0213333
R7437 VGND.n5608 VGND 0.0213333
R7438 VGND.n5590 VGND 0.0213333
R7439 VGND.n5499 VGND 0.0213333
R7440 VGND.n5465 VGND 0.0213333
R7441 VGND VGND.n5922 0.0213333
R7442 VGND.n2021 VGND.n2020 0.0213333
R7443 VGND.n6180 VGND 0.0213333
R7444 VGND.n6992 VGND.n6991 0.0213333
R7445 VGND.n6398 VGND.n6397 0.0213333
R7446 VGND.n362 VGND.n361 0.0213333
R7447 VGND.n504 VGND 0.0213333
R7448 VGND.n6337 VGND.n6336 0.0207703
R7449 VGND.n6453 VGND.n6452 0.0207703
R7450 VGND.n6898 VGND.n6896 0.0207703
R7451 VGND.n6821 VGND.n6820 0.0207703
R7452 VGND.n2249 VGND.n2248 0.0207703
R7453 VGND.n1032 VGND.n1031 0.0207703
R7454 VGND.n1076 VGND.n1075 0.0207703
R7455 VGND.n2271 VGND.n2267 0.0207703
R7456 VGND.n2269 VGND.n2268 0.0207703
R7457 VGND.n6300 VGND.n6299 0.0207703
R7458 VGND.n3523 VGND.n3522 0.0207703
R7459 VGND.n3530 VGND.n3524 0.0207703
R7460 VGND.n7482 VGND.n7481 0.0207703
R7461 VGND.n169 VGND.n168 0.0207703
R7462 VGND.n721 VGND.n720 0.0207703
R7463 VGND.n705 VGND.n704 0.0207703
R7464 VGND.n3310 VGND.n3309 0.0207703
R7465 VGND.n3317 VGND.n3311 0.0207703
R7466 VGND.n7537 VGND.n7536 0.0207703
R7467 VGND.n115 VGND.n114 0.0207703
R7468 VGND.n7730 VGND.n7729 0.0207703
R7469 VGND.n7741 VGND.n7740 0.0207703
R7470 VGND.n4015 VGND.n4014 0.0207703
R7471 VGND.n4089 VGND.n4016 0.0207703
R7472 VGND.n3111 VGND.n3110 0.0207703
R7473 VGND.n3136 VGND.n3135 0.0207703
R7474 VGND.n3784 VGND.n3783 0.0207703
R7475 VGND.n3795 VGND.n3794 0.0207703
R7476 VGND.n2949 VGND.n2948 0.0207703
R7477 VGND.n4667 VGND.n2950 0.0207703
R7478 VGND.n4303 VGND.n4302 0.0207703
R7479 VGND.n4347 VGND.n4346 0.0207703
R7480 VGND.n2882 VGND.n2881 0.0207703
R7481 VGND.n2894 VGND.n2893 0.0207703
R7482 VGND.n4330 VGND.n4329 0.0207703
R7483 VGND.n2725 VGND.n2724 0.0207703
R7484 VGND.n4803 VGND.n4802 0.0207703
R7485 VGND.n4814 VGND.n4813 0.0207703
R7486 VGND.n4944 VGND.n4943 0.0207703
R7487 VGND.n2750 VGND.n2749 0.0207703
R7488 VGND.n2825 VGND.n2751 0.0207703
R7489 VGND.n1541 VGND.n1540 0.0207703
R7490 VGND.n1549 VGND.n1542 0.0207703
R7491 VGND.n1689 VGND.n1688 0.0207703
R7492 VGND.n1686 VGND.n1685 0.0207703
R7493 VGND.n2527 VGND.n2526 0.0207703
R7494 VGND.n2559 VGND.n2558 0.0207703
R7495 VGND.n5344 VGND.n5343 0.0207703
R7496 VGND.n5361 VGND.n5345 0.0207703
R7497 VGND.n1435 VGND.n1434 0.0207703
R7498 VGND.n2368 VGND.n2367 0.0207703
R7499 VGND.n1860 VGND.n1859 0.0207703
R7500 VGND.n1383 VGND.n1382 0.0207703
R7501 VGND.n5643 VGND.n5642 0.0207703
R7502 VGND.n2325 VGND.n2324 0.0207703
R7503 VGND.n1952 VGND.n1951 0.0207703
R7504 VGND.n5733 VGND.n5732 0.0207703
R7505 VGND.n5681 VGND.n5680 0.0207703
R7506 VGND.n1336 VGND.n1335 0.0207703
R7507 VGND.n1299 VGND.n1298 0.0207703
R7508 VGND.n1303 VGND.n1300 0.0207703
R7509 VGND.n6125 VGND.n6040 0.0207703
R7510 VGND.n6653 VGND.n6652 0.0207703
R7511 VGND.n6715 VGND.n6654 0.0207703
R7512 VGND.n932 VGND.n931 0.0207703
R7513 VGND.n7309 VGND.n933 0.0207703
R7514 VGND.n24 VGND.n23 0.0207703
R7515 VGND.n7901 VGND.n25 0.0207703
R7516 VGND.n7152 VGND.n7151 0.0207703
R7517 VGND.n598 VGND.n597 0.0207703
R7518 VGND.n8006 VGND.n8005 0.0207703
R7519 VGND.n7994 VGND.n7993 0.0207703
R7520 VGND.n6978 VGND.n6977 0.0207703
R7521 VGND.n7029 VGND.n7028 0.0207703
R7522 VGND.n350 VGND.n349 0.0207703
R7523 VGND.n298 VGND.n297 0.0207703
R7524 VGND.n7605 VGND.n7604 0.0204349
R7525 VGND.n4374 VGND.n4373 0.0204349
R7526 VGND.n2170 VGND.n2169 0.0202124
R7527 VGND.n1028 VGND.n1027 0.0202124
R7528 VGND.n1098 VGND.n1097 0.0202124
R7529 VGND.n1084 VGND.n1083 0.0202124
R7530 VGND.n2142 VGND.n2141 0.0202124
R7531 VGND.n2264 VGND.n2263 0.0202124
R7532 VGND.n2013 VGND.n2012 0.0202124
R7533 VGND.n6327 VGND.n6326 0.0202124
R7534 VGND.n3455 VGND.n3454 0.0202124
R7535 VGND.n3526 VGND.n3525 0.0202124
R7536 VGND.n7408 VGND.n7407 0.0202124
R7537 VGND.n165 VGND.n164 0.0202124
R7538 VGND.n260 VGND.n259 0.0202124
R7539 VGND.n698 VGND.n697 0.0202124
R7540 VGND.n42 VGND.n41 0.0202124
R7541 VGND.n7874 VGND.n7873 0.0202124
R7542 VGND.n3338 VGND.n3337 0.0202124
R7543 VGND.n3313 VGND.n3312 0.0202124
R7544 VGND.n7521 VGND.n7520 0.0202124
R7545 VGND.n119 VGND.n118 0.0202124
R7546 VGND.n91 VGND.n90 0.0202124
R7547 VGND.n86 VGND.n85 0.0202124
R7548 VGND.n7856 VGND.n7855 0.0202124
R7549 VGND.n63 VGND.n62 0.0202124
R7550 VGND.n3157 VGND.n3156 0.0202124
R7551 VGND.n4011 VGND.n4010 0.0202124
R7552 VGND.n3095 VGND.n3094 0.0202124
R7553 VGND.n3132 VGND.n3131 0.0202124
R7554 VGND.n3735 VGND.n3734 0.0202124
R7555 VGND.n3670 VGND.n3669 0.0202124
R7556 VGND.n3648 VGND.n3647 0.0202124
R7557 VGND.n3905 VGND.n3904 0.0202124
R7558 VGND.n4632 VGND.n4631 0.0202124
R7559 VGND.n2952 VGND.n2951 0.0202124
R7560 VGND.n4287 VGND.n4286 0.0202124
R7561 VGND.n4343 VGND.n4342 0.0202124
R7562 VGND.n4224 VGND.n4223 0.0202124
R7563 VGND.n2889 VGND.n2888 0.0202124
R7564 VGND.n4507 VGND.n4506 0.0202124
R7565 VGND.n3090 VGND.n3089 0.0202124
R7566 VGND.n4314 VGND.n4313 0.0202124
R7567 VGND.n2721 VGND.n2720 0.0202124
R7568 VGND.n4698 VGND.n4697 0.0202124
R7569 VGND.n2876 VGND.n2875 0.0202124
R7570 VGND.n2859 VGND.n2858 0.0202124
R7571 VGND.n2863 VGND.n2862 0.0202124
R7572 VGND.n2837 VGND.n2836 0.0202124
R7573 VGND.n5050 VGND.n5049 0.0202124
R7574 VGND.n5219 VGND.n5218 0.0202124
R7575 VGND.n1476 VGND.n1475 0.0202124
R7576 VGND.n2383 VGND.n2382 0.0202124
R7577 VGND.n2459 VGND.n2458 0.0202124
R7578 VGND.n1466 VGND.n1465 0.0202124
R7579 VGND.n5347 VGND.n5346 0.0202124
R7580 VGND.n1418 VGND.n1417 0.0202124
R7581 VGND.n1443 VGND.n1442 0.0202124
R7582 VGND.n1695 VGND.n1694 0.0202124
R7583 VGND.n1864 VGND.n1863 0.0202124
R7584 VGND.n2437 VGND.n2436 0.0202124
R7585 VGND.n5657 VGND.n5656 0.0202124
R7586 VGND.n1908 VGND.n1907 0.0202124
R7587 VGND.n1956 VGND.n1955 0.0202124
R7588 VGND.n5663 VGND.n5662 0.0202124
R7589 VGND.n5688 VGND.n5687 0.0202124
R7590 VGND.n1331 VGND.n1330 0.0202124
R7591 VGND.n1325 VGND.n1324 0.0202124
R7592 VGND.n5994 VGND.n5993 0.0202124
R7593 VGND.n6022 VGND.n6021 0.0202124
R7594 VGND.n1186 VGND.n1185 0.0202124
R7595 VGND.n1205 VGND.n1204 0.0202124
R7596 VGND.n6155 VGND.n6154 0.0202124
R7597 VGND.n6145 VGND.n6144 0.0202124
R7598 VGND.n1049 VGND.n1048 0.0202124
R7599 VGND.n6649 VGND.n6648 0.0202124
R7600 VGND.n7264 VGND.n7263 0.0202124
R7601 VGND.n7303 VGND.n7302 0.0202124
R7602 VGND.n462 VGND.n461 0.0202124
R7603 VGND.n34 VGND.n33 0.0202124
R7604 VGND.n965 VGND.n964 0.0202124
R7605 VGND.n7146 VGND.n7145 0.0202124
R7606 VGND.n588 VGND.n587 0.0202124
R7607 VGND.n426 VGND.n425 0.0202124
R7608 VGND.n7414 VGND.n7413 0.0202124
R7609 VGND.n8013 VGND.n8012 0.0202124
R7610 VGND.n6818 VGND.n6817 0.0202124
R7611 VGND.n6981 VGND.n6980 0.0202124
R7612 VGND.n7021 VGND.n7020 0.0202124
R7613 VGND.n274 VGND.n273 0.0202124
R7614 VGND.n385 VGND.n384 0.0202124
R7615 VGND.n1111 VGND.n1110 0.0202124
R7616 VGND.n6 VGND.n5 0.0200989
R7617 VGND.n782 VGND 0.0200312
R7618 VGND VGND.n816 0.0200312
R7619 VGND VGND.n3423 0.0200312
R7620 VGND.n3464 VGND.n3463 0.0200312
R7621 VGND.n3540 VGND.n3539 0.0200312
R7622 VGND VGND.n7666 0.0200312
R7623 VGND VGND.n7756 0.0200312
R7624 VGND.n7831 VGND 0.0200312
R7625 VGND.n7832 VGND.n7831 0.0200312
R7626 VGND.n3332 VGND.n3331 0.0200312
R7627 VGND.n3327 VGND.n3326 0.0200312
R7628 VGND.n4153 VGND 0.0200312
R7629 VGND.n4108 VGND.n4107 0.0200312
R7630 VGND.n4129 VGND.n4128 0.0200312
R7631 VGND.n4019 VGND.n4018 0.0200312
R7632 VGND.n4652 VGND.n4651 0.0200312
R7633 VGND.n4680 VGND.n4679 0.0200312
R7634 VGND.n4675 VGND.n4674 0.0200312
R7635 VGND VGND.n5101 0.0200312
R7636 VGND VGND.n4914 0.0200312
R7637 VGND.n5060 VGND.n5059 0.0200312
R7638 VGND.n2754 VGND.n2753 0.0200312
R7639 VGND.n5185 VGND 0.0200312
R7640 VGND.n5309 VGND.n1574 0.0200312
R7641 VGND.n1559 VGND.n1558 0.0200312
R7642 VGND.n5339 VGND.n5338 0.0200312
R7643 VGND.n5427 VGND.n5426 0.0200312
R7644 VGND VGND.n1875 0.0200312
R7645 VGND VGND.n5714 0.0200312
R7646 VGND.n5988 VGND.n1317 0.0200312
R7647 VGND.n1313 VGND.n1312 0.0200312
R7648 VGND.n6321 VGND 0.0200312
R7649 VGND.n6305 VGND.n6304 0.0200312
R7650 VGND.n6233 VGND.n6232 0.0200312
R7651 VGND.n6111 VGND.n6110 0.0200312
R7652 VGND.n6116 VGND.n6115 0.0200312
R7653 VGND VGND.n6853 0.0200312
R7654 VGND.n7123 VGND.n7122 0.0200312
R7655 VGND.n7324 VGND.n7323 0.0200312
R7656 VGND.n7319 VGND.n7318 0.0200312
R7657 VGND.n891 VGND 0.0200312
R7658 VGND VGND.n2191 0.0200312
R7659 VGND.n6738 VGND.n6737 0.0200312
R7660 VGND.n6758 VGND.n6757 0.0200312
R7661 VGND.n552 VGND 0.0200312
R7662 VGND.n7965 VGND.n7964 0.0200312
R7663 VGND.n7960 VGND.n7959 0.0200312
R7664 VGND.n818 VGND 0.0199818
R7665 VGND.n7513 VGND.n7512 0.0195896
R7666 VGND.n7612 VGND.n7611 0.0195896
R7667 VGND.n4216 VGND.n4215 0.0195896
R7668 VGND.n4382 VGND.n4381 0.0195896
R7669 VGND.n5157 VGND.n5156 0.0195896
R7670 VGND.n2344 VGND.n2342 0.0195896
R7671 VGND.n2300 VGND.n2298 0.0195896
R7672 VGND.n8000 VGND.n7999 0.0195896
R7673 VGND.n6904 VGND.n6903 0.0193669
R7674 VGND.n6338 VGND.n6337 0.0190811
R7675 VGND.n6437 VGND.n6436 0.0190811
R7676 VGND.n6811 VGND.n6810 0.0190811
R7677 VGND.n6832 VGND.n6831 0.0190811
R7678 VGND.n6885 VGND.n6884 0.0190811
R7679 VGND.n6898 VGND.n6897 0.0190811
R7680 VGND.n2208 VGND.n2207 0.0190811
R7681 VGND.n2174 VGND.n2173 0.0190811
R7682 VGND.n2241 VGND.n2240 0.0190811
R7683 VGND.n2248 VGND.n2247 0.0190811
R7684 VGND.n2154 VGND.n2153 0.0190811
R7685 VGND.n2158 VGND.n2157 0.0190811
R7686 VGND.n2285 VGND.n2147 0.0190811
R7687 VGND.n2271 VGND.n2270 0.0190811
R7688 VGND.n2017 VGND.n1993 0.0190811
R7689 VGND.n2005 VGND.n2004 0.0190811
R7690 VGND.n6324 VGND.n1119 0.0190811
R7691 VGND.n3524 VGND.n3523 0.0190811
R7692 VGND.n158 VGND.n157 0.0190811
R7693 VGND.n7405 VGND.n7397 0.0190811
R7694 VGND.n7495 VGND.n7494 0.0190811
R7695 VGND.n7481 VGND.n7480 0.0190811
R7696 VGND.n722 VGND.n721 0.0190811
R7697 VGND.n264 VGND.n263 0.0190811
R7698 VGND.n737 VGND.n736 0.0190811
R7699 VGND.n814 VGND.n43 0.0190811
R7700 VGND.n3360 VGND.n3359 0.0190811
R7701 VGND.n3311 VGND.n3310 0.0190811
R7702 VGND.n7551 VGND.n7550 0.0190811
R7703 VGND.n7525 VGND.n7524 0.0190811
R7704 VGND.n7529 VGND.n7528 0.0190811
R7705 VGND.n7536 VGND.n7535 0.0190811
R7706 VGND.n7731 VGND.n7730 0.0190811
R7707 VGND.n95 VGND.n94 0.0190811
R7708 VGND.n7717 VGND.n105 0.0190811
R7709 VGND.n7859 VGND.n7858 0.0190811
R7710 VGND.n59 VGND.n58 0.0190811
R7711 VGND.n4016 VGND.n4015 0.0190811
R7712 VGND.n3125 VGND.n3124 0.0190811
R7713 VGND.n3099 VGND.n3098 0.0190811
R7714 VGND.n3103 VGND.n3102 0.0190811
R7715 VGND.n3110 VGND.n3109 0.0190811
R7716 VGND.n3785 VGND.n3784 0.0190811
R7717 VGND.n3739 VGND.n3738 0.0190811
R7718 VGND.n3756 VGND.n3755 0.0190811
R7719 VGND.n3651 VGND.n3650 0.0190811
R7720 VGND.n3640 VGND.n3639 0.0190811
R7721 VGND.n2950 VGND.n2949 0.0190811
R7722 VGND.n4284 VGND.n4283 0.0190811
R7723 VGND.n4291 VGND.n4290 0.0190811
R7724 VGND.n4295 VGND.n4294 0.0190811
R7725 VGND.n4302 VGND.n4301 0.0190811
R7726 VGND.n2883 VGND.n2882 0.0190811
R7727 VGND.n4228 VGND.n4227 0.0190811
R7728 VGND.n4489 VGND.n4238 0.0190811
R7729 VGND.n4510 VGND.n4509 0.0190811
R7730 VGND.n3086 VGND.n3085 0.0190811
R7731 VGND.n5118 VGND.n5117 0.0190811
R7732 VGND.n4318 VGND.n4317 0.0190811
R7733 VGND.n4322 VGND.n4321 0.0190811
R7734 VGND.n4329 VGND.n4328 0.0190811
R7735 VGND.n4804 VGND.n4803 0.0190811
R7736 VGND.n4702 VGND.n4701 0.0190811
R7737 VGND.n4790 VGND.n4712 0.0190811
R7738 VGND.n4912 VGND.n2857 0.0190811
R7739 VGND.n4931 VGND.n4930 0.0190811
R7740 VGND.n2751 VGND.n2750 0.0190811
R7741 VGND.n5226 VGND.n5225 0.0190811
R7742 VGND.n5247 VGND.n5246 0.0190811
R7743 VGND.n1542 VGND.n1541 0.0190811
R7744 VGND.n2399 VGND.n2398 0.0190811
R7745 VGND.n2714 VGND.n2389 0.0190811
R7746 VGND.n1688 VGND.n1687 0.0190811
R7747 VGND.n2527 VGND.n2525 0.0190811
R7748 VGND.n1670 VGND.n1669 0.0190811
R7749 VGND.n2548 VGND.n2547 0.0190811
R7750 VGND.n5345 VGND.n5344 0.0190811
R7751 VGND.n1433 VGND.n1432 0.0190811
R7752 VGND.n1422 VGND.n1421 0.0190811
R7753 VGND.n1725 VGND.n1724 0.0190811
R7754 VGND.n1746 VGND.n1745 0.0190811
R7755 VGND.n2360 VGND.n1698 0.0190811
R7756 VGND.n2367 VGND.n2366 0.0190811
R7757 VGND.n1384 VGND.n1383 0.0190811
R7758 VGND.n2441 VGND.n2440 0.0190811
R7759 VGND.n5654 VGND.n1394 0.0190811
R7760 VGND.n1901 VGND.n1900 0.0190811
R7761 VGND.n1919 VGND.n1918 0.0190811
R7762 VGND.n2317 VGND.n1910 0.0190811
R7763 VGND.n2324 VGND.n2323 0.0190811
R7764 VGND.n5733 VGND.n5731 0.0190811
R7765 VGND.n5673 VGND.n5672 0.0190811
R7766 VGND.n5707 VGND.n5706 0.0190811
R7767 VGND.n1334 VGND.n1333 0.0190811
R7768 VGND.n1344 VGND.n1343 0.0190811
R7769 VGND.n1300 VGND.n1299 0.0190811
R7770 VGND.n1192 VGND.n1191 0.0190811
R7771 VGND.n1212 VGND.n1211 0.0190811
R7772 VGND.n6040 VGND.n6039 0.0190811
R7773 VGND.n6654 VGND.n6653 0.0190811
R7774 VGND.n933 VGND.n932 0.0190811
R7775 VGND.n25 VGND.n24 0.0190811
R7776 VGND.n951 VGND.n950 0.0190811
R7777 VGND.n948 VGND.n947 0.0190811
R7778 VGND.n596 VGND.n595 0.0190811
R7779 VGND.n7423 VGND.n7422 0.0190811
R7780 VGND.n7464 VGND.n7426 0.0190811
R7781 VGND.n7466 VGND.n1 0.0190811
R7782 VGND.n8005 VGND.n2 0.0190811
R7783 VGND.n6984 VGND.n6978 0.0190811
R7784 VGND.n986 VGND.n985 0.0190811
R7785 VGND.n7018 VGND.n1002 0.0190811
R7786 VGND.n354 VGND.n350 0.0190811
R7787 VGND.n283 VGND.n282 0.0190811
R7788 VGND.n3366 VGND 0.0188432
R7789 VGND.n7401 VGND.n7398 0.0187292
R7790 VGND.n255 VGND.n254 0.0187292
R7791 VGND.n816 VGND 0.0187292
R7792 VGND.n7881 VGND.n45 0.0187292
R7793 VGND.n3370 VGND.n3368 0.0187292
R7794 VGND.n7596 VGND.n7592 0.0187292
R7795 VGND.n7710 VGND.n7709 0.0187292
R7796 VGND.n7840 VGND.n7839 0.0187292
R7797 VGND.n3176 VGND.n69 0.0187292
R7798 VGND VGND.n3177 0.0187292
R7799 VGND.n4194 VGND.n4192 0.0187292
R7800 VGND VGND.n3876 0.0187292
R7801 VGND.n3885 VGND.n3884 0.0187292
R7802 VGND.n3922 VGND.n3921 0.0187292
R7803 VGND.n4280 VGND 0.0187292
R7804 VGND.n4365 VGND.n4363 0.0187292
R7805 VGND.n4481 VGND.n4480 0.0187292
R7806 VGND.n4534 VGND.n4533 0.0187292
R7807 VGND.n4548 VGND.n4546 0.0187292
R7808 VGND.n4549 VGND 0.0187292
R7809 VGND.n5135 VGND.n5132 0.0187292
R7810 VGND.n4782 VGND.n4781 0.0187292
R7811 VGND.n4914 VGND 0.0187292
R7812 VGND.n4964 VGND.n4962 0.0187292
R7813 VGND.n2393 VGND.n2391 0.0187292
R7814 VGND.n2543 VGND.n2541 0.0187292
R7815 VGND.n5264 VGND.n5263 0.0187292
R7816 VGND.n5279 VGND.n5278 0.0187292
R7817 VGND.n1731 VGND 0.0187292
R7818 VGND.n1741 VGND.n1699 0.0187292
R7819 VGND.n1766 VGND.n1395 0.0187292
R7820 VGND.n5537 VGND.n5536 0.0187292
R7821 VGND.n5528 VGND.n5526 0.0187292
R7822 VGND.n5524 VGND 0.0187292
R7823 VGND.n1914 VGND.n1911 0.0187292
R7824 VGND.n5713 VGND.n5711 0.0187292
R7825 VGND.n5885 VGND.n5884 0.0187292
R7826 VGND.n5899 VGND.n5897 0.0187292
R7827 VGND VGND.n5901 0.0187292
R7828 VGND.n2151 VGND.n2149 0.0187292
R7829 VGND.n6241 VGND.n6240 0.0187292
R7830 VGND.n6227 VGND.n6226 0.0187292
R7831 VGND.n6224 VGND 0.0187292
R7832 VGND.n6871 VGND.n6869 0.0187292
R7833 VGND.n7012 VGND.n7010 0.0187292
R7834 VGND.n7166 VGND.n7164 0.0187292
R7835 VGND.n2220 VGND.n2218 0.0187292
R7836 VGND.n6418 VGND.n6416 0.0187292
R7837 VGND.n6563 VGND.n6562 0.0187292
R7838 VGND.n6579 VGND.n6578 0.0187292
R7839 VGND VGND.n6580 0.0187292
R7840 VGND.n7460 VGND.n7458 0.0187292
R7841 VGND.n381 VGND.n380 0.0187292
R7842 VGND.n571 VGND.n570 0.0187292
R7843 VGND.n562 VGND.n561 0.0187292
R7844 VGND.n558 VGND 0.0187292
R7845 VGND.n2415 VGND 0.0179232
R7846 VGND.n7830 VGND.n7828 0.0174271
R7847 VGND.n3875 VGND.n3873 0.0174271
R7848 VGND.n2972 VGND.n2971 0.0174271
R7849 VGND.n4916 VGND.n4915 0.0174271
R7850 VGND.n2631 VGND.n2630 0.0174271
R7851 VGND.n5561 VGND.n5559 0.0174271
R7852 VGND.n1358 VGND.n1357 0.0174271
R7853 VGND.n6231 VGND.n6229 0.0174271
R7854 VGND.n7126 VGND.n7125 0.0174271
R7855 VGND.n6538 VGND.n6537 0.0174271
R7856 VGND.n415 VGND.n414 0.0174271
R7857 VGND.n6436 VGND.n6435 0.0173919
R7858 VGND.n6833 VGND.n6832 0.0173919
R7859 VGND.n2175 VGND.n2174 0.0173919
R7860 VGND.n2158 VGND.n2146 0.0173919
R7861 VGND.n2004 VGND.n2003 0.0173919
R7862 VGND.n3452 VGND.n3451 0.0173919
R7863 VGND.n7406 VGND.n7405 0.0173919
R7864 VGND.n263 VGND.n262 0.0173919
R7865 VGND.n3166 VGND.n3165 0.0173919
R7866 VGND.n7526 VGND.n7525 0.0173919
R7867 VGND.n94 VGND.n93 0.0173919
R7868 VGND.n3617 VGND.n3616 0.0173919
R7869 VGND.n3100 VGND.n3099 0.0173919
R7870 VGND.n3738 VGND.n3737 0.0173919
R7871 VGND.n4625 VGND.n4624 0.0173919
R7872 VGND.n4292 VGND.n4291 0.0173919
R7873 VGND.n4227 VGND.n4226 0.0173919
R7874 VGND.n4319 VGND.n4318 0.0173919
R7875 VGND.n4701 VGND.n4700 0.0173919
R7876 VGND.n2831 VGND.n2830 0.0173919
R7877 VGND.n1480 VGND.n1479 0.0173919
R7878 VGND.n2399 VGND.n2388 0.0173919
R7879 VGND.n1669 VGND.n1668 0.0173919
R7880 VGND.n1463 VGND.n1462 0.0173919
R7881 VGND.n1746 VGND.n1696 0.0173919
R7882 VGND.n2440 VGND.n2439 0.0173919
R7883 VGND.n1919 VGND.n1909 0.0173919
R7884 VGND.n5672 VGND.n5671 0.0173919
R7885 VGND.n1251 VGND.n1250 0.0173919
R7886 VGND.n6100 VGND.n6099 0.0173919
R7887 VGND.n1054 VGND.n1053 0.0173919
R7888 VGND.n939 VGND.n938 0.0173919
R7889 VGND.n455 VGND.n454 0.0173919
R7890 VGND.n7465 VGND.n7464 0.0173919
R7891 VGND.n282 VGND.n281 0.0173919
R7892 VGND.n4655 VGND.n4653 0.017391
R7893 VGND.n2535 VGND.n2534 0.0173894
R7894 VGND.n7957 VGND.n18 0.0172667
R7895 VGND.n3564 VGND.n3563 0.0172634
R7896 VGND.n6731 VGND.n6730 0.0172634
R7897 VGND.n6314 VGND.n6313 0.0172616
R7898 VGND.n6760 VGND.n6759 0.0170064
R7899 VGND.n6760 VGND.n1044 0.0168883
R7900 VGND.n2211 VGND.n2210 0.0168788
R7901 VGND.n6802 VGND.n1029 0.0168788
R7902 VGND.n6549 VGND.n1099 0.0168788
R7903 VGND.n6554 VGND.n1085 0.0168788
R7904 VGND.n3571 VGND.n3341 0.0168788
R7905 VGND.n3529 VGND.n3527 0.0168788
R7906 VGND.n161 VGND.n160 0.0168788
R7907 VGND.n7516 VGND.n166 0.0168788
R7908 VGND.n724 VGND.n723 0.0168788
R7909 VGND.n716 VGND.n699 0.0168788
R7910 VGND.n824 VGND.n823 0.0168788
R7911 VGND.n3353 VGND.n3351 0.0168788
R7912 VGND.n3609 VGND.n3160 0.0168788
R7913 VGND.n3316 VGND.n3314 0.0168788
R7914 VGND.n7554 VGND.n7553 0.0168788
R7915 VGND.n7559 VGND.n120 0.0168788
R7916 VGND.n7733 VGND.n7732 0.0168788
R7917 VGND.n7738 VGND.n87 0.0168788
R7918 VGND.n7821 VGND.n7820 0.0168788
R7919 VGND.n7852 VGND.n66 0.0168788
R7920 VGND.n4095 VGND.n4094 0.0168788
R7921 VGND.n4090 VGND.n4012 0.0168788
R7922 VGND.n3128 VGND.n3127 0.0168788
R7923 VGND.n4219 VGND.n3133 0.0168788
R7924 VGND.n3787 VGND.n3786 0.0168788
R7925 VGND.n3792 VGND.n3671 0.0168788
R7926 VGND.n3866 VGND.n3865 0.0168788
R7927 VGND.n3899 VGND.n3896 0.0168788
R7928 VGND.n4662 VGND.n2958 0.0168788
R7929 VGND.n4666 VGND.n2953 0.0168788
R7930 VGND.n4356 VGND.n4355 0.0168788
R7931 VGND.n4351 VGND.n4344 0.0168788
R7932 VGND.n2885 VGND.n2884 0.0168788
R7933 VGND.n4693 VGND.n2890 0.0168788
R7934 VGND.n3075 VGND.n3074 0.0168788
R7935 VGND.n4523 VGND.n2968 0.0168788
R7936 VGND.n5121 VGND.n5120 0.0168788
R7937 VGND.n5160 VGND.n2722 0.0168788
R7938 VGND.n4806 VGND.n4805 0.0168788
R7939 VGND.n4811 VGND.n2877 0.0168788
R7940 VGND.n4924 VGND.n4923 0.0168788
R7941 VGND.n2870 VGND.n2864 0.0168788
R7942 VGND.n5045 VGND.n5044 0.0168788
R7943 VGND.n2826 VGND.n2748 0.0168788
R7944 VGND.n5356 VGND.n5352 0.0168788
R7945 VGND.n5360 VGND.n5348 0.0168788
R7946 VGND.n5554 VGND.n5553 0.0168788
R7947 VGND.n5549 VGND.n1444 0.0168788
R7948 VGND.n1728 VGND.n1727 0.0168788
R7949 VGND.n2339 VGND.n1865 0.0168788
R7950 VGND.n1386 VGND.n1385 0.0168788
R7951 VGND.n5640 VGND.n5638 0.0168788
R7952 VGND.n1904 VGND.n1903 0.0168788
R7953 VGND.n2295 VGND.n1957 0.0168788
R7954 VGND.n5730 VGND.n5729 0.0168788
R7955 VGND.n5691 VGND.n5689 0.0168788
R7956 VGND.n5869 VGND.n5868 0.0168788
R7957 VGND.n5874 VGND.n1326 0.0168788
R7958 VGND.n6016 VGND.n6015 0.0168788
R7959 VGND.n1302 VGND.n1301 0.0168788
R7960 VGND.n6721 VGND.n6720 0.0168788
R7961 VGND.n6716 VGND.n6650 0.0168788
R7962 VGND.n7266 VGND.n7265 0.0168788
R7963 VGND.n7308 VGND.n934 0.0168788
R7964 VGND.n489 VGND.n488 0.0168788
R7965 VGND.n7900 VGND.n35 0.0168788
R7966 VGND.n7136 VGND.n966 0.0168788
R7967 VGND.n7141 VGND.n7138 0.0168788
R7968 VGND.n608 VGND.n607 0.0168788
R7969 VGND.n584 VGND.n427 0.0168788
R7970 VGND.n7412 VGND.n7411 0.0168788
R7971 VGND.n8011 VGND.n8010 0.0168788
R7972 VGND.n6815 VGND.n6814 0.0168788
R7973 VGND.n6825 VGND.n6819 0.0168788
R7974 VGND.n6983 VGND.n6982 0.0168788
R7975 VGND.n7026 VGND.n981 0.0168788
R7976 VGND.n353 VGND.n352 0.0168788
R7977 VGND.n691 VGND.n294 0.0168788
R7978 VGND.n6341 VGND.n6340 0.0168788
R7979 VGND.n6450 VGND.n1112 0.0168788
R7980 VGND.n4672 VGND.n4670 0.0166396
R7981 VGND.n7958 VGND.n7957 0.016628
R7982 VGND.n3565 VGND.n3564 0.0166244
R7983 VGND.n6730 VGND.n1058 0.0166244
R7984 VGND.n6313 VGND.n6312 0.0166226
R7985 VGND.n6798 VGND 0.0166211
R7986 VGND.n4656 VGND.n4655 0.0164962
R7987 VGND.n2534 VGND.n2533 0.0164946
R7988 VGND.n233 VGND.n231 0.016464
R7989 VGND.n7688 VGND.n7686 0.016464
R7990 VGND.n3780 VGND.n3779 0.016464
R7991 VGND.n4461 VGND.n4239 0.016464
R7992 VGND.n4759 VGND.n4757 0.016464
R7993 VGND.n2516 VGND.n2515 0.016464
R7994 VGND.n1783 VGND.n1782 0.016464
R7995 VGND.n5740 VGND.n5739 0.016464
R7996 VGND.n2024 VGND.n2023 0.016464
R7997 VGND.n6989 VGND.n6987 0.016464
R7998 VGND.n6395 VGND.n6393 0.016464
R7999 VGND.n359 VGND.n357 0.016464
R8000 VGND.n4673 VGND.n4672 0.0162568
R8001 VGND.n7503 VGND.n7502 0.016125
R8002 VGND.n7506 VGND.n7505 0.016125
R8003 VGND.n706 VGND 0.016125
R8004 VGND.n712 VGND.n711 0.016125
R8005 VGND.n811 VGND.n809 0.016125
R8006 VGND.n3537 VGND.n3534 0.016125
R8007 VGND.n7607 VGND.n7606 0.016125
R8008 VGND.n7610 VGND.n7609 0.016125
R8009 VGND VGND.n7711 0.016125
R8010 VGND.n7745 VGND.n7744 0.016125
R8011 VGND.n7837 VGND.n7835 0.016125
R8012 VGND.n7841 VGND.n7840 0.016125
R8013 VGND.n3324 VGND.n3320 0.016125
R8014 VGND.n4210 VGND.n4209 0.016125
R8015 VGND.n4213 VGND.n4212 0.016125
R8016 VGND.n3731 VGND 0.016125
R8017 VGND.n3799 VGND.n3798 0.016125
R8018 VGND.n3882 VGND.n3880 0.016125
R8019 VGND.n4025 VGND.n4024 0.016125
R8020 VGND.n4087 VGND 0.016125
R8021 VGND.n4376 VGND.n4375 0.016125
R8022 VGND.n4379 VGND.n4378 0.016125
R8023 VGND VGND.n4484 0.016125
R8024 VGND.n4689 VGND.n4688 0.016125
R8025 VGND.n4531 VGND.n4529 0.016125
R8026 VGND.n4535 VGND.n4534 0.016125
R8027 VGND.n5128 VGND 0.016125
R8028 VGND.n5151 VGND.n5150 0.016125
R8029 VGND.n5154 VGND.n5153 0.016125
R8030 VGND VGND.n4785 0.016125
R8031 VGND.n4819 VGND.n4817 0.016125
R8032 VGND VGND.n4950 0.016125
R8033 VGND.n4952 VGND.n4951 0.016125
R8034 VGND.n2760 VGND.n2759 0.016125
R8035 VGND VGND.n2760 0.016125
R8036 VGND.n2703 VGND.n2701 0.016125
R8037 VGND.n2699 VGND.n2698 0.016125
R8038 VGND.n2544 VGND 0.016125
R8039 VGND.n2564 VGND.n2562 0.016125
R8040 VGND.n5262 VGND.n5261 0.016125
R8041 VGND.n5265 VGND.n5264 0.016125
R8042 VGND.n1556 VGND.n1552 0.016125
R8043 VGND.n2350 VGND.n2348 0.016125
R8044 VGND.n2346 VGND.n2345 0.016125
R8045 VGND VGND.n5648 0.016125
R8046 VGND.n5635 VGND.n5634 0.016125
R8047 VGND.n5534 VGND.n5532 0.016125
R8048 VGND.n5538 VGND.n5537 0.016125
R8049 VGND.n5424 VGND.n5420 0.016125
R8050 VGND.n5420 VGND 0.016125
R8051 VGND.n2302 VGND.n2301 0.016125
R8052 VGND.n5697 VGND 0.016125
R8053 VGND.n5684 VGND.n5683 0.016125
R8054 VGND.n5882 VGND.n5880 0.016125
R8055 VGND.n5886 VGND.n5885 0.016125
R8056 VGND.n1310 VGND.n1307 0.016125
R8057 VGND.n2162 VGND.n2161 0.016125
R8058 VGND.n6291 VGND.n6290 0.016125
R8059 VGND.n6238 VGND.n6236 0.016125
R8060 VGND.n6242 VGND.n6241 0.016125
R8061 VGND.n6122 VGND.n6120 0.016125
R8062 VGND.n7016 VGND 0.016125
R8063 VGND.n7033 VGND.n7032 0.016125
R8064 VGND.n7120 VGND.n7117 0.016125
R8065 VGND.n7115 VGND 0.016125
R8066 VGND.n7154 VGND.n7153 0.016125
R8067 VGND.n7316 VGND.n7312 0.016125
R8068 VGND VGND.n2176 0.016125
R8069 VGND.n2230 VGND.n2228 0.016125
R8070 VGND.n2226 VGND.n1035 0.016125
R8071 VGND VGND.n6422 0.016125
R8072 VGND.n6458 VGND.n6456 0.016125
R8073 VGND.n6561 VGND.n6560 0.016125
R8074 VGND.n6564 VGND.n6563 0.016125
R8075 VGND.n687 VGND.n686 0.016125
R8076 VGND.n568 VGND.n566 0.016125
R8077 VGND.n572 VGND.n571 0.016125
R8078 VGND.n1069 VGND.n1068 0.0157027
R8079 VGND.n3359 VGND.n3358 0.0157027
R8080 VGND.n58 VGND.n57 0.0157027
R8081 VGND.n3639 VGND.n3638 0.0157027
R8082 VGND.n3085 VGND.n3084 0.0157027
R8083 VGND.n5246 VGND.n5245 0.0157027
R8084 VGND.n1211 VGND.n1210 0.0157027
R8085 VGND.n947 VGND.n946 0.0157027
R8086 VGND.n430 VGND.n429 0.0157027
R8087 VGND.n7404 VGND.n7402 0.0148229
R8088 VGND.n7496 VGND 0.0148229
R8089 VGND.n7504 VGND.n7503 0.0148229
R8090 VGND.n240 VGND.n239 0.0148229
R8091 VGND.n738 VGND.n256 0.0148229
R8092 VGND.n713 VGND.n707 0.0148229
R8093 VGND.n813 VGND.n812 0.0148229
R8094 VGND.n3362 VGND.n3361 0.0148229
R8095 VGND.n3559 VGND 0.0148229
R8096 VGND.n3538 VGND.n3537 0.0148229
R8097 VGND.n7598 VGND.n7597 0.0148229
R8098 VGND.n7601 VGND.n7600 0.0148229
R8099 VGND.n7608 VGND.n7607 0.0148229
R8100 VGND.n7695 VGND.n7694 0.0148229
R8101 VGND.n7716 VGND.n7712 0.0148229
R8102 VGND.n7743 VGND.n81 0.0148229
R8103 VGND.n7833 VGND.n7832 0.0148229
R8104 VGND.n7845 VGND.n7844 0.0148229
R8105 VGND.n3592 VGND 0.0148229
R8106 VGND.n3325 VGND.n3324 0.0148229
R8107 VGND.n4196 VGND.n4195 0.0148229
R8108 VGND.n4199 VGND.n4198 0.0148229
R8109 VGND.n4211 VGND.n4210 0.0148229
R8110 VGND.n3772 VGND.n3771 0.0148229
R8111 VGND.n3757 VGND.n3731 0.0148229
R8112 VGND.n3797 VGND.n3667 0.0148229
R8113 VGND.n3878 VGND.n3877 0.0148229
R8114 VGND.n3913 VGND.n3912 0.0148229
R8115 VGND VGND.n4110 0.0148229
R8116 VGND.n4024 VGND.n4020 0.0148229
R8117 VGND.n4367 VGND.n4366 0.0148229
R8118 VGND.n4370 VGND.n4369 0.0148229
R8119 VGND.n4377 VGND.n4376 0.0148229
R8120 VGND.n4468 VGND.n4467 0.0148229
R8121 VGND.n4488 VGND.n4485 0.0148229
R8122 VGND.n4690 VGND.n2895 0.0148229
R8123 VGND.n4527 VGND.n4526 0.0148229
R8124 VGND.n4539 VGND.n4538 0.0148229
R8125 VGND.n4649 VGND 0.0148229
R8126 VGND.n5137 VGND.n5136 0.0148229
R8127 VGND.n5140 VGND.n5139 0.0148229
R8128 VGND.n5152 VGND.n5151 0.0148229
R8129 VGND.n4766 VGND.n4765 0.0148229
R8130 VGND.n4789 VGND.n4786 0.0148229
R8131 VGND.n4816 VGND.n2873 0.0148229
R8132 VGND.n4911 VGND.n4910 0.0148229
R8133 VGND.n4956 VGND.n4955 0.0148229
R8134 VGND.n2844 VGND 0.0148229
R8135 VGND.n2759 VGND.n2755 0.0148229
R8136 VGND.n2400 VGND.n2394 0.0148229
R8137 VGND VGND.n2713 0.0148229
R8138 VGND.n2701 VGND.n2700 0.0148229
R8139 VGND.n2532 VGND.n2531 0.0148229
R8140 VGND.n2546 VGND.n2544 0.0148229
R8141 VGND.n2561 VGND.n2551 0.0148229
R8142 VGND.n5259 VGND.n5258 0.0148229
R8143 VGND.n5269 VGND.n5268 0.0148229
R8144 VGND.n1582 VGND 0.0148229
R8145 VGND.n1557 VGND.n1556 0.0148229
R8146 VGND.n1747 VGND.n1742 0.0148229
R8147 VGND VGND.n2359 0.0148229
R8148 VGND.n2348 VGND.n2347 0.0148229
R8149 VGND.n1776 VGND.n1775 0.0148229
R8150 VGND.n5653 VGND.n5649 0.0148229
R8151 VGND.n5646 VGND.n5645 0.0148229
R8152 VGND.n5530 VGND.n5529 0.0148229
R8153 VGND.n5542 VGND.n5541 0.0148229
R8154 VGND.n5441 VGND 0.0148229
R8155 VGND.n5425 VGND.n5424 0.0148229
R8156 VGND.n1920 VGND.n1915 0.0148229
R8157 VGND VGND.n2316 0.0148229
R8158 VGND.n2304 VGND.n2303 0.0148229
R8159 VGND.n5674 VGND.n5669 0.0148229
R8160 VGND.n5709 VGND.n5697 0.0148229
R8161 VGND.n5685 VGND.n5682 0.0148229
R8162 VGND.n5878 VGND.n5877 0.0148229
R8163 VGND.n5890 VGND.n5889 0.0148229
R8164 VGND.n6001 VGND 0.0148229
R8165 VGND.n1311 VGND.n1310 0.0148229
R8166 VGND.n2159 VGND.n2152 0.0148229
R8167 VGND VGND.n2284 0.0148229
R8168 VGND.n2272 VGND.n2163 0.0148229
R8169 VGND.n6311 VGND.n6310 0.0148229
R8170 VGND.n6323 VGND.n6305 0.0148229
R8171 VGND.n6303 VGND.n6302 0.0148229
R8172 VGND.n6234 VGND.n6233 0.0148229
R8173 VGND.n6246 VGND.n6245 0.0148229
R8174 VGND VGND.n6102 0.0148229
R8175 VGND.n6120 VGND.n6117 0.0148229
R8176 VGND.n6873 VGND.n6872 0.0148229
R8177 VGND.n6876 VGND.n6875 0.0148229
R8178 VGND.n6899 VGND.n1020 0.0148229
R8179 VGND.n6996 VGND.n6995 0.0148229
R8180 VGND.n7017 VGND.n7016 0.0148229
R8181 VGND.n7031 VGND.n978 0.0148229
R8182 VGND.n7122 VGND.n7121 0.0148229
R8183 VGND.n7158 VGND.n7157 0.0148229
R8184 VGND VGND.n7281 0.0148229
R8185 VGND.n7317 VGND.n7316 0.0148229
R8186 VGND.n2222 VGND.n2221 0.0148229
R8187 VGND.n2225 VGND.n2224 0.0148229
R8188 VGND.n2228 VGND.n2227 0.0148229
R8189 VGND.n6402 VGND.n6401 0.0148229
R8190 VGND.n6425 VGND.n6423 0.0148229
R8191 VGND.n6455 VGND.n1108 0.0148229
R8192 VGND.n6558 VGND.n6557 0.0148229
R8193 VGND.n6568 VGND.n6567 0.0148229
R8194 VGND.n7463 VGND.n7461 0.0148229
R8195 VGND VGND.n8021 0.0148229
R8196 VGND.n8004 VGND.n8003 0.0148229
R8197 VGND.n366 VGND.n365 0.0148229
R8198 VGND.n392 VGND.n391 0.0148229
R8199 VGND.n688 VGND.n397 0.0148229
R8200 VGND.n564 VGND.n563 0.0148229
R8201 VGND.n576 VGND.n575 0.0148229
R8202 VGND.n473 VGND 0.0148229
R8203 VGND.n2255 VGND.n2254 0.0145155
R8204 VGND.n2254 VGND.n2253 0.0145155
R8205 VGND.n1073 VGND.n1072 0.0145155
R8206 VGND.n2144 VGND.n2143 0.0145155
R8207 VGND.n1115 VGND.n1114 0.0145155
R8208 VGND.n3554 VGND.n3553 0.0145155
R8209 VGND.n3553 VGND.n3552 0.0145155
R8210 VGND.n7488 VGND.n7487 0.0145155
R8211 VGND.n7487 VGND.n7486 0.0145155
R8212 VGND.n731 VGND.n730 0.0145155
R8213 VGND.n732 VGND.n731 0.0145155
R8214 VGND.n7888 VGND.n7887 0.0145155
R8215 VGND.n3587 VGND.n3586 0.0145155
R8216 VGND.n3586 VGND.n3585 0.0145155
R8217 VGND.n7543 VGND.n7542 0.0145155
R8218 VGND.n7542 VGND.n7541 0.0145155
R8219 VGND.n7723 VGND.n7722 0.0145155
R8220 VGND.n7722 VGND.n7721 0.0145155
R8221 VGND.n7866 VGND.n7865 0.0145155
R8222 VGND.n4118 VGND.n4117 0.0145155
R8223 VGND.n4119 VGND.n4118 0.0145155
R8224 VGND.n3117 VGND.n3116 0.0145155
R8225 VGND.n3116 VGND.n3115 0.0145155
R8226 VGND.n3750 VGND.n3749 0.0145155
R8227 VGND.n3751 VGND.n3750 0.0145155
R8228 VGND.n3892 VGND.n3891 0.0145155
R8229 VGND.n4644 VGND.n4643 0.0145155
R8230 VGND.n4643 VGND.n4642 0.0145155
R8231 VGND.n4309 VGND.n4308 0.0145155
R8232 VGND.n4308 VGND.n4307 0.0145155
R8233 VGND.n4495 VGND.n4494 0.0145155
R8234 VGND.n4494 VGND.n4493 0.0145155
R8235 VGND.n4517 VGND.n4516 0.0145155
R8236 VGND.n4336 VGND.n4335 0.0145155
R8237 VGND.n4335 VGND.n4334 0.0145155
R8238 VGND.n4796 VGND.n4795 0.0145155
R8239 VGND.n4795 VGND.n4794 0.0145155
R8240 VGND.n4938 VGND.n4937 0.0145155
R8241 VGND.n4937 VGND.n4936 0.0145155
R8242 VGND.n2839 VGND.n2838 0.0145155
R8243 VGND.n5222 VGND.n5221 0.0145155
R8244 VGND.n5221 VGND.n5220 0.0145155
R8245 VGND.n5317 VGND.n5316 0.0145155
R8246 VGND.n5316 VGND.n5315 0.0145155
R8247 VGND.n2386 VGND.n2385 0.0145155
R8248 VGND.n2385 VGND.n2384 0.0145155
R8249 VGND.n2433 VGND.n2432 0.0145155
R8250 VGND.n2434 VGND.n2433 0.0145155
R8251 VGND.n5436 VGND.n5435 0.0145155
R8252 VGND.n5435 VGND.n5434 0.0145155
R8253 VGND.n1429 VGND.n1428 0.0145155
R8254 VGND.n1428 VGND.n1427 0.0145155
R8255 VGND.n2374 VGND.n2373 0.0145155
R8256 VGND.n2373 VGND.n2372 0.0145155
R8257 VGND.n2449 VGND.n2448 0.0145155
R8258 VGND.n2331 VGND.n2330 0.0145155
R8259 VGND.n2330 VGND.n2329 0.0145155
R8260 VGND.n5701 VGND.n5700 0.0145155
R8261 VGND.n5702 VGND.n5701 0.0145155
R8262 VGND.n1351 VGND.n1350 0.0145155
R8263 VGND.n1350 VGND.n1349 0.0145155
R8264 VGND.n5996 VGND.n5995 0.0145155
R8265 VGND.n1188 VGND.n1187 0.0145155
R8266 VGND.n6151 VGND.n6150 0.0145155
R8267 VGND.n6747 VGND.n6746 0.0145155
R8268 VGND.n6748 VGND.n6747 0.0145155
R8269 VGND.n7289 VGND.n7288 0.0145155
R8270 VGND.n7290 VGND.n7289 0.0145155
R8271 VGND.n468 VGND.n467 0.0145155
R8272 VGND.n467 VGND.n466 0.0145155
R8273 VGND.n958 VGND.n957 0.0145155
R8274 VGND.n959 VGND.n958 0.0145155
R8275 VGND.n592 VGND.n591 0.0145155
R8276 VGND.n591 VGND.n590 0.0145155
R8277 VGND.n7416 VGND.n7415 0.0145155
R8278 VGND.n6891 VGND.n6890 0.0145155
R8279 VGND.n6892 VGND.n6891 0.0145155
R8280 VGND.n995 VGND.n994 0.0145155
R8281 VGND.n996 VGND.n995 0.0145155
R8282 VGND.n278 VGND.n277 0.0145155
R8283 VGND.n277 VGND.n276 0.0145155
R8284 VGND.n6432 VGND.n6431 0.0145155
R8285 VGND.n6431 VGND.n6430 0.0145155
R8286 VGND.n710 VGND.n709 0.014042
R8287 VGND.n7747 VGND.n7746 0.014042
R8288 VGND.n3801 VGND.n3800 0.014042
R8289 VGND.n5633 VGND.n5632 0.014042
R8290 VGND.n1369 VGND.n1368 0.014042
R8291 VGND.n6289 VGND.n1120 0.014042
R8292 VGND.n7036 VGND.n7035 0.014042
R8293 VGND.n685 VGND.n684 0.014042
R8294 VGND.n6444 VGND.n6438 0.0140135
R8295 VGND.n6444 VGND.n6443 0.0140135
R8296 VGND.n6427 VGND.n6345 0.0140135
R8297 VGND.n6887 VGND.n6886 0.0140135
R8298 VGND.n6884 VGND.n6883 0.0140135
R8299 VGND.n6895 VGND.n1023 0.0140135
R8300 VGND.n2243 VGND.n2242 0.0140135
R8301 VGND.n2240 VGND.n2239 0.0140135
R8302 VGND.n2250 VGND.n2246 0.0140135
R8303 VGND.n1093 VGND.n1092 0.0140135
R8304 VGND.n1081 VGND.n1078 0.0140135
R8305 VGND.n2287 VGND.n2286 0.0140135
R8306 VGND.n2282 VGND.n2147 0.0140135
R8307 VGND.n2266 VGND.n2166 0.0140135
R8308 VGND.n2010 VGND.n2006 0.0140135
R8309 VGND.n2010 VGND.n2009 0.0140135
R8310 VGND.n6325 VGND.n1117 0.0140135
R8311 VGND.n3557 VGND.n3453 0.0140135
R8312 VGND.n3545 VGND.n3544 0.0140135
R8313 VGND.n3549 VGND.n3545 0.0140135
R8314 VGND.n7492 VGND.n7491 0.0140135
R8315 VGND.n7494 VGND.n7493 0.0140135
R8316 VGND.n7483 VGND.n7479 0.0140135
R8317 VGND.n271 VGND.n265 0.0140135
R8318 VGND.n271 VGND.n270 0.0140135
R8319 VGND.n735 VGND.n258 0.0140135
R8320 VGND.n7886 VGND.n7885 0.0140135
R8321 VGND.n7877 VGND.n7876 0.0140135
R8322 VGND.n3590 VGND.n3336 0.0140135
R8323 VGND.n3578 VGND.n3577 0.0140135
R8324 VGND.n3582 VGND.n3578 0.0140135
R8325 VGND.n7531 VGND.n7530 0.0140135
R8326 VGND.n7528 VGND.n7527 0.0140135
R8327 VGND.n7538 VGND.n7534 0.0140135
R8328 VGND.n102 VGND.n96 0.0140135
R8329 VGND.n102 VGND.n101 0.0140135
R8330 VGND.n7718 VGND.n104 0.0140135
R8331 VGND.n7864 VGND.n7863 0.0140135
R8332 VGND.n61 VGND.n55 0.0140135
R8333 VGND.n4114 VGND.n4113 0.0140135
R8334 VGND.n3155 VGND.n3154 0.0140135
R8335 VGND.n4122 VGND.n3155 0.0140135
R8336 VGND.n3105 VGND.n3104 0.0140135
R8337 VGND.n3102 VGND.n3101 0.0140135
R8338 VGND.n3112 VGND.n3108 0.0140135
R8339 VGND.n3746 VGND.n3740 0.0140135
R8340 VGND.n3746 VGND.n3745 0.0140135
R8341 VGND.n3754 VGND.n3733 0.0140135
R8342 VGND.n3890 VGND.n3889 0.0140135
R8343 VGND.n3908 VGND.n3907 0.0140135
R8344 VGND.n4647 VGND.n4630 0.0140135
R8345 VGND.n4635 VGND.n4634 0.0140135
R8346 VGND.n4639 VGND.n4635 0.0140135
R8347 VGND.n4297 VGND.n4296 0.0140135
R8348 VGND.n4294 VGND.n4293 0.0140135
R8349 VGND.n4304 VGND.n4300 0.0140135
R8350 VGND.n4235 VGND.n4229 0.0140135
R8351 VGND.n4235 VGND.n4234 0.0140135
R8352 VGND.n4490 VGND.n4237 0.0140135
R8353 VGND.n4515 VGND.n4514 0.0140135
R8354 VGND.n3088 VGND.n3082 0.0140135
R8355 VGND.n4324 VGND.n4323 0.0140135
R8356 VGND.n4321 VGND.n4320 0.0140135
R8357 VGND.n4331 VGND.n4327 0.0140135
R8358 VGND.n4709 VGND.n4703 0.0140135
R8359 VGND.n4709 VGND.n4708 0.0140135
R8360 VGND.n4791 VGND.n4711 0.0140135
R8361 VGND.n4942 VGND.n4941 0.0140135
R8362 VGND.n4933 VGND.n4929 0.0140135
R8363 VGND.n2842 VGND.n2835 0.0140135
R8364 VGND.n2743 VGND.n2742 0.0140135
R8365 VGND.n5052 VGND.n2743 0.0140135
R8366 VGND.n5231 VGND.n5230 0.0140135
R8367 VGND.n5249 VGND.n5243 0.0140135
R8368 VGND.n5314 VGND.n5313 0.0140135
R8369 VGND.n1563 VGND.n1562 0.0140135
R8370 VGND.n1567 VGND.n1563 0.0140135
R8371 VGND.n2716 VGND.n2715 0.0140135
R8372 VGND.n2711 VGND.n2389 0.0140135
R8373 VGND.n1690 VGND.n1684 0.0140135
R8374 VGND.n1675 VGND.n1671 0.0140135
R8375 VGND.n1675 VGND.n1674 0.0140135
R8376 VGND.n2461 VGND.n2431 0.0140135
R8377 VGND.n5439 VGND.n1464 0.0140135
R8378 VGND.n5327 VGND.n5326 0.0140135
R8379 VGND.n5431 VGND.n5327 0.0140135
R8380 VGND.n1439 VGND.n1438 0.0140135
R8381 VGND.n1424 VGND.n1420 0.0140135
R8382 VGND.n2362 VGND.n2361 0.0140135
R8383 VGND.n1698 VGND.n1697 0.0140135
R8384 VGND.n2369 VGND.n2365 0.0140135
R8385 VGND.n2447 VGND.n2442 0.0140135
R8386 VGND.n2447 VGND.n2446 0.0140135
R8387 VGND.n5655 VGND.n1393 0.0140135
R8388 VGND.n2319 VGND.n2318 0.0140135
R8389 VGND.n2314 VGND.n1910 0.0140135
R8390 VGND.n2326 VGND.n2322 0.0140135
R8391 VGND.n5724 VGND.n5665 0.0140135
R8392 VGND.n5724 VGND.n5723 0.0140135
R8393 VGND.n5705 VGND.n5699 0.0140135
R8394 VGND.n1340 VGND.n1339 0.0140135
R8395 VGND.n1346 VGND.n1342 0.0140135
R8396 VGND.n5999 VGND.n5992 0.0140135
R8397 VGND.n6026 VGND.n6025 0.0140135
R8398 VGND.n6031 VGND.n6026 0.0140135
R8399 VGND.n1197 VGND.n1196 0.0140135
R8400 VGND.n1214 VGND.n1208 0.0140135
R8401 VGND.n6103 VGND.n1239 0.0140135
R8402 VGND.n6137 VGND.n6136 0.0140135
R8403 VGND.n6143 VGND.n6137 0.0140135
R8404 VGND.n6743 VGND.n6742 0.0140135
R8405 VGND.n1047 VGND.n1046 0.0140135
R8406 VGND.n6751 VGND.n1047 0.0140135
R8407 VGND.n7285 VGND.n7284 0.0140135
R8408 VGND.n7296 VGND.n7295 0.0140135
R8409 VGND.n7301 VGND.n7296 0.0140135
R8410 VGND.n471 VGND.n460 0.0140135
R8411 VGND.n28 VGND.n27 0.0140135
R8412 VGND.n31 VGND.n28 0.0140135
R8413 VGND.n954 VGND.n953 0.0140135
R8414 VGND.n7149 VGND.n7148 0.0140135
R8415 VGND.n602 VGND.n601 0.0140135
R8416 VGND.n423 VGND.n420 0.0140135
R8417 VGND.n7468 VGND.n7467 0.0140135
R8418 VGND.n8019 VGND.n1 0.0140135
R8419 VGND.n8016 VGND.n8015 0.0140135
R8420 VGND.n991 VGND.n987 0.0140135
R8421 VGND.n991 VGND.n990 0.0140135
R8422 VGND.n7019 VGND.n1001 0.0140135
R8423 VGND.n290 VGND.n284 0.0140135
R8424 VGND.n290 VGND.n289 0.0140135
R8425 VGND.n387 VGND.n383 0.0140135
R8426 VGND.n7404 VGND.n7403 0.0135208
R8427 VGND.n239 VGND.n238 0.0135208
R8428 VGND.n246 VGND.n244 0.0135208
R8429 VGND.n708 VGND 0.0135208
R8430 VGND.n3561 VGND.n3560 0.0135208
R8431 VGND.n7599 VGND.n7598 0.0135208
R8432 VGND.n7694 VGND.n7693 0.0135208
R8433 VGND.n7701 VGND.n7699 0.0135208
R8434 VGND VGND.n7748 0.0135208
R8435 VGND.n3594 VGND.n3593 0.0135208
R8436 VGND.n4197 VGND.n4196 0.0135208
R8437 VGND.n3773 VGND.n3772 0.0135208
R8438 VGND.n3768 VGND.n3766 0.0135208
R8439 VGND VGND.n3802 0.0135208
R8440 VGND.n4109 VGND.n4108 0.0135208
R8441 VGND VGND.n4361 0.0135208
R8442 VGND.n4368 VGND.n4367 0.0135208
R8443 VGND.n4467 VGND.n4466 0.0135208
R8444 VGND.n4471 VGND.n4470 0.0135208
R8445 VGND VGND.n2979 0.0135208
R8446 VGND.n5138 VGND.n5137 0.0135208
R8447 VGND.n4765 VGND.n4764 0.0135208
R8448 VGND.n4772 VGND.n4770 0.0135208
R8449 VGND VGND.n4823 0.0135208
R8450 VGND.n2846 VGND.n2845 0.0135208
R8451 VGND.n2401 VGND.n2400 0.0135208
R8452 VGND.n2531 VGND.n2530 0.0135208
R8453 VGND VGND.n2567 0.0135208
R8454 VGND.n1584 VGND.n1583 0.0135208
R8455 VGND.n1733 VGND 0.0135208
R8456 VGND.n1748 VGND.n1747 0.0135208
R8457 VGND.n1777 VGND.n1776 0.0135208
R8458 VGND.n1773 VGND.n1772 0.0135208
R8459 VGND.n5443 VGND.n5442 0.0135208
R8460 VGND.n5669 VGND.n5668 0.0135208
R8461 VGND.n5679 VGND.n5678 0.0135208
R8462 VGND.n1367 VGND 0.0135208
R8463 VGND.n6003 VGND.n6002 0.0135208
R8464 VGND.n6310 VGND.n6309 0.0135208
R8465 VGND VGND.n1125 0.0135208
R8466 VGND.n6095 VGND.n6094 0.0135208
R8467 VGND.n6874 VGND.n6873 0.0135208
R8468 VGND.n6995 VGND.n6994 0.0135208
R8469 VGND.n7002 VGND.n7000 0.0135208
R8470 VGND.n7034 VGND 0.0135208
R8471 VGND.n7280 VGND.n7279 0.0135208
R8472 VGND VGND.n2216 0.0135208
R8473 VGND.n2223 VGND.n2222 0.0135208
R8474 VGND.n6401 VGND.n6400 0.0135208
R8475 VGND.n6408 VGND.n6406 0.0135208
R8476 VGND VGND.n6461 0.0135208
R8477 VGND.n6734 VGND.n6733 0.0135208
R8478 VGND.n7463 VGND.n7462 0.0135208
R8479 VGND.n365 VGND.n364 0.0135208
R8480 VGND.n372 VGND.n370 0.0135208
R8481 VGND.n683 VGND 0.0135208
R8482 VGND.n475 VGND.n474 0.0135208
R8483 VGND.n1029 VGND.n1028 0.0130912
R8484 VGND.n1099 VGND.n1098 0.0130912
R8485 VGND.n1085 VGND.n1084 0.0130912
R8486 VGND.n2141 VGND.n2140 0.0130912
R8487 VGND.n2014 VGND.n2013 0.0130912
R8488 VGND.n3527 VGND.n3526 0.0130912
R8489 VGND.n166 VGND.n165 0.0130912
R8490 VGND.n699 VGND.n698 0.0130912
R8491 VGND.n3314 VGND.n3313 0.0130912
R8492 VGND.n120 VGND.n119 0.0130912
R8493 VGND.n87 VGND.n86 0.0130912
R8494 VGND.n4012 VGND.n4011 0.0130912
R8495 VGND.n3133 VGND.n3132 0.0130912
R8496 VGND.n3671 VGND.n3670 0.0130912
R8497 VGND.n2953 VGND.n2952 0.0130912
R8498 VGND.n4344 VGND.n4343 0.0130912
R8499 VGND.n2890 VGND.n2889 0.0130912
R8500 VGND.n2722 VGND.n2721 0.0130912
R8501 VGND.n2877 VGND.n2876 0.0130912
R8502 VGND.n2864 VGND.n2863 0.0130912
R8503 VGND.n5218 VGND.n5217 0.0130912
R8504 VGND.n1652 VGND.n1651 0.0130912
R8505 VGND.n1475 VGND.n1474 0.0130912
R8506 VGND.n1544 VGND.n1543 0.0130912
R8507 VGND.n2382 VGND.n2381 0.0130912
R8508 VGND.n1679 VGND.n1678 0.0130912
R8509 VGND.n2522 VGND.n2521 0.0130912
R8510 VGND.n2458 VGND.n2457 0.0130912
R8511 VGND.n5348 VGND.n5347 0.0130912
R8512 VGND.n1444 VGND.n1443 0.0130912
R8513 VGND.n1865 VGND.n1864 0.0130912
R8514 VGND.n1957 VGND.n1956 0.0130912
R8515 VGND.n5689 VGND.n5688 0.0130912
R8516 VGND.n1326 VGND.n1325 0.0130912
R8517 VGND.n6156 VGND.n6155 0.0130912
R8518 VGND.n6650 VGND.n6649 0.0130912
R8519 VGND.n7265 VGND.n7264 0.0130912
R8520 VGND.n35 VGND.n34 0.0130912
R8521 VGND.n966 VGND.n965 0.0130912
R8522 VGND.n427 VGND.n426 0.0130912
R8523 VGND.n7413 VGND.n7412 0.0130912
R8524 VGND.n8012 VGND.n8011 0.0130912
R8525 VGND.n6814 VGND.n6813 0.0130912
R8526 VGND.n6819 VGND.n6818 0.0130912
R8527 VGND.n6982 VGND.n6981 0.0130912
R8528 VGND.n384 VGND.n294 0.0130912
R8529 VGND.n6340 VGND.n6339 0.0130912
R8530 VGND.n1112 VGND.n1111 0.0130912
R8531 VGND.n2139 VGND.n2138 0.0126061
R8532 VGND.n2016 VGND.n2015 0.0126061
R8533 VGND.n2639 VGND.n1653 0.0126061
R8534 VGND.n5255 VGND.n5253 0.0126061
R8535 VGND.n1598 VGND.n1597 0.0126061
R8536 VGND.n1548 VGND.n1545 0.0126061
R8537 VGND.n5207 VGND.n5206 0.0126061
R8538 VGND.n2411 VGND.n1680 0.0126061
R8539 VGND.n2524 VGND.n2523 0.0126061
R8540 VGND.n2556 VGND.n2554 0.0126061
R8541 VGND.n6158 VGND.n6157 0.0126061
R8542 VGND.n6443 VGND.n6442 0.0123243
R8543 VGND.n1077 VGND.n1076 0.0123243
R8544 VGND.n1081 VGND.n1080 0.0123243
R8545 VGND.n2155 VGND.n2154 0.0123243
R8546 VGND.n2009 VGND.n2008 0.0123243
R8547 VGND.n270 VGND.n269 0.0123243
R8548 VGND.n7878 VGND.n46 0.0123243
R8549 VGND.n7876 VGND.n47 0.0123243
R8550 VGND.n101 VGND.n100 0.0123243
R8551 VGND.n54 VGND.n53 0.0123243
R8552 VGND.n61 VGND.n60 0.0123243
R8553 VGND.n3745 VGND.n3744 0.0123243
R8554 VGND.n3909 VGND.n3636 0.0123243
R8555 VGND.n3907 VGND.n3641 0.0123243
R8556 VGND.n4234 VGND.n4233 0.0123243
R8557 VGND.n3081 VGND.n3080 0.0123243
R8558 VGND.n3088 VGND.n3087 0.0123243
R8559 VGND.n4708 VGND.n4707 0.0123243
R8560 VGND.n4933 VGND.n4932 0.0123243
R8561 VGND.n5242 VGND.n5241 0.0123243
R8562 VGND.n5249 VGND.n5248 0.0123243
R8563 VGND.n2396 VGND.n2395 0.0123243
R8564 VGND.n1674 VGND.n1673 0.0123243
R8565 VGND.n1424 VGND.n1423 0.0123243
R8566 VGND.n2446 VGND.n2445 0.0123243
R8567 VGND.n5723 VGND.n5722 0.0123243
R8568 VGND.n1346 VGND.n1345 0.0123243
R8569 VGND.n1207 VGND.n1206 0.0123243
R8570 VGND.n1214 VGND.n1213 0.0123243
R8571 VGND.n7151 VGND.n7150 0.0123243
R8572 VGND.n7148 VGND.n949 0.0123243
R8573 VGND.n423 VGND.n422 0.0123243
R8574 VGND.n7424 VGND.n7423 0.0123243
R8575 VGND.n990 VGND.n989 0.0123243
R8576 VGND.n289 VGND.n288 0.0123243
R8577 VGND.n7502 VGND.n7501 0.0122188
R8578 VGND.n3364 VGND.n3362 0.0122188
R8579 VGND.n7847 VGND.n7845 0.0122188
R8580 VGND.n4209 VGND.n4207 0.0122188
R8581 VGND VGND.n3774 0.0122188
R8582 VGND.n3918 VGND.n3913 0.0122188
R8583 VGND VGND.n4084 0.0122188
R8584 VGND.n2978 VGND.n2896 0.0122188
R8585 VGND.n4542 VGND.n4539 0.0122188
R8586 VGND.n5150 VGND.n5148 0.0122188
R8587 VGND.n4821 VGND.n4820 0.0122188
R8588 VGND.n4958 VGND.n4956 0.0122188
R8589 VGND VGND.n2820 0.0122188
R8590 VGND.n2705 VGND.n2703 0.0122188
R8591 VGND.n2529 VGND 0.0122188
R8592 VGND.n2566 VGND.n2565 0.0122188
R8593 VGND.n5275 VGND.n5269 0.0122188
R8594 VGND.n2352 VGND.n2350 0.0122188
R8595 VGND.n5544 VGND.n5542 0.0122188
R8596 VGND.n5415 VGND 0.0122188
R8597 VGND.n2308 VGND.n2306 0.0122188
R8598 VGND VGND.n2304 0.0122188
R8599 VGND.n5667 VGND 0.0122188
R8600 VGND.n5893 VGND.n5890 0.0122188
R8601 VGND.n2276 VGND.n2274 0.0122188
R8602 VGND VGND.n2272 0.0122188
R8603 VGND.n6248 VGND.n6246 0.0122188
R8604 VGND.n6900 VGND.n1018 0.0122188
R8605 VGND VGND.n6899 0.0122188
R8606 VGND.n6993 VGND 0.0122188
R8607 VGND.n7160 VGND.n7158 0.0122188
R8608 VGND.n2232 VGND.n2230 0.0122188
R8609 VGND.n6460 VGND.n6459 0.0122188
R8610 VGND.n6575 VGND.n6568 0.0122188
R8611 VGND VGND.n6710 0.0122188
R8612 VGND.n8004 VGND 0.0122188
R8613 VGND.n363 VGND 0.0122188
R8614 VGND.n579 VGND.n576 0.0122188
R8615 VGND.n2101 VGND.n2100 0.0118576
R8616 VGND.n6297 VGND.n6295 0.0118576
R8617 VGND.n6127 VGND.n6126 0.0118576
R8618 VGND.n6259 VGND.n6258 0.0118576
R8619 VGND.n6255 VGND.n6253 0.0118576
R8620 VGND.n5322 VGND.n5321 0.0117818
R8621 VGND.n5216 VGND.n5215 0.0117818
R8622 VGND.n2380 VGND.n2379 0.0117818
R8623 VGND.n2455 VGND.n2454 0.0117818
R8624 VGND.n6 VGND.n4 0.0115273
R8625 VGND.n148 VGND.n147 0.0114169
R8626 VGND.n7586 VGND.n7585 0.0114169
R8627 VGND.n5196 VGND.n5195 0.0114169
R8628 VGND.n4185 VGND.n4184 0.0114169
R8629 VGND.n4281 VGND.n4278 0.0114169
R8630 VGND.n5126 VGND.n5116 0.0114169
R8631 VGND.n1737 VGND.n1723 0.0114169
R8632 VGND.n1891 VGND.n1890 0.0114169
R8633 VGND.n2129 VGND.n2128 0.0114169
R8634 VGND.n6862 VGND.n6861 0.0114169
R8635 VGND.n2205 VGND.n2202 0.0114169
R8636 VGND.n7451 VGND.n7450 0.0114169
R8637 VGND.n7606 VGND.n7605 0.0111911
R8638 VGND.n4375 VGND.n4374 0.0111911
R8639 VGND.n7497 VGND.n7496 0.0109167
R8640 VGND.n7500 VGND.n7499 0.0109167
R8641 VGND.n7879 VGND 0.0109167
R8642 VGND.n3562 VGND 0.0109167
R8643 VGND.n7602 VGND.n7601 0.0109167
R8644 VGND.n3601 VGND.n3599 0.0109167
R8645 VGND.n3599 VGND.n3597 0.0109167
R8646 VGND.n3595 VGND 0.0109167
R8647 VGND.n4200 VGND.n4199 0.0109167
R8648 VGND.n4205 VGND.n4203 0.0109167
R8649 VGND VGND.n3910 0.0109167
R8650 VGND.n4104 VGND.n4102 0.0109167
R8651 VGND.n4106 VGND.n4104 0.0109167
R8652 VGND.n4085 VGND 0.0109167
R8653 VGND.n4371 VGND.n4370 0.0109167
R8654 VGND VGND.n4650 0.0109167
R8655 VGND.n5141 VGND.n5140 0.0109167
R8656 VGND.n5146 VGND.n5144 0.0109167
R8657 VGND.n2853 VGND.n2851 0.0109167
R8658 VGND.n2851 VGND.n2849 0.0109167
R8659 VGND.n2847 VGND 0.0109167
R8660 VGND.n2821 VGND 0.0109167
R8661 VGND.n2713 VGND.n2712 0.0109167
R8662 VGND.n2708 VGND.n2707 0.0109167
R8663 VGND.n2513 VGND 0.0109167
R8664 VGND.n2528 VGND 0.0109167
R8665 VGND.n1591 VGND.n1589 0.0109167
R8666 VGND.n1589 VGND.n1587 0.0109167
R8667 VGND.n1585 VGND 0.0109167
R8668 VGND.n2359 VGND.n2358 0.0109167
R8669 VGND.n2355 VGND.n2354 0.0109167
R8670 VGND.n5450 VGND.n5448 0.0109167
R8671 VGND.n5448 VGND.n5446 0.0109167
R8672 VGND.n5444 VGND 0.0109167
R8673 VGND VGND.n5362 0.0109167
R8674 VGND.n2316 VGND.n2315 0.0109167
R8675 VGND.n2311 VGND.n2310 0.0109167
R8676 VGND.n5735 VGND 0.0109167
R8677 VGND VGND.n5734 0.0109167
R8678 VGND.n6008 VGND.n6007 0.0109167
R8679 VGND.n6007 VGND.n6006 0.0109167
R8680 VGND.n6004 VGND 0.0109167
R8681 VGND.n2284 VGND.n2283 0.0109167
R8682 VGND.n2279 VGND.n2278 0.0109167
R8683 VGND VGND.n6243 0.0109167
R8684 VGND.n6090 VGND.n6088 0.0109167
R8685 VGND.n6092 VGND.n6090 0.0109167
R8686 VGND VGND.n6093 0.0109167
R8687 VGND.n6882 VGND.n6876 0.0109167
R8688 VGND.n6879 VGND.n6878 0.0109167
R8689 VGND VGND.n7155 0.0109167
R8690 VGND.n7275 VGND.n7273 0.0109167
R8691 VGND.n7277 VGND.n7275 0.0109167
R8692 VGND VGND.n7278 0.0109167
R8693 VGND.n2238 VGND.n2225 0.0109167
R8694 VGND.n2235 VGND.n2234 0.0109167
R8695 VGND VGND.n6797 0.0109167
R8696 VGND VGND.n6732 0.0109167
R8697 VGND.n6711 VGND 0.0109167
R8698 VGND.n8021 VGND.n8020 0.0109167
R8699 VGND.n482 VGND.n480 0.0109167
R8700 VGND.n480 VGND.n478 0.0109167
R8701 VGND.n476 VGND 0.0109167
R8702 VGND.n6442 VGND.n6441 0.0106351
R8703 VGND.n6451 VGND.n1109 0.0106351
R8704 VGND.n1080 VGND.n1079 0.0106351
R8705 VGND.n1070 VGND.n1069 0.0106351
R8706 VGND.n2008 VGND.n2007 0.0106351
R8707 VGND.n6298 VGND.n6293 0.0106351
R8708 VGND.n3569 VGND.n3568 0.0106351
R8709 VGND.n3548 VGND.n3547 0.0106351
R8710 VGND.n3522 VGND.n3521 0.0106351
R8711 VGND.n269 VGND.n268 0.0106351
R8712 VGND.n715 VGND.n703 0.0106351
R8713 VGND.n3360 VGND.n47 0.0106351
R8714 VGND.n3358 VGND.n3357 0.0106351
R8715 VGND.n3607 VGND.n3606 0.0106351
R8716 VGND.n3581 VGND.n3580 0.0106351
R8717 VGND.n3309 VGND.n3308 0.0106351
R8718 VGND.n100 VGND.n99 0.0106351
R8719 VGND.n7739 VGND.n84 0.0106351
R8720 VGND.n60 VGND.n59 0.0106351
R8721 VGND.n57 VGND.n56 0.0106351
R8722 VGND.n4005 VGND.n4004 0.0106351
R8723 VGND.n4125 VGND.n4124 0.0106351
R8724 VGND.n4014 VGND.n4013 0.0106351
R8725 VGND.n4083 VGND.n4017 0.0106351
R8726 VGND.n3744 VGND.n3743 0.0106351
R8727 VGND.n3793 VGND.n3668 0.0106351
R8728 VGND.n3641 VGND.n3640 0.0106351
R8729 VGND.n3638 VGND.n3637 0.0106351
R8730 VGND.n4660 VGND.n4659 0.0106351
R8731 VGND.n4638 VGND.n4637 0.0106351
R8732 VGND.n2948 VGND.n2947 0.0106351
R8733 VGND.n4233 VGND.n4232 0.0106351
R8734 VGND.n4692 VGND.n2892 0.0106351
R8735 VGND.n3087 VGND.n3086 0.0106351
R8736 VGND.n3084 VGND.n3083 0.0106351
R8737 VGND.n4707 VGND.n4706 0.0106351
R8738 VGND.n4812 VGND.n2874 0.0106351
R8739 VGND.n4932 VGND.n4931 0.0106351
R8740 VGND.n2867 VGND.n2866 0.0106351
R8741 VGND.n5042 VGND.n5041 0.0106351
R8742 VGND.n5056 VGND.n5055 0.0106351
R8743 VGND.n2819 VGND.n2752 0.0106351
R8744 VGND.n5248 VGND.n5247 0.0106351
R8745 VGND.n5245 VGND.n5244 0.0106351
R8746 VGND.n1595 VGND.n1594 0.0106351
R8747 VGND.n1571 VGND.n1570 0.0106351
R8748 VGND.n1673 VGND.n1672 0.0106351
R8749 VGND.n2557 VGND.n2553 0.0106351
R8750 VGND.n5354 VGND.n5353 0.0106351
R8751 VGND.n5430 VGND.n5329 0.0106351
R8752 VGND.n5343 VGND.n5342 0.0106351
R8753 VGND.n5417 VGND.n5416 0.0106351
R8754 VGND.n1423 VGND.n1422 0.0106351
R8755 VGND.n1446 VGND.n1445 0.0106351
R8756 VGND.n2445 VGND.n2444 0.0106351
R8757 VGND.n5641 VGND.n5637 0.0106351
R8758 VGND.n5722 VGND.n5666 0.0106351
R8759 VGND.n5693 VGND.n5692 0.0106351
R8760 VGND.n1345 VGND.n1344 0.0106351
R8761 VGND.n1322 VGND.n1321 0.0106351
R8762 VGND.n6013 VGND.n6012 0.0106351
R8763 VGND.n6030 VGND.n6029 0.0106351
R8764 VGND.n1213 VGND.n1212 0.0106351
R8765 VGND.n1210 VGND.n1209 0.0106351
R8766 VGND.n6142 VGND.n6141 0.0106351
R8767 VGND.n6139 VGND.n6138 0.0106351
R8768 VGND.n6645 VGND.n6644 0.0106351
R8769 VGND.n6754 VGND.n6753 0.0106351
R8770 VGND.n6652 VGND.n6651 0.0106351
R8771 VGND.n6709 VGND.n6655 0.0106351
R8772 VGND.n7261 VGND.n7260 0.0106351
R8773 VGND.n7300 VGND.n7299 0.0106351
R8774 VGND.n486 VGND.n485 0.0106351
R8775 VGND.n30 VGND.n29 0.0106351
R8776 VGND.n23 VGND.n22 0.0106351
R8777 VGND.n949 VGND.n948 0.0106351
R8778 VGND.n946 VGND.n945 0.0106351
R8779 VGND.n422 VGND.n421 0.0106351
R8780 VGND.n431 VGND.n430 0.0106351
R8781 VGND.n989 VGND.n988 0.0106351
R8782 VGND.n7027 VGND.n980 0.0106351
R8783 VGND.n288 VGND.n287 0.0106351
R8784 VGND.n690 VGND.n296 0.0106351
R8785 VGND.n819 VGND.n818 0.0103319
R8786 VGND.n6323 VGND.n6322 0.0102388
R8787 VGND.n3758 VGND.n3757 0.00990278
R8788 VGND.n2257 VGND.n2170 0.00975758
R8789 VGND.n2256 VGND.n2255 0.00975758
R8790 VGND.n2253 VGND.n2252 0.00975758
R8791 VGND.n1097 VGND.n1096 0.00975758
R8792 VGND.n1095 VGND.n1094 0.00975758
R8793 VGND.n1074 VGND.n1073 0.00975758
R8794 VGND.n1083 VGND.n1082 0.00975758
R8795 VGND.n2288 VGND.n2142 0.00975758
R8796 VGND.n2145 VGND.n2144 0.00975758
R8797 VGND.n2168 VGND.n2167 0.00975758
R8798 VGND.n2265 VGND.n2264 0.00975758
R8799 VGND.n2012 VGND.n2011 0.00975758
R8800 VGND.n2000 VGND.n1999 0.00975758
R8801 VGND.n1116 VGND.n1115 0.00975758
R8802 VGND.n6328 VGND.n6327 0.00975758
R8803 VGND.n3556 VGND.n3455 0.00975758
R8804 VGND.n3555 VGND.n3554 0.00975758
R8805 VGND.n3552 VGND.n3551 0.00975758
R8806 VGND.n7490 VGND.n7408 0.00975758
R8807 VGND.n7489 VGND.n7488 0.00975758
R8808 VGND.n7486 VGND.n7485 0.00975758
R8809 VGND.n728 VGND.n260 0.00975758
R8810 VGND.n730 VGND.n729 0.00975758
R8811 VGND.n733 VGND.n732 0.00975758
R8812 VGND.n7890 VGND.n42 0.00975758
R8813 VGND.n7889 VGND.n7888 0.00975758
R8814 VGND.n49 VGND.n48 0.00975758
R8815 VGND.n7875 VGND.n7874 0.00975758
R8816 VGND.n3589 VGND.n3338 0.00975758
R8817 VGND.n3588 VGND.n3587 0.00975758
R8818 VGND.n3585 VGND.n3584 0.00975758
R8819 VGND.n7545 VGND.n7521 0.00975758
R8820 VGND.n7544 VGND.n7543 0.00975758
R8821 VGND.n7541 VGND.n7540 0.00975758
R8822 VGND.n7725 VGND.n91 0.00975758
R8823 VGND.n7724 VGND.n7723 0.00975758
R8824 VGND.n7721 VGND.n7720 0.00975758
R8825 VGND.n7868 VGND.n7856 0.00975758
R8826 VGND.n7867 VGND.n7866 0.00975758
R8827 VGND.n52 VGND.n51 0.00975758
R8828 VGND.n64 VGND.n63 0.00975758
R8829 VGND.n4115 VGND.n3157 0.00975758
R8830 VGND.n4117 VGND.n4116 0.00975758
R8831 VGND.n4120 VGND.n4119 0.00975758
R8832 VGND.n3119 VGND.n3095 0.00975758
R8833 VGND.n3118 VGND.n3117 0.00975758
R8834 VGND.n3115 VGND.n3114 0.00975758
R8835 VGND.n3747 VGND.n3735 0.00975758
R8836 VGND.n3749 VGND.n3748 0.00975758
R8837 VGND.n3752 VGND.n3751 0.00975758
R8838 VGND.n3894 VGND.n3648 0.00975758
R8839 VGND.n3893 VGND.n3892 0.00975758
R8840 VGND.n3643 VGND.n3642 0.00975758
R8841 VGND.n3906 VGND.n3905 0.00975758
R8842 VGND.n4646 VGND.n4632 0.00975758
R8843 VGND.n4645 VGND.n4644 0.00975758
R8844 VGND.n4642 VGND.n4641 0.00975758
R8845 VGND.n4311 VGND.n4287 0.00975758
R8846 VGND.n4310 VGND.n4309 0.00975758
R8847 VGND.n4307 VGND.n4306 0.00975758
R8848 VGND.n4497 VGND.n4224 0.00975758
R8849 VGND.n4496 VGND.n4495 0.00975758
R8850 VGND.n4493 VGND.n4492 0.00975758
R8851 VGND.n4519 VGND.n4507 0.00975758
R8852 VGND.n4518 VGND.n4517 0.00975758
R8853 VGND.n3079 VGND.n3078 0.00975758
R8854 VGND.n3091 VGND.n3090 0.00975758
R8855 VGND.n4338 VGND.n4314 0.00975758
R8856 VGND.n4337 VGND.n4336 0.00975758
R8857 VGND.n4334 VGND.n4333 0.00975758
R8858 VGND.n4798 VGND.n4698 0.00975758
R8859 VGND.n4797 VGND.n4796 0.00975758
R8860 VGND.n4794 VGND.n4793 0.00975758
R8861 VGND.n4940 VGND.n2859 0.00975758
R8862 VGND.n4939 VGND.n4938 0.00975758
R8863 VGND.n4936 VGND.n4935 0.00975758
R8864 VGND.n2841 VGND.n2837 0.00975758
R8865 VGND.n2840 VGND.n2839 0.00975758
R8866 VGND.n2745 VGND.n2744 0.00975758
R8867 VGND.n5051 VGND.n5050 0.00975758
R8868 VGND.n5232 VGND.n5219 0.00975758
R8869 VGND.n5223 VGND.n5222 0.00975758
R8870 VGND.n5251 VGND.n5250 0.00975758
R8871 VGND.n5319 VGND.n1476 0.00975758
R8872 VGND.n5318 VGND.n5317 0.00975758
R8873 VGND.n1566 VGND.n1565 0.00975758
R8874 VGND.n2717 VGND.n2383 0.00975758
R8875 VGND.n2387 VGND.n2386 0.00975758
R8876 VGND.n1692 VGND.n1691 0.00975758
R8877 VGND.n1676 VGND.n1665 0.00975758
R8878 VGND.n2435 VGND.n2434 0.00975758
R8879 VGND.n2460 VGND.n2459 0.00975758
R8880 VGND.n5438 VGND.n1466 0.00975758
R8881 VGND.n5437 VGND.n5436 0.00975758
R8882 VGND.n5434 VGND.n5433 0.00975758
R8883 VGND.n1440 VGND.n1418 0.00975758
R8884 VGND.n1430 VGND.n1429 0.00975758
R8885 VGND.n1427 VGND.n1426 0.00975758
R8886 VGND.n2376 VGND.n1695 0.00975758
R8887 VGND.n2375 VGND.n2374 0.00975758
R8888 VGND.n2372 VGND.n2371 0.00975758
R8889 VGND.n2451 VGND.n2437 0.00975758
R8890 VGND.n2450 VGND.n2449 0.00975758
R8891 VGND.n1390 VGND.n1389 0.00975758
R8892 VGND.n5658 VGND.n5657 0.00975758
R8893 VGND.n2333 VGND.n1908 0.00975758
R8894 VGND.n2332 VGND.n2331 0.00975758
R8895 VGND.n2329 VGND.n2328 0.00975758
R8896 VGND.n5725 VGND.n5663 0.00975758
R8897 VGND.n5700 VGND.n5664 0.00975758
R8898 VGND.n5703 VGND.n5702 0.00975758
R8899 VGND.n1353 VGND.n1331 0.00975758
R8900 VGND.n1352 VGND.n1351 0.00975758
R8901 VGND.n1349 VGND.n1348 0.00975758
R8902 VGND.n5998 VGND.n5994 0.00975758
R8903 VGND.n5997 VGND.n5996 0.00975758
R8904 VGND.n6020 VGND.n6019 0.00975758
R8905 VGND.n6032 VGND.n6022 0.00975758
R8906 VGND.n1198 VGND.n1186 0.00975758
R8907 VGND.n1189 VGND.n1188 0.00975758
R8908 VGND.n1203 VGND.n1202 0.00975758
R8909 VGND.n1215 VGND.n1205 0.00975758
R8910 VGND.n6154 VGND.n6153 0.00975758
R8911 VGND.n6152 VGND.n6151 0.00975758
R8912 VGND.n6132 VGND.n6131 0.00975758
R8913 VGND.n6146 VGND.n6145 0.00975758
R8914 VGND.n6744 VGND.n1049 0.00975758
R8915 VGND.n6746 VGND.n6745 0.00975758
R8916 VGND.n6749 VGND.n6748 0.00975758
R8917 VGND.n7288 VGND.n7287 0.00975758
R8918 VGND.n7291 VGND.n7290 0.00975758
R8919 VGND.n7304 VGND.n7303 0.00975758
R8920 VGND.n470 VGND.n462 0.00975758
R8921 VGND.n469 VGND.n468 0.00975758
R8922 VGND.n466 VGND.n465 0.00975758
R8923 VGND.n33 VGND.n32 0.00975758
R8924 VGND.n957 VGND.n956 0.00975758
R8925 VGND.n960 VGND.n959 0.00975758
R8926 VGND.n7147 VGND.n7146 0.00975758
R8927 VGND.n603 VGND.n588 0.00975758
R8928 VGND.n593 VGND.n592 0.00975758
R8929 VGND.n590 VGND.n589 0.00975758
R8930 VGND.n425 VGND.n424 0.00975758
R8931 VGND.n7469 VGND.n7414 0.00975758
R8932 VGND.n7417 VGND.n7416 0.00975758
R8933 VGND.n8008 VGND.n8007 0.00975758
R8934 VGND.n8014 VGND.n8013 0.00975758
R8935 VGND.n6888 VGND.n1024 0.00975758
R8936 VGND.n6890 VGND.n6889 0.00975758
R8937 VGND.n6893 VGND.n6892 0.00975758
R8938 VGND.n994 VGND.n993 0.00975758
R8939 VGND.n997 VGND.n996 0.00975758
R8940 VGND.n7022 VGND.n7021 0.00975758
R8941 VGND.n291 VGND.n274 0.00975758
R8942 VGND.n279 VGND.n278 0.00975758
R8943 VGND.n276 VGND.n275 0.00975758
R8944 VGND.n386 VGND.n385 0.00975758
R8945 VGND.n6445 VGND.n6343 0.00975758
R8946 VGND.n6433 VGND.n6432 0.00975758
R8947 VGND.n6430 VGND.n6429 0.00975758
R8948 VGND.n147 VGND.n145 0.00961458
R8949 VGND.n248 VGND.n246 0.00961458
R8950 VGND VGND.n7880 0.00961458
R8951 VGND.n7880 VGND.n7879 0.00961458
R8952 VGND VGND.n3561 0.00961458
R8953 VGND.n7585 VGND.n7584 0.00961458
R8954 VGND.n7592 VGND.n7591 0.00961458
R8955 VGND.n7703 VGND.n7701 0.00961458
R8956 VGND.n7842 VGND.n7841 0.00961458
R8957 VGND.n3603 VGND.n3601 0.00961458
R8958 VGND VGND.n3594 0.00961458
R8959 VGND.n4184 VGND.n4182 0.00961458
R8960 VGND.n4192 VGND.n4191 0.00961458
R8961 VGND.n3766 VGND.n3764 0.00961458
R8962 VGND VGND.n3635 0.00961458
R8963 VGND.n3910 VGND.n3635 0.00961458
R8964 VGND.n4102 VGND.n4100 0.00961458
R8965 VGND.n4278 VGND.n4276 0.00961458
R8966 VGND.n4363 VGND.n4362 0.00961458
R8967 VGND.n4473 VGND.n4471 0.00961458
R8968 VGND.n4536 VGND.n4535 0.00961458
R8969 VGND.n5116 VGND.n5114 0.00961458
R8970 VGND VGND.n5127 0.00961458
R8971 VGND.n5132 VGND.n5131 0.00961458
R8972 VGND.n4775 VGND.n4772 0.00961458
R8973 VGND.n4953 VGND.n4952 0.00961458
R8974 VGND.n5038 VGND.n2853 0.00961458
R8975 VGND VGND.n2846 0.00961458
R8976 VGND.n5195 VGND.n5193 0.00961458
R8977 VGND.n2391 VGND.n2390 0.00961458
R8978 VGND VGND.n2406 0.00961458
R8979 VGND.n5266 VGND.n5265 0.00961458
R8980 VGND.n1593 VGND.n1591 0.00961458
R8981 VGND VGND.n1584 0.00961458
R8982 VGND.n1723 VGND.n1721 0.00961458
R8983 VGND.n1732 VGND.n1699 0.00961458
R8984 VGND.n1772 VGND.n1771 0.00961458
R8985 VGND.n5539 VGND.n5538 0.00961458
R8986 VGND.n5452 VGND.n5450 0.00961458
R8987 VGND VGND.n5443 0.00961458
R8988 VGND.n1890 VGND.n1888 0.00961458
R8989 VGND VGND.n5679 0.00961458
R8990 VGND.n5887 VGND.n5886 0.00961458
R8991 VGND.n6009 VGND.n6008 0.00961458
R8992 VGND VGND.n6003 0.00961458
R8993 VGND.n2128 VGND.n2126 0.00961458
R8994 VGND.n2149 VGND.n2148 0.00961458
R8995 VGND.n6243 VGND.n6242 0.00961458
R8996 VGND.n6088 VGND.n1236 0.00961458
R8997 VGND.n6094 VGND 0.00961458
R8998 VGND.n6861 VGND.n6859 0.00961458
R8999 VGND.n6869 VGND.n6868 0.00961458
R9000 VGND.n7004 VGND.n7002 0.00961458
R9001 VGND.n7155 VGND.n7154 0.00961458
R9002 VGND.n7273 VGND.n7271 0.00961458
R9003 VGND.n7279 VGND 0.00961458
R9004 VGND.n2202 VGND.n2200 0.00961458
R9005 VGND.n2204 VGND 0.00961458
R9006 VGND.n2218 VGND.n2217 0.00961458
R9007 VGND.n6410 VGND.n6408 0.00961458
R9008 VGND.n6565 VGND.n6564 0.00961458
R9009 VGND.n6733 VGND 0.00961458
R9010 VGND.n7450 VGND.n7448 0.00961458
R9011 VGND.n7458 VGND.n7457 0.00961458
R9012 VGND.n374 VGND.n372 0.00961458
R9013 VGND.n573 VGND.n572 0.00961458
R9014 VGND.n484 VGND.n482 0.00961458
R9015 VGND VGND.n475 0.00961458
R9016 VGND.n6338 VGND.n6335 0.00894595
R9017 VGND.n6435 VGND.n6434 0.00894595
R9018 VGND.n6438 VGND.n6437 0.00894595
R9019 VGND.n6454 VGND.n6451 0.00894595
R9020 VGND.n6824 VGND.n1015 0.00894595
R9021 VGND.n6801 VGND.n6800 0.00894595
R9022 VGND.n6548 VGND.n6543 0.00894595
R9023 VGND.n6548 VGND.n6547 0.00894595
R9024 VGND.n1091 VGND.n1090 0.00894595
R9025 VGND.n6556 VGND.n6555 0.00894595
R9026 VGND.n2099 VGND.n2098 0.00894595
R9027 VGND.n2018 VGND.n2017 0.00894595
R9028 VGND.n2003 VGND.n2002 0.00894595
R9029 VGND.n2006 VGND.n2005 0.00894595
R9030 VGND.n6301 VGND.n6298 0.00894595
R9031 VGND.n3570 VGND.n3567 0.00894595
R9032 VGND.n3544 VGND.n3457 0.00894595
R9033 VGND.n3547 VGND.n3546 0.00894595
R9034 VGND.n3531 VGND.n3530 0.00894595
R9035 VGND.n7515 VGND.n7514 0.00894595
R9036 VGND.n722 VGND.n719 0.00894595
R9037 VGND.n262 VGND.n261 0.00894595
R9038 VGND.n265 VGND.n264 0.00894595
R9039 VGND.n715 VGND.n714 0.00894595
R9040 VGND.n826 VGND.n825 0.00894595
R9041 VGND.n825 VGND.n821 0.00894595
R9042 VGND.n7884 VGND.n7883 0.00894595
R9043 VGND.n3355 VGND.n3354 0.00894595
R9044 VGND.n3608 VGND.n3605 0.00894595
R9045 VGND.n3577 VGND.n3576 0.00894595
R9046 VGND.n3580 VGND.n3579 0.00894595
R9047 VGND.n3318 VGND.n3317 0.00894595
R9048 VGND.n7561 VGND.n7560 0.00894595
R9049 VGND.n7731 VGND.n7728 0.00894595
R9050 VGND.n93 VGND.n92 0.00894595
R9051 VGND.n96 VGND.n95 0.00894595
R9052 VGND.n7742 VGND.n7739 0.00894595
R9053 VGND.n7823 VGND.n7822 0.00894595
R9054 VGND.n7822 VGND.n7819 0.00894595
R9055 VGND.n7862 VGND.n7861 0.00894595
R9056 VGND.n7851 VGND.n7850 0.00894595
R9057 VGND.n4097 VGND.n4096 0.00894595
R9058 VGND.n3154 VGND.n3153 0.00894595
R9059 VGND.n4124 VGND.n4123 0.00894595
R9060 VGND.n4089 VGND.n4088 0.00894595
R9061 VGND.n4218 VGND.n4217 0.00894595
R9062 VGND.n3785 VGND.n3782 0.00894595
R9063 VGND.n3737 VGND.n3736 0.00894595
R9064 VGND.n3740 VGND.n3739 0.00894595
R9065 VGND.n3796 VGND.n3793 0.00894595
R9066 VGND.n3868 VGND.n3867 0.00894595
R9067 VGND.n3867 VGND.n3864 0.00894595
R9068 VGND.n3888 VGND.n3887 0.00894595
R9069 VGND.n3898 VGND.n3634 0.00894595
R9070 VGND.n4661 VGND.n4658 0.00894595
R9071 VGND.n4634 VGND.n4633 0.00894595
R9072 VGND.n4637 VGND.n4636 0.00894595
R9073 VGND.n4668 VGND.n4667 0.00894595
R9074 VGND.n4350 VGND.n4251 0.00894595
R9075 VGND.n2883 VGND.n2880 0.00894595
R9076 VGND.n4226 VGND.n4225 0.00894595
R9077 VGND.n4229 VGND.n4228 0.00894595
R9078 VGND.n4692 VGND.n4691 0.00894595
R9079 VGND.n3073 VGND.n3070 0.00894595
R9080 VGND.n3073 VGND.n3072 0.00894595
R9081 VGND.n4513 VGND.n4512 0.00894595
R9082 VGND.n4525 VGND.n4524 0.00894595
R9083 VGND.n5159 VGND.n5158 0.00894595
R9084 VGND.n4804 VGND.n4801 0.00894595
R9085 VGND.n4700 VGND.n4699 0.00894595
R9086 VGND.n4703 VGND.n4702 0.00894595
R9087 VGND.n4815 VGND.n4812 0.00894595
R9088 VGND.n4922 VGND.n4919 0.00894595
R9089 VGND.n4922 VGND.n4921 0.00894595
R9090 VGND.n4946 VGND.n4945 0.00894595
R9091 VGND.n2869 VGND.n2856 0.00894595
R9092 VGND.n5043 VGND.n5040 0.00894595
R9093 VGND.n2742 VGND.n2741 0.00894595
R9094 VGND.n5055 VGND.n5054 0.00894595
R9095 VGND.n2825 VGND.n2824 0.00894595
R9096 VGND.n2641 VGND.n2640 0.00894595
R9097 VGND.n2640 VGND.n2636 0.00894595
R9098 VGND.n5229 VGND.n5228 0.00894595
R9099 VGND.n5257 VGND.n5256 0.00894595
R9100 VGND.n1600 VGND.n1599 0.00894595
R9101 VGND.n1562 VGND.n1561 0.00894595
R9102 VGND.n1570 VGND.n1569 0.00894595
R9103 VGND.n1550 VGND.n1549 0.00894595
R9104 VGND.n2413 VGND.n2412 0.00894595
R9105 VGND.n2525 VGND.n2518 0.00894595
R9106 VGND.n1668 VGND.n1667 0.00894595
R9107 VGND.n1671 VGND.n1670 0.00894595
R9108 VGND.n2560 VGND.n2557 0.00894595
R9109 VGND.n5355 VGND.n1459 0.00894595
R9110 VGND.n5326 VGND.n5325 0.00894595
R9111 VGND.n5329 VGND.n5328 0.00894595
R9112 VGND.n5418 VGND.n5361 0.00894595
R9113 VGND.n5556 VGND.n5555 0.00894595
R9114 VGND.n5555 VGND.n1413 0.00894595
R9115 VGND.n1437 VGND.n1436 0.00894595
R9116 VGND.n5548 VGND.n5547 0.00894595
R9117 VGND.n2341 VGND.n2340 0.00894595
R9118 VGND.n1384 VGND.n1381 0.00894595
R9119 VGND.n2439 VGND.n2438 0.00894595
R9120 VGND.n2442 VGND.n2441 0.00894595
R9121 VGND.n5644 VGND.n5641 0.00894595
R9122 VGND.n2297 VGND.n2296 0.00894595
R9123 VGND.n5731 VGND.n1378 0.00894595
R9124 VGND.n5671 VGND.n5670 0.00894595
R9125 VGND.n5673 VGND.n5665 0.00894595
R9126 VGND.n5692 VGND.n5686 0.00894595
R9127 VGND.n5867 VGND.n5864 0.00894595
R9128 VGND.n5867 VGND.n5866 0.00894595
R9129 VGND.n1338 VGND.n1337 0.00894595
R9130 VGND.n5876 VGND.n5875 0.00894595
R9131 VGND.n6014 VGND.n6011 0.00894595
R9132 VGND.n6025 VGND.n6024 0.00894595
R9133 VGND.n6029 VGND.n6028 0.00894595
R9134 VGND.n1304 VGND.n1303 0.00894595
R9135 VGND.n6261 VGND.n6260 0.00894595
R9136 VGND.n6260 VGND.n1183 0.00894595
R9137 VGND.n1195 VGND.n1194 0.00894595
R9138 VGND.n6252 VGND.n6251 0.00894595
R9139 VGND.n6160 VGND.n6159 0.00894595
R9140 VGND.n6136 VGND.n6135 0.00894595
R9141 VGND.n6141 VGND.n6140 0.00894595
R9142 VGND.n6125 VGND.n6124 0.00894595
R9143 VGND.n6723 VGND.n6722 0.00894595
R9144 VGND.n1046 VGND.n1045 0.00894595
R9145 VGND.n6753 VGND.n6752 0.00894595
R9146 VGND.n6715 VGND.n6714 0.00894595
R9147 VGND.n7268 VGND.n7267 0.00894595
R9148 VGND.n7295 VGND.n7294 0.00894595
R9149 VGND.n7299 VGND.n7298 0.00894595
R9150 VGND.n7310 VGND.n7309 0.00894595
R9151 VGND.n491 VGND.n490 0.00894595
R9152 VGND.n27 VGND.n26 0.00894595
R9153 VGND.n7902 VGND.n7901 0.00894595
R9154 VGND.n7135 VGND.n7131 0.00894595
R9155 VGND.n7135 VGND.n7134 0.00894595
R9156 VGND.n7140 VGND.n943 0.00894595
R9157 VGND.n610 VGND.n609 0.00894595
R9158 VGND.n609 VGND.n418 0.00894595
R9159 VGND.n600 VGND.n599 0.00894595
R9160 VGND.n583 VGND.n582 0.00894595
R9161 VGND.n7998 VGND.n7997 0.00894595
R9162 VGND.n6985 VGND.n6984 0.00894595
R9163 VGND.n6976 VGND.n6975 0.00894595
R9164 VGND.n987 VGND.n986 0.00894595
R9165 VGND.n7030 VGND.n7027 0.00894595
R9166 VGND.n355 VGND.n354 0.00894595
R9167 VGND.n281 VGND.n280 0.00894595
R9168 VGND.n284 VGND.n283 0.00894595
R9169 VGND.n690 VGND.n689 0.00894595
R9170 VGND.n1960 VGND.n1959 0.00837842
R9171 VGND.n1962 VGND.n1961 0.00837842
R9172 VGND.n5212 VGND.n5211 0.00837842
R9173 VGND.n1965 VGND.n1964 0.00837842
R9174 VGND.n234 VGND.n233 0.0083125
R9175 VGND.n244 VGND.n242 0.0083125
R9176 VGND.n249 VGND.n248 0.0083125
R9177 VGND.n709 VGND.n708 0.0083125
R9178 VGND.n3361 VGND.n3356 0.0083125
R9179 VGND.n3365 VGND.n3364 0.0083125
R9180 VGND.n3542 VGND.n3541 0.0083125
R9181 VGND.n3539 VGND.n3538 0.0083125
R9182 VGND.n7689 VGND.n7688 0.0083125
R9183 VGND.n7699 VGND.n7697 0.0083125
R9184 VGND.n7704 VGND.n7703 0.0083125
R9185 VGND.n7748 VGND.n7747 0.0083125
R9186 VGND.n7844 VGND.n7843 0.0083125
R9187 VGND.n7848 VGND.n7847 0.0083125
R9188 VGND.n3329 VGND.n3328 0.0083125
R9189 VGND.n3326 VGND.n3325 0.0083125
R9190 VGND.n3779 VGND.n3777 0.0083125
R9191 VGND.n3770 VGND.n3768 0.0083125
R9192 VGND.n3764 VGND.n3762 0.0083125
R9193 VGND.n3802 VGND.n3801 0.0083125
R9194 VGND.n3912 VGND.n3911 0.0083125
R9195 VGND.n3919 VGND.n3918 0.0083125
R9196 VGND.n4126 VGND.n3152 0.0083125
R9197 VGND.n4020 VGND.n4019 0.0083125
R9198 VGND.n4086 VGND.n4085 0.0083125
R9199 VGND.n4462 VGND.n4461 0.0083125
R9200 VGND.n4470 VGND.n4469 0.0083125
R9201 VGND.n4474 VGND.n4473 0.0083125
R9202 VGND.n2979 VGND.n2978 0.0083125
R9203 VGND.n4538 VGND.n4537 0.0083125
R9204 VGND.n4543 VGND.n4542 0.0083125
R9205 VGND.n4677 VGND.n4676 0.0083125
R9206 VGND.n4674 VGND.n4673 0.0083125
R9207 VGND.n4760 VGND.n4759 0.0083125
R9208 VGND.n4770 VGND.n4768 0.0083125
R9209 VGND.n4776 VGND.n4775 0.0083125
R9210 VGND.n4823 VGND.n4821 0.0083125
R9211 VGND.n4955 VGND.n4954 0.0083125
R9212 VGND.n4959 VGND.n4958 0.0083125
R9213 VGND.n5057 VGND.n2739 0.0083125
R9214 VGND.n2755 VGND.n2754 0.0083125
R9215 VGND.n2822 VGND.n2821 0.0083125
R9216 VGND.n2697 VGND.n2402 0.0083125
R9217 VGND.n2515 VGND.n2514 0.0083125
R9218 VGND.n2536 VGND.n2535 0.0083125
R9219 VGND.n2567 VGND.n2566 0.0083125
R9220 VGND.n5268 VGND.n5267 0.0083125
R9221 VGND.n5276 VGND.n5275 0.0083125
R9222 VGND.n1572 VGND.n1560 0.0083125
R9223 VGND.n1558 VGND.n1557 0.0083125
R9224 VGND.n1782 VGND.n1781 0.0083125
R9225 VGND.n1774 VGND.n1773 0.0083125
R9226 VGND.n1771 VGND.n1770 0.0083125
R9227 VGND.n5632 VGND.n5631 0.0083125
R9228 VGND.n5541 VGND.n5540 0.0083125
R9229 VGND.n5545 VGND.n5544 0.0083125
R9230 VGND.n5429 VGND.n5428 0.0083125
R9231 VGND.n5426 VGND.n5425 0.0083125
R9232 VGND.n5362 VGND.n5341 0.0083125
R9233 VGND.n5739 VGND.n5736 0.0083125
R9234 VGND.n5678 VGND.n5676 0.0083125
R9235 VGND VGND.n5719 0.0083125
R9236 VGND.n1368 VGND.n1367 0.0083125
R9237 VGND.n5889 VGND.n5888 0.0083125
R9238 VGND.n5894 VGND.n5893 0.0083125
R9239 VGND.n1315 VGND.n1314 0.0083125
R9240 VGND.n1312 VGND.n1311 0.0083125
R9241 VGND.n2097 VGND.n1974 0.0083125
R9242 VGND.n2023 VGND.n2022 0.0083125
R9243 VGND.n6315 VGND.n6314 0.0083125
R9244 VGND.n1125 VGND.n1120 0.0083125
R9245 VGND.n6245 VGND.n6244 0.0083125
R9246 VGND.n6249 VGND.n6248 0.0083125
R9247 VGND.n6114 VGND.n6113 0.0083125
R9248 VGND.n6117 VGND.n6116 0.0083125
R9249 VGND.n1019 VGND 0.0083125
R9250 VGND VGND.n1016 0.0083125
R9251 VGND.n6990 VGND.n6989 0.0083125
R9252 VGND.n7000 VGND.n6998 0.0083125
R9253 VGND.n7005 VGND.n7004 0.0083125
R9254 VGND.n7035 VGND.n7034 0.0083125
R9255 VGND.n7157 VGND.n7156 0.0083125
R9256 VGND.n7161 VGND.n7160 0.0083125
R9257 VGND.n7321 VGND.n7320 0.0083125
R9258 VGND.n7318 VGND.n7317 0.0083125
R9259 VGND.n6796 VGND.n6795 0.0083125
R9260 VGND.n6396 VGND.n6395 0.0083125
R9261 VGND.n6406 VGND.n6404 0.0083125
R9262 VGND.n6411 VGND.n6410 0.0083125
R9263 VGND.n6461 VGND.n6460 0.0083125
R9264 VGND.n6567 VGND.n6566 0.0083125
R9265 VGND.n6576 VGND.n6575 0.0083125
R9266 VGND.n6756 VGND.n6755 0.0083125
R9267 VGND.n6759 VGND.n6758 0.0083125
R9268 VGND.n6712 VGND.n6711 0.0083125
R9269 VGND.n8002 VGND 0.0083125
R9270 VGND VGND.n8001 0.0083125
R9271 VGND.n360 VGND.n359 0.0083125
R9272 VGND.n370 VGND.n368 0.0083125
R9273 VGND.n375 VGND.n374 0.0083125
R9274 VGND.n684 VGND.n683 0.0083125
R9275 VGND.n575 VGND.n574 0.0083125
R9276 VGND.n580 VGND.n579 0.0083125
R9277 VGND.n7962 VGND.n7961 0.0083125
R9278 VGND.n7959 VGND.n7958 0.0083125
R9279 VGND.n1658 VGND.n1657 0.00803709
R9280 VGND.n1655 VGND.n1654 0.00803709
R9281 VGND.n2638 VGND.n2637 0.00762121
R9282 VGND.n1547 VGND.n1546 0.00762121
R9283 VGND.n2410 VGND.n2409 0.00762121
R9284 VGND.n2520 VGND.n2519 0.00762121
R9285 VGND.n6036 VGND.n6035 0.00735251
R9286 VGND.n1328 VGND.n1327 0.00735251
R9287 VGND.n2291 VGND.n2290 0.00735251
R9288 VGND.n1997 VGND.n1996 0.00735251
R9289 VGND.n6809 VGND.n6808 0.00725676
R9290 VGND.n2214 VGND.n2213 0.00725676
R9291 VGND.n2136 VGND.n2135 0.00725676
R9292 VGND.n3459 VGND.n3458 0.00725676
R9293 VGND.n156 VGND.n155 0.00725676
R9294 VGND.n3168 VGND.n3167 0.00725676
R9295 VGND.n7549 VGND.n7548 0.00725676
R9296 VGND.n3620 VGND.n3619 0.00725676
R9297 VGND.n3123 VGND.n3122 0.00725676
R9298 VGND.n4627 VGND.n4626 0.00725676
R9299 VGND.n4359 VGND.n4358 0.00725676
R9300 VGND.n5124 VGND.n5123 0.00725676
R9301 VGND.n1483 VGND.n1482 0.00725676
R9302 VGND.n5203 VGND.n5202 0.00725676
R9303 VGND.n5331 VGND.n5330 0.00725676
R9304 VGND.n1735 VGND.n1730 0.00725676
R9305 VGND.n1899 VGND.n1898 0.00725676
R9306 VGND.n6134 VGND.n6133 0.00725676
R9307 VGND.n1057 VGND.n1056 0.00725676
R9308 VGND.n7293 VGND.n7292 0.00725676
R9309 VGND.n457 VGND.n456 0.00725676
R9310 VGND.n7420 VGND.n7419 0.00725676
R9311 VGND.n7501 VGND.n7500 0.00701042
R9312 VGND.n238 VGND.n237 0.00701042
R9313 VGND.n242 VGND.n240 0.00701042
R9314 VGND.n809 VGND.n45 0.00701042
R9315 VGND.n7881 VGND 0.00701042
R9316 VGND.n3543 VGND 0.00701042
R9317 VGND.n3541 VGND.n3540 0.00701042
R9318 VGND.n7693 VGND.n7692 0.00701042
R9319 VGND.n7697 VGND.n7695 0.00701042
R9320 VGND.n7839 VGND.n7837 0.00701042
R9321 VGND.n3331 VGND.n3330 0.00701042
R9322 VGND.n3330 VGND 0.00701042
R9323 VGND.n3328 VGND.n3327 0.00701042
R9324 VGND.n4207 VGND.n4205 0.00701042
R9325 VGND.n3774 VGND.n3773 0.00701042
R9326 VGND.n3771 VGND.n3770 0.00701042
R9327 VGND.n3884 VGND.n3882 0.00701042
R9328 VGND.n3885 VGND 0.00701042
R9329 VGND.n4128 VGND.n4127 0.00701042
R9330 VGND.n4127 VGND 0.00701042
R9331 VGND.n4018 VGND.n3152 0.00701042
R9332 VGND VGND.n4025 0.00701042
R9333 VGND VGND.n4253 0.00701042
R9334 VGND.n4466 VGND.n4465 0.00701042
R9335 VGND.n4469 VGND.n4468 0.00701042
R9336 VGND.n4533 VGND.n4531 0.00701042
R9337 VGND.n4679 VGND.n4678 0.00701042
R9338 VGND.n4678 VGND 0.00701042
R9339 VGND.n4676 VGND.n4675 0.00701042
R9340 VGND.n5148 VGND.n5146 0.00701042
R9341 VGND.n4764 VGND.n4763 0.00701042
R9342 VGND.n4768 VGND.n4766 0.00701042
R9343 VGND.n4950 VGND.n4948 0.00701042
R9344 VGND.n5059 VGND.n5058 0.00701042
R9345 VGND.n5058 VGND 0.00701042
R9346 VGND.n2753 VGND.n2739 0.00701042
R9347 VGND.n2823 VGND 0.00701042
R9348 VGND.n2707 VGND.n2705 0.00701042
R9349 VGND.n2530 VGND.n2529 0.00701042
R9350 VGND.n2533 VGND.n2532 0.00701042
R9351 VGND.n5263 VGND.n5262 0.00701042
R9352 VGND.n1574 VGND.n1573 0.00701042
R9353 VGND.n1573 VGND 0.00701042
R9354 VGND.n1560 VGND.n1559 0.00701042
R9355 VGND.n1552 VGND 0.00701042
R9356 VGND.n1738 VGND 0.00701042
R9357 VGND.n2354 VGND.n2352 0.00701042
R9358 VGND.n1778 VGND.n1777 0.00701042
R9359 VGND.n1775 VGND.n1774 0.00701042
R9360 VGND.n5536 VGND.n5534 0.00701042
R9361 VGND.n5340 VGND.n5339 0.00701042
R9362 VGND VGND.n5340 0.00701042
R9363 VGND.n5428 VGND.n5427 0.00701042
R9364 VGND VGND.n5419 0.00701042
R9365 VGND VGND.n1920 0.00701042
R9366 VGND.n1921 VGND 0.00701042
R9367 VGND.n2310 VGND.n2308 0.00701042
R9368 VGND.n5668 VGND.n5667 0.00701042
R9369 VGND.n5676 VGND.n5674 0.00701042
R9370 VGND.n5884 VGND.n5882 0.00701042
R9371 VGND.n1317 VGND.n1316 0.00701042
R9372 VGND.n1316 VGND 0.00701042
R9373 VGND.n1314 VGND.n1313 0.00701042
R9374 VGND VGND.n2159 0.00701042
R9375 VGND.n2160 VGND 0.00701042
R9376 VGND.n2278 VGND.n2276 0.00701042
R9377 VGND.n6309 VGND.n6308 0.00701042
R9378 VGND.n6312 VGND.n6311 0.00701042
R9379 VGND.n6240 VGND.n6238 0.00701042
R9380 VGND.n6112 VGND.n6111 0.00701042
R9381 VGND VGND.n6112 0.00701042
R9382 VGND.n6115 VGND.n6114 0.00701042
R9383 VGND.n6878 VGND.n1018 0.00701042
R9384 VGND.n6994 VGND.n6993 0.00701042
R9385 VGND.n6998 VGND.n6996 0.00701042
R9386 VGND.n7117 VGND.n7115 0.00701042
R9387 VGND.n7323 VGND.n7322 0.00701042
R9388 VGND.n7322 VGND 0.00701042
R9389 VGND.n7320 VGND.n7319 0.00701042
R9390 VGND.n2234 VGND.n2232 0.00701042
R9391 VGND.n6400 VGND.n6399 0.00701042
R9392 VGND.n6404 VGND.n6402 0.00701042
R9393 VGND.n6562 VGND.n6561 0.00701042
R9394 VGND.n6737 VGND.n6736 0.00701042
R9395 VGND.n6736 VGND 0.00701042
R9396 VGND.n6757 VGND.n6756 0.00701042
R9397 VGND VGND.n1044 0.00701042
R9398 VGND.n6713 VGND 0.00701042
R9399 VGND.n364 VGND.n363 0.00701042
R9400 VGND.n368 VGND.n366 0.00701042
R9401 VGND.n570 VGND.n568 0.00701042
R9402 VGND.n7964 VGND.n7963 0.00701042
R9403 VGND.n7963 VGND 0.00701042
R9404 VGND.n7961 VGND.n7960 0.00701042
R9405 VGND.n1656 VGND.n1655 0.00696227
R9406 VGND.n1959 VGND.n1958 0.00696227
R9407 VGND.n5211 VGND.n5210 0.00657697
R9408 VGND.n5213 VGND.n1658 0.00657697
R9409 VGND.n1966 VGND.n1965 0.00657697
R9410 VGND.n1963 VGND.n1962 0.00657697
R9411 VGND.n2101 VGND.n1969 0.00648266
R9412 VGND.n6295 VGND.n6294 0.00648266
R9413 VGND.n6258 VGND.n6257 0.00648266
R9414 VGND.n6255 VGND.n6254 0.00648266
R9415 VGND.n6127 VGND.n6037 0.00648266
R9416 VGND.n2257 VGND.n2256 0.00619697
R9417 VGND.n2252 VGND.n2251 0.00619697
R9418 VGND.n1096 VGND.n1095 0.00619697
R9419 VGND.n1082 VGND.n1074 0.00619697
R9420 VGND.n2288 VGND.n2145 0.00619697
R9421 VGND.n2265 VGND.n2168 0.00619697
R9422 VGND.n2011 VGND.n2000 0.00619697
R9423 VGND.n6328 VGND.n1116 0.00619697
R9424 VGND.n3556 VGND.n3555 0.00619697
R9425 VGND.n3551 VGND.n3550 0.00619697
R9426 VGND.n7490 VGND.n7489 0.00619697
R9427 VGND.n7485 VGND.n7484 0.00619697
R9428 VGND.n729 VGND.n728 0.00619697
R9429 VGND.n734 VGND.n733 0.00619697
R9430 VGND.n7890 VGND.n7889 0.00619697
R9431 VGND.n7875 VGND.n49 0.00619697
R9432 VGND.n3589 VGND.n3588 0.00619697
R9433 VGND.n3584 VGND.n3583 0.00619697
R9434 VGND.n7545 VGND.n7544 0.00619697
R9435 VGND.n7540 VGND.n7539 0.00619697
R9436 VGND.n7725 VGND.n7724 0.00619697
R9437 VGND.n7720 VGND.n7719 0.00619697
R9438 VGND.n7868 VGND.n7867 0.00619697
R9439 VGND.n64 VGND.n52 0.00619697
R9440 VGND.n4116 VGND.n4115 0.00619697
R9441 VGND.n4121 VGND.n4120 0.00619697
R9442 VGND.n3119 VGND.n3118 0.00619697
R9443 VGND.n3114 VGND.n3113 0.00619697
R9444 VGND.n3748 VGND.n3747 0.00619697
R9445 VGND.n3753 VGND.n3752 0.00619697
R9446 VGND.n3894 VGND.n3893 0.00619697
R9447 VGND.n3906 VGND.n3643 0.00619697
R9448 VGND.n4646 VGND.n4645 0.00619697
R9449 VGND.n4641 VGND.n4640 0.00619697
R9450 VGND.n4311 VGND.n4310 0.00619697
R9451 VGND.n4306 VGND.n4305 0.00619697
R9452 VGND.n4497 VGND.n4496 0.00619697
R9453 VGND.n4492 VGND.n4491 0.00619697
R9454 VGND.n4519 VGND.n4518 0.00619697
R9455 VGND.n3091 VGND.n3079 0.00619697
R9456 VGND.n4338 VGND.n4337 0.00619697
R9457 VGND.n4333 VGND.n4332 0.00619697
R9458 VGND.n4798 VGND.n4797 0.00619697
R9459 VGND.n4793 VGND.n4792 0.00619697
R9460 VGND.n4940 VGND.n4939 0.00619697
R9461 VGND.n4935 VGND.n4934 0.00619697
R9462 VGND.n2841 VGND.n2840 0.00619697
R9463 VGND.n5051 VGND.n2745 0.00619697
R9464 VGND.n5232 VGND.n5223 0.00619697
R9465 VGND.n5251 VGND.n5240 0.00619697
R9466 VGND.n5319 VGND.n5318 0.00619697
R9467 VGND.n1566 VGND.n1564 0.00619697
R9468 VGND.n2717 VGND.n2387 0.00619697
R9469 VGND.n1692 VGND.n1681 0.00619697
R9470 VGND.n1676 VGND.n1666 0.00619697
R9471 VGND.n2460 VGND.n2435 0.00619697
R9472 VGND.n5438 VGND.n5437 0.00619697
R9473 VGND.n5433 VGND.n5432 0.00619697
R9474 VGND.n1440 VGND.n1430 0.00619697
R9475 VGND.n1426 VGND.n1425 0.00619697
R9476 VGND.n2376 VGND.n2375 0.00619697
R9477 VGND.n2371 VGND.n2370 0.00619697
R9478 VGND.n2451 VGND.n2450 0.00619697
R9479 VGND.n5658 VGND.n1390 0.00619697
R9480 VGND.n2333 VGND.n2332 0.00619697
R9481 VGND.n2328 VGND.n2327 0.00619697
R9482 VGND.n5725 VGND.n5664 0.00619697
R9483 VGND.n5704 VGND.n5703 0.00619697
R9484 VGND.n1353 VGND.n1352 0.00619697
R9485 VGND.n1348 VGND.n1347 0.00619697
R9486 VGND.n5998 VGND.n5997 0.00619697
R9487 VGND.n6032 VGND.n6020 0.00619697
R9488 VGND.n1198 VGND.n1189 0.00619697
R9489 VGND.n1215 VGND.n1203 0.00619697
R9490 VGND.n6153 VGND.n6152 0.00619697
R9491 VGND.n6146 VGND.n6132 0.00619697
R9492 VGND.n6745 VGND.n6744 0.00619697
R9493 VGND.n6750 VGND.n6749 0.00619697
R9494 VGND.n7287 VGND.n7286 0.00619697
R9495 VGND.n7304 VGND.n7291 0.00619697
R9496 VGND.n470 VGND.n469 0.00619697
R9497 VGND.n956 VGND.n955 0.00619697
R9498 VGND.n7147 VGND.n960 0.00619697
R9499 VGND.n603 VGND.n593 0.00619697
R9500 VGND.n7469 VGND.n7417 0.00619697
R9501 VGND.n8014 VGND.n8008 0.00619697
R9502 VGND.n6889 VGND.n6888 0.00619697
R9503 VGND.n6894 VGND.n6893 0.00619697
R9504 VGND.n993 VGND.n992 0.00619697
R9505 VGND.n7022 VGND.n997 0.00619697
R9506 VGND.n291 VGND.n279 0.00619697
R9507 VGND.n6445 VGND.n6433 0.00619697
R9508 VGND.n6429 VGND.n6428 0.00619697
R9509 VGND.n6149 VGND.n6036 0.00590801
R9510 VGND.n6147 VGND.n6130 0.00590801
R9511 VGND.n2262 VGND.n2261 0.00590801
R9512 VGND.n6330 VGND.n6329 0.00590801
R9513 VGND.n154 VGND.n153 0.00570833
R9514 VGND.n7403 VGND 0.00570833
R9515 VGND.n3463 VGND.n3462 0.00570833
R9516 VGND.n7590 VGND.n7589 0.00570833
R9517 VGND.n7828 VGND.n7826 0.00570833
R9518 VGND VGND.n7830 0.00570833
R9519 VGND.n3333 VGND.n3332 0.00570833
R9520 VGND.n4190 VGND.n4189 0.00570833
R9521 VGND.n3873 VGND.n3871 0.00570833
R9522 VGND.n4129 VGND.n3151 0.00570833
R9523 VGND.n4361 VGND.n4360 0.00570833
R9524 VGND.n3068 VGND.n2972 0.00570833
R9525 VGND.n4680 VGND.n2899 0.00570833
R9526 VGND.n5130 VGND.n5129 0.00570833
R9527 VGND.n4917 VGND.n4916 0.00570833
R9528 VGND.n4915 VGND 0.00570833
R9529 VGND.n5060 VGND.n2738 0.00570833
R9530 VGND.n5201 VGND.n5200 0.00570833
R9531 VGND VGND.n2401 0.00570833
R9532 VGND.n2634 VGND.n2631 0.00570833
R9533 VGND.n5310 VGND.n5309 0.00570833
R9534 VGND.n1734 VGND.n1733 0.00570833
R9535 VGND.n5563 VGND.n5561 0.00570833
R9536 VGND.n5338 VGND.n5334 0.00570833
R9537 VGND.n1897 VGND.n1896 0.00570833
R9538 VGND.n5862 VGND.n1358 0.00570833
R9539 VGND.n5989 VGND.n5988 0.00570833
R9540 VGND.n2134 VGND.n2133 0.00570833
R9541 VGND.n6229 VGND.n1181 0.00570833
R9542 VGND.n6110 VGND.n6106 0.00570833
R9543 VGND.n6867 VGND.n6866 0.00570833
R9544 VGND.n7129 VGND.n7126 0.00570833
R9545 VGND.n7324 VGND.n878 0.00570833
R9546 VGND.n2216 VGND.n2215 0.00570833
R9547 VGND.n6541 VGND.n6538 0.00570833
R9548 VGND.n6739 VGND.n6738 0.00570833
R9549 VGND.n7456 VGND.n7455 0.00570833
R9550 VGND.n7462 VGND 0.00570833
R9551 VGND.n416 VGND.n415 0.00570833
R9552 VGND.n7965 VGND.n17 0.00570833
R9553 VGND.n1968 VGND.n1967 0.005649
R9554 VGND.n6335 VGND.n6334 0.00556757
R9555 VGND.n6454 VGND.n6453 0.00556757
R9556 VGND.n6808 VGND.n6807 0.00556757
R9557 VGND.n6887 VGND.n6833 0.00556757
R9558 VGND.n2214 VGND.n2206 0.00556757
R9559 VGND.n2243 VGND.n2175 0.00556757
R9560 VGND.n6800 VGND.n6799 0.00556757
R9561 VGND.n2135 VGND.n2104 0.00556757
R9562 VGND.n2287 VGND.n2146 0.00556757
R9563 VGND.n2270 VGND.n2269 0.00556757
R9564 VGND.n2098 VGND.n1973 0.00556757
R9565 VGND.n2019 VGND.n2018 0.00556757
R9566 VGND.n6301 VGND.n6300 0.00556757
R9567 VGND.n155 VGND.n122 0.00556757
R9568 VGND.n7491 VGND.n7406 0.00556757
R9569 VGND.n719 VGND.n718 0.00556757
R9570 VGND.n714 VGND.n705 0.00556757
R9571 VGND.n7548 VGND.n7547 0.00556757
R9572 VGND.n7531 VGND.n7526 0.00556757
R9573 VGND.n7728 VGND.n7727 0.00556757
R9574 VGND.n7742 VGND.n7741 0.00556757
R9575 VGND.n4088 VGND.n4017 0.00556757
R9576 VGND.n3122 VGND.n3121 0.00556757
R9577 VGND.n3105 VGND.n3100 0.00556757
R9578 VGND.n3782 VGND.n3781 0.00556757
R9579 VGND.n3796 VGND.n3795 0.00556757
R9580 VGND.n4359 VGND.n4282 0.00556757
R9581 VGND.n4297 VGND.n4292 0.00556757
R9582 VGND.n2880 VGND.n2879 0.00556757
R9583 VGND.n4691 VGND.n2894 0.00556757
R9584 VGND.n5125 VGND.n5124 0.00556757
R9585 VGND.n4324 VGND.n4319 0.00556757
R9586 VGND.n4801 VGND.n4800 0.00556757
R9587 VGND.n4815 VGND.n4814 0.00556757
R9588 VGND.n2824 VGND.n2752 0.00556757
R9589 VGND.n5202 VGND.n5170 0.00556757
R9590 VGND.n2716 VGND.n2388 0.00556757
R9591 VGND.n1687 VGND.n1686 0.00556757
R9592 VGND.n2414 VGND.n2413 0.00556757
R9593 VGND.n2518 VGND.n2517 0.00556757
R9594 VGND.n2560 VGND.n2559 0.00556757
R9595 VGND.n5418 VGND.n5417 0.00556757
R9596 VGND.n1736 VGND.n1735 0.00556757
R9597 VGND.n2362 VGND.n1696 0.00556757
R9598 VGND.n1381 VGND.n1380 0.00556757
R9599 VGND.n5644 VGND.n5643 0.00556757
R9600 VGND.n1898 VGND.n1866 0.00556757
R9601 VGND.n2319 VGND.n1909 0.00556757
R9602 VGND.n1378 VGND.n1377 0.00556757
R9603 VGND.n5686 VGND.n5681 0.00556757
R9604 VGND.n6714 VGND.n6655 0.00556757
R9605 VGND.n7419 VGND.n7418 0.00556757
R9606 VGND.n7468 VGND.n7465 0.00556757
R9607 VGND.n7993 VGND.n2 0.00556757
R9608 VGND.n6986 VGND.n6985 0.00556757
R9609 VGND.n7030 VGND.n7029 0.00556757
R9610 VGND.n356 VGND.n355 0.00556757
R9611 VGND.n689 VGND.n298 0.00556757
R9612 VGND.n2290 VGND.n2289 0.00554564
R9613 VGND.n1998 VGND.n1997 0.00554564
R9614 VGND.n1216 VGND.n1201 0.00500002
R9615 VGND.n1327 VGND.n1199 0.00500002
R9616 VGND VGND.n2095 0.00490236
R9617 VGND.n5321 VGND.n5320 0.00482801
R9618 VGND.n5233 VGND.n5216 0.00482801
R9619 VGND.n2718 VGND.n2380 0.00482801
R9620 VGND.n2456 VGND.n2455 0.00482801
R9621 VGND.n2140 VGND.n2139 0.00477273
R9622 VGND.n2015 VGND.n2014 0.00477273
R9623 VGND.n5253 VGND.n1652 0.00477273
R9624 VGND.n1545 VGND.n1544 0.00477273
R9625 VGND.n1680 VGND.n1679 0.00477273
R9626 VGND.n2523 VGND.n2522 0.00477273
R9627 VGND.n6157 VGND.n6156 0.00477273
R9628 VGND.n464 VGND.n463 0.00460158
R9629 VGND.n7305 VGND.n937 0.00460158
R9630 VGND.n604 VGND.n586 0.00460158
R9631 VGND.n7892 VGND.n7891 0.00460158
R9632 VGND.n7870 VGND.n7869 0.00460158
R9633 VGND.n3895 VGND.n3646 0.00460158
R9634 VGND.n4520 VGND.n4505 0.00460158
R9635 VGND.n4927 VGND.n2860 0.00460158
R9636 VGND.n1415 VGND.n1354 0.00460158
R9637 VGND.n7144 VGND.n961 0.00460158
R9638 VGND.n7470 VGND.n7409 0.00460158
R9639 VGND.n7476 VGND.n7475 0.00460158
R9640 VGND.n7546 VGND.n7519 0.00460158
R9641 VGND.n3120 VGND.n3093 0.00460158
R9642 VGND.n4312 VGND.n4285 0.00460158
R9643 VGND.n4340 VGND.n4339 0.00460158
R9644 VGND.n2378 VGND.n2377 0.00460158
R9645 VGND.n2335 VGND.n2334 0.00460158
R9646 VGND.n2259 VGND.n2258 0.00460158
R9647 VGND.n292 VGND.n272 0.00460158
R9648 VGND.n727 VGND.n695 0.00460158
R9649 VGND.n7726 VGND.n89 0.00460158
R9650 VGND.n3674 VGND.n3673 0.00460158
R9651 VGND.n4499 VGND.n4498 0.00460158
R9652 VGND.n4799 VGND.n4696 0.00460158
R9653 VGND.n2453 VGND.n2452 0.00460158
R9654 VGND.n5726 VGND.n5661 0.00460158
R9655 VGND.n7023 VGND.n984 0.00460158
R9656 VGND.n154 VGND.n151 0.00440625
R9657 VGND.n7505 VGND.n7504 0.00440625
R9658 VGND.n235 VGND.n234 0.00440625
R9659 VGND.n738 VGND.n255 0.00440625
R9660 VGND VGND.n256 0.00440625
R9661 VGND.n713 VGND.n712 0.00440625
R9662 VGND.n3372 VGND.n3370 0.00440625
R9663 VGND.n3543 VGND 0.00440625
R9664 VGND VGND.n3542 0.00440625
R9665 VGND.n7589 VGND.n7588 0.00440625
R9666 VGND.n7609 VGND.n7608 0.00440625
R9667 VGND.n7690 VGND.n7689 0.00440625
R9668 VGND.n7716 VGND.n7710 0.00440625
R9669 VGND.n7712 VGND 0.00440625
R9670 VGND.n7744 VGND.n7743 0.00440625
R9671 VGND.n3177 VGND.n3176 0.00440625
R9672 VGND VGND.n3329 0.00440625
R9673 VGND.n4189 VGND.n4188 0.00440625
R9674 VGND.n4212 VGND.n4211 0.00440625
R9675 VGND.n3777 VGND.n3776 0.00440625
R9676 VGND VGND.n3730 0.00440625
R9677 VGND.n3798 VGND.n3797 0.00440625
R9678 VGND.n3923 VGND.n3922 0.00440625
R9679 VGND VGND.n4126 0.00440625
R9680 VGND.n4087 VGND.n4086 0.00440625
R9681 VGND.n4360 VGND.n4253 0.00440625
R9682 VGND.n4378 VGND.n4377 0.00440625
R9683 VGND.n4463 VGND.n4462 0.00440625
R9684 VGND.n4488 VGND.n4481 0.00440625
R9685 VGND.n4485 VGND 0.00440625
R9686 VGND.n4690 VGND.n4689 0.00440625
R9687 VGND.n4549 VGND.n4548 0.00440625
R9688 VGND VGND.n4677 0.00440625
R9689 VGND.n5129 VGND.n5128 0.00440625
R9690 VGND.n5153 VGND.n5152 0.00440625
R9691 VGND.n4761 VGND.n4760 0.00440625
R9692 VGND.n4789 VGND.n4782 0.00440625
R9693 VGND.n4786 VGND 0.00440625
R9694 VGND.n4817 VGND.n4816 0.00440625
R9695 VGND.n4965 VGND.n4964 0.00440625
R9696 VGND VGND.n5057 0.00440625
R9697 VGND.n2823 VGND.n2822 0.00440625
R9698 VGND.n5201 VGND.n5199 0.00440625
R9699 VGND.n2700 VGND.n2699 0.00440625
R9700 VGND.n2406 VGND.n2402 0.00440625
R9701 VGND.n2514 VGND.n2513 0.00440625
R9702 VGND.n2546 VGND.n2543 0.00440625
R9703 VGND.n2550 VGND 0.00440625
R9704 VGND.n2562 VGND.n2561 0.00440625
R9705 VGND.n5280 VGND.n5279 0.00440625
R9706 VGND VGND.n1572 0.00440625
R9707 VGND.n1734 VGND.n1731 0.00440625
R9708 VGND.n2347 VGND.n2346 0.00440625
R9709 VGND.n1781 VGND.n1780 0.00440625
R9710 VGND.n5653 VGND.n1395 0.00440625
R9711 VGND.n5649 VGND 0.00440625
R9712 VGND.n5645 VGND.n5635 0.00440625
R9713 VGND.n5526 VGND.n5524 0.00440625
R9714 VGND.n5429 VGND 0.00440625
R9715 VGND.n5419 VGND.n5341 0.00440625
R9716 VGND.n1897 VGND.n1894 0.00440625
R9717 VGND.n2306 VGND 0.00440625
R9718 VGND.n2303 VGND.n2302 0.00440625
R9719 VGND.n5736 VGND.n5735 0.00440625
R9720 VGND.n5715 VGND 0.00440625
R9721 VGND.n5711 VGND.n5709 0.00440625
R9722 VGND VGND.n5696 0.00440625
R9723 VGND.n5685 VGND.n5684 0.00440625
R9724 VGND.n5901 VGND.n5899 0.00440625
R9725 VGND VGND.n1315 0.00440625
R9726 VGND.n2134 VGND.n2132 0.00440625
R9727 VGND.n2274 VGND 0.00440625
R9728 VGND.n2163 VGND.n2162 0.00440625
R9729 VGND.n2097 VGND.n2096 0.00440625
R9730 VGND.n2022 VGND.n2021 0.00440625
R9731 VGND VGND.n6320 0.00440625
R9732 VGND.n6302 VGND.n6291 0.00440625
R9733 VGND.n6226 VGND.n6224 0.00440625
R9734 VGND.n6113 VGND 0.00440625
R9735 VGND.n6866 VGND.n6865 0.00440625
R9736 VGND.n6900 VGND 0.00440625
R9737 VGND.n1020 VGND.n1019 0.00440625
R9738 VGND.n6991 VGND.n6990 0.00440625
R9739 VGND.n7017 VGND.n7012 0.00440625
R9740 VGND VGND.n7015 0.00440625
R9741 VGND.n7032 VGND.n7031 0.00440625
R9742 VGND.n7168 VGND.n7166 0.00440625
R9743 VGND VGND.n7321 0.00440625
R9744 VGND.n2215 VGND.n2176 0.00440625
R9745 VGND.n2227 VGND.n2226 0.00440625
R9746 VGND.n6797 VGND.n6796 0.00440625
R9747 VGND.n6397 VGND.n6396 0.00440625
R9748 VGND.n6425 VGND.n6418 0.00440625
R9749 VGND.n6423 VGND 0.00440625
R9750 VGND.n6456 VGND.n6455 0.00440625
R9751 VGND.n6580 VGND.n6579 0.00440625
R9752 VGND.n6755 VGND 0.00440625
R9753 VGND.n6713 VGND.n6712 0.00440625
R9754 VGND.n7455 VGND.n7454 0.00440625
R9755 VGND.n4 VGND 0.00440625
R9756 VGND.n8003 VGND.n8002 0.00440625
R9757 VGND.n361 VGND.n360 0.00440625
R9758 VGND.n391 VGND.n381 0.00440625
R9759 VGND VGND.n392 0.00440625
R9760 VGND.n396 VGND 0.00440625
R9761 VGND.n688 VGND.n687 0.00440625
R9762 VGND.n561 VGND.n558 0.00440625
R9763 VGND VGND.n7962 0.00440625
R9764 VGND.n6802 VGND.n1030 0.00406061
R9765 VGND.n6549 VGND.n1088 0.00406061
R9766 VGND.n6554 VGND.n6553 0.00406061
R9767 VGND.n2100 VGND.n1970 0.00406061
R9768 VGND.n6297 VGND.n6296 0.00406061
R9769 VGND.n3571 VGND.n3340 0.00406061
R9770 VGND.n7516 VGND.n167 0.00406061
R9771 VGND.n716 VGND.n700 0.00406061
R9772 VGND.n3609 VGND.n3159 0.00406061
R9773 VGND.n7559 VGND.n7558 0.00406061
R9774 VGND.n7738 VGND.n7737 0.00406061
R9775 VGND.n4095 VGND.n4006 0.00406061
R9776 VGND.n4219 VGND.n3134 0.00406061
R9777 VGND.n3792 VGND.n3791 0.00406061
R9778 VGND.n4662 VGND.n2957 0.00406061
R9779 VGND.n4351 VGND.n4345 0.00406061
R9780 VGND.n4693 VGND.n2891 0.00406061
R9781 VGND.n5160 VGND.n2723 0.00406061
R9782 VGND.n4811 VGND.n4810 0.00406061
R9783 VGND.n2870 VGND.n2865 0.00406061
R9784 VGND.n2639 VGND.n2638 0.00406061
R9785 VGND.n5255 VGND.n5254 0.00406061
R9786 VGND.n1598 VGND.n1596 0.00406061
R9787 VGND.n1548 VGND.n1547 0.00406061
R9788 VGND.n5206 VGND.n5169 0.00406061
R9789 VGND.n2411 VGND.n2410 0.00406061
R9790 VGND.n2524 VGND.n2520 0.00406061
R9791 VGND.n2556 VGND.n2555 0.00406061
R9792 VGND.n5356 VGND.n5351 0.00406061
R9793 VGND.n5554 VGND.n1414 0.00406061
R9794 VGND.n2339 VGND.n2338 0.00406061
R9795 VGND.n2295 VGND.n2294 0.00406061
R9796 VGND.n5691 VGND.n5690 0.00406061
R9797 VGND.n5874 VGND.n5873 0.00406061
R9798 VGND.n6259 VGND.n1184 0.00406061
R9799 VGND.n6253 VGND.n1217 0.00406061
R9800 VGND.n6126 VGND.n6038 0.00406061
R9801 VGND.n6721 VGND.n6646 0.00406061
R9802 VGND.n7266 VGND.n7262 0.00406061
R9803 VGND.n7900 VGND.n7899 0.00406061
R9804 VGND.n7136 VGND.n963 0.00406061
R9805 VGND.n584 VGND.n428 0.00406061
R9806 VGND.n8010 VGND.n8009 0.00406061
R9807 VGND.n6815 VGND.n6806 0.00406061
R9808 VGND.n6983 VGND.n6979 0.00406061
R9809 VGND.n691 VGND.n295 0.00406061
R9810 VGND.n6341 VGND.n6333 0.00406061
R9811 VGND.n3456 VGND.n37 0.00393497
R9812 VGND.n3573 VGND.n3572 0.00393497
R9813 VGND.n3575 VGND.n3574 0.00393497
R9814 VGND.n3611 VGND.n3610 0.00393497
R9815 VGND.n3613 VGND.n3612 0.00393497
R9816 VGND.n4093 VGND.n4009 0.00393497
R9817 VGND.n4007 VGND.n2954 0.00393497
R9818 VGND.n4663 VGND.n2956 0.00393497
R9819 VGND.n5048 VGND.n2746 0.00393497
R9820 VGND.n5324 VGND.n5323 0.00393497
R9821 VGND.n5357 VGND.n5350 0.00393497
R9822 VGND.n6034 VGND.n6033 0.00393497
R9823 VGND.n6128 VGND.n1050 0.00393497
R9824 VGND.n6719 VGND.n6647 0.00393497
R9825 VGND.n7898 VGND.n7897 0.00393497
R9826 VGND.n936 VGND.n935 0.00393497
R9827 VGND.n2955 VGND.n2747 0.00393497
R9828 VGND.n5349 VGND.n1240 0.00393497
R9829 VGND.n5214 VGND.n1441 0.00393497
R9830 VGND.n5552 VGND.n1416 0.00393497
R9831 VGND.n5872 VGND.n1329 0.00393497
R9832 VGND.n6552 VGND.n1086 0.00393497
R9833 VGND.n585 VGND.n39 0.00393497
R9834 VGND.n7137 VGND.n962 0.00393497
R9835 VGND.n2871 VGND.n2861 0.00393497
R9836 VGND.n3092 VGND.n3077 0.00393497
R9837 VGND.n3903 VGND.n3902 0.00393497
R9838 VGND.n3645 VGND.n65 0.00393497
R9839 VGND.n7872 VGND.n7871 0.00393497
R9840 VGND.n6550 VGND.n1087 0.00393497
R9841 VGND.n7518 VGND.n7517 0.00393497
R9842 VGND.n7557 VGND.n121 0.00393497
R9843 VGND.n4221 VGND.n4220 0.00393497
R9844 VGND.n4352 VGND.n4341 0.00393497
R9845 VGND.n5162 VGND.n5161 0.00393497
R9846 VGND.n2337 VGND.n2336 0.00393497
R9847 VGND.n2293 VGND.n2292 0.00393497
R9848 VGND.n6804 VGND.n6803 0.00393497
R9849 VGND.n6828 VGND.n1025 0.00393497
R9850 VGND.n7473 VGND.n7472 0.00393497
R9851 VGND.n6816 VGND.n6805 0.00393497
R9852 VGND.n717 VGND.n696 0.00393497
R9853 VGND.n7736 VGND.n88 0.00393497
R9854 VGND.n3790 VGND.n3672 0.00393497
R9855 VGND.n4695 VGND.n4694 0.00393497
R9856 VGND.n4809 VGND.n2878 0.00393497
R9857 VGND.n6447 VGND.n6446 0.00393497
R9858 VGND.n693 VGND.n692 0.00393497
R9859 VGND.n983 VGND.n982 0.00393497
R9860 VGND.n1995 VGND.n1379 0.00393497
R9861 VGND.n5660 VGND.n5659 0.00393497
R9862 VGND.n6342 VGND.n6332 0.00393497
R9863 VGND.n150 VGND.n148 0.00360244
R9864 VGND.n7587 VGND.n7586 0.00360244
R9865 VGND.n5198 VGND.n5196 0.00360244
R9866 VGND.n4187 VGND.n4185 0.00360244
R9867 VGND.n4281 VGND.n4280 0.00360244
R9868 VGND.n5127 VGND.n5126 0.00360244
R9869 VGND.n1738 VGND.n1737 0.00360244
R9870 VGND.n1893 VGND.n1891 0.00360244
R9871 VGND.n2131 VGND.n2129 0.00360244
R9872 VGND.n6864 VGND.n6862 0.00360244
R9873 VGND.n2205 VGND.n2204 0.00360244
R9874 VGND.n7453 VGND.n7451 0.00360244
R9875 VGND.n6130 VGND.n6129 0.00358437
R9876 VGND.n1201 VGND.n1200 0.00358437
R9877 VGND.n2261 VGND.n2260 0.00358437
R9878 VGND.n6331 VGND.n6330 0.00358437
R9879 VGND.n2138 VGND.n2103 0.0033671
R9880 VGND.n2016 VGND.n1994 0.0033671
R9881 VGND.n6158 VGND.n1238 0.0033671
R9882 VGND.n1471 VGND.n1470 0.0032017
R9883 VGND.n1470 VGND.n1469 0.0032017
R9884 VGND.n5237 VGND.n5236 0.0032017
R9885 VGND.n5238 VGND.n5237 0.0032017
R9886 VGND.n5167 VGND.n5166 0.0032017
R9887 VGND.n5166 VGND.n5165 0.0032017
R9888 VGND.n1662 VGND.n1661 0.0032017
R9889 VGND.n1663 VGND.n1662 0.0032017
R9890 VGND.n935 VGND 0.00314375
R9891 VGND.n962 VGND 0.00314375
R9892 VGND.n1025 VGND 0.00314375
R9893 VGND.n982 VGND 0.00314375
R9894 VGND VGND.n3464 0.00310417
R9895 VGND.n4688 VGND.n2896 0.00310417
R9896 VGND.n4651 VGND 0.00310417
R9897 VGND.n4820 VGND.n4819 0.00310417
R9898 VGND.n4951 VGND 0.00310417
R9899 VGND.n2565 VGND.n2564 0.00310417
R9900 VGND VGND.n1748 0.00310417
R9901 VGND.n5631 VGND 0.00310417
R9902 VGND.n7153 VGND 0.00310417
R9903 VGND.n6459 VGND.n6458 0.00310417
R9904 VGND.n464 VGND.n36 0.0028004
R9905 VGND.n7306 VGND.n7305 0.0028004
R9906 VGND.n605 VGND.n604 0.0028004
R9907 VGND.n7144 VGND.n7143 0.0028004
R9908 VGND.n5871 VGND.n1354 0.0028004
R9909 VGND.n4521 VGND.n4520 0.0028004
R9910 VGND.n3901 VGND.n3895 0.0028004
R9911 VGND.n7869 VGND.n7854 0.0028004
R9912 VGND.n7891 VGND.n40 0.0028004
R9913 VGND.n4927 VGND.n4926 0.0028004
R9914 VGND.n7476 VGND.n163 0.0028004
R9915 VGND.n7556 VGND.n7546 0.0028004
R9916 VGND.n3130 VGND.n3120 0.0028004
R9917 VGND.n4353 VGND.n4312 0.0028004
R9918 VGND.n4339 VGND.n2719 0.0028004
R9919 VGND.n2377 VGND.n1693 0.0028004
R9920 VGND.n2334 VGND.n1906 0.0028004
R9921 VGND.n2258 VGND.n1026 0.0028004
R9922 VGND.n7471 VGND.n7470 0.0028004
R9923 VGND.n293 VGND.n292 0.0028004
R9924 VGND.n7024 VGND.n7023 0.0028004
R9925 VGND.n4808 VGND.n4799 0.0028004
R9926 VGND.n4498 VGND.n2887 0.0028004
R9927 VGND.n3789 VGND.n3674 0.0028004
R9928 VGND.n7735 VGND.n7726 0.0028004
R9929 VGND.n727 VGND.n726 0.0028004
R9930 VGND.n2452 VGND.n1388 0.0028004
R9931 VGND.n5727 VGND.n5726 0.0028004
R9932 VGND.n162 VGND.n161 0.00251462
R9933 VGND.n725 VGND.n724 0.00251462
R9934 VGND.n824 VGND.n822 0.00251462
R9935 VGND.n7555 VGND.n7554 0.00251462
R9936 VGND.n7734 VGND.n7733 0.00251462
R9937 VGND.n7821 VGND.n50 0.00251462
R9938 VGND.n3129 VGND.n3128 0.00251462
R9939 VGND.n3788 VGND.n3787 0.00251462
R9940 VGND.n3866 VGND.n3644 0.00251462
R9941 VGND.n4356 VGND.n4354 0.00251462
R9942 VGND.n2886 VGND.n2885 0.00251462
R9943 VGND.n3076 VGND.n3075 0.00251462
R9944 VGND.n5121 VGND.n5119 0.00251462
R9945 VGND.n4807 VGND.n4806 0.00251462
R9946 VGND.n4925 VGND.n4924 0.00251462
R9947 VGND.n5046 VGND.n5045 0.00251462
R9948 VGND.n1728 VGND.n1726 0.00251462
R9949 VGND.n1387 VGND.n1386 0.00251462
R9950 VGND.n1905 VGND.n1904 0.00251462
R9951 VGND.n5730 VGND.n5728 0.00251462
R9952 VGND.n5870 VGND.n5869 0.00251462
R9953 VGND.n6017 VGND.n6016 0.00251462
R9954 VGND.n2827 VGND.n2826 0.00251462
R9955 VGND.n1302 VGND.n1241 0.00251462
R9956 VGND.n4523 VGND.n4522 0.00251462
R9957 VGND.n3900 VGND.n3899 0.00251462
R9958 VGND.n7853 VGND.n7852 0.00251462
R9959 VGND.n3353 VGND.n3352 0.00251462
R9960 VGND.n5640 VGND.n5639 0.00251462
R9961 VGND.n7026 VGND.n7025 0.00251462
R9962 VGND.n7898 VGND.n36 0.00246749
R9963 VGND.n5047 VGND.n2747 0.00246749
R9964 VGND.n6018 VGND.n1240 0.00246749
R9965 VGND.n7306 VGND.n936 0.00246749
R9966 VGND.n6719 VGND.n6718 0.00246749
R9967 VGND.n3572 VGND.n3339 0.00246749
R9968 VGND.n3610 VGND.n3158 0.00246749
R9969 VGND.n4093 VGND.n4092 0.00246749
R9970 VGND.n4664 VGND.n4663 0.00246749
R9971 VGND.n4664 VGND.n2954 0.00246749
R9972 VGND.n4092 VGND.n3613 0.00246749
R9973 VGND.n3575 VGND.n3158 0.00246749
R9974 VGND.n3456 VGND.n3339 0.00246749
R9975 VGND.n5048 VGND.n5047 0.00246749
R9976 VGND.n5358 VGND.n5357 0.00246749
R9977 VGND.n5358 VGND.n5324 0.00246749
R9978 VGND.n6718 VGND.n1050 0.00246749
R9979 VGND.n6033 VGND.n6018 0.00246749
R9980 VGND.n605 VGND.n585 0.00246749
R9981 VGND.n7872 VGND.n40 0.00246749
R9982 VGND.n7854 VGND.n65 0.00246749
R9983 VGND.n3903 VGND.n3901 0.00246749
R9984 VGND.n4521 VGND.n3092 0.00246749
R9985 VGND.n4926 VGND.n2871 0.00246749
R9986 VGND.n6551 VGND.n6550 0.00246749
R9987 VGND.n7143 VGND.n7137 0.00246749
R9988 VGND.n5872 VGND.n5871 0.00246749
R9989 VGND.n5552 VGND.n5551 0.00246749
R9990 VGND.n5551 VGND.n1441 0.00246749
R9991 VGND.n6552 VGND.n6551 0.00246749
R9992 VGND.n7472 VGND.n7471 0.00246749
R9993 VGND.n6827 VGND.n6816 0.00246749
R9994 VGND.n7517 VGND.n163 0.00246749
R9995 VGND.n7557 VGND.n7556 0.00246749
R9996 VGND.n4220 VGND.n3130 0.00246749
R9997 VGND.n4353 VGND.n4352 0.00246749
R9998 VGND.n5161 VGND.n2719 0.00246749
R9999 VGND.n2337 VGND.n1693 0.00246749
R10000 VGND.n2293 VGND.n1906 0.00246749
R10001 VGND.n6803 VGND.n1026 0.00246749
R10002 VGND.n6828 VGND.n6827 0.00246749
R10003 VGND.n692 VGND.n293 0.00246749
R10004 VGND.n5659 VGND.n1388 0.00246749
R10005 VGND.n5727 VGND.n1379 0.00246749
R10006 VGND.n6448 VGND.n6342 0.00246749
R10007 VGND.n7024 VGND.n983 0.00246749
R10008 VGND.n4809 VGND.n4808 0.00246749
R10009 VGND.n4694 VGND.n2887 0.00246749
R10010 VGND.n3790 VGND.n3789 0.00246749
R10011 VGND.n7736 VGND.n7735 0.00246749
R10012 VGND.n726 VGND.n717 0.00246749
R10013 VGND.n6448 VGND.n6447 0.00246749
R10014 VGND.n3800 VGND.n3799 0.00228056
R10015 VGND.n5683 VGND.n1369 0.00228056
R10016 VGND.n7036 VGND.n7033 0.00228056
R10017 VGND.n686 VGND.n685 0.00228056
R10018 VGND.n711 VGND.n710 0.00228056
R10019 VGND.n7746 VGND.n7745 0.00228056
R10020 VGND.n5634 VGND.n5633 0.00228056
R10021 VGND.n6290 VGND.n6289 0.00228056
R10022 VGND.n6440 VGND.n6439 0.00218919
R10023 VGND.n6812 VGND.n6809 0.00218919
R10024 VGND.n6831 VGND.n6830 0.00218919
R10025 VGND.n1022 VGND.n1021 0.00218919
R10026 VGND.n6896 VGND.n6895 0.00218919
R10027 VGND.n6824 VGND.n6823 0.00218919
R10028 VGND.n2213 VGND.n2212 0.00218919
R10029 VGND.n2173 VGND.n2172 0.00218919
R10030 VGND.n2245 VGND.n2244 0.00218919
R10031 VGND.n2250 VGND.n2249 0.00218919
R10032 VGND.n6801 VGND.n1034 0.00218919
R10033 VGND.n2137 VGND.n2136 0.00218919
R10034 VGND.n2157 VGND.n2156 0.00218919
R10035 VGND.n2165 VGND.n2164 0.00218919
R10036 VGND.n2267 VGND.n2266 0.00218919
R10037 VGND.n2099 VGND.n1972 0.00218919
R10038 VGND.n6318 VGND.n6317 0.00218919
R10039 VGND.n3450 VGND.n3449 0.00218919
R10040 VGND.n3558 VGND.n3452 0.00218919
R10041 VGND.n159 VGND.n156 0.00218919
R10042 VGND.n7397 VGND.n7396 0.00218919
R10043 VGND.n7478 VGND.n7477 0.00218919
R10044 VGND.n7483 VGND.n7482 0.00218919
R10045 VGND.n7515 VGND.n171 0.00218919
R10046 VGND.n267 VGND.n266 0.00218919
R10047 VGND.n3164 VGND.n3163 0.00218919
R10048 VGND.n3591 VGND.n3166 0.00218919
R10049 VGND.n7552 VGND.n7549 0.00218919
R10050 VGND.n7524 VGND.n7523 0.00218919
R10051 VGND.n7533 VGND.n7532 0.00218919
R10052 VGND.n7538 VGND.n7537 0.00218919
R10053 VGND.n7560 VGND.n117 0.00218919
R10054 VGND.n98 VGND.n97 0.00218919
R10055 VGND.n3615 VGND.n3614 0.00218919
R10056 VGND.n3618 VGND.n3617 0.00218919
R10057 VGND.n3126 VGND.n3123 0.00218919
R10058 VGND.n3098 VGND.n3097 0.00218919
R10059 VGND.n3107 VGND.n3106 0.00218919
R10060 VGND.n3112 VGND.n3111 0.00218919
R10061 VGND.n4218 VGND.n3138 0.00218919
R10062 VGND.n3742 VGND.n3741 0.00218919
R10063 VGND.n4623 VGND.n4622 0.00218919
R10064 VGND.n4648 VGND.n4625 0.00218919
R10065 VGND.n4358 VGND.n4357 0.00218919
R10066 VGND.n4290 VGND.n4289 0.00218919
R10067 VGND.n4299 VGND.n4298 0.00218919
R10068 VGND.n4304 VGND.n4303 0.00218919
R10069 VGND.n4350 VGND.n4349 0.00218919
R10070 VGND.n4231 VGND.n4230 0.00218919
R10071 VGND.n5123 VGND.n5122 0.00218919
R10072 VGND.n4317 VGND.n4316 0.00218919
R10073 VGND.n4326 VGND.n4325 0.00218919
R10074 VGND.n4331 VGND.n4330 0.00218919
R10075 VGND.n5159 VGND.n2727 0.00218919
R10076 VGND.n4705 VGND.n4704 0.00218919
R10077 VGND.n2829 VGND.n2828 0.00218919
R10078 VGND.n2843 VGND.n2831 0.00218919
R10079 VGND.n1478 VGND.n1477 0.00218919
R10080 VGND.n1481 VGND.n1480 0.00218919
R10081 VGND.n5205 VGND.n5203 0.00218919
R10082 VGND.n2398 VGND.n2397 0.00218919
R10083 VGND.n1683 VGND.n1682 0.00218919
R10084 VGND.n1690 VGND.n1689 0.00218919
R10085 VGND.n2412 VGND.n2408 0.00218919
R10086 VGND.n2429 VGND.n2428 0.00218919
R10087 VGND.n1461 VGND.n1460 0.00218919
R10088 VGND.n5440 VGND.n1463 0.00218919
R10089 VGND.n1730 VGND.n1729 0.00218919
R10090 VGND.n1745 VGND.n1744 0.00218919
R10091 VGND.n2364 VGND.n2363 0.00218919
R10092 VGND.n2369 VGND.n2368 0.00218919
R10093 VGND.n2340 VGND.n1862 0.00218919
R10094 VGND.n1902 VGND.n1899 0.00218919
R10095 VGND.n1918 VGND.n1917 0.00218919
R10096 VGND.n2321 VGND.n2320 0.00218919
R10097 VGND.n2326 VGND.n2325 0.00218919
R10098 VGND.n2296 VGND.n1954 0.00218919
R10099 VGND.n5717 VGND.n5716 0.00218919
R10100 VGND.n1249 VGND.n1248 0.00218919
R10101 VGND.n6000 VGND.n1251 0.00218919
R10102 VGND.n6098 VGND.n6097 0.00218919
R10103 VGND.n6101 VGND.n6100 0.00218919
R10104 VGND.n1052 VGND.n1051 0.00218919
R10105 VGND.n1055 VGND.n1054 0.00218919
R10106 VGND.n7259 VGND.n7258 0.00218919
R10107 VGND.n940 VGND.n939 0.00218919
R10108 VGND.n453 VGND.n452 0.00218919
R10109 VGND.n472 VGND.n455 0.00218919
R10110 VGND.n7421 VGND.n7420 0.00218919
R10111 VGND.n7426 VGND.n7425 0.00218919
R10112 VGND.n8018 VGND.n8017 0.00218919
R10113 VGND.n8015 VGND.n8006 0.00218919
R10114 VGND.n7997 VGND.n7996 0.00218919
R10115 VGND.n999 VGND.n998 0.00218919
R10116 VGND.n286 VGND.n285 0.00218919
R10117 VGND.n2211 VGND.n2209 0.00218193
R10118 VGND.n6717 VGND.n6716 0.00218193
R10119 VGND.n7308 VGND.n7307 0.00218193
R10120 VGND.n489 VGND.n487 0.00218193
R10121 VGND.n4666 VGND.n4665 0.00218193
R10122 VGND.n4091 VGND.n4090 0.00218193
R10123 VGND.n3316 VGND.n3315 0.00218193
R10124 VGND.n3529 VGND.n3528 0.00218193
R10125 VGND.n5360 VGND.n5359 0.00218193
R10126 VGND.n7142 VGND.n7141 0.00218193
R10127 VGND.n608 VGND.n606 0.00218193
R10128 VGND.n5550 VGND.n5549 0.00218193
R10129 VGND.n7411 VGND.n7410 0.00218193
R10130 VGND.n6826 VGND.n6825 0.00218193
R10131 VGND.n353 VGND.n351 0.00218193
R10132 VGND.n6450 VGND.n6449 0.00218193
R10133 VGND.n2289 VGND.n2102 0.00185526
R10134 VGND.n7402 VGND.n7401 0.00180208
R10135 VGND.n7499 VGND.n7498 0.00180208
R10136 VGND.n251 VGND.n250 0.00180208
R10137 VGND VGND.n813 0.00180208
R10138 VGND.n3563 VGND.n3562 0.00180208
R10139 VGND.n3560 VGND.n3559 0.00180208
R10140 VGND.n7597 VGND.n7596 0.00180208
R10141 VGND.n7604 VGND.n7603 0.00180208
R10142 VGND.n7706 VGND.n7705 0.00180208
R10143 VGND.n3597 VGND.n3595 0.00180208
R10144 VGND.n3593 VGND.n3592 0.00180208
R10145 VGND.n4195 VGND.n4194 0.00180208
R10146 VGND.n4203 VGND.n4202 0.00180208
R10147 VGND.n3761 VGND.n3760 0.00180208
R10148 VGND.n3877 VGND 0.00180208
R10149 VGND.n4107 VGND.n4106 0.00180208
R10150 VGND.n4110 VGND.n4109 0.00180208
R10151 VGND.n4366 VGND.n4365 0.00180208
R10152 VGND.n4373 VGND.n4372 0.00180208
R10153 VGND.n4476 VGND.n4475 0.00180208
R10154 VGND.n4653 VGND.n4652 0.00180208
R10155 VGND.n4650 VGND.n4649 0.00180208
R10156 VGND.n5136 VGND.n5135 0.00180208
R10157 VGND.n5144 VGND.n5143 0.00180208
R10158 VGND.n4778 VGND.n4777 0.00180208
R10159 VGND VGND.n4911 0.00180208
R10160 VGND.n2849 VGND.n2847 0.00180208
R10161 VGND.n2845 VGND.n2844 0.00180208
R10162 VGND.n2394 VGND.n2393 0.00180208
R10163 VGND.n2710 VGND.n2708 0.00180208
R10164 VGND.n2538 VGND.n2537 0.00180208
R10165 VGND.n1587 VGND.n1585 0.00180208
R10166 VGND.n1583 VGND.n1582 0.00180208
R10167 VGND.n1742 VGND.n1741 0.00180208
R10168 VGND.n2357 VGND.n2355 0.00180208
R10169 VGND.n1769 VGND.n1768 0.00180208
R10170 VGND.n5446 VGND.n5444 0.00180208
R10171 VGND.n5442 VGND.n5441 0.00180208
R10172 VGND.n1915 VGND.n1914 0.00180208
R10173 VGND.n2313 VGND.n2311 0.00180208
R10174 VGND.n5718 VGND.n5715 0.00180208
R10175 VGND.n6006 VGND.n6004 0.00180208
R10176 VGND.n6002 VGND.n6001 0.00180208
R10177 VGND.n2152 VGND.n2151 0.00180208
R10178 VGND.n2281 VGND.n2279 0.00180208
R10179 VGND.n6320 VGND.n6319 0.00180208
R10180 VGND.n6093 VGND.n6092 0.00180208
R10181 VGND.n6102 VGND.n6095 0.00180208
R10182 VGND.n6872 VGND.n6871 0.00180208
R10183 VGND.n6881 VGND.n6879 0.00180208
R10184 VGND.n7007 VGND.n7006 0.00180208
R10185 VGND.n7278 VGND.n7277 0.00180208
R10186 VGND.n7281 VGND.n7280 0.00180208
R10187 VGND.n2221 VGND.n2220 0.00180208
R10188 VGND.n2237 VGND.n2235 0.00180208
R10189 VGND.n6413 VGND.n6412 0.00180208
R10190 VGND.n6732 VGND.n6731 0.00180208
R10191 VGND.n6735 VGND.n6734 0.00180208
R10192 VGND.n7461 VGND.n7460 0.00180208
R10193 VGND.n5 VGND.n0 0.00180208
R10194 VGND.n377 VGND.n376 0.00180208
R10195 VGND.n478 VGND.n476 0.00180208
R10196 VGND.n474 VGND.n473 0.00180208
R10197 VGND.n6148 VGND.n6147 0.0014919
R10198 VGND.n6149 VGND.n6148 0.0014919
R10199 VGND.n2262 VGND.n2102 0.0014919
R10200 VGND.n6329 VGND.n1113 0.0014919
R10201 VGND.n5320 VGND.n1473 0.00142658
R10202 VGND.n5252 VGND.n5233 0.00142658
R10203 VGND.n5208 VGND.n2718 0.00142658
R10204 VGND.n2456 VGND.n1677 0.00142658
R10205 VGND.n6256 VGND.n1199 0.00140106
R10206 VGND.n6256 VGND.n1216 0.00140106
R10207 VGND.n1472 VGND.n1471 0.00107355
R10208 VGND.n5239 VGND.n5238 0.00107355
R10209 VGND.n5168 VGND.n5167 0.00107355
R10210 VGND.n1664 VGND.n1663 0.00107355
R10211 VGND.n1469 VGND.n1468 0.00107344
R10212 VGND.n1468 VGND.n1467 0.00107344
R10213 VGND.n5235 VGND.n5234 0.00107344
R10214 VGND.n5236 VGND.n5235 0.00107344
R10215 VGND.n5165 VGND.n5164 0.00107344
R10216 VGND.n5164 VGND.n5163 0.00107344
R10217 VGND.n1661 VGND.n1660 0.00107344
R10218 VGND.n1660 VGND.n1659 0.00107344
R10219 VGND.n1473 VGND.n1472 0.00107332
R10220 VGND.n5252 VGND.n5239 0.00107332
R10221 VGND.n5208 VGND.n5168 0.00107332
R10222 VGND.n1677 VGND.n1664 0.00107332
R10223 VPWR.n6043 VPWR 2228.5
R10224 VPWR.n6708 VPWR 1881.54
R10225 VPWR.n954 VPWR 1727.12
R10226 VPWR.n3680 VPWR.n3643 1409.47
R10227 VPWR.n4865 VPWR 1263.87
R10228 VPWR VPWR.n5734 1139.41
R10229 VPWR.n6045 VPWR 1139.41
R10230 VPWR.n2930 VPWR 1052.39
R10231 VPWR.n7274 VPWR 897.968
R10232 VPWR.n6853 VPWR 646.202
R10233 VPWR.n1095 VPWR 646.202
R10234 VPWR VPWR.n2121 646.202
R10235 VPWR VPWR.n5748 597.819
R10236 VPWR.n3118 VPWR 491.784
R10237 VPWR.n5058 VPWR 491.784
R10238 VPWR.n5142 VPWR 491.784
R10239 VPWR VPWR.n6707 491.784
R10240 VPWR.n7584 VPWR 491.784
R10241 VPWR VPWR.n7274 491.784
R10242 VPWR.n953 VPWR 491.784
R10243 VPWR.n442 VPWR 491.784
R10244 VPWR VPWR.n1431 491.784
R10245 VPWR VPWR.n3866 491.784
R10246 VPWR.n1646 VPWR 491.784
R10247 VPWR VPWR.n1481 491.784
R10248 VPWR.n2123 VPWR 491.784
R10249 VPWR.n2122 VPWR 491.784
R10250 VPWR VPWR.n3284 339.046
R10251 VPWR.n45 VPWR 339.046
R10252 VPWR.n955 VPWR 339.046
R10253 VPWR VPWR.n1091 339.046
R10254 VPWR.n1096 VPWR 339.046
R10255 VPWR.n4075 VPWR 339.046
R10256 VPWR.n1734 VPWR 339.046
R10257 VPWR.n1571 VPWR 339.046
R10258 VPWR.n3439 VPWR 339.046
R10259 VPWR.n2560 VPWR 337.368
R10260 VPWR.n5056 VPWR 337.368
R10261 VPWR.n6044 VPWR 316.668
R10262 VPWR.n5468 VPWR 308.834
R10263 VPWR.n4074 VPWR 281.979
R10264 VPWR.n5159 VPWR.t251 252.238
R10265 VPWR.n6481 VPWR.t37 252.238
R10266 VPWR.n6506 VPWR.t31 252.006
R10267 VPWR.n6413 VPWR.t78 251.977
R10268 VPWR.n5669 VPWR.t35 251.977
R10269 VPWR.n5593 VPWR.t203 251.946
R10270 VPWR.n2510 VPWR.t49 236.891
R10271 VPWR.n1342 VPWR.t183 236.891
R10272 VPWR.n5741 VPWR.t253 230.734
R10273 VPWR.n6342 VPWR.t176 230.734
R10274 VPWR.n6175 VPWR.t114 230.734
R10275 VPWR.n3073 VPWR.t207 230.734
R10276 VPWR.n2513 VPWR.t101 230.734
R10277 VPWR.n3167 VPWR.t56 230.734
R10278 VPWR.n3130 VPWR.t65 230.734
R10279 VPWR.n3254 VPWR.t42 230.734
R10280 VPWR.n3226 VPWR.t230 230.734
R10281 VPWR.n3297 VPWR.t69 230.734
R10282 VPWR.n3296 VPWR.t240 230.734
R10283 VPWR.n2639 VPWR.t83 230.734
R10284 VPWR.n6465 VPWR.t44 230.734
R10285 VPWR.n6391 VPWR.t87 230.734
R10286 VPWR.n6490 VPWR.t93 230.734
R10287 VPWR.n6515 VPWR.t155 230.734
R10288 VPWR.n6542 VPWR.t21 230.734
R10289 VPWR.n4976 VPWR.t190 230.734
R10290 VPWR.n4996 VPWR.t30 230.734
R10291 VPWR.n6718 VPWR.t171 230.734
R10292 VPWR.n7592 VPWR.t196 230.734
R10293 VPWR.n7527 VPWR.t1 230.734
R10294 VPWR.n7541 VPWR.t184 230.734
R10295 VPWR.n6641 VPWR.t241 230.734
R10296 VPWR.n5150 VPWR.t123 230.734
R10297 VPWR.n5177 VPWR.t4 230.734
R10298 VPWR.n5196 VPWR.t10 230.734
R10299 VPWR.n6935 VPWR.t38 230.734
R10300 VPWR.n5515 VPWR.t149 230.734
R10301 VPWR.n5540 VPWR.t153 230.734
R10302 VPWR.n5567 VPWR.t164 230.734
R10303 VPWR.n5451 VPWR.t174 230.734
R10304 VPWR.n7101 VPWR.t191 230.734
R10305 VPWR.n5257 VPWR.t175 230.734
R10306 VPWR.n5281 VPWR.t165 230.734
R10307 VPWR.n1192 VPWR.t116 230.734
R10308 VPWR.n4670 VPWR.t154 230.734
R10309 VPWR.n4649 VPWR.t91 230.734
R10310 VPWR.n4547 VPWR.t124 230.734
R10311 VPWR.n4516 VPWR.t34 230.734
R10312 VPWR.n1168 VPWR.t106 230.734
R10313 VPWR.n1017 VPWR.t122 230.734
R10314 VPWR.n3885 VPWR.t152 230.734
R10315 VPWR.n3881 VPWR.t161 230.734
R10316 VPWR.n4336 VPWR.t215 230.734
R10317 VPWR.n1351 VPWR.t232 230.734
R10318 VPWR.n1315 VPWR.t194 230.734
R10319 VPWR.n1970 VPWR.t159 230.734
R10320 VPWR.n2135 VPWR.t67 230.734
R10321 VPWR.n3546 VPWR.t142 230.734
R10322 VPWR.n1776 VPWR.t72 230.734
R10323 VPWR.n3666 VPWR.t226 230.734
R10324 VPWR.n2307 VPWR.t90 230.734
R10325 VPWR.n2307 VPWR.t227 230.734
R10326 VPWR.n3426 VPWR.t150 230.734
R10327 VPWR.n2253 VPWR.t177 230.734
R10328 VPWR.n2877 VPWR.t108 230.734
R10329 VPWR.n2959 VPWR.t213 230.734
R10330 VPWR.n2229 VPWR.t206 230.734
R10331 VPWR.n2908 VPWR.t131 230.734
R10332 VPWR.n2209 VPWR.t229 230.734
R10333 VPWR.n5868 VPWR.t157 230.734
R10334 VPWR.n5734 VPWR 221.964
R10335 VPWR.n6045 VPWR 221.964
R10336 VPWR VPWR.n6044 221.964
R10337 VPWR VPWR.n6043 221.964
R10338 VPWR.n5748 VPWR 219.004
R10339 VPWR VPWR.n3117 182.952
R10340 VPWR.n3285 VPWR 182.952
R10341 VPWR.n6854 VPWR 182.952
R10342 VPWR.n7275 VPWR 182.952
R10343 VPWR.n376 VPWR 182.952
R10344 VPWR VPWR.n4074 181.273
R10345 VPWR.n1476 VPWR.t16 179.971
R10346 VPWR.n5063 VPWR 179.595
R10347 VPWR.n5057 VPWR 179.595
R10348 VPWR VPWR.n5464 179.595
R10349 VPWR VPWR.n4921 179.595
R10350 VPWR.n5312 VPWR 179.595
R10351 VPWR.n5311 VPWR 179.595
R10352 VPWR.n956 VPWR 179.595
R10353 VPWR.n952 VPWR 179.595
R10354 VPWR.n377 VPWR 179.595
R10355 VPWR.n3867 VPWR 179.595
R10356 VPWR.n1645 VPWR 179.595
R10357 VPWR VPWR.n2805 179.595
R10358 VPWR.n2930 VPWR 179.595
R10359 VPWR.n2929 VPWR 179.595
R10360 VPWR.n3438 VPWR 179.595
R10361 VPWR.n3306 VPWR.t0 178.661
R10362 VPWR.n3306 VPWR.t205 178.661
R10363 VPWR.n2561 VPWR.t63 178.661
R10364 VPWR.n2415 VPWR.t163 178.661
R10365 VPWR.n2582 VPWR.t111 178.661
R10366 VPWR.n2582 VPWR.t46 178.661
R10367 VPWR.n54 VPWR.t29 178.661
R10368 VPWR.n54 VPWR.t228 178.661
R10369 VPWR.n50 VPWR.t245 178.661
R10370 VPWR.n6380 VPWR.t82 178.661
R10371 VPWR.n6380 VPWR.t9 178.661
R10372 VPWR.n6383 VPWR.t92 178.661
R10373 VPWR.n5004 VPWR.t141 178.661
R10374 VPWR.n5096 VPWR.t52 178.661
R10375 VPWR.n5095 VPWR.t102 178.661
R10376 VPWR.n5095 VPWR.t33 178.661
R10377 VPWR.n174 VPWR.t84 178.661
R10378 VPWR.n174 VPWR.t25 178.661
R10379 VPWR.n7444 VPWR.t20 178.661
R10380 VPWR.n7444 VPWR.t136 178.661
R10381 VPWR.n5467 VPWR.t208 178.661
R10382 VPWR.n6822 VPWR.t32 178.661
R10383 VPWR.n5429 VPWR.t238 178.661
R10384 VPWR.n5429 VPWR.t172 178.661
R10385 VPWR.n7329 VPWR.t133 178.661
R10386 VPWR.n7329 VPWR.t80 178.661
R10387 VPWR.n7071 VPWR.t120 178.661
R10388 VPWR.n7272 VPWR.t192 178.661
R10389 VPWR.n5353 VPWR.t125 178.661
R10390 VPWR.n5353 VPWR.t62 178.661
R10391 VPWR.n5347 VPWR.t70 178.661
R10392 VPWR.n4800 VPWR.t252 178.661
R10393 VPWR.n4800 VPWR.t198 178.661
R10394 VPWR.n583 VPWR.t40 178.661
R10395 VPWR.n639 VPWR.t218 178.661
R10396 VPWR.n479 VPWR.t8 178.661
R10397 VPWR.n479 VPWR.t200 178.661
R10398 VPWR.n477 VPWR.t156 178.661
R10399 VPWR.n342 VPWR.t118 178.661
R10400 VPWR.n342 VPWR.t58 178.661
R10401 VPWR.n1021 VPWR.t145 178.661
R10402 VPWR.n1021 VPWR.t81 178.661
R10403 VPWR.n3888 VPWR.t224 178.661
R10404 VPWR.n3888 VPWR.t162 178.661
R10405 VPWR.n1229 VPWR.t146 178.661
R10406 VPWR.n1229 VPWR.t95 178.661
R10407 VPWR.n431 VPWR.t236 178.661
R10408 VPWR.n1528 VPWR.t48 178.661
R10409 VPWR.n3998 VPWR.t160 178.661
R10410 VPWR.n3998 VPWR.t28 178.661
R10411 VPWR.n4197 VPWR.t166 178.661
R10412 VPWR.n1961 VPWR.t169 178.661
R10413 VPWR.n1848 VPWR.t15 178.661
R10414 VPWR.n1848 VPWR.t217 178.661
R10415 VPWR.n1675 VPWR.t128 178.661
R10416 VPWR.n1675 VPWR.t73 178.661
R10417 VPWR.n1579 VPWR.t64 178.661
R10418 VPWR.n1583 VPWR.t26 178.661
R10419 VPWR.n2126 VPWR.t247 178.661
R10420 VPWR.n3591 VPWR.t119 178.661
R10421 VPWR.n3648 VPWR.t27 178.661
R10422 VPWR.n3648 VPWR.t221 178.661
R10423 VPWR.n2292 VPWR.t137 178.661
R10424 VPWR.n2292 VPWR.t85 178.661
R10425 VPWR.n2693 VPWR.t243 178.661
R10426 VPWR.n2693 VPWR.t189 178.661
R10427 VPWR.n2696 VPWR.t195 178.661
R10428 VPWR.n2944 VPWR.t110 178.661
R10429 VPWR.n2435 VPWR.t43 178.406
R10430 VPWR.n3234 VPWR.t2 177.762
R10431 VPWR.n5173 VPWR.t36 177.762
R10432 VPWR.n6957 VPWR.t14 177.762
R10433 VPWR.n1142 VPWR.t212 177.762
R10434 VPWR VPWR.t170 177.762
R10435 VPWR.n3776 VPWR.t250 174.971
R10436 VPWR.n6402 VPWR.n6401 169.036
R10437 VPWR.n5110 VPWR.n5109 169.036
R10438 VPWR.n6286 VPWR.t201 166.282
R10439 VPWR.n6305 VPWR.t181 166.282
R10440 VPWR.n6059 VPWR.t100 166.282
R10441 VPWR.n2602 VPWR.t88 166.282
R10442 VPWR.n5897 VPWR.t168 166.282
R10443 VPWR.n5931 VPWR.t167 166.282
R10444 VPWR.n3777 VPWR.t185 143.667
R10445 VPWR.n2416 VPWR.t147 141.607
R10446 VPWR.n5184 VPWR.t86 141.607
R10447 VPWR.n4869 VPWR.t178 141.008
R10448 VPWR.n1139 VPWR.t117 140.364
R10449 VPWR.n1643 VPWR.t158 140.364
R10450 VPWR.n3230 VPWR.t75 138.72
R10451 VPWR.n1336 VPWR.t235 134.994
R10452 VPWR.n5738 VPWR.t182 134.964
R10453 VPWR.n6135 VPWR.t66 134.964
R10454 VPWR.n6054 VPWR.t138 134.964
R10455 VPWR.n2584 VPWR.t89 134.964
R10456 VPWR.n46 VPWR.t54 134.964
R10457 VPWR.n38 VPWR.t239 134.964
R10458 VPWR.n35 VPWR.t222 134.964
R10459 VPWR.n5020 VPWR.t214 134.964
R10460 VPWR.n7438 VPWR.t39 134.964
R10461 VPWR.n4923 VPWR.t45 134.964
R10462 VPWR.n6862 VPWR.t132 134.964
R10463 VPWR.n7336 VPWR.t210 134.964
R10464 VPWR.n5348 VPWR.t104 134.964
R10465 VPWR.n5378 VPWR.t144 134.964
R10466 VPWR.n319 VPWR.t211 134.964
R10467 VPWR.n903 VPWR.t233 134.964
R10468 VPWR.n896 VPWR.t7 134.964
R10469 VPWR.n808 VPWR.t50 134.964
R10470 VPWR.n755 VPWR.t6 134.964
R10471 VPWR.n508 VPWR.t231 134.964
R10472 VPWR.n4499 VPWR.t223 134.964
R10473 VPWR.n3995 VPWR.t180 134.964
R10474 VPWR.n1952 VPWR.t121 134.964
R10475 VPWR.n1863 VPWR.t151 134.964
R10476 VPWR.n1870 VPWR.t47 134.964
R10477 VPWR.n1877 VPWR.t109 134.964
R10478 VPWR.n2145 VPWR.t148 134.964
R10479 VPWR.n1602 VPWR.t129 134.964
R10480 VPWR.n2797 VPWR.t219 134.964
R10481 VPWR.n2706 VPWR.t220 134.964
R10482 VPWR.n2892 VPWR.t139 134.964
R10483 VPWR.n5853 VPWR.t94 134.964
R10484 VPWR VPWR.n5057 129.24
R10485 VPWR VPWR.n5056 129.24
R10486 VPWR VPWR.n4865 129.24
R10487 VPWR.n6148 VPWR.n5826 126.659
R10488 VPWR.n2560 VPWR 125.883
R10489 VPWR.n3118 VPWR 125.883
R10490 VPWR.n3284 VPWR 125.883
R10491 VPWR.n3285 VPWR 125.883
R10492 VPWR.n5063 VPWR 125.883
R10493 VPWR VPWR.n5058 125.883
R10494 VPWR VPWR.n45 125.883
R10495 VPWR.n5142 VPWR 125.883
R10496 VPWR.n6707 VPWR 125.883
R10497 VPWR.n6708 VPWR 125.883
R10498 VPWR.n7584 VPWR 125.883
R10499 VPWR VPWR.n7583 125.883
R10500 VPWR.n5464 VPWR 125.883
R10501 VPWR.n5468 VPWR 125.883
R10502 VPWR VPWR.n4921 125.883
R10503 VPWR.n6854 VPWR 125.883
R10504 VPWR VPWR.n6853 125.883
R10505 VPWR.n5312 VPWR 125.883
R10506 VPWR.n956 VPWR 125.883
R10507 VPWR VPWR.n955 125.883
R10508 VPWR VPWR.n954 125.883
R10509 VPWR VPWR.n953 125.883
R10510 VPWR VPWR.n952 125.883
R10511 VPWR.n1091 VPWR 125.883
R10512 VPWR.n1096 VPWR 125.883
R10513 VPWR VPWR.n1095 125.883
R10514 VPWR VPWR.n377 125.883
R10515 VPWR VPWR.n376 125.883
R10516 VPWR.n442 VPWR 125.883
R10517 VPWR.n3867 VPWR 125.883
R10518 VPWR.n1646 VPWR 125.883
R10519 VPWR VPWR.n1645 125.883
R10520 VPWR VPWR.n1481 125.883
R10521 VPWR.n4075 VPWR 125.883
R10522 VPWR.n1734 VPWR 125.883
R10523 VPWR.n2123 VPWR 125.883
R10524 VPWR VPWR.n2122 125.883
R10525 VPWR VPWR.n1571 125.883
R10526 VPWR VPWR.n2929 125.883
R10527 VPWR.n3439 VPWR 125.883
R10528 VPWR VPWR.n3438 125.883
R10529 VPWR.n3117 VPWR 124.206
R10530 VPWR VPWR.n5311 124.206
R10531 VPWR.n7275 VPWR 124.206
R10532 VPWR.n1430 VPWR 124.206
R10533 VPWR.n1431 VPWR 124.206
R10534 VPWR.n3866 VPWR 124.206
R10535 VPWR.n2121 VPWR 124.206
R10536 VPWR.n2805 VPWR 124.206
R10537 VPWR.n7583 VPWR.n7582 120.481
R10538 VPWR.n6853 VPWR.n6852 120.481
R10539 VPWR.n7276 VPWR.n7275 120.481
R10540 VPWR.n952 VPWR.n951 120.481
R10541 VPWR.n953 VPWR.n577 120.481
R10542 VPWR.n4074 VPWR.n1521 120.481
R10543 VPWR.n2121 VPWR.n2120 120.481
R10544 VPWR.n3438 VPWR.n3437 120.481
R10545 VPWR.n6044 VPWR.n5830 120.481
R10546 VPWR.n6046 VPWR.n6045 120.481
R10547 VPWR.n6219 VPWR.n5748 120.481
R10548 VPWR.n6264 VPWR.n5734 120.481
R10549 VPWR.n6709 VPWR.n6708 120.481
R10550 VPWR.n5500 VPWR.n5468 120.481
R10551 VPWR.n5313 VPWR.n5312 120.481
R10552 VPWR.n957 VPWR.n956 120.481
R10553 VPWR.n1647 VPWR.n1646 120.481
R10554 VPWR.n2122 VPWR.n1578 120.481
R10555 VPWR.n2929 VPWR.n2928 120.481
R10556 VPWR.n6043 VPWR.n6042 120.481
R10557 VPWR.n4197 VPWR.n1481 119.094
R10558 VPWR.n3119 VPWR.n3118 118.513
R10559 VPWR.n3868 VPWR.n3867 117.906
R10560 VPWR.n2561 VPWR.n2560 117.627
R10561 VPWR.n3286 VPWR.n3285 116.73
R10562 VPWR.n6523 VPWR.n5058 116.73
R10563 VPWR.n5056 VPWR.n31 116.73
R10564 VPWR.n7674 VPWR.n45 116.73
R10565 VPWR.n5057 VPWR.n5055 116.73
R10566 VPWR.n6707 VPWR.n6706 116.73
R10567 VPWR.n7585 VPWR.n7584 116.73
R10568 VPWR.n5189 VPWR.n5142 116.73
R10569 VPWR.n6855 VPWR.n6854 116.73
R10570 VPWR.n6953 VPWR.n4921 116.73
R10571 VPWR.n5560 VPWR.n5464 116.73
R10572 VPWR.n5311 VPWR.n5310 116.73
R10573 VPWR.n7274 VPWR.n7273 116.73
R10574 VPWR.n7098 VPWR.n4865 116.73
R10575 VPWR.n955 VPWR.n575 116.73
R10576 VPWR.n954 VPWR.n576 116.73
R10577 VPWR.n1134 VPWR.n1096 116.73
R10578 VPWR.n376 VPWR.n367 116.73
R10579 VPWR.n4622 VPWR.n377 116.73
R10580 VPWR.n1095 VPWR.n395 116.73
R10581 VPWR.n1430 VPWR.n1429 116.73
R10582 VPWR.n3866 VPWR.n3865 116.73
R10583 VPWR.n4359 VPWR.n1431 116.73
R10584 VPWR.n1645 VPWR.n1641 116.73
R10585 VPWR.n4076 VPWR.n4075 116.73
R10586 VPWR.n3636 VPWR.n1571 116.73
R10587 VPWR.n2124 VPWR.n2123 116.73
R10588 VPWR.n1735 VPWR.n1734 116.73
R10589 VPWR.n2931 VPWR.n2930 116.73
R10590 VPWR.n3440 VPWR.n3439 116.73
R10591 VPWR.n2805 VPWR.n2796 116.73
R10592 VPWR.n5064 VPWR.n5063 116.728
R10593 VPWR.n1189 VPWR.n1091 116.728
R10594 VPWR.n1324 VPWR.n442 116.728
R10595 VPWR.n6147 VPWR.n6146 114.165
R10596 VPWR.n7668 VPWR.t249 95.6157
R10597 VPWR.n5476 VPWR.t143 95.615
R10598 VPWR.n2430 VPWR.t188 95.5078
R10599 VPWR.n7722 VPWR.t199 95.5078
R10600 VPWR.n7520 VPWR.t197 95.5078
R10601 VPWR.n5091 VPWR.t41 95.5078
R10602 VPWR.n277 VPWR.t22 95.5078
R10603 VPWR.n4868 VPWR.t68 95.5078
R10604 VPWR.n5237 VPWR.t103 95.5078
R10605 VPWR.n645 VPWR.t5 95.5078
R10606 VPWR.n4487 VPWR.t3 95.5078
R10607 VPWR.n4065 VPWR.t244 95.5078
R10608 VPWR.n1531 VPWR.t13 95.5078
R10609 VPWR.n1733 VPWR.t24 95.5078
R10610 VPWR.n1569 VPWR.t96 95.5078
R10611 VPWR.n7232 VPWR.t193 95.5071
R10612 VPWR.n642 VPWR.t254 95.5071
R10613 VPWR.n337 VPWR.t23 95.5071
R10614 VPWR.n374 VPWR.t130 95.5071
R10615 VPWR.n1225 VPWR.t204 95.5071
R10616 VPWR.n3302 VPWR.t113 95.034
R10617 VPWR.n2431 VPWR.t242 93.6187
R10618 VPWR.n6401 VPWR.t57 93.6187
R10619 VPWR.n5109 VPWR.t18 93.6187
R10620 VPWR.n6686 VPWR.t11 93.5832
R10621 VPWR.n3313 VPWR.t17 93.2069
R10622 VPWR.n5062 VPWR.t98 93.0776
R10623 VPWR.n5144 VPWR.t53 93.0776
R10624 VPWR.n7681 VPWR.t248 91.34
R10625 VPWR.n170 VPWR.t71 91.34
R10626 VPWR.n7359 VPWR.t134 91.34
R10627 VPWR.n683 VPWR.t60 91.34
R10628 VPWR.n4657 VPWR.t74 91.34
R10629 VPWR.n1374 VPWR.t246 91.34
R10630 VPWR.n4213 VPWR.t225 91.34
R10631 VPWR.n3628 VPWR.t97 91.34
R10632 VPWR.n2238 VPWR.t107 91.34
R10633 VPWR.n2858 VPWR.t115 91.34
R10634 VPWR.n7598 VPWR.t51 91.34
R10635 VPWR.n4918 VPWR.t127 91.34
R10636 VPWR.n5305 VPWR.t76 91.34
R10637 VPWR.n1026 VPWR.t126 91.34
R10638 VPWR.n4073 VPWR.t61 91.34
R10639 VPWR.n2001 VPWR.t79 91.34
R10640 VPWR.n2722 VPWR.t140 91.34
R10641 VPWR.n2328 VPWR.t237 91.34
R10642 VPWR.n5046 VPWR.t186 91.2541
R10643 VPWR.n6827 VPWR.t59 91.2541
R10644 VPWR.n7104 VPWR.t112 91.2541
R10645 VPWR.n2423 VPWR.t12 91.2541
R10646 VPWR.n3276 VPWR.t55 91.2541
R10647 VPWR.n7228 VPWR.t216 91.2541
R10648 VPWR.n3876 VPWR.t19 91.2541
R10649 VPWR.n3604 VPWR.t173 91.2541
R10650 VPWR.n3674 VPWR.t135 89.7
R10651 VPWR.n4510 VPWR.t77 88.7695
R10652 VPWR.n7082 VPWR.t202 88.005
R10653 VPWR.n3273 VPWR.t234 86.1982
R10654 VPWR.n6149 VPWR.n6148 76.0005
R10655 VPWR.n3146 VPWR.n3145 76.0005
R10656 VPWR.n5551 VPWR.n5550 76.0005
R10657 VPWR.n7132 VPWR.n7131 76.0005
R10658 VPWR.n6034 VPWR.n6033 76.0005
R10659 VPWR.n3284 VPWR.n3283 60.2417
R10660 VPWR.n3117 VPWR.n3116 60.2417
R10661 VPWR.n6147 VPWR.t99 50.5057
R10662 VPWR.n3144 VPWR.t187 50.5057
R10663 VPWR.n5549 VPWR.t209 50.5057
R10664 VPWR.n7130 VPWR.t179 50.5057
R10665 VPWR.n6032 VPWR.t105 50.5057
R10666 VPWR.n6855 VPWR.n6798 34.6358
R10667 VPWR.n6961 VPWR.n4920 34.6358
R10668 VPWR.n7346 VPWR.n7345 34.6358
R10669 VPWR.n1858 VPWR.n1845 34.6358
R10670 VPWR.n3625 VPWR.n1575 34.6358
R10671 VPWR.n2701 VPWR.n2692 34.6358
R10672 VPWR.n3440 VPWR.n2212 34.6358
R10673 VPWR.n2931 VPWR.n2804 34.6358
R10674 VPWR.n6298 VPWR.n6297 34.6358
R10675 VPWR.n6299 VPWR.n6298 34.6358
R10676 VPWR.n6122 VPWR.n6121 34.6358
R10677 VPWR.n3235 VPWR.n3234 34.6358
R10678 VPWR.n67 VPWR.n48 34.6358
R10679 VPWR.n63 VPWR.n48 34.6358
R10680 VPWR.n7686 VPWR.n7685 34.6358
R10681 VPWR.n5055 VPWR.n4980 34.6358
R10682 VPWR.n5032 VPWR.n5031 34.6358
R10683 VPWR.n7458 VPWR.n7439 34.6358
R10684 VPWR.n6839 VPWR.n6838 34.6358
R10685 VPWR.n6805 VPWR.n6798 34.6358
R10686 VPWR.n6973 VPWR.n6972 34.6358
R10687 VPWR.n6953 VPWR.n6952 34.6358
R10688 VPWR.n5440 VPWR.n5427 34.6358
R10689 VPWR.n7350 VPWR.n7326 34.6358
R10690 VPWR.n7280 VPWR.n290 34.6358
R10691 VPWR.n7124 VPWR.n4863 34.6358
R10692 VPWR.n5361 VPWR.n5360 34.6358
R10693 VPWR.n5376 VPWR.n5346 34.6358
R10694 VPWR.n4821 VPWR.n4820 34.6358
R10695 VPWR.n4830 VPWR.n4829 34.6358
R10696 VPWR.n658 VPWR.n657 34.6358
R10697 VPWR.n784 VPWR.n576 34.6358
R10698 VPWR.n638 VPWR.n575 34.6358
R10699 VPWR.n4623 VPWR.n4622 34.6358
R10700 VPWR.n4485 VPWR.n398 34.6358
R10701 VPWR.n1134 VPWR.n1097 34.6358
R10702 VPWR.n1135 VPWR.n1134 34.6358
R10703 VPWR.n1146 VPWR.n1145 34.6358
R10704 VPWR.n3858 VPWR.n3816 34.6358
R10705 VPWR.n3854 VPWR.n3816 34.6358
R10706 VPWR.n3859 VPWR.n3858 34.6358
R10707 VPWR.n3865 VPWR.n3780 34.6358
R10708 VPWR.n4359 VPWR.n1432 34.6358
R10709 VPWR.n4360 VPWR.n4359 34.6358
R10710 VPWR.n4106 VPWR.n4105 34.6358
R10711 VPWR.n4113 VPWR.n4112 34.6358
R10712 VPWR.n4119 VPWR.n1520 34.6358
R10713 VPWR.n4177 VPWR.n4176 34.6358
R10714 VPWR.n4176 VPWR.n1484 34.6358
R10715 VPWR.n4227 VPWR.n4226 34.6358
R10716 VPWR.n2012 VPWR.n2011 34.6358
R10717 VPWR.n2011 VPWR.n1641 34.6358
R10718 VPWR.n1701 VPWR.n1700 34.6358
R10719 VPWR.n1749 VPWR.n1748 34.6358
R10720 VPWR.n1789 VPWR.n1735 34.6358
R10721 VPWR.n3637 VPWR.n3636 34.6358
R10722 VPWR.n2976 VPWR.n2796 34.6358
R10723 VPWR.n2697 VPWR.n2692 34.6358
R10724 VPWR.n2987 VPWR.n2793 34.6358
R10725 VPWR.n2982 VPWR.n2794 34.6358
R10726 VPWR.n2816 VPWR.n2804 34.6358
R10727 VPWR.n2932 VPWR.n2931 34.6358
R10728 VPWR.n5891 VPWR.n5832 34.6358
R10729 VPWR.n5943 VPWR.n5926 34.6358
R10730 VPWR.n767 VPWR.n766 33.6462
R10731 VPWR.n3837 VPWR.n3819 33.6462
R10732 VPWR.n4379 VPWR.n4378 33.6462
R10733 VPWR.n4383 VPWR.n4382 33.6462
R10734 VPWR.n4006 VPWR.n4005 32.377
R10735 VPWR.n1129 VPWR.n1098 32.0005
R10736 VPWR.n1696 VPWR.n1673 32.0005
R10737 VPWR.n2016 VPWR.n2015 30.8711
R10738 VPWR.n4120 VPWR.n4119 30.4946
R10739 VPWR.n5055 VPWR.n4981 30.1181
R10740 VPWR.n2943 VPWR.n2801 30.1181
R10741 VPWR.n490 VPWR.n476 29.0829
R10742 VPWR.n6739 VPWR.n6738 28.9887
R10743 VPWR.n4460 VPWR 28.6123
R10744 VPWR.n7583 VPWR 28.5341
R10745 VPWR VPWR.n1430 28.5341
R10746 VPWR VPWR.n6256 28.2358
R10747 VPWR.n2595 VPWR 28.2358
R10748 VPWR VPWR.n7697 28.2358
R10749 VPWR.n662 VPWR 28.2358
R10750 VPWR.n1858 VPWR 28.2358
R10751 VPWR.n2526 VPWR 28.2358
R10752 VPWR.n3235 VPWR 28.2358
R10753 VPWR.n3865 VPWR.n3781 28.2358
R10754 VPWR.n7273 VPWR.n292 27.8593
R10755 VPWR.n817 VPWR 27.8593
R10756 VPWR.n1744 VPWR.n1586 27.8593
R10757 VPWR.n5944 VPWR.n5943 27.8593
R10758 VPWR.n4663 VPWR.n4662 27.2962
R10759 VPWR.n7080 VPWR.n4867 27.2033
R10760 VPWR.n6215 VPWR.n6214 27.0566
R10761 VPWR.n5444 VPWR.n5427 27.0566
R10762 VPWR.n4347 VPWR.n4346 27.0566
R10763 VPWR.n1787 VPWR.n1786 27.0566
R10764 VPWR.n3433 VPWR.n2213 27.0566
R10765 VPWR.n2221 VPWR.n2220 27.0566
R10766 VPWR.n3441 VPWR.n3440 26.7859
R10767 VPWR.n4622 VPWR.n378 26.7859
R10768 VPWR.n6229 VPWR.n5745 26.7859
R10769 VPWR.n6161 VPWR.n6160 26.7859
R10770 VPWR.n5012 VPWR.n5011 26.7859
R10771 VPWR.n6735 VPWR.n6734 26.7859
R10772 VPWR.n6627 VPWR.n6626 26.7859
R10773 VPWR.n6920 VPWR.n4926 26.7859
R10774 VPWR.n1987 VPWR.n1986 26.7859
R10775 VPWR.n2530 VPWR.n2529 26.7299
R10776 VPWR.n1242 VPWR.n1241 26.7299
R10777 VPWR.n3123 VPWR.n2416 26.2083
R10778 VPWR.n5185 VPWR.n5184 26.2083
R10779 VPWR.n6292 VPWR.n6291 25.6005
R10780 VPWR.n6303 VPWR.n6280 25.6005
R10781 VPWR.n6156 VPWR.n6155 25.6005
R10782 VPWR.n6128 VPWR.n6127 25.6005
R10783 VPWR.n1234 VPWR.n1233 25.6005
R10784 VPWR.n1857 VPWR.n1846 25.6005
R10785 VPWR.n5955 VPWR.n5922 25.6005
R10786 VPWR.n5945 VPWR.n5924 25.6005
R10787 VPWR.n5937 VPWR.n5936 25.6005
R10788 VPWR.n6297 VPWR.n6282 25.224
R10789 VPWR.n6122 VPWR.n6051 25.224
R10790 VPWR.n2436 VPWR.n2428 25.224
R10791 VPWR.n2531 VPWR.n2517 25.224
R10792 VPWR.n2531 VPWR.n2530 25.224
R10793 VPWR.n1243 VPWR.n1242 25.224
R10794 VPWR.n1852 VPWR.n1847 25.224
R10795 VPWR.n2713 VPWR.n2691 25.224
R10796 VPWR.n5951 VPWR.n5950 25.224
R10797 VPWR.n5927 VPWR.n5926 25.224
R10798 VPWR.n7710 VPWR.n7709 25.1912
R10799 VPWR.n6856 VPWR.n6855 25.1912
R10800 VPWR.n4493 VPWR.n395 25.1912
R10801 VPWR.n4020 VPWR.n4019 25.1912
R10802 VPWR.n1793 VPWR.n1735 25.1912
R10803 VPWR.n3636 VPWR.n1574 25.1912
R10804 VPWR.n6256 VPWR.n5736 25.1912
R10805 VPWR.n6121 VPWR.n6052 25.1912
R10806 VPWR.n6115 VPWR.n6055 25.1912
R10807 VPWR.n76 VPWR.n75 25.1912
R10808 VPWR.n7685 VPWR.n42 25.1912
R10809 VPWR.n7691 VPWR.n7690 25.1912
R10810 VPWR.n7697 VPWR.n37 25.1912
R10811 VPWR.n7716 VPWR.n7715 25.1912
R10812 VPWR.n5031 VPWR.n5019 25.1912
R10813 VPWR.n5025 VPWR.n5022 25.1912
R10814 VPWR.n192 VPWR.n171 25.1912
R10815 VPWR.n7465 VPWR.n7464 25.1912
R10816 VPWR.n6838 VPWR.n6803 25.1912
R10817 VPWR.n6983 VPWR.n6982 25.1912
R10818 VPWR.n6972 VPWR.n4919 25.1912
R10819 VPWR.n6952 VPWR.n4922 25.1912
R10820 VPWR.n7351 VPWR.n7350 25.1912
R10821 VPWR.n7239 VPWR.n7238 25.1912
R10822 VPWR.n7258 VPWR.n7257 25.1912
R10823 VPWR.n5360 VPWR.n5351 25.1912
R10824 VPWR.n681 VPWR.n638 25.1912
R10825 VPWR.n1951 VPWR.n1648 25.1912
R10826 VPWR.n1862 VPWR.n1845 25.1912
R10827 VPWR.n2859 VPWR.n2856 25.1912
R10828 VPWR.n2988 VPWR.n2987 25.1912
R10829 VPWR.n2925 VPWR.n2924 25.1912
R10830 VPWR.n5854 VPWR.n5850 25.1912
R10831 VPWR.n6307 VPWR.n6304 24.8476
R10832 VPWR.n3239 VPWR.n3238 24.8476
R10833 VPWR.n5014 VPWR.n4980 24.8476
R10834 VPWR.n1247 VPWR.n1246 24.8476
R10835 VPWR.n4354 VPWR.n4353 24.8476
R10836 VPWR.n3621 VPWR.n1575 24.8476
R10837 VPWR.n2796 VPWR.n2795 24.8476
R10838 VPWR.n6154 VPWR.n5824 24.7608
R10839 VPWR.n7125 VPWR.n7124 24.7608
R10840 VPWR.n1154 VPWR.n1153 24.5271
R10841 VPWR.n752 VPWR.n751 24.5034
R10842 VPWR.n781 VPWR.n576 24.4711
R10843 VPWR.n6293 VPWR.n6292 24.4711
R10844 VPWR.n6127 VPWR.n6126 24.4711
R10845 VPWR.n7453 VPWR.n7440 24.4711
R10846 VPWR.n4813 VPWR.n4812 24.4711
R10847 VPWR.n3852 VPWR.n3851 24.4711
R10848 VPWR.n4365 VPWR.n435 24.4711
R10849 VPWR.n4085 VPWR.n1530 24.4711
R10850 VPWR.n1853 VPWR.n1846 24.4711
R10851 VPWR.n1682 VPWR.n1681 24.4711
R10852 VPWR.n5949 VPWR.n5924 24.4711
R10853 VPWR.n5938 VPWR.n5937 24.4711
R10854 VPWR.n657 VPWR.n644 24.4333
R10855 VPWR.n3871 VPWR.n3776 24.4327
R10856 VPWR.n6222 VPWR.n5746 24.0946
R10857 VPWR.n6299 VPWR.n6280 24.0946
R10858 VPWR.n6155 VPWR.n6154 24.0946
R10859 VPWR.n4471 VPWR.n4470 24.0946
R10860 VPWR.n3813 VPWR.n3780 24.0946
R10861 VPWR.n4347 VPWR.n1436 24.0946
R10862 VPWR.n5951 VPWR.n5922 24.0946
R10863 VPWR.n4498 VPWR.n395 24.0757
R10864 VPWR.n7081 VPWR.n7080 23.8912
R10865 VPWR.n3314 VPWR.n3301 23.7181
R10866 VPWR.n7273 VPWR.n7272 23.7181
R10867 VPWR.n639 VPWR.n575 23.7181
R10868 VPWR.n4486 VPWR.n4485 23.7181
R10869 VPWR.n2007 VPWR.n1641 23.7181
R10870 VPWR.n2124 VPWR.n1583 23.7181
R10871 VPWR.n6220 VPWR.n6219 23.7181
R10872 VPWR.n6219 VPWR.n5747 23.7181
R10873 VPWR.n5846 VPWR.n5830 23.7181
R10874 VPWR.n2436 VPWR.n2435 23.7181
R10875 VPWR.n3116 VPWR.n2419 23.7181
R10876 VPWR.n3116 VPWR.n2420 23.7181
R10877 VPWR.n6852 VPWR.n6800 23.7181
R10878 VPWR.n7276 VPWR.n290 23.7181
R10879 VPWR.n7069 VPWR.n4872 23.7181
R10880 VPWR.n5313 VPWR.n5233 23.7181
R10881 VPWR.n5314 VPWR.n5313 23.7181
R10882 VPWR.n5361 VPWR.n5347 23.7181
R10883 VPWR.n5365 VPWR.n5347 23.7181
R10884 VPWR.n957 VPWR.n573 23.7181
R10885 VPWR.n646 VPWR.n573 23.7181
R10886 VPWR.n479 VPWR.n478 23.7181
R10887 VPWR.n485 VPWR.n477 23.7181
R10888 VPWR.n505 VPWR.n475 23.7181
R10889 VPWR.n358 VPWR.n357 23.7181
R10890 VPWR.n4623 VPWR.n375 23.7181
R10891 VPWR.n1249 VPWR.n1226 23.7181
R10892 VPWR.n4085 VPWR.n4084 23.7181
R10893 VPWR.n4112 VPWR.n1521 23.7181
R10894 VPWR.n4197 VPWR.n1480 23.7181
R10895 VPWR.n4197 VPWR.n1479 23.7181
R10896 VPWR.n1848 VPWR.n1847 23.7181
R10897 VPWR.n3639 VPWR.n1570 23.7181
R10898 VPWR.n3437 VPWR.n2213 23.7181
R10899 VPWR.n2697 VPWR.n2696 23.7181
R10900 VPWR.n5850 VPWR.n5830 23.7181
R10901 VPWR.n506 VPWR.n505 23.6811
R10902 VPWR.n5379 VPWR.n5376 23.6784
R10903 VPWR.n363 VPWR.n362 23.3565
R10904 VPWR.n4383 VPWR.n431 23.0405
R10905 VPWR.n6817 VPWR.n6816 22.9652
R10906 VPWR.n7342 VPWR.n7341 22.9652
R10907 VPWR.n5366 VPWR.n5365 22.9652
R10908 VPWR.n490 VPWR.n489 22.9652
R10909 VPWR.n1485 VPWR.n1484 22.9652
R10910 VPWR.n2718 VPWR.n2690 22.9652
R10911 VPWR.n813 VPWR.n601 22.9323
R10912 VPWR.n6962 VPWR.n6961 22.9184
R10913 VPWR.n3851 VPWR.n3817 22.5887
R10914 VPWR.n4366 VPWR.n4365 22.5887
R10915 VPWR.n4767 VPWR.n4766 22.5559
R10916 VPWR.n6056 VPWR.n6055 22.2123
R10917 VPWR.n6110 VPWR.n6056 22.2123
R10918 VPWR.n2421 VPWR.n2419 22.2123
R10919 VPWR.n2592 VPWR.n2591 22.2123
R10920 VPWR.n7070 VPWR.n7069 22.2123
R10921 VPWR.n7120 VPWR.n4863 22.2123
R10922 VPWR.n482 VPWR.n478 22.2123
R10923 VPWR.n483 VPWR.n482 22.2123
R10924 VPWR.n358 VPWR.n336 22.2123
R10925 VPWR.n4636 VPWR.n4635 22.2123
R10926 VPWR.n4108 VPWR.n1522 22.2123
R10927 VPWR.n1482 VPWR.n1480 22.2123
R10928 VPWR.n4200 VPWR.n1479 22.2123
R10929 VPWR.n4201 VPWR.n4200 22.2123
R10930 VPWR.n1744 VPWR.n1742 22.2123
R10931 VPWR.n1748 VPWR.n1742 22.2123
R10932 VPWR.n2714 VPWR.n2713 22.2123
R10933 VPWR.n2714 VPWR.n2690 22.2123
R10934 VPWR.n3593 VPWR.n3591 21.7466
R10935 VPWR.n1034 VPWR.n1033 21.5933
R10936 VPWR.n2596 VPWR.n2595 21.4593
R10937 VPWR.n5434 VPWR.n5433 21.4593
R10938 VPWR.n7281 VPWR.n7280 21.4593
R10939 VPWR.n1753 VPWR.n1752 21.4593
R10940 VPWR.n1762 VPWR.n1761 21.0952
R10941 VPWR.n1425 VPWR.n438 21.0829
R10942 VPWR.n1740 VPWR.n1739 21.0829
R10943 VPWR.n744 VPWR.n743 20.7415
R10944 VPWR.n6293 VPWR.n6282 20.7064
R10945 VPWR.n6126 VPWR.n6051 20.7064
R10946 VPWR.n1853 VPWR.n1852 20.7064
R10947 VPWR.n5950 VPWR.n5949 20.7064
R10948 VPWR.n5938 VPWR.n5927 20.7064
R10949 VPWR.n2517 VPWR.n2516 20.3859
R10950 VPWR.n3142 VPWR.n3141 20.0749
R10951 VPWR.n5555 VPWR.n5548 20.0749
R10952 VPWR.n6291 VPWR.n6284 19.9534
R10953 VPWR.n6128 VPWR.n6049 19.9534
R10954 VPWR.n5022 VPWR.n26 19.9534
R10955 VPWR.n5433 VPWR.n5428 19.9534
R10956 VPWR.n7223 VPWR.n292 19.9534
R10957 VPWR.n3813 VPWR.n3812 19.9534
R10958 VPWR.n4218 VPWR.n4217 19.9534
R10959 VPWR.n3602 VPWR.n1577 19.9534
R10960 VPWR.n5945 VPWR.n5944 19.9534
R10961 VPWR.n5936 VPWR.n5929 19.9534
R10962 VPWR.n3606 VPWR.n3602 19.9057
R10963 VPWR.n6304 VPWR.n6303 19.577
R10964 VPWR.n6156 VPWR.n5822 19.577
R10965 VPWR.n3317 VPWR.n3300 19.577
R10966 VPWR.n57 VPWR.n52 19.577
R10967 VPWR.n7724 VPWR.n7723 19.577
R10968 VPWR.n177 VPWR.n172 19.577
R10969 VPWR.n951 VPWR.n580 19.577
R10970 VPWR.n5956 VPWR.n5955 19.577
R10971 VPWR.n947 VPWR.n578 19.5441
R10972 VPWR.n348 VPWR.n339 19.5347
R10973 VPWR.n5526 VPWR.n5525 19.2067
R10974 VPWR.n5272 VPWR.n5236 19.2067
R10975 VPWR.n3911 VPWR.n3910 19.2067
R10976 VPWR.n6477 VPWR.n5062 18.9594
R10977 VPWR.n5164 VPWR.n5144 18.9594
R10978 VPWR.n5101 VPWR.n5092 18.824
R10979 VPWR VPWR.n6306 18.7912
R10980 VPWR VPWR.n6109 18.7912
R10981 VPWR.n5038 VPWR.n5037 18.7912
R10982 VPWR.n3626 VPWR 18.7912
R10983 VPWR.n2702 VPWR 18.7912
R10984 VPWR.n2709 VPWR.n2691 18.7912
R10985 VPWR VPWR.n6228 18.4476
R10986 VPWR.n5822 VPWR 18.4476
R10987 VPWR VPWR.n7449 18.4476
R10988 VPWR VPWR.n4805 18.4476
R10989 VPWR.n888 VPWR.n887 18.4476
R10990 VPWR VPWR.n347 18.4476
R10991 VPWR.n5892 VPWR 18.4476
R10992 VPWR VPWR.n5956 18.4476
R10993 VPWR.n6287 VPWR.n6284 18.4147
R10994 VPWR.n6049 VPWR.n6048 18.4147
R10995 VPWR.n5930 VPWR.n5929 18.4147
R10996 VPWR.n7450 VPWR.n7441 18.0711
R10997 VPWR.n4806 VPWR.n4797 18.0711
R10998 VPWR.n662 VPWR.n643 18.0711
R10999 VPWR VPWR.n4186 18.0711
R11000 VPWR.n1528 VPWR.n1527 17.6946
R11001 VPWR.n6313 VPWR.n6312 17.612
R11002 VPWR.n6946 VPWR.n6945 17.612
R11003 VPWR.n2869 VPWR.n2868 17.612
R11004 VPWR.n2919 VPWR.n2918 17.612
R11005 VPWR.n5860 VPWR.n5859 17.612
R11006 VPWR.n6250 VPWR.n5739 17.612
R11007 VPWR.n2610 VPWR.n2609 17.612
R11008 VPWR.n2970 VPWR.n2969 17.612
R11009 VPWR.n5097 VPWR.n5096 17.3181
R11010 VPWR.n1140 VPWR.n1139 17.3181
R11011 VPWR.n1139 VPWR.n1138 17.3181
R11012 VPWR.n2428 VPWR.n2427 17.2853
R11013 VPWR.n2152 VPWR.n1580 17.2339
R11014 VPWR.n7216 VPWR 17.1239
R11015 VPWR.n5429 VPWR.n5428 16.9417
R11016 VPWR.n1230 VPWR.n1229 16.9417
R11017 VPWR.n1676 VPWR.n1675 16.9417
R11018 VPWR.n3648 VPWR.n3647 16.9417
R11019 VPWR.n1201 VPWR.n1090 16.8979
R11020 VPWR.n4526 VPWR.n391 16.6514
R11021 VPWR.n3654 VPWR.n3653 16.6212
R11022 VPWR.n5885 VPWR.n5884 16.6212
R11023 VPWR.n2007 VPWR.n2006 16.6183
R11024 VPWR.n1371 VPWR.n1370 16.5652
R11025 VPWR.n5249 VPWR.n5248 16.4496
R11026 VPWR.n3124 VPWR.n3123 16.3211
R11027 VPWR.n5185 VPWR.n5183 16.3211
R11028 VPWR.n4663 VPWR.n367 16.3211
R11029 VPWR.n4530 VPWR.n391 16.3211
R11030 VPWR.n2244 VPWR.n2217 16.2403
R11031 VPWR.n2126 VPWR.n2124 16.2176
R11032 VPWR.n6384 VPWR.n6383 16.139
R11033 VPWR.n6710 VPWR.n6709 16.139
R11034 VPWR.n1962 VPWR.n1961 16.139
R11035 VPWR.n2127 VPWR.n2126 16.139
R11036 VPWR.n2317 VPWR.n2316 15.995
R11037 VPWR.n6265 VPWR.n6264 15.8683
R11038 VPWR.n3283 VPWR.n2385 15.8683
R11039 VPWR.n2562 VPWR.n2561 15.8683
R11040 VPWR.n7582 VPWR.n7581 15.8683
R11041 VPWR.n3889 VPWR.n3888 15.8683
R11042 VPWR.n1331 VPWR.n1330 15.8683
R11043 VPWR.n3437 VPWR.n2214 15.8683
R11044 VPWR.n2928 VPWR.n2806 15.8683
R11045 VPWR.n2945 VPWR.n2944 15.8683
R11046 VPWR.n336 VPWR 15.8123
R11047 VPWR.n7675 VPWR.n7674 15.7465
R11048 VPWR.n4077 VPWR.n4076 15.7465
R11049 VPWR.n1871 VPWR.n1868 15.7465
R11050 VPWR.n756 VPWR.n752 15.7306
R11051 VPWR.n7276 VPWR.n291 15.4358
R11052 VPWR.n3290 VPWR.n3289 15.3068
R11053 VPWR.n3314 VPWR.n3313 15.1382
R11054 VPWR.n5501 VPWR.n5500 15.0923
R11055 VPWR.n6863 VPWR.n6796 15.0265
R11056 VPWR.n909 VPWR.n908 15.0265
R11057 VPWR.n3824 VPWR.n3823 14.9948
R11058 VPWR.n6652 VPWR.n6651 14.9474
R11059 VPWR.n2120 VPWR.n1585 14.6829
R11060 VPWR.n1429 VPWR.n438 14.65
R11061 VPWR.n4205 VPWR.n4204 14.65
R11062 VPWR.n3620 VPWR.n3619 14.65
R11063 VPWR.n5899 VPWR.n5898 14.65
R11064 VPWR.n3111 VPWR.n2421 14.6331
R11065 VPWR.n3838 VPWR.n3837 14.6291
R11066 VPWR.n2293 VPWR.n2292 14.5851
R11067 VPWR.n3872 VPWR.n3871 14.5729
R11068 VPWR.n5105 VPWR.n5092 14.3064
R11069 VPWR.n7218 VPWR.n7216 14.3064
R11070 VPWR.n4353 VPWR.n1434 14.3064
R11071 VPWR.n6139 VPWR.n6046 14.2735
R11072 VPWR.n6136 VPWR.n6046 14.2735
R11073 VPWR.n2583 VPWR.n2582 14.2735
R11074 VPWR.n7330 VPWR.n7329 14.2735
R11075 VPWR.n5354 VPWR.n5353 14.2735
R11076 VPWR.n897 VPWR.n577 14.2735
R11077 VPWR.n671 VPWR.n670 14.2735
R11078 VPWR.n1025 VPWR.n1020 14.2735
R11079 VPWR.n3999 VPWR.n3998 14.2735
R11080 VPWR.n4067 VPWR.n4066 14.2735
R11081 VPWR.n1953 VPWR.n1647 14.2735
R11082 VPWR.n1596 VPWR.n1583 14.2735
R11083 VPWR.n6042 VPWR.n5831 14.2735
R11084 VPWR.n431 VPWR.n430 14.2634
R11085 VPWR.n3321 VPWR.n3300 13.9299
R11086 VPWR.n6822 VPWR.n6821 13.9299
R11087 VPWR.n762 VPWR.n761 13.902
R11088 VPWR.n3826 VPWR.n3824 13.8976
R11089 VPWR.n6042 VPWR.n6041 13.8432
R11090 VPWR.n3140 VPWR.n3139 13.6753
R11091 VPWR.n5547 VPWR.n5466 13.6753
R11092 VPWR.n50 VPWR.n49 13.5534
R11093 VPWR.n890 VPWR.n583 13.5534
R11094 VPWR.n3598 VPWR.n1577 13.5534
R11095 VPWR.n2983 VPWR.n2982 13.5534
R11096 VPWR.n182 VPWR.n181 13.5206
R11097 VPWR.n4634 VPWR.n4633 13.5206
R11098 VPWR.n2245 VPWR.n2244 13.4744
R11099 VPWR VPWR.n3306 13.41
R11100 VPWR.n6264 VPWR.n5733 13.177
R11101 VPWR.n54 VPWR.n53 13.177
R11102 VPWR.n174 VPWR.n173 13.177
R11103 VPWR.n7444 VPWR.n7443 13.177
R11104 VPWR.n4800 VPWR.n4799 13.177
R11105 VPWR.n342 VPWR.n341 13.177
R11106 VPWR.n1436 VPWR.n1435 13.177
R11107 VPWR.n4642 VPWR.n4641 13.0915
R11108 VPWR.n6480 VPWR.n5062 13.0319
R11109 VPWR.n5145 VPWR.n5144 13.0319
R11110 VPWR.n3283 VPWR.n2384 12.8005
R11111 VPWR.n2591 VPWR.n2590 12.8005
R11112 VPWR.n6383 VPWR.n6380 12.8005
R11113 VPWR.n5096 VPWR.n5095 12.8005
R11114 VPWR.n7582 VPWR.n160 12.8005
R11115 VPWR.n5477 VPWR.n5467 12.8005
R11116 VPWR.n6852 VPWR.n6799 12.8005
R11117 VPWR.n7071 VPWR.n4869 12.8005
R11118 VPWR.n5238 VPWR.n5233 12.8005
R11119 VPWR.n583 VPWR.n577 12.8005
R11120 VPWR.n489 VPWR.n477 12.8005
R11121 VPWR.n1021 VPWR.n1020 12.8005
R11122 VPWR.n3868 VPWR.n3778 12.8005
R11123 VPWR.n1961 VPWR.n1647 12.8005
R11124 VPWR.n1579 VPWR.n1578 12.8005
R11125 VPWR.n3591 VPWR.n1578 12.8005
R11126 VPWR.n2696 VPWR.n2693 12.8005
R11127 VPWR.n36 VPWR 12.424
R11128 VPWR.n7443 VPWR.n7442 12.424
R11129 VPWR.n4799 VPWR.n4798 12.424
R11130 VPWR.n341 VPWR.n340 12.424
R11131 VPWR.n3621 VPWR.n3620 12.424
R11132 VPWR.n51 VPWR.n50 12.0476
R11133 VPWR.n5500 VPWR.n5467 12.0476
R11134 VPWR.n7341 VPWR.n7327 12.0476
R11135 VPWR.n2719 VPWR.n2718 12.0147
R11136 VPWR.n3265 VPWR.n3264 11.9246
R11137 VPWR.n3240 VPWR.n3239 11.7271
R11138 VPWR.n52 VPWR.n51 11.6711
R11139 VPWR.n181 VPWR.n172 11.6711
R11140 VPWR.n1373 VPWR.n1372 11.6382
R11141 VPWR.n2561 VPWR.n2507 11.5544
R11142 VPWR.n3230 VPWR.n2383 11.4546
R11143 VPWR.n3119 VPWR.n2418 11.4366
R11144 VPWR.n7071 VPWR.n7070 11.2946
R11145 VPWR.n7119 VPWR.n4864 11.2946
R11146 VPWR.n1522 VPWR.n1521 11.2946
R11147 VPWR.n2590 VPWR.n2589 11.2618
R11148 VPWR.n7337 VPWR.n7327 11.2618
R11149 VPWR.n2520 VPWR.n2519 10.9181
R11150 VPWR.n2604 VPWR 10.9181
R11151 VPWR.n1483 VPWR.n1482 10.9181
R11152 VPWR.n2604 VPWR.n2603 10.8853
R11153 VPWR.n5051 VPWR.n4981 10.8853
R11154 VPWR.n6823 VPWR.n6822 10.8853
R11155 VPWR.n7272 VPWR.n7230 10.8853
R11156 VPWR.n7704 VPWR.n7703 10.8646
R11157 VPWR.n2898 VPWR.n2897 10.5506
R11158 VPWR.n7233 VPWR.n7231 10.5417
R11159 VPWR.n951 VPWR.n578 10.5417
R11160 VPWR.n2897 VPWR.n2895 10.3589
R11161 VPWR.n6477 VPWR.n6476 10.3343
R11162 VPWR.n5466 VPWR.n5465 10.3343
R11163 VPWR.n3289 VPWR.n2383 9.90679
R11164 VPWR.n68 VPWR.n67 9.78874
R11165 VPWR.n193 VPWR.n192 9.78874
R11166 VPWR.n7120 VPWR.n7119 9.78874
R11167 VPWR.n1947 VPWR.n1946 9.78874
R11168 VPWR.n1688 VPWR.n1687 9.78874
R11169 VPWR.n6246 VPWR.n5739 9.73273
R11170 VPWR.n6246 VPWR.n6245 9.73273
R11171 VPWR.n6245 VPWR.n6244 9.73273
R11172 VPWR.n6241 VPWR.n6240 9.73273
R11173 VPWR.n6240 VPWR.n6239 9.73273
R11174 VPWR.n6239 VPWR.n5743 9.73273
R11175 VPWR.n6235 VPWR.n5743 9.73273
R11176 VPWR.n6235 VPWR.n6234 9.73273
R11177 VPWR.n6234 VPWR.n6233 9.73273
R11178 VPWR.n6233 VPWR.n5745 9.73273
R11179 VPWR.n2452 VPWR.n2451 9.73273
R11180 VPWR.n2538 VPWR.n2537 9.73273
R11181 VPWR.n2537 VPWR.n2536 9.73273
R11182 VPWR.n2536 VPWR.n2516 9.73273
R11183 VPWR.n2554 VPWR.n2508 9.73273
R11184 VPWR.n6390 VPWR.n6379 9.73273
R11185 VPWR.n6396 VPWR.n6395 9.73273
R11186 VPWR.n6476 VPWR.n5064 9.73273
R11187 VPWR.n7568 VPWR.n7567 9.73273
R11188 VPWR.n7585 VPWR.n159 9.73273
R11189 VPWR.n5171 VPWR.n5170 9.73273
R11190 VPWR.n6925 VPWR.n6924 9.73273
R11191 VPWR.n6924 VPWR.n4926 9.73273
R11192 VPWR.n5560 VPWR.n5465 9.73273
R11193 VPWR.n5445 VPWR.n5444 9.73273
R11194 VPWR.n5458 VPWR.n5426 9.73273
R11195 VPWR.n7094 VPWR.n4866 9.73273
R11196 VPWR.n7098 VPWR.n4866 9.73273
R11197 VPWR.n5255 VPWR.n5254 9.73273
R11198 VPWR.n5276 VPWR.n5236 9.73273
R11199 VPWR.n5277 VPWR.n5276 9.73273
R11200 VPWR.n5310 VPWR.n5235 9.73273
R11201 VPWR.n5310 VPWR.n5309 9.73273
R11202 VPWR.n4667 VPWR.n367 9.73273
R11203 VPWR.n4668 VPWR.n4667 9.73273
R11204 VPWR.n4648 VPWR.n371 9.73273
R11205 VPWR.n4654 VPWR.n370 9.73273
R11206 VPWR.n4531 VPWR.n4530 9.73273
R11207 VPWR.n4524 VPWR.n4523 9.73273
R11208 VPWR.n1190 VPWR.n1189 9.73273
R11209 VPWR.n1189 VPWR.n1092 9.73273
R11210 VPWR.n1185 VPWR.n1184 9.73273
R11211 VPWR.n1044 VPWR.n1043 9.73273
R11212 VPWR.n3910 VPWR.n3884 9.73273
R11213 VPWR.n3906 VPWR.n3884 9.73273
R11214 VPWR.n3906 VPWR.n3905 9.73273
R11215 VPWR.n3902 VPWR.n3901 9.73273
R11216 VPWR.n3901 VPWR.n3886 9.73273
R11217 VPWR.n3897 VPWR.n3886 9.73273
R11218 VPWR.n1366 VPWR.n1365 9.73273
R11219 VPWR.n1324 VPWR.n443 9.73273
R11220 VPWR.n1325 VPWR.n1324 9.73273
R11221 VPWR.n2142 VPWR.n1581 9.73273
R11222 VPWR.n3663 VPWR.n3644 9.73273
R11223 VPWR.n3659 VPWR.n3658 9.73273
R11224 VPWR.n3658 VPWR.n3645 9.73273
R11225 VPWR.n2882 VPWR.n2807 9.73273
R11226 VPWR.n2883 VPWR.n2882 9.73273
R11227 VPWR.n2902 VPWR.n2901 9.73273
R11228 VPWR.n958 VPWR.n957 9.67237
R11229 VPWR.n910 VPWR.n909 9.41227
R11230 VPWR.n675 VPWR.n639 9.41227
R11231 VPWR.n1700 VPWR.n1673 9.41227
R11232 VPWR.n234 VPWR.n233 9.30284
R11233 VPWR.n5668 VPWR.n5667 9.3005
R11234 VPWR.n5140 VPWR.n5139 9.3005
R11235 VPWR.n5666 VPWR.n5665 9.3005
R11236 VPWR.n206 VPWR.n205 9.3005
R11237 VPWR.n216 VPWR.n215 9.3005
R11238 VPWR.n208 VPWR.n207 9.3005
R11239 VPWR.n6756 VPWR.n6755 9.3005
R11240 VPWR.n6754 VPWR.n6753 9.3005
R11241 VPWR.n5592 VPWR.n5591 9.3005
R11242 VPWR.n5619 VPWR.n5618 9.3005
R11243 VPWR.n5601 VPWR.n5600 9.3005
R11244 VPWR.n5590 VPWR.n5589 9.3005
R11245 VPWR.n7421 VPWR.n7420 9.3005
R11246 VPWR.n7477 VPWR.n7476 9.3005
R11247 VPWR.n7411 VPWR.n7410 9.3005
R11248 VPWR.n7413 VPWR.n7412 9.3005
R11249 VPWR.n5334 VPWR.n5333 9.3005
R11250 VPWR.n5342 VPWR.n5341 9.3005
R11251 VPWR.n5332 VPWR.n5331 9.3005
R11252 VPWR.n7306 VPWR.n7305 9.3005
R11253 VPWR.n7367 VPWR.n7366 9.3005
R11254 VPWR.n7369 VPWR.n7368 9.3005
R11255 VPWR.n7309 VPWR.n7308 9.3005
R11256 VPWR.n4836 VPWR.n4835 9.3005
R11257 VPWR.n4838 VPWR.n4837 9.3005
R11258 VPWR.n4770 VPWR.n4769 9.3005
R11259 VPWR.n4772 VPWR.n4771 9.3005
R11260 VPWR.n520 VPWR.n519 9.3005
R11261 VPWR.n561 VPWR.n560 9.3005
R11262 VPWR.n1128 VPWR.n1127 9.3005
R11263 VPWR.n1056 VPWR.n1055 9.3005
R11264 VPWR.n1082 VPWR.n1081 9.3005
R11265 VPWR.n1084 VPWR.n1083 9.3005
R11266 VPWR.n4536 VPWR.n4535 9.3005
R11267 VPWR.n4704 VPWR.n4703 9.3005
R11268 VPWR.n4722 VPWR.n4721 9.3005
R11269 VPWR.n4720 VPWR.n4719 9.3005
R11270 VPWR.n4694 VPWR.n4693 9.3005
R11271 VPWR.n4696 VPWR.n4695 9.3005
R11272 VPWR.n4611 VPWR.n4610 9.3005
R11273 VPWR.n4608 VPWR.n4607 9.3005
R11274 VPWR.n4538 VPWR.n4537 9.3005
R11275 VPWR.n402 VPWR.n401 9.3005
R11276 VPWR.n1100 VPWR.n1099 9.3005
R11277 VPWR.n1125 VPWR.n1124 9.3005
R11278 VPWR.n1074 VPWR.n1073 9.3005
R11279 VPWR.n1058 VPWR.n1057 9.3005
R11280 VPWR.n1303 VPWR.n1302 9.3005
R11281 VPWR.n1439 VPWR.n1438 9.3005
R11282 VPWR.n3941 VPWR.n3940 9.3005
R11283 VPWR.n1441 VPWR.n1440 9.3005
R11284 VPWR.n1391 VPWR.n1390 9.3005
R11285 VPWR.n1393 VPWR.n1392 9.3005
R11286 VPWR.n1305 VPWR.n1304 9.3005
R11287 VPWR.n1258 VPWR.n1257 9.3005
R11288 VPWR.n2017 VPWR.n2016 9.3005
R11289 VPWR.n1939 VPWR.n1938 9.3005
R11290 VPWR.n4160 VPWR.n4159 9.3005
R11291 VPWR.n4121 VPWR.n4120 9.3005
R11292 VPWR.n4124 VPWR.n4123 9.3005
R11293 VPWR.n4162 VPWR.n4161 9.3005
R11294 VPWR.n2020 VPWR.n2019 9.3005
R11295 VPWR.n1941 VPWR.n1940 9.3005
R11296 VPWR.n1931 VPWR.n1930 9.3005
R11297 VPWR.n1928 VPWR.n1927 9.3005
R11298 VPWR.n3583 VPWR.n3582 9.3005
R11299 VPWR.n2114 VPWR.n2113 9.3005
R11300 VPWR.n3560 VPWR.n3559 9.3005
R11301 VPWR.n3580 VPWR.n3579 9.3005
R11302 VPWR.n3558 VPWR.n3557 9.3005
R11303 VPWR.n2087 VPWR.n2086 9.3005
R11304 VPWR.n2089 VPWR.n2088 9.3005
R11305 VPWR.n2111 VPWR.n2110 9.3005
R11306 VPWR.n2821 VPWR.n2820 9.3005
R11307 VPWR.n2788 VPWR.n2787 9.3005
R11308 VPWR.n3452 VPWR.n3451 9.3005
R11309 VPWR.n2332 VPWR.n2331 9.3005
R11310 VPWR.n3422 VPWR.n3421 9.3005
R11311 VPWR.n3420 VPWR.n3419 9.3005
R11312 VPWR.n3455 VPWR.n3454 9.3005
R11313 VPWR.n3475 VPWR.n3474 9.3005
R11314 VPWR.n3477 VPWR.n3476 9.3005
R11315 VPWR.n2824 VPWR.n2823 9.3005
R11316 VPWR.n2790 VPWR.n2789 9.3005
R11317 VPWR.n2764 VPWR.n2763 9.3005
R11318 VPWR.n6530 VPWR.n6529 9.3005
R11319 VPWR.n6412 VPWR.n6411 9.3005
R11320 VPWR.n6429 VPWR.n6428 9.3005
R11321 VPWR.n6410 VPWR.n6409 9.3005
R11322 VPWR.n6533 VPWR.n6532 9.3005
R11323 VPWR.n6554 VPWR.n6553 9.3005
R11324 VPWR.n6556 VPWR.n6555 9.3005
R11325 VPWR.n7725 VPWR.n7724 9.3005
R11326 VPWR.n7728 VPWR.n7727 9.3005
R11327 VPWR.n2618 VPWR.n2617 9.3005
R11328 VPWR.n2645 VPWR.n2644 9.3005
R11329 VPWR.n3110 VPWR.n3109 9.3005
R11330 VPWR.n3216 VPWR.n3215 9.3005
R11331 VPWR.n3350 VPWR.n3349 9.3005
R11332 VPWR.n3358 VPWR.n3357 9.3005
R11333 VPWR.n3332 VPWR.n3331 9.3005
R11334 VPWR.n3360 VPWR.n3359 9.3005
R11335 VPWR.n3213 VPWR.n3212 9.3005
R11336 VPWR.n3107 VPWR.n3106 9.3005
R11337 VPWR.n3085 VPWR.n3084 9.3005
R11338 VPWR.n3087 VPWR.n3086 9.3005
R11339 VPWR.n2634 VPWR.n2633 9.3005
R11340 VPWR.n2643 VPWR.n2642 9.3005
R11341 VPWR.n2616 VPWR.n2615 9.3005
R11342 VPWR.n6212 VPWR.n6211 9.3005
R11343 VPWR.n6321 VPWR.n6320 9.3005
R11344 VPWR.n6346 VPWR.n6345 9.3005
R11345 VPWR.n6319 VPWR.n6318 9.3005
R11346 VPWR.n6337 VPWR.n6336 9.3005
R11347 VPWR.n6348 VPWR.n6347 9.3005
R11348 VPWR.n6209 VPWR.n6208 9.3005
R11349 VPWR.n6189 VPWR.n6188 9.3005
R11350 VPWR.n6187 VPWR.n6186 9.3005
R11351 VPWR.n5963 VPWR.n5962 9.3005
R11352 VPWR.n5971 VPWR.n5970 9.3005
R11353 VPWR.n5961 VPWR.n5960 9.3005
R11354 VPWR.n5989 VPWR.n5988 9.3005
R11355 VPWR.n3264 VPWR.n3228 9.20592
R11356 VPWR.n601 VPWR 9.03579
R11357 VPWR.n4635 VPWR.n4634 9.03579
R11358 VPWR.n1372 VPWR.n1371 9.03579
R11359 VPWR.n2120 VPWR.n1586 9.03579
R11360 VPWR.n2944 VPWR.n2943 9.03579
R11361 VPWR.n7405 VPWR.n7404 9.02415
R11362 VPWR.n5325 VPWR.n5324 9.02415
R11363 VPWR.n4764 VPWR.n4763 9.02415
R11364 VPWR.n971 VPWR.n970 9.02415
R11365 VPWR.n4687 VPWR.n4686 9.02415
R11366 VPWR.n1205 VPWR.n1204 9.02415
R11367 VPWR.n4059 VPWR.n4058 9.02415
R11368 VPWR.n2991 VPWR.n2990 9.02415
R11369 VPWR.n6655 VPWR.n6654 9.00388
R11370 VPWR.n5664 VPWR.n5663 9.0005
R11371 VPWR.n5671 VPWR.n5670 9.0005
R11372 VPWR.n5136 VPWR.n5135 9.0005
R11373 VPWR.n6764 VPWR.n6763 9.0005
R11374 VPWR.n6758 VPWR.n6757 9.0005
R11375 VPWR.n6752 VPWR.n6751 9.0005
R11376 VPWR.n162 VPWR.n161 9.0005
R11377 VPWR.n230 VPWR.n229 9.0005
R11378 VPWR.n221 VPWR.n220 9.0005
R11379 VPWR.n210 VPWR.n209 9.0005
R11380 VPWR.n7616 VPWR.n7615 9.0005
R11381 VPWR.n6611 VPWR.n6610 9.0005
R11382 VPWR.n5588 VPWR.n5587 9.0005
R11383 VPWR.n5595 VPWR.n5594 9.0005
R11384 VPWR.n5615 VPWR.n5614 9.0005
R11385 VPWR.n5606 VPWR.n5605 9.0005
R11386 VPWR.n6911 VPWR.n6910 9.0005
R11387 VPWR.n7409 VPWR.n7408 9.0005
R11388 VPWR.n7415 VPWR.n7414 9.0005
R11389 VPWR.n7426 VPWR.n7425 9.0005
R11390 VPWR.n7482 VPWR.n7481 9.0005
R11391 VPWR.n5330 VPWR.n5329 9.0005
R11392 VPWR.n5336 VPWR.n5335 9.0005
R11393 VPWR.n5399 VPWR.n5398 9.0005
R11394 VPWR.n5402 VPWR.n5401 9.0005
R11395 VPWR.n7181 VPWR.n7180 9.0005
R11396 VPWR.n7159 VPWR.n7158 9.0005
R11397 VPWR.n7311 VPWR.n7310 9.0005
R11398 VPWR.n7372 VPWR.n7371 9.0005
R11399 VPWR.n4768 VPWR.n4767 9.0005
R11400 VPWR.n4774 VPWR.n4773 9.0005
R11401 VPWR.n4841 VPWR.n4840 9.0005
R11402 VPWR.n525 VPWR.n524 9.0005
R11403 VPWR.n557 VPWR.n556 9.0005
R11404 VPWR.n1086 VPWR.n1085 9.0005
R11405 VPWR.n1070 VPWR.n1069 9.0005
R11406 VPWR.n1080 VPWR.n1079 9.0005
R11407 VPWR.n4540 VPWR.n4539 9.0005
R11408 VPWR.n4534 VPWR.n4533 9.0005
R11409 VPWR.n4692 VPWR.n4691 9.0005
R11410 VPWR.n4698 VPWR.n4697 9.0005
R11411 VPWR.n4709 VPWR.n4708 9.0005
R11412 VPWR.n4717 VPWR.n4716 9.0005
R11413 VPWR.n4606 VPWR.n4605 9.0005
R11414 VPWR.n1061 VPWR.n1060 9.0005
R11415 VPWR.n1123 VPWR.n1122 9.0005
R11416 VPWR.n1102 VPWR.n1101 9.0005
R11417 VPWR.n4459 VPWR.n4458 9.0005
R11418 VPWR.n1307 VPWR.n1306 9.0005
R11419 VPWR.n1263 VPWR.n1262 9.0005
R11420 VPWR.n1301 VPWR.n1300 9.0005
R11421 VPWR.n1443 VPWR.n1442 9.0005
R11422 VPWR.n3784 VPWR.n3783 9.0005
R11423 VPWR.n3937 VPWR.n3936 9.0005
R11424 VPWR.n1272 VPWR.n1271 9.0005
R11425 VPWR.n1395 VPWR.n1394 9.0005
R11426 VPWR.n1389 VPWR.n1388 9.0005
R11427 VPWR.n1943 VPWR.n1942 9.0005
R11428 VPWR.n4164 VPWR.n4163 9.0005
R11429 VPWR.n4158 VPWR.n4157 9.0005
R11430 VPWR VPWR.n1518 9.0005
R11431 VPWR.n4126 VPWR.n4125 9.0005
R11432 VPWR.n1937 VPWR.n1936 9.0005
R11433 VPWR.n1892 VPWR.n1891 9.0005
R11434 VPWR.n1926 VPWR.n1925 9.0005
R11435 VPWR.n2022 VPWR.n2021 9.0005
R11436 VPWR.n3578 VPWR.n3577 9.0005
R11437 VPWR.n3689 VPWR.n3688 9.0005
R11438 VPWR.n3556 VPWR.n3555 9.0005
R11439 VPWR.n3562 VPWR.n3561 9.0005
R11440 VPWR.n2109 VPWR.n2107 9.0005
R11441 VPWR.n2109 VPWR.n2108 9.0005
R11442 VPWR.n2091 VPWR.n2090 9.0005
R11443 VPWR.n2085 VPWR.n2084 9.0005
R11444 VPWR.n2792 VPWR.n2791 9.0005
R11445 VPWR.n3424 VPWR.n3423 9.0005
R11446 VPWR.n3418 VPWR.n3417 9.0005
R11447 VPWR.n2337 VPWR.n2336 9.0005
R11448 VPWR.n3457 VPWR.n3456 9.0005
R11449 VPWR.n3479 VPWR.n3478 9.0005
R11450 VPWR.n3473 VPWR.n3472 9.0005
R11451 VPWR.n2786 VPWR.n2785 9.0005
R11452 VPWR.n2751 VPWR.n2750 9.0005
R11453 VPWR.n2760 VPWR.n2759 9.0005
R11454 VPWR.n2826 VPWR.n2825 9.0005
R11455 VPWR.n6535 VPWR.n6534 9.0005
R11456 VPWR.n6552 VPWR.n6551 9.0005
R11457 VPWR.n6558 VPWR.n6557 9.0005
R11458 VPWR.n7730 VPWR.n7729 9.0005
R11459 VPWR VPWR.n7737 9.0005
R11460 VPWR.n87 VPWR.n86 9.0005
R11461 VPWR.n5066 VPWR.n5065 9.0005
R11462 VPWR.n6415 VPWR.n6414 9.0005
R11463 VPWR.n6434 VPWR.n6433 9.0005
R11464 VPWR.n3105 VPWR.n3104 9.0005
R11465 VPWR.n3089 VPWR.n3088 9.0005
R11466 VPWR.n3083 VPWR.n3082 9.0005
R11467 VPWR.n3211 VPWR.n3210 9.0005
R11468 VPWR.n3192 VPWR.n3191 9.0005
R11469 VPWR.n2647 VPWR.n2646 9.0005
R11470 VPWR.n2641 VPWR.n2640 9.0005
R11471 VPWR.n2630 VPWR.n2629 9.0005
R11472 VPWR.n2621 VPWR.n2620 9.0005
R11473 VPWR.n3362 VPWR.n3361 9.0005
R11474 VPWR.n3356 VPWR.n3355 9.0005
R11475 VPWR.n3346 VPWR.n3345 9.0005
R11476 VPWR.n3337 VPWR.n3336 9.0005
R11477 VPWR.n5906 VPWR.n5905 9.0005
R11478 VPWR.n6207 VPWR.n6206 9.0005
R11479 VPWR.n6350 VPWR.n6349 9.0005
R11480 VPWR.n6344 VPWR.n6343 9.0005
R11481 VPWR.n6324 VPWR.n6323 9.0005
R11482 VPWR.n6333 VPWR.n6332 9.0005
R11483 VPWR.n6191 VPWR.n6190 9.0005
R11484 VPWR.n6185 VPWR.n6184 9.0005
R11485 VPWR.n5976 VPWR.n5975 9.0005
R11486 VPWR.n5965 VPWR.n5964 9.0005
R11487 VPWR.n5985 VPWR.n5984 9.0005
R11488 VPWR.n6706 VPWR.n4941 8.99224
R11489 VPWR.n5189 VPWR.n5143 8.93934
R11490 VPWR.n3586 VPWR.n1579 8.93934
R11491 VPWR.n3593 VPWR.n3592 8.72346
R11492 VPWR.n3111 VPWR.n3110 8.67488
R11493 VPWR.n1527 VPWR.n1526 8.65932
R11494 VPWR.n4005 VPWR.n3996 8.62646
R11495 VPWR.n1603 VPWR.n1593 8.62646
R11496 VPWR VPWR.n5164 8.53595
R11497 VPWR.n6686 VPWR.n4941 8.49384
R11498 VPWR.n6524 VPWR.n6523 8.49383
R11499 VPWR.n5459 VPWR.n5458 8.49383
R11500 VPWR.n2538 VPWR.n2514 8.44958
R11501 VPWR.n3244 VPWR.n3243 8.44958
R11502 VPWR.n6472 VPWR.n5064 8.44958
R11503 VPWR.n6523 VPWR.n5060 8.44958
R11504 VPWR.n4997 VPWR.n4995 8.44958
R11505 VPWR.n6706 VPWR.n4940 8.44958
R11506 VPWR.n5190 VPWR.n5189 8.44958
R11507 VPWR.n5561 VPWR.n5560 8.44958
R11508 VPWR.n1360 VPWR.n1359 8.44958
R11509 VPWR.n6400 VPWR.n6378 8.35119
R11510 VPWR VPWR.n2554 7.93438
R11511 VPWR.n5254 VPWR 7.93438
R11512 VPWR.n7449 VPWR.n7442 7.90638
R11513 VPWR.n4805 VPWR.n4798 7.90638
R11514 VPWR.n347 VPWR.n340 7.90638
R11515 VPWR.n3147 VPWR.n3146 7.87742
R11516 VPWR.n5554 VPWR.n5551 7.87742
R11517 VPWR.n2153 VPWR 7.8286
R11518 VPWR.n3322 VPWR.n3321 7.76772
R11519 VPWR.n2451 VPWR.n2425 7.75995
R11520 VPWR.n7586 VPWR.n7585 7.75995
R11521 VPWR.n7099 VPWR.n7098 7.75995
R11522 VPWR.n5309 VPWR.n5286 7.75995
R11523 VPWR.n4655 VPWR.n4654 7.75995
R11524 VPWR.n4523 VPWR.n394 7.75995
R11525 VPWR.n3917 VPWR.n3916 7.75995
R11526 VPWR.n2146 VPWR.n2142 7.75995
R11527 VPWR.n3664 VPWR.n3663 7.75995
R11528 VPWR.n2235 VPWR.n2234 7.75995
R11529 VPWR.n494 VPWR.n493 7.71815
R11530 VPWR.n3286 VPWR.n2383 7.60924
R11531 VPWR.n3272 VPWR.n2384 7.56696
R11532 VPWR.n3868 VPWR.n3776 7.52685
R11533 VPWR.n7459 VPWR.n7458 7.49348
R11534 VPWR.n3139 VPWR.n2414 7.26653
R11535 VPWR.n6499 VPWR.n6498 7.21067
R11536 VPWR.n4991 VPWR.n4989 7.21067
R11537 VPWR.n4095 VPWR.n1528 7.15344
R11538 VPWR.n6148 VPWR.n6147 7.11866
R11539 VPWR.n3145 VPWR.n3144 7.11866
R11540 VPWR.n5550 VPWR.n5549 7.11866
R11541 VPWR.n7131 VPWR.n7130 7.11866
R11542 VPWR.n6033 VPWR.n6032 7.11866
R11543 VPWR.n7115 VPWR.n4864 7.07809
R11544 VPWR.n3778 VPWR.n3777 7.05764
R11545 VPWR.n6687 VPWR.n6686 6.9375
R11546 VPWR.n3231 VPWR.n3230 6.77697
R11547 VPWR VPWR.n816 6.77697
R11548 VPWR.n3135 VPWR.n2414 6.66496
R11549 VPWR.n5006 VPWR.n5005 6.66496
R11550 VPWR.n1047 VPWR.n1046 6.66488
R11551 VPWR.n6529 VPWR.n6528 6.59529
R11552 VPWR.n6286 VPWR.n6285 6.58925
R11553 VPWR.n5932 VPWR.n5931 6.58194
R11554 VPWR.n6229 VPWR 6.4005
R11555 VPWR.n6257 VPWR 6.4005
R11556 VPWR.n6307 VPWR 6.4005
R11557 VPWR.n6160 VPWR 6.4005
R11558 VPWR.n6110 VPWR 6.4005
R11559 VPWR.n2529 VPWR 6.4005
R11560 VPWR.n3238 VPWR 6.4005
R11561 VPWR.n2592 VPWR 6.4005
R11562 VPWR.n7698 VPWR 6.4005
R11563 VPWR.n7450 VPWR 6.4005
R11564 VPWR.n4806 VPWR 6.4005
R11565 VPWR VPWR.n661 6.4005
R11566 VPWR.n348 VPWR 6.4005
R11567 VPWR.n362 VPWR 6.4005
R11568 VPWR.n4187 VPWR 6.4005
R11569 VPWR VPWR.n1857 6.4005
R11570 VPWR VPWR.n3625 6.4005
R11571 VPWR VPWR.n2701 6.4005
R11572 VPWR VPWR.n5891 6.4005
R11573 VPWR.n5957 VPWR 6.4005
R11574 VPWR.n762 VPWR.n602 6.21764
R11575 VPWR.n2432 VPWR.n2431 6.158
R11576 VPWR.n6401 VPWR.n6400 6.158
R11577 VPWR.n5109 VPWR.n5108 6.158
R11578 VPWR.n7698 VPWR.n36 6.02403
R11579 VPWR.n7533 VPWR.n7532 5.97806
R11580 VPWR.n1179 VPWR.n1178 5.97806
R11581 VPWR.n3823 VPWR.n3822 5.85193
R11582 VPWR.n2418 VPWR.n2417 5.76367
R11583 VPWR.n2417 VPWR.n2416 5.75665
R11584 VPWR.n5184 VPWR.n5143 5.75665
R11585 VPWR.n2432 VPWR.n2430 5.70476
R11586 VPWR.n5108 VPWR.n5091 5.70476
R11587 VPWR.n2550 VPWR.n2549 5.66204
R11588 VPWR.n2549 VPWR.n2548 5.66204
R11589 VPWR.n2548 VPWR.n2511 5.66204
R11590 VPWR.n2544 VPWR.n2543 5.66204
R11591 VPWR.n2543 VPWR.n2542 5.66204
R11592 VPWR.n2542 VPWR.n2514 5.66204
R11593 VPWR.n3228 VPWR.n3227 5.66204
R11594 VPWR.n6483 VPWR.n6482 5.66204
R11595 VPWR.n6498 VPWR.n6497 5.66204
R11596 VPWR.n6505 VPWR.n5061 5.66204
R11597 VPWR.n5060 VPWR.n5059 5.66204
R11598 VPWR.n6528 VPWR.n4979 5.66204
R11599 VPWR.n4991 VPWR.n4990 5.66204
R11600 VPWR.n4940 VPWR.n4939 5.66204
R11601 VPWR.n1344 VPWR.n1343 5.66204
R11602 VPWR.n2316 VPWR.n2290 5.66204
R11603 VPWR.n3278 VPWR.n3273 5.48841
R11604 VPWR.n1337 VPWR.n1336 5.41234
R11605 VPWR.n580 VPWR.n579 5.27109
R11606 VPWR.n809 VPWR.n805 5.23701
R11607 VPWR.n6244 VPWR.n5741 5.18397
R11608 VPWR.n6391 VPWR.n6390 5.18397
R11609 VPWR.n4997 VPWR.n4996 5.18397
R11610 VPWR.n5178 VPWR.n5177 5.18397
R11611 VPWR.n5281 VPWR.n5280 5.18397
R11612 VPWR.n4649 VPWR.n4648 5.18397
R11613 VPWR.n4548 VPWR.n4547 5.18397
R11614 VPWR.n1040 VPWR.n1017 5.18397
R11615 VPWR.n3905 VPWR.n3885 5.18397
R11616 VPWR.n3547 VPWR.n3546 5.18397
R11617 VPWR.n3427 VPWR.n3426 5.18397
R11618 VPWR.n2210 VPWR.n2209 5.18397
R11619 VPWR.n2510 VPWR.n2508 5.03171
R11620 VPWR.n1342 VPWR.n1341 5.03171
R11621 VPWR.n752 VPWR.n603 4.91172
R11622 VPWR.n1619 VPWR.n1618 4.91172
R11623 VPWR.n763 VPWR.n762 4.89665
R11624 VPWR.n5005 VPWR 4.86662
R11625 VPWR.n1607 VPWR.n1606 4.84444
R11626 VPWR.n1338 VPWR.n1337 4.76083
R11627 VPWR.n2428 VPWR 4.73093
R11628 VPWR.n6252 VPWR.n6251 4.67352
R11629 VPWR.n6141 VPWR.n5828 4.67352
R11630 VPWR.n6141 VPWR.n6140 4.67352
R11631 VPWR.n6134 VPWR.n6133 4.67352
R11632 VPWR.n6117 VPWR.n6116 4.67352
R11633 VPWR.n3309 VPWR.n3308 4.67352
R11634 VPWR.n2442 VPWR.n2426 4.67352
R11635 VPWR.n2585 VPWR.n2579 4.67352
R11636 VPWR.n7670 VPWR.n47 4.67352
R11637 VPWR.n44 VPWR.n43 4.67352
R11638 VPWR.n40 VPWR.n39 4.67352
R11639 VPWR.n34 VPWR.n33 4.67352
R11640 VPWR.n7721 VPWR.n31 4.67352
R11641 VPWR.n7717 VPWR.n31 4.67352
R11642 VPWR.n5026 VPWR.n5021 4.67352
R11643 VPWR.n170 VPWR.n169 4.67352
R11644 VPWR.n4918 VPWR.n4917 4.67352
R11645 VPWR.n4925 VPWR.n4924 4.67352
R11646 VPWR.n6861 VPWR.n6860 4.67352
R11647 VPWR.n7335 VPWR.n7334 4.67352
R11648 VPWR.n7235 VPWR.n7234 4.67352
R11649 VPWR.n7076 VPWR.n7075 4.67352
R11650 VPWR.n7076 VPWR.n4867 4.67352
R11651 VPWR.n7084 VPWR.n7083 4.67352
R11652 VPWR.n5350 VPWR.n5349 4.67352
R11653 VPWR.n895 VPWR.n894 4.67352
R11654 VPWR.n807 VPWR.n806 4.67352
R11655 VPWR.n641 VPWR.n640 4.67352
R11656 VPWR.n354 VPWR.n353 4.67352
R11657 VPWR.n353 VPWR.n352 4.67352
R11658 VPWR.n4502 VPWR.n4500 4.67352
R11659 VPWR.n4488 VPWR.n396 4.67352
R11660 VPWR.n4492 VPWR.n396 4.67352
R11661 VPWR.n1028 VPWR.n1026 4.67352
R11662 VPWR.n1027 VPWR.n1018 4.67352
R11663 VPWR.n1376 VPWR.n1374 4.67352
R11664 VPWR.n1376 VPWR.n1375 4.67352
R11665 VPWR.n1375 VPWR.n437 4.67352
R11666 VPWR.n3994 VPWR.n3993 4.67352
R11667 VPWR.n4073 VPWR.n4072 4.67352
R11668 VPWR.n4072 VPWR.n1536 4.67352
R11669 VPWR.n1538 VPWR.n1536 4.67352
R11670 VPWR.n4213 VPWR.n4212 4.67352
R11671 VPWR.n4212 VPWR.n4211 4.67352
R11672 VPWR.n2006 VPWR.n1644 4.67352
R11673 VPWR.n1955 VPWR.n1954 4.67352
R11674 VPWR.n1865 VPWR.n1864 4.67352
R11675 VPWR.n1869 VPWR.n1843 4.67352
R11676 VPWR.n1796 VPWR.n1795 4.67352
R11677 VPWR.n1795 VPWR.n1794 4.67352
R11678 VPWR.n1573 VPWR.n1572 4.67352
R11679 VPWR.n2858 VPWR.n2857 4.67352
R11680 VPWR.n2799 VPWR.n2798 4.67352
R11681 VPWR.n2708 VPWR.n2707 4.67352
R11682 VPWR.n2894 VPWR.n2893 4.67352
R11683 VPWR.n5852 VPWR.n5851 4.67352
R11684 VPWR.n6251 VPWR.n6250 4.67352
R11685 VPWR.n6312 VPWR.n6278 4.67352
R11686 VPWR.n6140 VPWR.n6139 4.67352
R11687 VPWR.n6133 VPWR.n6048 4.67352
R11688 VPWR.n6116 VPWR.n6115 4.67352
R11689 VPWR.n3308 VPWR.n3307 4.67352
R11690 VPWR.n2427 VPWR.n2426 4.67352
R11691 VPWR.n2609 VPWR.n2576 4.67352
R11692 VPWR.n2589 VPWR.n2579 4.67352
R11693 VPWR.n7681 VPWR.n42 4.67352
R11694 VPWR.n7675 VPWR.n44 4.67352
R11695 VPWR.n7691 VPWR.n40 4.67352
R11696 VPWR.n7717 VPWR.n7716 4.67352
R11697 VPWR.n5018 VPWR.n5017 4.67352
R11698 VPWR.n5038 VPWR.n5018 4.67352
R11699 VPWR.n5026 VPWR.n5025 4.67352
R11700 VPWR.n171 VPWR.n170 4.67352
R11701 VPWR.n6652 VPWR.n6612 4.67352
R11702 VPWR.n7437 VPWR.n7436 4.67352
R11703 VPWR.n6802 VPWR.n6801 4.67352
R11704 VPWR.n6803 VPWR.n6802 4.67352
R11705 VPWR.n4919 VPWR.n4918 4.67352
R11706 VPWR.n6946 VPWR.n4925 4.67352
R11707 VPWR.n7239 VPWR.n7235 4.67352
R11708 VPWR.n7230 VPWR.n7229 4.67352
R11709 VPWR.n5351 VPWR.n5350 4.67352
R11710 VPWR.n321 VPWR.n320 4.67352
R11711 VPWR.n4766 VPWR.n321 4.67352
R11712 VPWR.n908 VPWR.n582 4.67352
R11713 VPWR.n683 VPWR.n681 4.67352
R11714 VPWR.n670 VPWR.n641 4.67352
R11715 VPWR.n352 VPWR.n339 4.67352
R11716 VPWR.n4502 VPWR.n4501 4.67352
R11717 VPWR.n4493 VPWR.n4492 4.67352
R11718 VPWR.n1026 VPWR.n1025 4.67352
R11719 VPWR.n1033 VPWR.n1018 4.67352
R11720 VPWR.n1374 VPWR.n1373 4.67352
R11721 VPWR.n1429 VPWR.n437 4.67352
R11722 VPWR.n1534 VPWR.n1533 4.67352
R11723 VPWR.n4077 VPWR.n1534 4.67352
R11724 VPWR.n4076 VPWR.n4073 4.67352
R11725 VPWR.n4067 VPWR.n1538 4.67352
R11726 VPWR.n4213 VPWR.n1478 4.67352
R11727 VPWR.n2001 VPWR.n2000 4.67352
R11728 VPWR.n1954 VPWR.n1953 4.67352
R11729 VPWR.n1794 VPWR.n1793 4.67352
R11730 VPWR.n1601 VPWR.n1600 4.67352
R11731 VPWR.n3606 VPWR.n3605 4.67352
R11732 VPWR.n1574 VPWR.n1573 4.67352
R11733 VPWR.n3681 VPWR.n3680 4.67352
R11734 VPWR.n2859 VPWR.n2858 4.67352
R11735 VPWR.n2970 VPWR.n2799 4.67352
R11736 VPWR.n2709 VPWR.n2708 4.67352
R11737 VPWR.n2919 VPWR.n2894 4.67352
R11738 VPWR.n5896 VPWR.n5831 4.67352
R11739 VPWR.n7093 VPWR.n7092 4.65596
R11740 VPWR.n5250 VPWR.n5249 4.65519
R11741 VPWR.n754 VPWR.n753 4.65505
R11742 VPWR.n5502 VPWR.n5501 4.6532
R11743 VPWR.n655 VPWR.n644 4.65151
R11744 VPWR.n6963 VPWR.n6962 4.65148
R11745 VPWR.n5380 VPWR.n5379 4.65148
R11746 VPWR.n5203 VPWR.n5141 4.6505
R11747 VPWR.n5098 VPWR.n5097 4.6505
R11748 VPWR.n5100 VPWR.n5099 4.6505
R11749 VPWR.n5102 VPWR.n5101 4.6505
R11750 VPWR.n5103 VPWR.n5092 4.6505
R11751 VPWR.n5202 VPWR.n5201 4.6505
R11752 VPWR.n5200 VPWR.n5199 4.6505
R11753 VPWR.n5198 VPWR.n5197 4.6505
R11754 VPWR.n5195 VPWR.n5194 4.6505
R11755 VPWR.n5193 VPWR.n5192 4.6505
R11756 VPWR.n5191 VPWR.n5190 4.6505
R11757 VPWR.n5189 VPWR.n5188 4.6505
R11758 VPWR.n5186 VPWR.n5185 4.6505
R11759 VPWR.n5179 VPWR.n5178 4.6505
R11760 VPWR.n5176 VPWR.n5175 4.6505
R11761 VPWR.n5174 VPWR.n5173 4.6505
R11762 VPWR.n5172 VPWR.n5171 4.6505
R11763 VPWR.n5168 VPWR.n5167 4.6505
R11764 VPWR.n5161 VPWR.n5160 4.6505
R11765 VPWR.n5158 VPWR.n5157 4.6505
R11766 VPWR.n5156 VPWR.n5155 4.6505
R11767 VPWR.n5154 VPWR.n5153 4.6505
R11768 VPWR.n5152 VPWR.n5151 4.6505
R11769 VPWR.n5149 VPWR.n5148 4.6505
R11770 VPWR.n5146 VPWR.n4940 4.6505
R11771 VPWR.n6706 VPWR.n6705 4.6505
R11772 VPWR.n6746 VPWR.n6745 4.6505
R11773 VPWR.n6742 VPWR.n6741 4.6505
R11774 VPWR.n6738 VPWR.n6737 4.6505
R11775 VPWR.n6709 VPWR.n4938 4.6505
R11776 VPWR.n6618 VPWR.n6615 4.6505
R11777 VPWR.n6619 VPWR.n6614 4.6505
R11778 VPWR.n6624 VPWR.n6613 4.6505
R11779 VPWR.n6651 VPWR.n6650 4.6505
R11780 VPWR.n6711 VPWR.n6710 4.6505
R11781 VPWR.n6713 VPWR.n6712 4.6505
R11782 VPWR.n6715 VPWR.n6714 4.6505
R11783 VPWR.n6717 VPWR.n6716 4.6505
R11784 VPWR.n6720 VPWR.n6719 4.6505
R11785 VPWR.n6722 VPWR.n6721 4.6505
R11786 VPWR.n6724 VPWR.n6723 4.6505
R11787 VPWR.n6726 VPWR.n6725 4.6505
R11788 VPWR.n6728 VPWR.n6727 4.6505
R11789 VPWR.n6730 VPWR.n6729 4.6505
R11790 VPWR.n6732 VPWR.n6731 4.6505
R11791 VPWR.n6734 VPWR.n6733 4.6505
R11792 VPWR.n7585 VPWR.n158 4.6505
R11793 VPWR.n7582 VPWR.n7526 4.6505
R11794 VPWR.n7524 VPWR.n160 4.6505
R11795 VPWR.n7523 VPWR.n160 4.6505
R11796 VPWR.n201 VPWR.n168 4.6505
R11797 VPWR.n181 VPWR.n180 4.6505
R11798 VPWR.n179 VPWR.n172 4.6505
R11799 VPWR.n176 VPWR.n173 4.6505
R11800 VPWR.n200 VPWR.n199 4.6505
R11801 VPWR.n198 VPWR.n197 4.6505
R11802 VPWR.n196 VPWR.n195 4.6505
R11803 VPWR.n194 VPWR.n193 4.6505
R11804 VPWR.n192 VPWR.n191 4.6505
R11805 VPWR.n190 VPWR.n171 4.6505
R11806 VPWR.n187 VPWR.n186 4.6505
R11807 VPWR.n185 VPWR.n184 4.6505
R11808 VPWR.n183 VPWR.n182 4.6505
R11809 VPWR.n178 VPWR.n177 4.6505
R11810 VPWR.n7599 VPWR.n7598 4.6505
R11811 VPWR.n7594 VPWR.n7593 4.6505
R11812 VPWR.n7591 VPWR.n7590 4.6505
R11813 VPWR.n7589 VPWR.n7588 4.6505
R11814 VPWR.n7587 VPWR.n7586 4.6505
R11815 VPWR.n7528 VPWR.n159 4.6505
R11816 VPWR.n7530 VPWR.n7529 4.6505
R11817 VPWR.n7532 VPWR.n7531 4.6505
R11818 VPWR.n7534 VPWR.n7533 4.6505
R11819 VPWR.n7536 VPWR.n7535 4.6505
R11820 VPWR.n7538 VPWR.n7537 4.6505
R11821 VPWR.n7540 VPWR.n7539 4.6505
R11822 VPWR.n7543 VPWR.n7542 4.6505
R11823 VPWR.n7545 VPWR.n7544 4.6505
R11824 VPWR.n7547 VPWR.n7546 4.6505
R11825 VPWR.n7549 VPWR.n7548 4.6505
R11826 VPWR.n7551 VPWR.n7550 4.6505
R11827 VPWR.n7553 VPWR.n7552 4.6505
R11828 VPWR.n7555 VPWR.n7554 4.6505
R11829 VPWR.n7557 VPWR.n7556 4.6505
R11830 VPWR.n7559 VPWR.n7558 4.6505
R11831 VPWR.n7561 VPWR.n7560 4.6505
R11832 VPWR.n7563 VPWR.n7562 4.6505
R11833 VPWR.n7565 VPWR.n7564 4.6505
R11834 VPWR.n7567 VPWR.n7566 4.6505
R11835 VPWR.n7569 VPWR.n7568 4.6505
R11836 VPWR.n7571 VPWR.n7570 4.6505
R11837 VPWR.n7573 VPWR.n7572 4.6505
R11838 VPWR.n7575 VPWR.n7574 4.6505
R11839 VPWR.n7577 VPWR.n7576 4.6505
R11840 VPWR.n7579 VPWR.n7578 4.6505
R11841 VPWR.n7581 VPWR.n7580 4.6505
R11842 VPWR.n7522 VPWR.n7521 4.6505
R11843 VPWR.n203 VPWR.n202 4.6505
R11844 VPWR.n6744 VPWR.n6743 4.6505
R11845 VPWR.n6740 VPWR.n6739 4.6505
R11846 VPWR.n6736 VPWR.n6735 4.6505
R11847 VPWR.n6617 VPWR.n6616 4.6505
R11848 VPWR.n6621 VPWR.n6620 4.6505
R11849 VPWR.n6623 VPWR.n6622 4.6505
R11850 VPWR.n6626 VPWR.n6625 4.6505
R11851 VPWR.n6628 VPWR.n6627 4.6505
R11852 VPWR.n6630 VPWR.n6629 4.6505
R11853 VPWR.n6632 VPWR.n6631 4.6505
R11854 VPWR.n6634 VPWR.n6633 4.6505
R11855 VPWR.n6636 VPWR.n6635 4.6505
R11856 VPWR.n6638 VPWR.n6637 4.6505
R11857 VPWR.n6640 VPWR.n6639 4.6505
R11858 VPWR.n6643 VPWR.n6642 4.6505
R11859 VPWR.n6645 VPWR.n6644 4.6505
R11860 VPWR.n6647 VPWR.n6646 4.6505
R11861 VPWR.n6649 VPWR.n6648 4.6505
R11862 VPWR.n6653 VPWR.n6652 4.6505
R11863 VPWR.n5166 VPWR.n5165 4.6505
R11864 VPWR.n5170 VPWR.n5169 4.6505
R11865 VPWR.n5181 VPWR.n5180 4.6505
R11866 VPWR.n5183 VPWR.n5182 4.6505
R11867 VPWR.n5111 VPWR.n5110 4.6505
R11868 VPWR.n5116 VPWR.n5115 4.6505
R11869 VPWR.n5574 VPWR.n5463 4.6505
R11870 VPWR.n5500 VPWR.n5499 4.6505
R11871 VPWR.n5431 VPWR.n5428 4.6505
R11872 VPWR.n5435 VPWR.n5434 4.6505
R11873 VPWR.n5573 VPWR.n5572 4.6505
R11874 VPWR.n5571 VPWR.n5570 4.6505
R11875 VPWR.n5569 VPWR.n5568 4.6505
R11876 VPWR.n5566 VPWR.n5565 4.6505
R11877 VPWR.n5564 VPWR.n5563 4.6505
R11878 VPWR.n5562 VPWR.n5561 4.6505
R11879 VPWR.n5560 VPWR.n5559 4.6505
R11880 VPWR.n5556 VPWR.n5555 4.6505
R11881 VPWR.n5544 VPWR.n5543 4.6505
R11882 VPWR.n5542 VPWR.n5541 4.6505
R11883 VPWR.n5539 VPWR.n5538 4.6505
R11884 VPWR.n5527 VPWR.n5526 4.6505
R11885 VPWR.n5523 VPWR.n5522 4.6505
R11886 VPWR.n6865 VPWR.n6796 4.6505
R11887 VPWR.n6855 VPWR.n6797 4.6505
R11888 VPWR.n6810 VPWR.n6809 4.6505
R11889 VPWR.n6812 VPWR.n6811 4.6505
R11890 VPWR.n6814 VPWR.n6813 4.6505
R11891 VPWR.n6818 VPWR.n6817 4.6505
R11892 VPWR.n6842 VPWR.n6841 4.6505
R11893 VPWR.n6844 VPWR.n6843 4.6505
R11894 VPWR.n6848 VPWR.n6847 4.6505
R11895 VPWR.n7455 VPWR.n7440 4.6505
R11896 VPWR.n7452 VPWR.n7441 4.6505
R11897 VPWR.n7449 VPWR.n7448 4.6505
R11898 VPWR.n7447 VPWR.n7442 4.6505
R11899 VPWR.n7446 VPWR.n7443 4.6505
R11900 VPWR.n7470 VPWR.n7469 4.6505
R11901 VPWR.n7468 VPWR.n7467 4.6505
R11902 VPWR.n7466 VPWR.n7465 4.6505
R11903 VPWR.n7464 VPWR.n7463 4.6505
R11904 VPWR.n7460 VPWR.n7459 4.6505
R11905 VPWR.n7458 VPWR.n7457 4.6505
R11906 VPWR.n7456 VPWR.n7439 4.6505
R11907 VPWR.n7454 VPWR.n7453 4.6505
R11908 VPWR.n7451 VPWR.n7450 4.6505
R11909 VPWR.n7472 VPWR.n7471 4.6505
R11910 VPWR.n6864 VPWR.n6863 4.6505
R11911 VPWR.n6857 VPWR.n6856 4.6505
R11912 VPWR.n6804 VPWR.n6798 4.6505
R11913 VPWR.n6806 VPWR.n6805 4.6505
R11914 VPWR.n6808 VPWR.n6807 4.6505
R11915 VPWR.n6816 VPWR.n6815 4.6505
R11916 VPWR.n6824 VPWR.n6823 4.6505
R11917 VPWR.n6826 VPWR.n6825 4.6505
R11918 VPWR.n6829 VPWR.n6828 4.6505
R11919 VPWR.n6831 VPWR.n6830 4.6505
R11920 VPWR.n6833 VPWR.n6832 4.6505
R11921 VPWR.n6836 VPWR.n6803 4.6505
R11922 VPWR.n6838 VPWR.n6837 4.6505
R11923 VPWR.n6840 VPWR.n6839 4.6505
R11924 VPWR.n6846 VPWR.n6845 4.6505
R11925 VPWR.n6849 VPWR.n6800 4.6505
R11926 VPWR.n6852 VPWR.n6851 4.6505
R11927 VPWR.n7407 VPWR.n7406 4.6505
R11928 VPWR.n6990 VPWR.n6989 4.6505
R11929 VPWR.n6988 VPWR.n6987 4.6505
R11930 VPWR.n6986 VPWR.n6985 4.6505
R11931 VPWR.n6984 VPWR.n6983 4.6505
R11932 VPWR.n6982 VPWR.n6981 4.6505
R11933 VPWR.n6980 VPWR.n6979 4.6505
R11934 VPWR.n6978 VPWR.n6977 4.6505
R11935 VPWR.n6976 VPWR.n6975 4.6505
R11936 VPWR.n6974 VPWR.n6973 4.6505
R11937 VPWR.n6972 VPWR.n6971 4.6505
R11938 VPWR.n6970 VPWR.n4919 4.6505
R11939 VPWR.n6967 VPWR.n6966 4.6505
R11940 VPWR.n6965 VPWR.n6964 4.6505
R11941 VPWR.n6961 VPWR.n6960 4.6505
R11942 VPWR.n6959 VPWR.n4920 4.6505
R11943 VPWR.n6958 VPWR.n6957 4.6505
R11944 VPWR.n6956 VPWR.n6955 4.6505
R11945 VPWR.n6954 VPWR.n6953 4.6505
R11946 VPWR.n6952 VPWR.n6951 4.6505
R11947 VPWR.n6950 VPWR.n4922 4.6505
R11948 VPWR.n6947 VPWR.n6946 4.6505
R11949 VPWR.n6945 VPWR.n6944 4.6505
R11950 VPWR.n6943 VPWR.n6942 4.6505
R11951 VPWR.n6941 VPWR.n6940 4.6505
R11952 VPWR.n6939 VPWR.n6938 4.6505
R11953 VPWR.n6937 VPWR.n6936 4.6505
R11954 VPWR.n6934 VPWR.n6933 4.6505
R11955 VPWR.n6932 VPWR.n6931 4.6505
R11956 VPWR.n6930 VPWR.n6929 4.6505
R11957 VPWR.n6928 VPWR.n6927 4.6505
R11958 VPWR.n6926 VPWR.n6925 4.6505
R11959 VPWR.n6924 VPWR.n6923 4.6505
R11960 VPWR.n6922 VPWR.n4926 4.6505
R11961 VPWR.n6921 VPWR.n6920 4.6505
R11962 VPWR.n5497 VPWR.n5467 4.6505
R11963 VPWR.n5504 VPWR.n5503 4.6505
R11964 VPWR.n5506 VPWR.n5505 4.6505
R11965 VPWR.n5508 VPWR.n5507 4.6505
R11966 VPWR.n5510 VPWR.n5509 4.6505
R11967 VPWR.n5512 VPWR.n5511 4.6505
R11968 VPWR.n5514 VPWR.n5513 4.6505
R11969 VPWR.n5517 VPWR.n5516 4.6505
R11970 VPWR.n5519 VPWR.n5518 4.6505
R11971 VPWR.n5521 VPWR.n5520 4.6505
R11972 VPWR.n5525 VPWR.n5524 4.6505
R11973 VPWR.n5529 VPWR.n5528 4.6505
R11974 VPWR.n5531 VPWR.n5530 4.6505
R11975 VPWR.n5533 VPWR.n5532 4.6505
R11976 VPWR.n5535 VPWR.n5534 4.6505
R11977 VPWR.n5537 VPWR.n5536 4.6505
R11978 VPWR.n5558 VPWR.n5465 4.6505
R11979 VPWR.n5433 VPWR.n5432 4.6505
R11980 VPWR.n5437 VPWR.n5436 4.6505
R11981 VPWR.n5439 VPWR.n5438 4.6505
R11982 VPWR.n5441 VPWR.n5440 4.6505
R11983 VPWR.n5442 VPWR.n5427 4.6505
R11984 VPWR.n5444 VPWR.n5443 4.6505
R11985 VPWR.n5446 VPWR.n5445 4.6505
R11986 VPWR.n5448 VPWR.n5447 4.6505
R11987 VPWR.n5450 VPWR.n5449 4.6505
R11988 VPWR.n5453 VPWR.n5452 4.6505
R11989 VPWR.n5455 VPWR.n5454 4.6505
R11990 VPWR.n5456 VPWR.n5426 4.6505
R11991 VPWR.n5458 VPWR.n5457 4.6505
R11992 VPWR.n5460 VPWR.n5459 4.6505
R11993 VPWR.n5462 VPWR.n5461 4.6505
R11994 VPWR.n5323 VPWR.n5231 4.6505
R11995 VPWR.n5318 VPWR.n5232 4.6505
R11996 VPWR.n5313 VPWR.n5234 4.6505
R11997 VPWR.n5310 VPWR.n5285 4.6505
R11998 VPWR.n5367 VPWR.n5366 4.6505
R11999 VPWR.n5371 VPWR.n5370 4.6505
R12000 VPWR.n5373 VPWR.n5372 4.6505
R12001 VPWR.n5242 VPWR.n5241 4.6505
R12002 VPWR.n5244 VPWR.n5243 4.6505
R12003 VPWR.n5246 VPWR.n5245 4.6505
R12004 VPWR.n5248 VPWR.n5247 4.6505
R12005 VPWR.n5252 VPWR.n5251 4.6505
R12006 VPWR.n5254 VPWR.n5253 4.6505
R12007 VPWR.n5256 VPWR.n5255 4.6505
R12008 VPWR.n5259 VPWR.n5258 4.6505
R12009 VPWR.n5261 VPWR.n5260 4.6505
R12010 VPWR.n5263 VPWR.n5262 4.6505
R12011 VPWR.n5265 VPWR.n5264 4.6505
R12012 VPWR.n5267 VPWR.n5266 4.6505
R12013 VPWR.n5269 VPWR.n5268 4.6505
R12014 VPWR.n5271 VPWR.n5270 4.6505
R12015 VPWR.n5273 VPWR.n5272 4.6505
R12016 VPWR.n5274 VPWR.n5236 4.6505
R12017 VPWR.n5276 VPWR.n5275 4.6505
R12018 VPWR.n5278 VPWR.n5277 4.6505
R12019 VPWR.n5280 VPWR.n5279 4.6505
R12020 VPWR.n5283 VPWR.n5282 4.6505
R12021 VPWR.n5284 VPWR.n5235 4.6505
R12022 VPWR.n5309 VPWR.n5308 4.6505
R12023 VPWR.n5307 VPWR.n5286 4.6505
R12024 VPWR.n5306 VPWR.n5305 4.6505
R12025 VPWR.n7069 VPWR 4.6505
R12026 VPWR.n7070 VPWR.n4871 4.6505
R12027 VPWR.n7072 VPWR.n7071 4.6505
R12028 VPWR.n7117 VPWR.n4864 4.6505
R12029 VPWR.n7119 VPWR.n7118 4.6505
R12030 VPWR.n7121 VPWR.n7120 4.6505
R12031 VPWR.n7222 VPWR.n7221 4.6505
R12032 VPWR.n7225 VPWR.n292 4.6505
R12033 VPWR.n7273 VPWR.n7226 4.6505
R12034 VPWR.n7247 VPWR.n7231 4.6505
R12035 VPWR.n7246 VPWR.n7233 4.6505
R12036 VPWR.n7236 VPWR.n291 4.6505
R12037 VPWR.n7278 VPWR.n290 4.6505
R12038 VPWR.n7282 VPWR.n7281 4.6505
R12039 VPWR.n7339 VPWR.n7327 4.6505
R12040 VPWR.n7341 VPWR.n7340 4.6505
R12041 VPWR.n7360 VPWR.n7359 4.6505
R12042 VPWR.n7358 VPWR.n7357 4.6505
R12043 VPWR.n7356 VPWR.n7355 4.6505
R12044 VPWR.n7354 VPWR.n7353 4.6505
R12045 VPWR.n7352 VPWR.n7351 4.6505
R12046 VPWR.n7347 VPWR.n7346 4.6505
R12047 VPWR.n7331 VPWR.n7330 4.6505
R12048 VPWR.n7338 VPWR.n7337 4.6505
R12049 VPWR.n7343 VPWR.n7342 4.6505
R12050 VPWR.n7345 VPWR.n7344 4.6505
R12051 VPWR.n7348 VPWR.n7326 4.6505
R12052 VPWR.n7350 VPWR.n7349 4.6505
R12053 VPWR.n7362 VPWR.n7361 4.6505
R12054 VPWR.n7224 VPWR.n7223 4.6505
R12055 VPWR.n7270 VPWR.n7230 4.6505
R12056 VPWR.n7267 VPWR.n7266 4.6505
R12057 VPWR.n7265 VPWR.n7264 4.6505
R12058 VPWR.n7263 VPWR.n7262 4.6505
R12059 VPWR.n7261 VPWR.n7260 4.6505
R12060 VPWR.n7259 VPWR.n7258 4.6505
R12061 VPWR.n7257 VPWR.n7256 4.6505
R12062 VPWR.n7255 VPWR.n7254 4.6505
R12063 VPWR.n7253 VPWR.n7252 4.6505
R12064 VPWR.n7251 VPWR.n7250 4.6505
R12065 VPWR.n7249 VPWR.n7248 4.6505
R12066 VPWR.n7244 VPWR.n7243 4.6505
R12067 VPWR.n7240 VPWR.n7239 4.6505
R12068 VPWR.n7238 VPWR.n7237 4.6505
R12069 VPWR.n7277 VPWR.n7276 4.6505
R12070 VPWR.n7280 VPWR.n7279 4.6505
R12071 VPWR.n7284 VPWR.n7283 4.6505
R12072 VPWR.n7286 VPWR.n7285 4.6505
R12073 VPWR.n7219 VPWR.n7218 4.6505
R12074 VPWR.n7075 VPWR.n7074 4.6505
R12075 VPWR.n7077 VPWR.n7076 4.6505
R12076 VPWR.n7080 VPWR.n7079 4.6505
R12077 VPWR.n7087 VPWR.n7086 4.6505
R12078 VPWR.n7091 VPWR.n7090 4.6505
R12079 VPWR.n7095 VPWR.n7094 4.6505
R12080 VPWR.n7096 VPWR.n4866 4.6505
R12081 VPWR.n7098 VPWR.n7097 4.6505
R12082 VPWR.n7100 VPWR.n7099 4.6505
R12083 VPWR.n7103 VPWR.n7102 4.6505
R12084 VPWR.n7106 VPWR.n7105 4.6505
R12085 VPWR.n7108 VPWR.n7107 4.6505
R12086 VPWR.n7110 VPWR.n7109 4.6505
R12087 VPWR.n7116 VPWR.n7115 4.6505
R12088 VPWR.n7122 VPWR.n4863 4.6505
R12089 VPWR.n7124 VPWR.n7123 4.6505
R12090 VPWR.n7126 VPWR.n7125 4.6505
R12091 VPWR.n7129 VPWR.n7128 4.6505
R12092 VPWR.n7134 VPWR.n7133 4.6505
R12093 VPWR.n7137 VPWR.n7136 4.6505
R12094 VPWR.n7139 VPWR.n7138 4.6505
R12095 VPWR.n5239 VPWR.n5233 4.6505
R12096 VPWR.n5315 VPWR.n5314 4.6505
R12097 VPWR.n5320 VPWR.n5319 4.6505
R12098 VPWR.n5322 VPWR.n5321 4.6505
R12099 VPWR.n5355 VPWR.n5354 4.6505
R12100 VPWR.n5358 VPWR.n5351 4.6505
R12101 VPWR.n5360 VPWR.n5359 4.6505
R12102 VPWR.n5362 VPWR.n5361 4.6505
R12103 VPWR.n5365 VPWR.n5364 4.6505
R12104 VPWR.n5369 VPWR.n5368 4.6505
R12105 VPWR.n5374 VPWR.n5346 4.6505
R12106 VPWR.n5376 VPWR.n5375 4.6505
R12107 VPWR.n969 VPWR.n571 4.6505
R12108 VPWR.n968 VPWR.n572 4.6505
R12109 VPWR.n957 VPWR.n574 4.6505
R12110 VPWR.n672 VPWR.n671 4.6505
R12111 VPWR.n676 VPWR.n675 4.6505
R12112 VPWR.n678 VPWR.n575 4.6505
R12113 VPWR.n482 VPWR.n481 4.6505
R12114 VPWR.n489 VPWR.n488 4.6505
R12115 VPWR.n503 VPWR.n475 4.6505
R12116 VPWR.n963 VPWR.n962 4.6505
R12117 VPWR.n961 VPWR.n960 4.6505
R12118 VPWR.n650 VPWR.n649 4.6505
R12119 VPWR.n652 VPWR.n651 4.6505
R12120 VPWR.n654 VPWR.n653 4.6505
R12121 VPWR.n659 VPWR.n658 4.6505
R12122 VPWR.n681 VPWR.n680 4.6505
R12123 VPWR.n684 VPWR.n683 4.6505
R12124 VPWR.n776 VPWR.n775 4.6505
R12125 VPWR.n778 VPWR.n777 4.6505
R12126 VPWR.n782 VPWR.n781 4.6505
R12127 VPWR.n783 VPWR.n576 4.6505
R12128 VPWR.n793 VPWR.n792 4.6505
R12129 VPWR.n797 VPWR.n796 4.6505
R12130 VPWR.n891 VPWR.n890 4.6505
R12131 VPWR.n898 VPWR.n897 4.6505
R12132 VPWR.n909 VPWR.n581 4.6505
R12133 VPWR.n911 VPWR.n910 4.6505
R12134 VPWR.n925 VPWR.n924 4.6505
R12135 VPWR.n931 VPWR.n930 4.6505
R12136 VPWR.n933 VPWR.n932 4.6505
R12137 VPWR.n935 VPWR.n934 4.6505
R12138 VPWR.n943 VPWR.n942 4.6505
R12139 VPWR.n945 VPWR.n580 4.6505
R12140 VPWR.n949 VPWR.n578 4.6505
R12141 VPWR.n4802 VPWR.n4799 4.6505
R12142 VPWR.n4803 VPWR.n4798 4.6505
R12143 VPWR.n4805 VPWR.n4804 4.6505
R12144 VPWR.n4808 VPWR.n4797 4.6505
R12145 VPWR.n4812 VPWR.n4811 4.6505
R12146 VPWR.n4825 VPWR.n4796 4.6505
R12147 VPWR.n4807 VPWR.n4806 4.6505
R12148 VPWR.n4810 VPWR.n4809 4.6505
R12149 VPWR.n4814 VPWR.n4813 4.6505
R12150 VPWR.n4816 VPWR.n4815 4.6505
R12151 VPWR.n4818 VPWR.n4817 4.6505
R12152 VPWR.n4820 VPWR.n4819 4.6505
R12153 VPWR.n4822 VPWR.n4821 4.6505
R12154 VPWR.n4824 VPWR.n4823 4.6505
R12155 VPWR.n4827 VPWR.n4826 4.6505
R12156 VPWR.n4829 VPWR.n4828 4.6505
R12157 VPWR.n4831 VPWR.n4830 4.6505
R12158 VPWR.n889 VPWR.n888 4.6505
R12159 VPWR.n893 VPWR.n577 4.6505
R12160 VPWR.n902 VPWR.n901 4.6505
R12161 VPWR.n905 VPWR.n904 4.6505
R12162 VPWR.n908 VPWR.n907 4.6505
R12163 VPWR.n913 VPWR.n912 4.6505
R12164 VPWR.n915 VPWR.n914 4.6505
R12165 VPWR.n917 VPWR.n916 4.6505
R12166 VPWR.n919 VPWR.n918 4.6505
R12167 VPWR.n921 VPWR.n920 4.6505
R12168 VPWR.n923 VPWR.n922 4.6505
R12169 VPWR.n927 VPWR.n926 4.6505
R12170 VPWR.n929 VPWR.n928 4.6505
R12171 VPWR.n937 VPWR.n936 4.6505
R12172 VPWR.n939 VPWR.n938 4.6505
R12173 VPWR.n941 VPWR.n940 4.6505
R12174 VPWR.n951 VPWR.n950 4.6505
R12175 VPWR.n948 VPWR.n947 4.6505
R12176 VPWR.n4766 VPWR.n4765 4.6505
R12177 VPWR.n747 VPWR.n746 4.6505
R12178 VPWR.n749 VPWR.n748 4.6505
R12179 VPWR.n751 VPWR.n750 4.6505
R12180 VPWR.n757 VPWR.n756 4.6505
R12181 VPWR.n761 VPWR.n760 4.6505
R12182 VPWR.n766 VPWR.n765 4.6505
R12183 VPWR.n768 VPWR.n767 4.6505
R12184 VPWR.n770 VPWR.n769 4.6505
R12185 VPWR.n772 VPWR.n771 4.6505
R12186 VPWR.n774 VPWR.n773 4.6505
R12187 VPWR.n780 VPWR.n779 4.6505
R12188 VPWR.n785 VPWR.n784 4.6505
R12189 VPWR.n787 VPWR.n786 4.6505
R12190 VPWR.n789 VPWR.n788 4.6505
R12191 VPWR.n791 VPWR.n790 4.6505
R12192 VPWR.n795 VPWR.n794 4.6505
R12193 VPWR.n799 VPWR.n798 4.6505
R12194 VPWR.n801 VPWR.n800 4.6505
R12195 VPWR.n803 VPWR.n802 4.6505
R12196 VPWR.n805 VPWR.n804 4.6505
R12197 VPWR.n810 VPWR.n809 4.6505
R12198 VPWR.n814 VPWR.n813 4.6505
R12199 VPWR.n816 VPWR.n815 4.6505
R12200 VPWR.n818 VPWR.n817 4.6505
R12201 VPWR.n820 VPWR.n819 4.6505
R12202 VPWR.n745 VPWR.n744 4.6505
R12203 VPWR.n679 VPWR.n638 4.6505
R12204 VPWR.n674 VPWR.n673 4.6505
R12205 VPWR.n670 VPWR.n669 4.6505
R12206 VPWR.n666 VPWR.n665 4.6505
R12207 VPWR.n663 VPWR.n662 4.6505
R12208 VPWR.n661 VPWR.n660 4.6505
R12209 VPWR.n657 VPWR.n656 4.6505
R12210 VPWR.n647 VPWR.n573 4.6505
R12211 VPWR.n959 VPWR.n958 4.6505
R12212 VPWR.n965 VPWR.n964 4.6505
R12213 VPWR.n967 VPWR.n966 4.6505
R12214 VPWR VPWR.n478 4.6505
R12215 VPWR.n484 VPWR.n483 4.6505
R12216 VPWR.n486 VPWR.n485 4.6505
R12217 VPWR.n491 VPWR.n490 4.6505
R12218 VPWR.n493 VPWR.n492 4.6505
R12219 VPWR.n498 VPWR.n497 4.6505
R12220 VPWR.n500 VPWR.n499 4.6505
R12221 VPWR.n502 VPWR.n501 4.6505
R12222 VPWR.n505 VPWR.n504 4.6505
R12223 VPWR.n507 VPWR.n506 4.6505
R12224 VPWR.n510 VPWR.n509 4.6505
R12225 VPWR.n1203 VPWR.n1090 4.6505
R12226 VPWR.n1153 VPWR.n1152 4.6505
R12227 VPWR.n1149 VPWR.n1093 4.6505
R12228 VPWR.n1148 VPWR.n1094 4.6505
R12229 VPWR.n1131 VPWR.n1098 4.6505
R12230 VPWR.n1196 VPWR.n1195 4.6505
R12231 VPWR.n1191 VPWR.n1190 4.6505
R12232 VPWR.n1189 VPWR.n1188 4.6505
R12233 VPWR.n1182 VPWR.n1181 4.6505
R12234 VPWR.n1145 VPWR.n1144 4.6505
R12235 VPWR.n1143 VPWR.n1142 4.6505
R12236 VPWR.n1141 VPWR.n1140 4.6505
R12237 VPWR.n1138 VPWR.n1137 4.6505
R12238 VPWR.n1134 VPWR.n1133 4.6505
R12239 VPWR.n4472 VPWR.n4471 4.6505
R12240 VPWR.n4482 VPWR.n4481 4.6505
R12241 VPWR.n4634 VPWR.n373 4.6505
R12242 VPWR.n344 VPWR.n341 4.6505
R12243 VPWR.n345 VPWR.n340 4.6505
R12244 VPWR.n347 VPWR.n346 4.6505
R12245 VPWR.n360 VPWR.n336 4.6505
R12246 VPWR.n349 VPWR.n348 4.6505
R12247 VPWR.n350 VPWR.n339 4.6505
R12248 VPWR.n352 VPWR.n351 4.6505
R12249 VPWR.n353 VPWR.n338 4.6505
R12250 VPWR.n355 VPWR.n354 4.6505
R12251 VPWR.n359 VPWR.n358 4.6505
R12252 VPWR.n362 VPWR.n361 4.6505
R12253 VPWR.n364 VPWR.n363 4.6505
R12254 VPWR.n366 VPWR.n365 4.6505
R12255 VPWR.n4613 VPWR.n4612 4.6505
R12256 VPWR.n4615 VPWR.n4614 4.6505
R12257 VPWR.n4617 VPWR.n4616 4.6505
R12258 VPWR.n4619 VPWR.n4618 4.6505
R12259 VPWR.n4620 VPWR.n378 4.6505
R12260 VPWR.n4622 VPWR.n4621 4.6505
R12261 VPWR.n4624 VPWR.n4623 4.6505
R12262 VPWR.n4627 VPWR.n4626 4.6505
R12263 VPWR.n4629 VPWR.n4628 4.6505
R12264 VPWR.n4631 VPWR.n4630 4.6505
R12265 VPWR.n4633 VPWR.n4632 4.6505
R12266 VPWR.n4637 VPWR.n4636 4.6505
R12267 VPWR.n4639 VPWR.n4638 4.6505
R12268 VPWR.n4641 VPWR.n4640 4.6505
R12269 VPWR.n4643 VPWR.n4642 4.6505
R12270 VPWR.n4645 VPWR.n4644 4.6505
R12271 VPWR.n4646 VPWR.n371 4.6505
R12272 VPWR.n4648 VPWR.n4647 4.6505
R12273 VPWR.n4651 VPWR.n4650 4.6505
R12274 VPWR.n4652 VPWR.n370 4.6505
R12275 VPWR.n4654 VPWR.n4653 4.6505
R12276 VPWR.n4656 VPWR.n4655 4.6505
R12277 VPWR.n4658 VPWR.n4657 4.6505
R12278 VPWR.n4662 VPWR.n4661 4.6505
R12279 VPWR.n4664 VPWR.n4663 4.6505
R12280 VPWR.n4665 VPWR.n367 4.6505
R12281 VPWR.n4667 VPWR.n4666 4.6505
R12282 VPWR.n4669 VPWR.n4668 4.6505
R12283 VPWR.n4672 VPWR.n4671 4.6505
R12284 VPWR.n4674 VPWR.n4673 4.6505
R12285 VPWR.n4676 VPWR.n4675 4.6505
R12286 VPWR.n4464 VPWR.n4463 4.6505
R12287 VPWR.n4466 VPWR.n4465 4.6505
R12288 VPWR.n4468 VPWR.n4467 4.6505
R12289 VPWR.n4470 VPWR.n4469 4.6505
R12290 VPWR.n4474 VPWR.n4473 4.6505
R12291 VPWR.n4476 VPWR.n4475 4.6505
R12292 VPWR.n4478 VPWR.n4477 4.6505
R12293 VPWR.n4480 VPWR.n4479 4.6505
R12294 VPWR.n4483 VPWR.n398 4.6505
R12295 VPWR.n4485 VPWR.n4484 4.6505
R12296 VPWR.n4489 VPWR.n4488 4.6505
R12297 VPWR.n4492 VPWR.n4491 4.6505
R12298 VPWR.n4494 VPWR.n4493 4.6505
R12299 VPWR.n4495 VPWR.n395 4.6505
R12300 VPWR.n4498 VPWR.n4497 4.6505
R12301 VPWR.n4503 VPWR.n4502 4.6505
R12302 VPWR.n4507 VPWR.n4506 4.6505
R12303 VPWR.n4509 VPWR.n4508 4.6505
R12304 VPWR.n4513 VPWR.n4512 4.6505
R12305 VPWR.n4515 VPWR.n4514 4.6505
R12306 VPWR.n4518 VPWR.n4517 4.6505
R12307 VPWR.n4521 VPWR.n394 4.6505
R12308 VPWR.n4523 VPWR.n4522 4.6505
R12309 VPWR.n4525 VPWR.n4524 4.6505
R12310 VPWR.n4527 VPWR.n4526 4.6505
R12311 VPWR.n4528 VPWR.n391 4.6505
R12312 VPWR.n4530 VPWR.n4529 4.6505
R12313 VPWR.n4532 VPWR.n4531 4.6505
R12314 VPWR.n1130 VPWR.n1129 4.6505
R12315 VPWR.n1132 VPWR.n1097 4.6505
R12316 VPWR.n1136 VPWR.n1135 4.6505
R12317 VPWR.n1147 VPWR.n1146 4.6505
R12318 VPWR.n1151 VPWR.n1150 4.6505
R12319 VPWR.n1155 VPWR.n1154 4.6505
R12320 VPWR.n1157 VPWR.n1156 4.6505
R12321 VPWR.n1159 VPWR.n1158 4.6505
R12322 VPWR.n1161 VPWR.n1160 4.6505
R12323 VPWR.n1163 VPWR.n1162 4.6505
R12324 VPWR.n1165 VPWR.n1164 4.6505
R12325 VPWR.n1167 VPWR.n1166 4.6505
R12326 VPWR.n1170 VPWR.n1169 4.6505
R12327 VPWR.n1172 VPWR.n1171 4.6505
R12328 VPWR.n1174 VPWR.n1173 4.6505
R12329 VPWR.n1176 VPWR.n1175 4.6505
R12330 VPWR.n1178 VPWR.n1177 4.6505
R12331 VPWR.n1180 VPWR.n1179 4.6505
R12332 VPWR.n1184 VPWR.n1183 4.6505
R12333 VPWR.n1186 VPWR.n1185 4.6505
R12334 VPWR.n1187 VPWR.n1092 4.6505
R12335 VPWR.n1194 VPWR.n1193 4.6505
R12336 VPWR.n1198 VPWR.n1197 4.6505
R12337 VPWR.n1200 VPWR.n1199 4.6505
R12338 VPWR.n1202 VPWR.n1201 4.6505
R12339 VPWR.n1025 VPWR.n1024 4.6505
R12340 VPWR.n1026 VPWR.n1019 4.6505
R12341 VPWR.n1029 VPWR.n1028 4.6505
R12342 VPWR.n1033 VPWR.n1032 4.6505
R12343 VPWR.n1035 VPWR.n1034 4.6505
R12344 VPWR.n1037 VPWR.n1036 4.6505
R12345 VPWR.n1039 VPWR.n1038 4.6505
R12346 VPWR.n1041 VPWR.n1040 4.6505
R12347 VPWR.n1043 VPWR.n1042 4.6505
R12348 VPWR.n1045 VPWR.n1044 4.6505
R12349 VPWR.n1310 VPWR.n1309 4.6505
R12350 VPWR.n1370 VPWR.n1369 4.6505
R12351 VPWR.n1372 VPWR.n441 4.6505
R12352 VPWR.n1427 VPWR.n438 4.6505
R12353 VPWR.n1424 VPWR.n1380 4.6505
R12354 VPWR.n1231 VPWR.n1230 4.6505
R12355 VPWR.n1235 VPWR.n1234 4.6505
R12356 VPWR.n1242 VPWR.n1227 4.6505
R12357 VPWR.n1246 VPWR.n1245 4.6505
R12358 VPWR.n1321 VPWR.n1320 4.6505
R12359 VPWR.n1324 VPWR.n1323 4.6505
R12360 VPWR.n1328 VPWR.n1327 4.6505
R12361 VPWR.n1333 VPWR.n1332 4.6505
R12362 VPWR.n1335 VPWR.n1334 4.6505
R12363 VPWR.n1339 VPWR.n1338 4.6505
R12364 VPWR.n1341 VPWR.n1340 4.6505
R12365 VPWR.n1345 VPWR.n1344 4.6505
R12366 VPWR.n1348 VPWR.n1347 4.6505
R12367 VPWR.n1350 VPWR.n1349 4.6505
R12368 VPWR.n1353 VPWR.n1352 4.6505
R12369 VPWR.n1355 VPWR.n1354 4.6505
R12370 VPWR.n1357 VPWR.n1356 4.6505
R12371 VPWR.n1359 VPWR.n1358 4.6505
R12372 VPWR.n1361 VPWR.n1360 4.6505
R12373 VPWR.n1363 VPWR.n1362 4.6505
R12374 VPWR.n1365 VPWR.n1364 4.6505
R12375 VPWR.n1367 VPWR.n1366 4.6505
R12376 VPWR.n1377 VPWR.n1376 4.6505
R12377 VPWR.n1379 VPWR.n437 4.6505
R12378 VPWR.n1429 VPWR.n1428 4.6505
R12379 VPWR.n4387 VPWR.n429 4.6505
R12380 VPWR.n4386 VPWR.n430 4.6505
R12381 VPWR.n4372 VPWR.n432 4.6505
R12382 VPWR.n4371 VPWR.n433 4.6505
R12383 VPWR.n4368 VPWR.n434 4.6505
R12384 VPWR.n4365 VPWR.n4364 4.6505
R12385 VPWR.n4362 VPWR.n436 4.6505
R12386 VPWR.n4356 VPWR.n1433 4.6505
R12387 VPWR.n4353 VPWR.n4352 4.6505
R12388 VPWR.n4351 VPWR.n1434 4.6505
R12389 VPWR.n4350 VPWR.n1435 4.6505
R12390 VPWR.n4349 VPWR.n1436 4.6505
R12391 VPWR.n3814 VPWR.n3813 4.6505
R12392 VPWR.n3863 VPWR.n3781 4.6505
R12393 VPWR.n3851 VPWR.n3850 4.6505
R12394 VPWR.n3842 VPWR.n3818 4.6505
R12395 VPWR.n3832 VPWR.n3820 4.6505
R12396 VPWR.n3831 VPWR.n3821 4.6505
R12397 VPWR.n3829 VPWR.n3823 4.6505
R12398 VPWR.n3828 VPWR.n3824 4.6505
R12399 VPWR.n3923 VPWR.n3922 4.6505
R12400 VPWR.n3918 VPWR.n3917 4.6505
R12401 VPWR.n3916 VPWR.n3915 4.6505
R12402 VPWR.n3914 VPWR.n3913 4.6505
R12403 VPWR.n3912 VPWR.n3911 4.6505
R12404 VPWR.n3910 VPWR.n3909 4.6505
R12405 VPWR.n3908 VPWR.n3884 4.6505
R12406 VPWR.n3907 VPWR.n3906 4.6505
R12407 VPWR.n3905 VPWR.n3904 4.6505
R12408 VPWR.n3903 VPWR.n3902 4.6505
R12409 VPWR.n3901 VPWR.n3900 4.6505
R12410 VPWR.n3899 VPWR.n3886 4.6505
R12411 VPWR.n3898 VPWR.n3897 4.6505
R12412 VPWR.n3896 VPWR.n3895 4.6505
R12413 VPWR.n3894 VPWR.n3893 4.6505
R12414 VPWR.n3892 VPWR.n3891 4.6505
R12415 VPWR.n3890 VPWR.n3889 4.6505
R12416 VPWR.n3808 VPWR.n3807 4.6505
R12417 VPWR.n3810 VPWR.n3809 4.6505
R12418 VPWR.n3812 VPWR.n3811 4.6505
R12419 VPWR.n3815 VPWR.n3780 4.6505
R12420 VPWR.n3865 VPWR.n3864 4.6505
R12421 VPWR.n3862 VPWR.n3861 4.6505
R12422 VPWR.n3860 VPWR.n3859 4.6505
R12423 VPWR.n3858 VPWR.n3857 4.6505
R12424 VPWR.n3856 VPWR.n3816 4.6505
R12425 VPWR.n3855 VPWR.n3854 4.6505
R12426 VPWR.n3853 VPWR.n3852 4.6505
R12427 VPWR.n3849 VPWR.n3817 4.6505
R12428 VPWR.n3848 VPWR.n3847 4.6505
R12429 VPWR.n3846 VPWR.n3845 4.6505
R12430 VPWR.n3844 VPWR.n3843 4.6505
R12431 VPWR.n3841 VPWR.n3840 4.6505
R12432 VPWR.n3839 VPWR.n3838 4.6505
R12433 VPWR.n3837 VPWR.n3836 4.6505
R12434 VPWR.n3835 VPWR.n3819 4.6505
R12435 VPWR.n3834 VPWR.n3833 4.6505
R12436 VPWR.n3868 VPWR.n3779 4.6505
R12437 VPWR.n3869 VPWR.n3868 4.6505
R12438 VPWR.n3871 VPWR.n3870 4.6505
R12439 VPWR.n3873 VPWR.n3872 4.6505
R12440 VPWR.n3875 VPWR.n3874 4.6505
R12441 VPWR.n3883 VPWR.n3882 4.6505
R12442 VPWR.n4384 VPWR.n4383 4.6505
R12443 VPWR.n4382 VPWR.n4381 4.6505
R12444 VPWR.n4380 VPWR.n4379 4.6505
R12445 VPWR.n4378 VPWR.n4377 4.6505
R12446 VPWR.n4376 VPWR.n4375 4.6505
R12447 VPWR.n4374 VPWR.n4373 4.6505
R12448 VPWR.n4370 VPWR.n4369 4.6505
R12449 VPWR.n4367 VPWR.n4366 4.6505
R12450 VPWR.n4363 VPWR.n435 4.6505
R12451 VPWR.n4361 VPWR.n4360 4.6505
R12452 VPWR.n4359 VPWR.n4358 4.6505
R12453 VPWR.n4357 VPWR.n1432 4.6505
R12454 VPWR.n4355 VPWR.n4354 4.6505
R12455 VPWR.n4348 VPWR.n4347 4.6505
R12456 VPWR.n4346 VPWR.n4345 4.6505
R12457 VPWR.n4344 VPWR.n4343 4.6505
R12458 VPWR.n4342 VPWR.n4341 4.6505
R12459 VPWR.n4340 VPWR.n4339 4.6505
R12460 VPWR.n4338 VPWR.n4337 4.6505
R12461 VPWR.n4335 VPWR.n4334 4.6505
R12462 VPWR.n4333 VPWR.n4332 4.6505
R12463 VPWR.n4331 VPWR.n4330 4.6505
R12464 VPWR.n4329 VPWR.n4328 4.6505
R12465 VPWR.n4327 VPWR.n4326 4.6505
R12466 VPWR.n1426 VPWR.n1425 4.6505
R12467 VPWR.n1330 VPWR.n1329 4.6505
R12468 VPWR.n1326 VPWR.n1325 4.6505
R12469 VPWR.n1322 VPWR.n443 4.6505
R12470 VPWR.n1319 VPWR.n1318 4.6505
R12471 VPWR.n1317 VPWR.n1316 4.6505
R12472 VPWR.n1314 VPWR.n1313 4.6505
R12473 VPWR.n1312 VPWR.n1311 4.6505
R12474 VPWR.n1233 VPWR.n1232 4.6505
R12475 VPWR.n1237 VPWR.n1236 4.6505
R12476 VPWR.n1239 VPWR.n1238 4.6505
R12477 VPWR.n1241 VPWR.n1240 4.6505
R12478 VPWR.n1244 VPWR.n1243 4.6505
R12479 VPWR.n1248 VPWR.n1247 4.6505
R12480 VPWR.n1250 VPWR.n1249 4.6505
R12481 VPWR.n1253 VPWR.n1252 4.6505
R12482 VPWR.n1256 VPWR.n1255 4.6505
R12483 VPWR.n1946 VPWR.n1945 4.6505
R12484 VPWR.n1959 VPWR.n1647 4.6505
R12485 VPWR.n1994 VPWR.n1993 4.6505
R12486 VPWR.n1996 VPWR.n1995 4.6505
R12487 VPWR.n2008 VPWR.n2007 4.6505
R12488 VPWR.n2009 VPWR.n1641 4.6505
R12489 VPWR.n1852 VPWR.n1851 4.6505
R12490 VPWR.n1855 VPWR.n1846 4.6505
R12491 VPWR.n1951 VPWR.n1950 4.6505
R12492 VPWR.n1956 VPWR.n1955 4.6505
R12493 VPWR.n1963 VPWR.n1962 4.6505
R12494 VPWR.n1965 VPWR.n1964 4.6505
R12495 VPWR.n1967 VPWR.n1966 4.6505
R12496 VPWR.n1969 VPWR.n1968 4.6505
R12497 VPWR.n1972 VPWR.n1971 4.6505
R12498 VPWR.n1974 VPWR.n1973 4.6505
R12499 VPWR.n1976 VPWR.n1975 4.6505
R12500 VPWR.n1978 VPWR.n1977 4.6505
R12501 VPWR.n1980 VPWR.n1979 4.6505
R12502 VPWR.n1982 VPWR.n1981 4.6505
R12503 VPWR.n1984 VPWR.n1983 4.6505
R12504 VPWR.n1986 VPWR.n1985 4.6505
R12505 VPWR.n2002 VPWR.n2001 4.6505
R12506 VPWR.n2006 VPWR.n2005 4.6505
R12507 VPWR.n4229 VPWR.n1474 4.6505
R12508 VPWR.n4220 VPWR.n1475 4.6505
R12509 VPWR.n4215 VPWR.n1478 4.6505
R12510 VPWR.n4204 VPWR.n4203 4.6505
R12511 VPWR.n4200 VPWR.n4199 4.6505
R12512 VPWR.n4195 VPWR.n1480 4.6505
R12513 VPWR.n4194 VPWR.n1482 4.6505
R12514 VPWR.n4193 VPWR.n1483 4.6505
R12515 VPWR.n4186 VPWR.n4185 4.6505
R12516 VPWR.n4173 VPWR.n1485 4.6505
R12517 VPWR.n4109 VPWR.n1522 4.6505
R12518 VPWR.n4103 VPWR.n1523 4.6505
R12519 VPWR.n4102 VPWR.n1524 4.6505
R12520 VPWR.n4101 VPWR.n1525 4.6505
R12521 VPWR.n4099 VPWR.n1527 4.6505
R12522 VPWR.n4098 VPWR.n1528 4.6505
R12523 VPWR.n4090 VPWR.n1529 4.6505
R12524 VPWR.n4087 VPWR.n1530 4.6505
R12525 VPWR.n4076 VPWR.n1535 4.6505
R12526 VPWR.n4005 VPWR.n4004 4.6505
R12527 VPWR.n4017 VPWR.n4016 4.6505
R12528 VPWR.n4015 VPWR.n4014 4.6505
R12529 VPWR.n4013 VPWR.n4012 4.6505
R12530 VPWR.n4011 VPWR.n4010 4.6505
R12531 VPWR.n4009 VPWR.n4008 4.6505
R12532 VPWR.n4007 VPWR.n4006 4.6505
R12533 VPWR.n4003 VPWR.n3996 4.6505
R12534 VPWR.n4000 VPWR.n3999 4.6505
R12535 VPWR.n4027 VPWR.n4026 4.6505
R12536 VPWR.n4025 VPWR.n4024 4.6505
R12537 VPWR.n4023 VPWR.n4022 4.6505
R12538 VPWR.n4021 VPWR.n4020 4.6505
R12539 VPWR.n4019 VPWR.n4018 4.6505
R12540 VPWR.n4119 VPWR.n4118 4.6505
R12541 VPWR.n4117 VPWR.n1520 4.6505
R12542 VPWR.n4116 VPWR.n4115 4.6505
R12543 VPWR.n4114 VPWR.n4113 4.6505
R12544 VPWR.n4112 VPWR.n4111 4.6505
R12545 VPWR.n4110 VPWR.n1521 4.6505
R12546 VPWR VPWR.n4108 4.6505
R12547 VPWR.n4107 VPWR.n4106 4.6505
R12548 VPWR.n4105 VPWR.n4104 4.6505
R12549 VPWR.n4096 VPWR.n4095 4.6505
R12550 VPWR.n4094 VPWR.n4093 4.6505
R12551 VPWR.n4092 VPWR.n4091 4.6505
R12552 VPWR.n4089 VPWR.n4088 4.6505
R12553 VPWR.n4086 VPWR.n4085 4.6505
R12554 VPWR.n4082 VPWR.n4081 4.6505
R12555 VPWR.n4078 VPWR.n4077 4.6505
R12556 VPWR.n4072 VPWR.n4071 4.6505
R12557 VPWR.n4070 VPWR.n1536 4.6505
R12558 VPWR.n4068 VPWR.n4067 4.6505
R12559 VPWR.n4231 VPWR.n4230 4.6505
R12560 VPWR.n4228 VPWR.n4227 4.6505
R12561 VPWR.n4226 VPWR.n4225 4.6505
R12562 VPWR.n4224 VPWR.n4223 4.6505
R12563 VPWR.n4222 VPWR.n4221 4.6505
R12564 VPWR.n4219 VPWR.n4218 4.6505
R12565 VPWR.n4217 VPWR.n1477 4.6505
R12566 VPWR.n4217 VPWR.n4216 4.6505
R12567 VPWR.n4214 VPWR.n4213 4.6505
R12568 VPWR.n4208 VPWR.n4207 4.6505
R12569 VPWR.n4206 VPWR.n4205 4.6505
R12570 VPWR.n4202 VPWR.n4201 4.6505
R12571 VPWR VPWR.n1479 4.6505
R12572 VPWR.n4198 VPWR.n4197 4.6505
R12573 VPWR.n4192 VPWR.n4191 4.6505
R12574 VPWR.n4190 VPWR.n4189 4.6505
R12575 VPWR.n4188 VPWR.n4187 4.6505
R12576 VPWR.n4184 VPWR.n4183 4.6505
R12577 VPWR.n4182 VPWR.n4181 4.6505
R12578 VPWR.n4178 VPWR.n4177 4.6505
R12579 VPWR.n4176 VPWR.n4175 4.6505
R12580 VPWR.n4174 VPWR.n1484 4.6505
R12581 VPWR.n2015 VPWR.n2014 4.6505
R12582 VPWR.n2013 VPWR.n2012 4.6505
R12583 VPWR.n2011 VPWR.n2010 4.6505
R12584 VPWR.n2000 VPWR.n1999 4.6505
R12585 VPWR.n1998 VPWR.n1997 4.6505
R12586 VPWR.n1992 VPWR.n1991 4.6505
R12587 VPWR.n1990 VPWR.n1989 4.6505
R12588 VPWR.n1988 VPWR.n1987 4.6505
R12589 VPWR.n1949 VPWR.n1648 4.6505
R12590 VPWR.n1948 VPWR.n1947 4.6505
R12591 VPWR.n1850 VPWR.n1847 4.6505
R12592 VPWR.n1854 VPWR.n1853 4.6505
R12593 VPWR.n1857 VPWR.n1856 4.6505
R12594 VPWR.n1859 VPWR.n1858 4.6505
R12595 VPWR.n1860 VPWR.n1845 4.6505
R12596 VPWR.n1862 VPWR.n1861 4.6505
R12597 VPWR.n1864 VPWR.n1844 4.6505
R12598 VPWR.n1866 VPWR.n1865 4.6505
R12599 VPWR.n1868 VPWR.n1867 4.6505
R12600 VPWR.n1872 VPWR.n1871 4.6505
R12601 VPWR.n1874 VPWR.n1843 4.6505
R12602 VPWR.n1876 VPWR.n1875 4.6505
R12603 VPWR.n1879 VPWR.n1878 4.6505
R12604 VPWR.n1882 VPWR.n1881 4.6505
R12605 VPWR.n3589 VPWR.n1578 4.6505
R12606 VPWR.n3597 VPWR.n3596 4.6505
R12607 VPWR.n3599 VPWR.n3598 4.6505
R12608 VPWR.n3600 VPWR.n1577 4.6505
R12609 VPWR.n3620 VPWR.n1576 4.6505
R12610 VPWR.n3622 VPWR.n3621 4.6505
R12611 VPWR.n1605 VPWR.n1593 4.6505
R12612 VPWR.n1595 VPWR.n1583 4.6505
R12613 VPWR.n2124 VPWR.n1584 4.6505
R12614 VPWR.n1791 VPWR.n1735 4.6505
R12615 VPWR.n1759 VPWR.n1737 4.6505
R12616 VPWR.n1758 VPWR.n1738 4.6505
R12617 VPWR.n1757 VPWR.n1740 4.6505
R12618 VPWR.n1755 VPWR.n1741 4.6505
R12619 VPWR.n1752 VPWR.n1751 4.6505
R12620 VPWR.n1746 VPWR.n1742 4.6505
R12621 VPWR.n1743 VPWR.n1586 4.6505
R12622 VPWR.n2118 VPWR.n1585 4.6505
R12623 VPWR.n2117 VPWR.n1587 4.6505
R12624 VPWR.n1677 VPWR.n1676 4.6505
R12625 VPWR.n1679 VPWR.n1678 4.6505
R12626 VPWR.n1681 VPWR.n1680 4.6505
R12627 VPWR.n1797 VPWR.n1796 4.6505
R12628 VPWR.n1793 VPWR.n1792 4.6505
R12629 VPWR.n1786 VPWR.n1785 4.6505
R12630 VPWR.n1784 VPWR.n1783 4.6505
R12631 VPWR.n1782 VPWR.n1781 4.6505
R12632 VPWR.n1780 VPWR.n1779 4.6505
R12633 VPWR.n1778 VPWR.n1777 4.6505
R12634 VPWR.n1775 VPWR.n1774 4.6505
R12635 VPWR.n1773 VPWR.n1772 4.6505
R12636 VPWR.n1771 VPWR.n1770 4.6505
R12637 VPWR.n1769 VPWR.n1768 4.6505
R12638 VPWR.n1767 VPWR.n1766 4.6505
R12639 VPWR.n1765 VPWR.n1764 4.6505
R12640 VPWR.n1763 VPWR.n1762 4.6505
R12641 VPWR.n2116 VPWR.n2115 4.6505
R12642 VPWR.n1629 VPWR.n1628 4.6505
R12643 VPWR.n1627 VPWR.n1626 4.6505
R12644 VPWR.n1625 VPWR.n1624 4.6505
R12645 VPWR.n1623 VPWR.n1622 4.6505
R12646 VPWR.n1621 VPWR.n1620 4.6505
R12647 VPWR.n1617 VPWR.n1616 4.6505
R12648 VPWR.n1615 VPWR.n1614 4.6505
R12649 VPWR.n1613 VPWR.n1612 4.6505
R12650 VPWR.n1611 VPWR.n1610 4.6505
R12651 VPWR.n1609 VPWR.n1608 4.6505
R12652 VPWR.n1597 VPWR.n1596 4.6505
R12653 VPWR.n2126 VPWR.n2125 4.6505
R12654 VPWR.n2128 VPWR.n2127 4.6505
R12655 VPWR.n2130 VPWR.n2129 4.6505
R12656 VPWR.n2132 VPWR.n2131 4.6505
R12657 VPWR.n2134 VPWR.n2133 4.6505
R12658 VPWR.n2137 VPWR.n2136 4.6505
R12659 VPWR.n2139 VPWR.n2138 4.6505
R12660 VPWR.n2140 VPWR.n1581 4.6505
R12661 VPWR.n2142 VPWR.n2141 4.6505
R12662 VPWR.n2147 VPWR.n2146 4.6505
R12663 VPWR.n2150 VPWR.n1580 4.6505
R12664 VPWR.n3587 VPWR.n3586 4.6505
R12665 VPWR.n3607 VPWR.n3606 4.6505
R12666 VPWR.n3623 VPWR.n1575 4.6505
R12667 VPWR.n3627 VPWR.n3626 4.6505
R12668 VPWR.n3629 VPWR.n3628 4.6505
R12669 VPWR.n3631 VPWR.n3630 4.6505
R12670 VPWR.n3634 VPWR.n1574 4.6505
R12671 VPWR.n3636 VPWR.n3635 4.6505
R12672 VPWR.n3651 VPWR.n3646 4.6505
R12673 VPWR.n3650 VPWR.n3647 4.6505
R12674 VPWR.n3682 VPWR.n3681 4.6505
R12675 VPWR.n3680 VPWR.n3679 4.6505
R12676 VPWR.n3678 VPWR.n3677 4.6505
R12677 VPWR.n3670 VPWR.n3669 4.6505
R12678 VPWR.n3668 VPWR.n3667 4.6505
R12679 VPWR.n3665 VPWR.n3664 4.6505
R12680 VPWR.n3663 VPWR.n3662 4.6505
R12681 VPWR.n3661 VPWR.n3644 4.6505
R12682 VPWR.n3660 VPWR.n3659 4.6505
R12683 VPWR.n3658 VPWR.n3657 4.6505
R12684 VPWR.n3656 VPWR.n3645 4.6505
R12685 VPWR.n3655 VPWR.n3654 4.6505
R12686 VPWR.n3653 VPWR.n3652 4.6505
R12687 VPWR.n3640 VPWR.n3639 4.6505
R12688 VPWR.n3638 VPWR.n3637 4.6505
R12689 VPWR.n3625 VPWR.n3624 4.6505
R12690 VPWR.n3619 VPWR.n3618 4.6505
R12691 VPWR.n3617 VPWR.n3616 4.6505
R12692 VPWR.n3615 VPWR.n3614 4.6505
R12693 VPWR.n3613 VPWR.n3612 4.6505
R12694 VPWR.n3611 VPWR.n3610 4.6505
R12695 VPWR.n3602 VPWR.n3601 4.6505
R12696 VPWR.n3594 VPWR.n3593 4.6505
R12697 VPWR.n3585 VPWR.n3584 4.6505
R12698 VPWR.n2156 VPWR.n2155 4.6505
R12699 VPWR.n2154 VPWR.n2153 4.6505
R12700 VPWR.n2152 VPWR.n2151 4.6505
R12701 VPWR.n1604 VPWR.n1603 4.6505
R12702 VPWR.n2120 VPWR.n2119 4.6505
R12703 VPWR.n1745 VPWR.n1744 4.6505
R12704 VPWR.n1748 VPWR.n1747 4.6505
R12705 VPWR.n1750 VPWR.n1749 4.6505
R12706 VPWR.n1754 VPWR.n1753 4.6505
R12707 VPWR.n1761 VPWR.n1760 4.6505
R12708 VPWR.n1788 VPWR.n1787 4.6505
R12709 VPWR.n1790 VPWR.n1789 4.6505
R12710 VPWR.n1683 VPWR.n1682 4.6505
R12711 VPWR.n1685 VPWR.n1684 4.6505
R12712 VPWR.n1687 VPWR.n1686 4.6505
R12713 VPWR.n1689 VPWR.n1688 4.6505
R12714 VPWR.n1691 VPWR.n1690 4.6505
R12715 VPWR.n1693 VPWR.n1692 4.6505
R12716 VPWR.n1695 VPWR.n1694 4.6505
R12717 VPWR.n1697 VPWR.n1696 4.6505
R12718 VPWR.n1700 VPWR.n1699 4.6505
R12719 VPWR.n1702 VPWR.n1701 4.6505
R12720 VPWR.n1704 VPWR.n1703 4.6505
R12721 VPWR.n1706 VPWR.n1705 4.6505
R12722 VPWR.n1708 VPWR.n1707 4.6505
R12723 VPWR.n2854 VPWR.n2853 4.6505
R12724 VPWR.n2928 VPWR.n2927 4.6505
R12725 VPWR.n2979 VPWR.n2795 4.6505
R12726 VPWR.n2978 VPWR.n2796 4.6505
R12727 VPWR.n2941 VPWR.n2801 4.6505
R12728 VPWR.n2938 VPWR.n2802 4.6505
R12729 VPWR.n2931 VPWR.n2803 4.6505
R12730 VPWR.n2819 VPWR.n2818 4.6505
R12731 VPWR.n2711 VPWR.n2691 4.6505
R12732 VPWR.n2715 VPWR.n2714 4.6505
R12733 VPWR.n2718 VPWR.n2717 4.6505
R12734 VPWR.n2975 VPWR.n2974 4.6505
R12735 VPWR.n2971 VPWR.n2970 4.6505
R12736 VPWR.n2969 VPWR.n2968 4.6505
R12737 VPWR.n2967 VPWR.n2966 4.6505
R12738 VPWR.n2965 VPWR.n2964 4.6505
R12739 VPWR.n2963 VPWR.n2962 4.6505
R12740 VPWR.n2961 VPWR.n2960 4.6505
R12741 VPWR.n2958 VPWR.n2957 4.6505
R12742 VPWR.n2956 VPWR.n2955 4.6505
R12743 VPWR.n2954 VPWR.n2953 4.6505
R12744 VPWR.n2952 VPWR.n2951 4.6505
R12745 VPWR.n2950 VPWR.n2949 4.6505
R12746 VPWR.n2948 VPWR.n2947 4.6505
R12747 VPWR.n2946 VPWR.n2945 4.6505
R12748 VPWR.n2860 VPWR.n2859 4.6505
R12749 VPWR.n2864 VPWR.n2863 4.6505
R12750 VPWR.n2866 VPWR.n2865 4.6505
R12751 VPWR.n2868 VPWR.n2867 4.6505
R12752 VPWR.n2870 VPWR.n2869 4.6505
R12753 VPWR.n2872 VPWR.n2871 4.6505
R12754 VPWR.n2874 VPWR.n2873 4.6505
R12755 VPWR.n2876 VPWR.n2875 4.6505
R12756 VPWR.n2879 VPWR.n2878 4.6505
R12757 VPWR.n2880 VPWR.n2807 4.6505
R12758 VPWR.n2882 VPWR.n2881 4.6505
R12759 VPWR.n2884 VPWR.n2883 4.6505
R12760 VPWR.n2886 VPWR.n2885 4.6505
R12761 VPWR.n2888 VPWR.n2887 4.6505
R12762 VPWR.n2890 VPWR.n2889 4.6505
R12763 VPWR.n2891 VPWR.n2806 4.6505
R12764 VPWR.n2924 VPWR.n2923 4.6505
R12765 VPWR.n2920 VPWR.n2919 4.6505
R12766 VPWR.n2918 VPWR.n2917 4.6505
R12767 VPWR.n2916 VPWR.n2915 4.6505
R12768 VPWR.n2914 VPWR.n2913 4.6505
R12769 VPWR.n2912 VPWR.n2911 4.6505
R12770 VPWR.n2910 VPWR.n2909 4.6505
R12771 VPWR.n2907 VPWR.n2906 4.6505
R12772 VPWR.n2905 VPWR.n2904 4.6505
R12773 VPWR.n2903 VPWR.n2902 4.6505
R12774 VPWR.n2901 VPWR.n2900 4.6505
R12775 VPWR.n2899 VPWR.n2898 4.6505
R12776 VPWR.n3440 VPWR.n2211 4.6505
R12777 VPWR.n2246 VPWR.n2245 4.6505
R12778 VPWR.n3435 VPWR.n2213 4.6505
R12779 VPWR.n2329 VPWR.n2328 4.6505
R12780 VPWR.n2324 VPWR.n2323 4.6505
R12781 VPWR.n2322 VPWR.n2321 4.6505
R12782 VPWR.n2320 VPWR.n2319 4.6505
R12783 VPWR.n2318 VPWR.n2317 4.6505
R12784 VPWR.n2316 VPWR.n2315 4.6505
R12785 VPWR.n2313 VPWR.n2312 4.6505
R12786 VPWR.n2311 VPWR.n2310 4.6505
R12787 VPWR.n2309 VPWR.n2308 4.6505
R12788 VPWR.n2306 VPWR.n2305 4.6505
R12789 VPWR.n2304 VPWR.n2303 4.6505
R12790 VPWR.n2302 VPWR.n2301 4.6505
R12791 VPWR.n2300 VPWR.n2299 4.6505
R12792 VPWR.n2298 VPWR.n2297 4.6505
R12793 VPWR.n2296 VPWR.n2295 4.6505
R12794 VPWR.n2294 VPWR.n2293 4.6505
R12795 VPWR.n3448 VPWR.n3447 4.6505
R12796 VPWR.n3446 VPWR.n3445 4.6505
R12797 VPWR.n3444 VPWR.n3443 4.6505
R12798 VPWR.n3442 VPWR.n3441 4.6505
R12799 VPWR.n2218 VPWR.n2212 4.6505
R12800 VPWR.n2220 VPWR.n2219 4.6505
R12801 VPWR.n2222 VPWR.n2221 4.6505
R12802 VPWR.n2224 VPWR.n2223 4.6505
R12803 VPWR.n2226 VPWR.n2225 4.6505
R12804 VPWR.n2228 VPWR.n2227 4.6505
R12805 VPWR.n2231 VPWR.n2230 4.6505
R12806 VPWR.n2233 VPWR.n2232 4.6505
R12807 VPWR.n2236 VPWR.n2235 4.6505
R12808 VPWR.n2239 VPWR.n2238 4.6505
R12809 VPWR.n2242 VPWR.n2217 4.6505
R12810 VPWR.n2244 VPWR.n2243 4.6505
R12811 VPWR.n2248 VPWR.n2247 4.6505
R12812 VPWR.n2250 VPWR.n2249 4.6505
R12813 VPWR.n2252 VPWR.n2251 4.6505
R12814 VPWR.n2255 VPWR.n2254 4.6505
R12815 VPWR.n2257 VPWR.n2256 4.6505
R12816 VPWR.n2259 VPWR.n2258 4.6505
R12817 VPWR.n2261 VPWR.n2260 4.6505
R12818 VPWR.n2263 VPWR.n2262 4.6505
R12819 VPWR.n2265 VPWR.n2264 4.6505
R12820 VPWR.n2267 VPWR.n2266 4.6505
R12821 VPWR.n2268 VPWR.n2214 4.6505
R12822 VPWR.n3437 VPWR.n3436 4.6505
R12823 VPWR.n3434 VPWR.n3433 4.6505
R12824 VPWR.n3432 VPWR.n3431 4.6505
R12825 VPWR.n3430 VPWR.n3429 4.6505
R12826 VPWR.n3428 VPWR.n3427 4.6505
R12827 VPWR.n3450 VPWR.n3449 4.6505
R12828 VPWR.n2895 VPWR.n2208 4.6505
R12829 VPWR.n2926 VPWR.n2925 4.6505
R12830 VPWR.n2856 VPWR.n2855 4.6505
R12831 VPWR.n2817 VPWR.n2816 4.6505
R12832 VPWR.n2815 VPWR.n2804 4.6505
R12833 VPWR.n2933 VPWR.n2932 4.6505
R12834 VPWR.n2935 VPWR.n2934 4.6505
R12835 VPWR.n2937 VPWR.n2936 4.6505
R12836 VPWR.n2940 VPWR.n2939 4.6505
R12837 VPWR.n2943 VPWR.n2942 4.6505
R12838 VPWR.n2977 VPWR.n2976 4.6505
R12839 VPWR.n2980 VPWR.n2794 4.6505
R12840 VPWR.n2982 VPWR.n2981 4.6505
R12841 VPWR.n2984 VPWR.n2983 4.6505
R12842 VPWR.n2985 VPWR.n2793 4.6505
R12843 VPWR.n2987 VPWR.n2986 4.6505
R12844 VPWR.n2989 VPWR.n2988 4.6505
R12845 VPWR.n2698 VPWR.n2697 4.6505
R12846 VPWR.n2699 VPWR.n2692 4.6505
R12847 VPWR.n2701 VPWR.n2700 4.6505
R12848 VPWR.n2703 VPWR.n2702 4.6505
R12849 VPWR.n2710 VPWR.n2709 4.6505
R12850 VPWR.n2713 VPWR.n2712 4.6505
R12851 VPWR.n2716 VPWR.n2690 4.6505
R12852 VPWR.n2720 VPWR.n2719 4.6505
R12853 VPWR.n2723 VPWR.n2722 4.6505
R12854 VPWR.n5015 VPWR.n5014 4.6505
R12855 VPWR.n5053 VPWR.n4981 4.6505
R12856 VPWR.n5037 VPWR.n5036 4.6505
R12857 VPWR.n6460 VPWR.n6459 4.6505
R12858 VPWR.n6462 VPWR.n6461 4.6505
R12859 VPWR.n6464 VPWR.n6463 4.6505
R12860 VPWR.n6467 VPWR.n6466 4.6505
R12861 VPWR.n6469 VPWR.n6468 4.6505
R12862 VPWR.n6471 VPWR.n6470 4.6505
R12863 VPWR.n6473 VPWR.n6472 4.6505
R12864 VPWR.n6474 VPWR.n5064 4.6505
R12865 VPWR.n6484 VPWR.n6483 4.6505
R12866 VPWR.n6487 VPWR.n6486 4.6505
R12867 VPWR.n6489 VPWR.n6488 4.6505
R12868 VPWR.n6492 VPWR.n6491 4.6505
R12869 VPWR.n6494 VPWR.n6493 4.6505
R12870 VPWR.n6500 VPWR.n6499 4.6505
R12871 VPWR.n6502 VPWR.n6501 4.6505
R12872 VPWR.n6505 VPWR.n6504 4.6505
R12873 VPWR.n6508 VPWR.n6507 4.6505
R12874 VPWR.n6510 VPWR.n6509 4.6505
R12875 VPWR.n6512 VPWR.n6511 4.6505
R12876 VPWR.n6514 VPWR.n6513 4.6505
R12877 VPWR.n6517 VPWR.n6516 4.6505
R12878 VPWR.n6519 VPWR.n6518 4.6505
R12879 VPWR.n6521 VPWR.n5060 4.6505
R12880 VPWR.n6523 VPWR.n6522 4.6505
R12881 VPWR.n6525 VPWR.n6524 4.6505
R12882 VPWR.n6528 VPWR.n6527 4.6505
R12883 VPWR.n4978 VPWR.n4977 4.6505
R12884 VPWR.n4983 VPWR.n4982 4.6505
R12885 VPWR.n4985 VPWR.n4984 4.6505
R12886 VPWR.n4987 VPWR.n4986 4.6505
R12887 VPWR.n4989 VPWR.n4988 4.6505
R12888 VPWR.n4992 VPWR.n4991 4.6505
R12889 VPWR.n4995 VPWR.n4994 4.6505
R12890 VPWR.n5000 VPWR.n4999 4.6505
R12891 VPWR.n5055 VPWR.n5054 4.6505
R12892 VPWR.n5052 VPWR.n5051 4.6505
R12893 VPWR.n5050 VPWR.n5049 4.6505
R12894 VPWR.n5048 VPWR.n5047 4.6505
R12895 VPWR.n5045 VPWR.n5044 4.6505
R12896 VPWR.n5043 VPWR.n5042 4.6505
R12897 VPWR.n5039 VPWR.n5038 4.6505
R12898 VPWR.n5033 VPWR.n5032 4.6505
R12899 VPWR.n5027 VPWR.n5026 4.6505
R12900 VPWR.n5025 VPWR.n5024 4.6505
R12901 VPWR.n7669 VPWR.n7664 4.6505
R12902 VPWR.n62 VPWR.n49 4.6505
R12903 VPWR.n60 VPWR.n51 4.6505
R12904 VPWR.n59 VPWR.n52 4.6505
R12905 VPWR.n56 VPWR.n53 4.6505
R12906 VPWR.n73 VPWR.n72 4.6505
R12907 VPWR.n71 VPWR.n70 4.6505
R12908 VPWR.n69 VPWR.n68 4.6505
R12909 VPWR.n67 VPWR.n66 4.6505
R12910 VPWR.n65 VPWR.n48 4.6505
R12911 VPWR.n64 VPWR.n63 4.6505
R12912 VPWR.n58 VPWR.n57 4.6505
R12913 VPWR.n80 VPWR.n79 4.6505
R12914 VPWR.n77 VPWR.n76 4.6505
R12915 VPWR.n75 VPWR.n74 4.6505
R12916 VPWR.n7671 VPWR.n7670 4.6505
R12917 VPWR.n7683 VPWR.n42 4.6505
R12918 VPWR.n7682 VPWR.n7681 4.6505
R12919 VPWR.n7680 VPWR.n7679 4.6505
R12920 VPWR.n7676 VPWR.n7675 4.6505
R12921 VPWR.n7674 VPWR.n7673 4.6505
R12922 VPWR.n7685 VPWR.n7684 4.6505
R12923 VPWR.n7687 VPWR.n7686 4.6505
R12924 VPWR.n7688 VPWR.n41 4.6505
R12925 VPWR.n7695 VPWR.n37 4.6505
R12926 VPWR.n7692 VPWR.n7691 4.6505
R12927 VPWR.n7690 VPWR.n7689 4.6505
R12928 VPWR.n7697 VPWR.n7696 4.6505
R12929 VPWR.n7699 VPWR.n7698 4.6505
R12930 VPWR.n7701 VPWR.n7700 4.6505
R12931 VPWR.n7711 VPWR.n7710 4.6505
R12932 VPWR.n7709 VPWR.n7708 4.6505
R12933 VPWR.n7705 VPWR.n7704 4.6505
R12934 VPWR.n7703 VPWR.n7702 4.6505
R12935 VPWR.n7713 VPWR.n7712 4.6505
R12936 VPWR.n7721 VPWR.n7720 4.6505
R12937 VPWR.n7719 VPWR.n31 4.6505
R12938 VPWR.n7718 VPWR.n7717 4.6505
R12939 VPWR.n7715 VPWR.n7714 4.6505
R12940 VPWR.n5023 VPWR.n5022 4.6505
R12941 VPWR.n5031 VPWR.n5030 4.6505
R12942 VPWR.n5035 VPWR.n5034 4.6505
R12943 VPWR.n5016 VPWR.n4980 4.6505
R12944 VPWR.n5013 VPWR.n5012 4.6505
R12945 VPWR.n5011 VPWR.n5010 4.6505
R12946 VPWR.n5009 VPWR.n5008 4.6505
R12947 VPWR.n5007 VPWR.n5006 4.6505
R12948 VPWR.n5002 VPWR.n5001 4.6505
R12949 VPWR.n4998 VPWR.n4997 4.6505
R12950 VPWR.n6476 VPWR.n6475 4.6505
R12951 VPWR.n6385 VPWR.n6384 4.6505
R12952 VPWR.n6387 VPWR.n6386 4.6505
R12953 VPWR.n6388 VPWR.n6379 4.6505
R12954 VPWR.n6390 VPWR.n6389 4.6505
R12955 VPWR.n6393 VPWR.n6392 4.6505
R12956 VPWR.n6395 VPWR.n6394 4.6505
R12957 VPWR.n6397 VPWR.n6396 4.6505
R12958 VPWR.n6398 VPWR.n6378 4.6505
R12959 VPWR.n6403 VPWR.n6402 4.6505
R12960 VPWR.n6408 VPWR.n6407 4.6505
R12961 VPWR.n2590 VPWR.n2578 4.6505
R12962 VPWR.n2591 VPWR.n2577 4.6505
R12963 VPWR.n2597 VPWR.n2596 4.6505
R12964 VPWR.n2605 VPWR.n2604 4.6505
R12965 VPWR.n2561 VPWR.n2559 4.6505
R12966 VPWR.n2533 VPWR.n2517 4.6505
R12967 VPWR.n2530 VPWR.n2518 4.6505
R12968 VPWR.n2523 VPWR.n2519 4.6505
R12969 VPWR.n2522 VPWR.n2520 4.6505
R12970 VPWR.n3114 VPWR.n2419 4.6505
R12971 VPWR.n3113 VPWR.n2421 4.6505
R12972 VPWR.n2438 VPWR.n2428 4.6505
R12973 VPWR.n3239 VPWR.n3229 4.6505
R12974 VPWR.n3287 VPWR.n3286 4.6505
R12975 VPWR.n3316 VPWR.n3301 4.6505
R12976 VPWR.n3319 VPWR.n3300 4.6505
R12977 VPWR.n3327 VPWR.n3326 4.6505
R12978 VPWR.n3325 VPWR.n3324 4.6505
R12979 VPWR.n3323 VPWR.n3322 4.6505
R12980 VPWR.n3315 VPWR.n3314 4.6505
R12981 VPWR.n3310 VPWR.n3309 4.6505
R12982 VPWR.n3318 VPWR.n3317 4.6505
R12983 VPWR.n3321 VPWR.n3320 4.6505
R12984 VPWR.n3220 VPWR.n3219 4.6505
R12985 VPWR.n3222 VPWR.n3221 4.6505
R12986 VPWR.n3224 VPWR.n3223 4.6505
R12987 VPWR.n3225 VPWR.n2385 4.6505
R12988 VPWR.n3283 VPWR.n3282 4.6505
R12989 VPWR.n3280 VPWR.n3279 4.6505
R12990 VPWR.n3268 VPWR.n3267 4.6505
R12991 VPWR.n3266 VPWR.n3265 4.6505
R12992 VPWR.n3262 VPWR.n3228 4.6505
R12993 VPWR.n3260 VPWR.n3259 4.6505
R12994 VPWR.n3258 VPWR.n3257 4.6505
R12995 VPWR.n3256 VPWR.n3255 4.6505
R12996 VPWR.n3253 VPWR.n3252 4.6505
R12997 VPWR.n3251 VPWR.n3250 4.6505
R12998 VPWR.n3249 VPWR.n3248 4.6505
R12999 VPWR.n3247 VPWR.n3246 4.6505
R13000 VPWR.n3245 VPWR.n3244 4.6505
R13001 VPWR.n3243 VPWR.n3242 4.6505
R13002 VPWR.n3241 VPWR.n3240 4.6505
R13003 VPWR.n3238 VPWR.n3237 4.6505
R13004 VPWR.n3236 VPWR.n3235 4.6505
R13005 VPWR.n3234 VPWR.n3233 4.6505
R13006 VPWR.n3232 VPWR.n3231 4.6505
R13007 VPWR.n3289 VPWR.n3288 4.6505
R13008 VPWR.n3291 VPWR.n3290 4.6505
R13009 VPWR.n3293 VPWR.n3292 4.6505
R13010 VPWR.n3295 VPWR.n3294 4.6505
R13011 VPWR.n3299 VPWR.n3298 4.6505
R13012 VPWR.n3329 VPWR.n3328 4.6505
R13013 VPWR.n3218 VPWR.n3217 4.6505
R13014 VPWR.n2437 VPWR.n2436 4.6505
R13015 VPWR.n2435 VPWR.n2429 4.6505
R13016 VPWR.n3120 VPWR.n3119 4.6505
R13017 VPWR.n3123 VPWR.n3122 4.6505
R13018 VPWR.n3125 VPWR.n3124 4.6505
R13019 VPWR.n3127 VPWR.n3126 4.6505
R13020 VPWR.n3129 VPWR.n3128 4.6505
R13021 VPWR.n3132 VPWR.n3131 4.6505
R13022 VPWR.n3134 VPWR.n3133 4.6505
R13023 VPWR.n3136 VPWR.n3135 4.6505
R13024 VPWR.n3143 VPWR.n3142 4.6505
R13025 VPWR.n3149 VPWR.n3148 4.6505
R13026 VPWR.n3151 VPWR.n3150 4.6505
R13027 VPWR.n2453 VPWR.n2452 4.6505
R13028 VPWR.n2451 VPWR.n2450 4.6505
R13029 VPWR.n2449 VPWR.n2425 4.6505
R13030 VPWR.n2446 VPWR.n2445 4.6505
R13031 VPWR.n2444 VPWR.n2443 4.6505
R13032 VPWR.n2442 VPWR.n2441 4.6505
R13033 VPWR.n2557 VPWR.n2507 4.6505
R13034 VPWR.n2556 VPWR.n2555 4.6505
R13035 VPWR.n2554 VPWR.n2553 4.6505
R13036 VPWR.n2552 VPWR.n2508 4.6505
R13037 VPWR.n2551 VPWR.n2550 4.6505
R13038 VPWR.n2549 VPWR.n2509 4.6505
R13039 VPWR.n2548 VPWR.n2547 4.6505
R13040 VPWR.n2546 VPWR.n2511 4.6505
R13041 VPWR.n2545 VPWR.n2544 4.6505
R13042 VPWR.n2543 VPWR.n2512 4.6505
R13043 VPWR.n2542 VPWR.n2541 4.6505
R13044 VPWR.n2540 VPWR.n2514 4.6505
R13045 VPWR.n2539 VPWR.n2538 4.6505
R13046 VPWR.n2537 VPWR.n2515 4.6505
R13047 VPWR.n2536 VPWR.n2535 4.6505
R13048 VPWR.n2534 VPWR.n2516 4.6505
R13049 VPWR.n2532 VPWR.n2531 4.6505
R13050 VPWR.n2529 VPWR.n2528 4.6505
R13051 VPWR.n2527 VPWR.n2526 4.6505
R13052 VPWR.n2525 VPWR.n2524 4.6505
R13053 VPWR.n2521 VPWR.n2420 4.6505
R13054 VPWR.n3116 VPWR.n3115 4.6505
R13055 VPWR.n3112 VPWR.n3111 4.6505
R13056 VPWR.n2575 VPWR.n2574 4.6505
R13057 VPWR.n2573 VPWR.n2572 4.6505
R13058 VPWR.n2571 VPWR.n2570 4.6505
R13059 VPWR.n2569 VPWR.n2568 4.6505
R13060 VPWR.n2567 VPWR.n2566 4.6505
R13061 VPWR.n2565 VPWR.n2564 4.6505
R13062 VPWR.n2563 VPWR.n2562 4.6505
R13063 VPWR.n2583 VPWR.n2580 4.6505
R13064 VPWR.n2586 VPWR.n2585 4.6505
R13065 VPWR.n2587 VPWR.n2579 4.6505
R13066 VPWR.n2589 VPWR.n2588 4.6505
R13067 VPWR.n2593 VPWR.n2592 4.6505
R13068 VPWR.n2595 VPWR.n2594 4.6505
R13069 VPWR.n2599 VPWR.n2598 4.6505
R13070 VPWR.n2601 VPWR.n2600 4.6505
R13071 VPWR.n2609 VPWR.n2608 4.6505
R13072 VPWR.n2611 VPWR.n2610 4.6505
R13073 VPWR.n2613 VPWR.n2612 4.6505
R13074 VPWR.n5933 VPWR.n5930 4.6505
R13075 VPWR.n5841 VPWR.n5840 4.6505
R13076 VPWR.n5845 VPWR.n5844 4.6505
R13077 VPWR.n5886 VPWR.n5885 4.6505
R13078 VPWR.n5893 VPWR.n5892 4.6505
R13079 VPWR.n5900 VPWR.n5899 4.6505
R13080 VPWR.n6042 VPWR.n5904 4.6505
R13081 VPWR.n6173 VPWR.n5821 4.6505
R13082 VPWR.n6158 VPWR.n5822 4.6505
R13083 VPWR.n6155 VPWR.n5823 4.6505
R13084 VPWR.n6130 VPWR.n6049 4.6505
R13085 VPWR.n6127 VPWR.n6050 4.6505
R13086 VPWR.n6124 VPWR.n6051 4.6505
R13087 VPWR.n6112 VPWR.n6056 4.6505
R13088 VPWR.n6277 VPWR.n5732 4.6505
R13089 VPWR.n6262 VPWR.n5733 4.6505
R13090 VPWR.n6259 VPWR.n5735 4.6505
R13091 VPWR.n6228 VPWR.n6227 4.6505
R13092 VPWR.n6224 VPWR.n5746 4.6505
R13093 VPWR.n6289 VPWR.n6284 4.6505
R13094 VPWR.n6292 VPWR.n6283 4.6505
R13095 VPWR.n6295 VPWR.n6282 4.6505
R13096 VPWR.n6301 VPWR.n6280 4.6505
R13097 VPWR.n6304 VPWR.n6279 4.6505
R13098 VPWR.n6276 VPWR.n6275 4.6505
R13099 VPWR.n6274 VPWR.n6273 4.6505
R13100 VPWR.n6272 VPWR.n6271 4.6505
R13101 VPWR.n6270 VPWR.n6269 4.6505
R13102 VPWR.n6268 VPWR.n6267 4.6505
R13103 VPWR.n6266 VPWR.n6265 4.6505
R13104 VPWR.n6264 VPWR.n6263 4.6505
R13105 VPWR.n6254 VPWR.n5736 4.6505
R13106 VPWR.n6253 VPWR.n6252 4.6505
R13107 VPWR.n6251 VPWR.n5737 4.6505
R13108 VPWR.n6250 VPWR.n6249 4.6505
R13109 VPWR.n6248 VPWR.n5739 4.6505
R13110 VPWR.n6247 VPWR.n6246 4.6505
R13111 VPWR.n6245 VPWR.n5740 4.6505
R13112 VPWR.n6244 VPWR.n6243 4.6505
R13113 VPWR.n6242 VPWR.n6241 4.6505
R13114 VPWR.n6240 VPWR.n5742 4.6505
R13115 VPWR.n6239 VPWR.n6238 4.6505
R13116 VPWR.n6237 VPWR.n5743 4.6505
R13117 VPWR.n6236 VPWR.n6235 4.6505
R13118 VPWR.n6234 VPWR.n5744 4.6505
R13119 VPWR.n6233 VPWR.n6232 4.6505
R13120 VPWR.n6231 VPWR.n5745 4.6505
R13121 VPWR.n6219 VPWR.n6218 4.6505
R13122 VPWR.n6214 VPWR.n6213 4.6505
R13123 VPWR.n6172 VPWR.n6171 4.6505
R13124 VPWR.n6170 VPWR.n6169 4.6505
R13125 VPWR.n6168 VPWR.n6167 4.6505
R13126 VPWR.n6166 VPWR.n6165 4.6505
R13127 VPWR.n6164 VPWR.n6163 4.6505
R13128 VPWR.n6162 VPWR.n6161 4.6505
R13129 VPWR.n6152 VPWR.n5824 4.6505
R13130 VPWR.n6151 VPWR.n6150 4.6505
R13131 VPWR.n5827 VPWR.n5825 4.6505
R13132 VPWR.n6145 VPWR.n6144 4.6505
R13133 VPWR.n6143 VPWR.n5828 4.6505
R13134 VPWR.n6142 VPWR.n6141 4.6505
R13135 VPWR.n6140 VPWR.n5829 4.6505
R13136 VPWR.n6139 VPWR 4.6505
R13137 VPWR.n6138 VPWR.n6046 4.6505
R13138 VPWR.n6137 VPWR.n6136 4.6505
R13139 VPWR.n6134 VPWR.n6047 4.6505
R13140 VPWR.n6133 VPWR.n6132 4.6505
R13141 VPWR.n6131 VPWR.n6048 4.6505
R13142 VPWR.n6119 VPWR.n6052 4.6505
R13143 VPWR.n6118 VPWR.n6117 4.6505
R13144 VPWR.n6116 VPWR.n6053 4.6505
R13145 VPWR.n6115 VPWR.n6114 4.6505
R13146 VPWR.n5848 VPWR.n5830 4.6505
R13147 VPWR.n5855 VPWR.n5854 4.6505
R13148 VPWR.n5859 VPWR.n5858 4.6505
R13149 VPWR.n5861 VPWR.n5860 4.6505
R13150 VPWR.n5863 VPWR.n5862 4.6505
R13151 VPWR.n5865 VPWR.n5864 4.6505
R13152 VPWR.n5867 VPWR.n5866 4.6505
R13153 VPWR.n5870 VPWR.n5869 4.6505
R13154 VPWR.n5872 VPWR.n5871 4.6505
R13155 VPWR.n5874 VPWR.n5873 4.6505
R13156 VPWR.n5876 VPWR.n5875 4.6505
R13157 VPWR.n5878 VPWR.n5877 4.6505
R13158 VPWR.n5880 VPWR.n5879 4.6505
R13159 VPWR.n5882 VPWR.n5881 4.6505
R13160 VPWR.n5884 VPWR.n5883 4.6505
R13161 VPWR.n5903 VPWR.n5831 4.6505
R13162 VPWR.n6028 VPWR.n6027 4.6505
R13163 VPWR.n6031 VPWR.n6030 4.6505
R13164 VPWR.n6036 VPWR.n6035 4.6505
R13165 VPWR.n6039 VPWR.n6038 4.6505
R13166 VPWR.n6041 VPWR.n6040 4.6505
R13167 VPWR.n5895 VPWR.n5894 4.6505
R13168 VPWR.n5891 VPWR.n5890 4.6505
R13169 VPWR.n5889 VPWR.n5832 4.6505
R13170 VPWR.n5888 VPWR.n5887 4.6505
R13171 VPWR.n5850 VPWR.n5849 4.6505
R13172 VPWR.n5847 VPWR.n5846 4.6505
R13173 VPWR.n5843 VPWR.n5842 4.6505
R13174 VPWR.n5839 VPWR.n5838 4.6505
R13175 VPWR.n6111 VPWR.n6110 4.6505
R13176 VPWR.n6113 VPWR.n6055 4.6505
R13177 VPWR.n6121 VPWR.n6120 4.6505
R13178 VPWR.n6123 VPWR.n6122 4.6505
R13179 VPWR.n6126 VPWR.n6125 4.6505
R13180 VPWR.n6129 VPWR.n6128 4.6505
R13181 VPWR.n6154 VPWR.n6153 4.6505
R13182 VPWR.n6157 VPWR.n6156 4.6505
R13183 VPWR.n6160 VPWR.n6159 4.6505
R13184 VPWR.n6216 VPWR.n6215 4.6505
R13185 VPWR.n6217 VPWR.n5747 4.6505
R13186 VPWR.n6221 VPWR.n6220 4.6505
R13187 VPWR.n6223 VPWR.n6222 4.6505
R13188 VPWR.n6226 VPWR.n6225 4.6505
R13189 VPWR.n6230 VPWR.n6229 4.6505
R13190 VPWR.n6256 VPWR.n6255 4.6505
R13191 VPWR.n6258 VPWR.n6257 4.6505
R13192 VPWR.n6261 VPWR.n6260 4.6505
R13193 VPWR.n6288 VPWR.n6287 4.6505
R13194 VPWR.n6291 VPWR.n6290 4.6505
R13195 VPWR.n6294 VPWR.n6293 4.6505
R13196 VPWR.n6297 VPWR.n6296 4.6505
R13197 VPWR.n6298 VPWR.n6281 4.6505
R13198 VPWR.n6300 VPWR.n6299 4.6505
R13199 VPWR.n6303 VPWR.n6302 4.6505
R13200 VPWR.n6308 VPWR.n6307 4.6505
R13201 VPWR.n6312 VPWR.n6311 4.6505
R13202 VPWR.n6314 VPWR.n6313 4.6505
R13203 VPWR.n6316 VPWR.n6315 4.6505
R13204 VPWR.n5958 VPWR.n5957 4.6505
R13205 VPWR.n5956 VPWR.n5921 4.6505
R13206 VPWR.n5955 VPWR.n5954 4.6505
R13207 VPWR.n5953 VPWR.n5922 4.6505
R13208 VPWR.n5952 VPWR.n5951 4.6505
R13209 VPWR.n5950 VPWR.n5923 4.6505
R13210 VPWR.n5949 VPWR.n5948 4.6505
R13211 VPWR.n5947 VPWR.n5924 4.6505
R13212 VPWR.n5946 VPWR.n5945 4.6505
R13213 VPWR.n5944 VPWR.n5925 4.6505
R13214 VPWR.n5943 VPWR.n5942 4.6505
R13215 VPWR.n5941 VPWR.n5926 4.6505
R13216 VPWR.n5940 VPWR.n5927 4.6505
R13217 VPWR.n5939 VPWR.n5938 4.6505
R13218 VPWR.n5937 VPWR.n5928 4.6505
R13219 VPWR.n5936 VPWR.n5935 4.6505
R13220 VPWR.n5934 VPWR.n5929 4.6505
R13221 VPWR.n1717 VPWR.n1716 4.64677
R13222 VPWR.n1876 VPWR.n1843 4.59011
R13223 VPWR.n1728 VPWR.n1727 4.57445
R13224 VPWR.n7620 VPWR.n7619 4.57427
R13225 VPWR.n6749 VPWR.n6748 4.57427
R13226 VPWR.n6692 VPWR.n6691 4.57427
R13227 VPWR.n6612 VPWR.n6580 4.57427
R13228 VPWR.n6918 VPWR.n4928 4.57427
R13229 VPWR.n6791 VPWR.n6790 4.57427
R13230 VPWR.n7195 VPWR.n7194 4.57427
R13231 VPWR.n7163 VPWR.n7162 4.57427
R13232 VPWR.n7022 VPWR.n7021 4.57427
R13233 VPWR.n868 VPWR.n867 4.57427
R13234 VPWR.n839 VPWR.n838 4.57427
R13235 VPWR.n743 VPWR.n742 4.57427
R13236 VPWR.n701 VPWR.n700 4.57427
R13237 VPWR.n4549 VPWR.n4548 4.57427
R13238 VPWR.n4598 VPWR.n4597 4.57427
R13239 VPWR.n4461 VPWR.n4460 4.57427
R13240 VPWR.n1115 VPWR.n1114 4.57427
R13241 VPWR.n4324 VPWR.n4323 4.57427
R13242 VPWR.n3795 VPWR.n3794 4.57427
R13243 VPWR.n428 VPWR.n427 4.57427
R13244 VPWR.n1402 VPWR.n1381 4.57427
R13245 VPWR.n4171 VPWR.n1487 4.57427
R13246 VPWR.n1513 VPWR.n1512 4.57427
R13247 VPWR.n4233 VPWR.n1462 4.57427
R13248 VPWR.n1460 VPWR.n1459 4.57427
R13249 VPWR.n3570 VPWR.n3569 4.57427
R13250 VPWR.n3548 VPWR.n3547 4.57427
R13251 VPWR.n2077 VPWR.n2076 4.57427
R13252 VPWR.n2099 VPWR.n2098 4.57427
R13253 VPWR.n3486 VPWR.n2210 4.57427
R13254 VPWR.n3465 VPWR.n3464 4.57427
R13255 VPWR.n2834 VPWR.n2833 4.57427
R13256 VPWR.n2851 VPWR.n2850 4.57427
R13257 VPWR.n7782 VPWR.n26 4.57427
R13258 VPWR.n6544 VPWR.n6543 4.57427
R13259 VPWR.n6566 VPWR.n6565 4.57427
R13260 VPWR.n7741 VPWR.n7740 4.57427
R13261 VPWR.n3169 VPWR.n3168 4.57427
R13262 VPWR.n3188 VPWR.n3187 4.57427
R13263 VPWR.n3075 VPWR.n3074 4.57427
R13264 VPWR.n3097 VPWR.n3096 4.57427
R13265 VPWR.n6199 VPWR.n6198 4.57427
R13266 VPWR.n6177 VPWR.n6176 4.57427
R13267 VPWR.n6109 VPWR.n6108 4.57427
R13268 VPWR.n6091 VPWR.n6090 4.57427
R13269 VPWR.n4785 VPWR.n4784 4.57412
R13270 VPWR.n6869 VPWR.n6868 4.57282
R13271 VPWR.n7216 VPWR.n7215 4.57282
R13272 VPWR.n887 VPWR.n886 4.57282
R13273 VPWR.n3804 VPWR.n3803 4.57282
R13274 VPWR.n5835 VPWR.n5834 4.57282
R13275 VPWR.n6701 VPWR.n6700 4.57249
R13276 VPWR.n1421 VPWR.n1420 4.57249
R13277 VPWR.n6908 VPWR.n6907 4.57152
R13278 VPWR.n6241 VPWR.n5741 4.54926
R13279 VPWR.n6176 VPWR.n6175 4.54926
R13280 VPWR.n3074 VPWR.n3073 4.54926
R13281 VPWR.n3131 VPWR.n3130 4.54926
R13282 VPWR.n6392 VPWR.n6391 4.54926
R13283 VPWR.n6719 VPWR.n6718 4.54926
R13284 VPWR.n7567 VPWR.n7527 4.54926
R13285 VPWR.n7542 VPWR.n7541 4.54926
R13286 VPWR.n6642 VPWR.n6641 4.54926
R13287 VPWR.n5177 VPWR.n5176 4.54926
R13288 VPWR.n6936 VPWR.n6935 4.54926
R13289 VPWR.n5516 VPWR.n5515 4.54926
R13290 VPWR.n5452 VPWR.n5451 4.54926
R13291 VPWR.n5258 VPWR.n5257 4.54926
R13292 VPWR.n5282 VPWR.n5281 4.54926
R13293 VPWR.n4671 VPWR.n4670 4.54926
R13294 VPWR.n4650 VPWR.n4649 4.54926
R13295 VPWR.n1169 VPWR.n1168 4.54926
R13296 VPWR.n1193 VPWR.n1192 4.54926
R13297 VPWR.n1043 VPWR.n1017 4.54926
R13298 VPWR.n4337 VPWR.n4336 4.54926
R13299 VPWR.n1316 VPWR.n1315 4.54926
R13300 VPWR.n1971 VPWR.n1970 4.54926
R13301 VPWR.n2136 VPWR.n2135 4.54926
R13302 VPWR.n1777 VPWR.n1776 4.54926
R13303 VPWR.n2254 VPWR.n2253 4.54926
R13304 VPWR.n2878 VPWR.n2877 4.54926
R13305 VPWR.n2960 VPWR.n2959 4.54926
R13306 VPWR.n2230 VPWR.n2229 4.54926
R13307 VPWR.n2909 VPWR.n2908 4.54926
R13308 VPWR.n5869 VPWR.n5868 4.54926
R13309 VPWR.n7068 VPWR.n7067 4.53667
R13310 VPWR.n740 VPWR.n739 4.53667
R13311 VPWR.n517 VPWR.n516 4.50829
R13312 VPWR.n5991 VPWR.n5959 4.50829
R13313 VPWR.n236 VPWR.n204 4.50828
R13314 VPWR.n7474 VPWR.n7473 4.50828
R13315 VPWR.n7364 VPWR.n7363 4.50828
R13316 VPWR.n4833 VPWR.n4832 4.50828
R13317 VPWR VPWR.n5397 4.5005
R13318 VPWR.n4779 VPWR.n4778 4.5005
R13319 VPWR.n566 VPWR.n565 4.5005
R13320 VPWR VPWR.n1889 4.5005
R13321 VPWR.n2023 VPWR.n1640 4.5005
R13322 VPWR.n3415 VPWR.n3414 4.5005
R13323 VPWR.n2993 VPWR.n2689 4.5005
R13324 VPWR.n2604 VPWR 4.3525
R13325 VPWR.n7408 VPWR.n7407 4.31796
R13326 VPWR.n700 VPWR.n696 4.31796
R13327 VPWR.n2443 VPWR.n2442 4.29549
R13328 VPWR.n1681 VPWR 4.26717
R13329 VPWR.n434 VPWR 4.18512
R13330 VPWR.n6145 VPWR.n5828 4.18384
R13331 VPWR.n683 VPWR.n682 4.16558
R13332 VPWR.n7194 VPWR.n7193 4.16558
R13333 VPWR.n2435 VPWR.n2430 4.12386
R13334 VPWR.n7723 VPWR.n7722 4.12386
R13335 VPWR.n5105 VPWR.n5091 4.12386
R13336 VPWR.n6799 VPWR.n277 4.12386
R13337 VPWR.n7233 VPWR.n7232 4.12386
R13338 VPWR.n4869 VPWR.n4868 4.12386
R13339 VPWR.n5238 VPWR.n5237 4.12386
R13340 VPWR.n646 VPWR.n645 4.12386
R13341 VPWR.n643 VPWR.n642 4.12386
R13342 VPWR.n357 VPWR.n337 4.12386
R13343 VPWR.n375 VPWR.n374 4.12386
R13344 VPWR.n4487 VPWR.n4486 4.12386
R13345 VPWR.n1226 VPWR.n1225 4.12386
R13346 VPWR.n4066 VPWR.n4065 4.12386
R13347 VPWR.n4084 VPWR.n1531 4.12386
R13348 VPWR.n1733 VPWR.n1731 4.12386
R13349 VPWR.n1570 VPWR.n1569 4.12386
R13350 VPWR.n743 VPWR.n604 4.11479
R13351 VPWR.n6691 VPWR.n6690 4.06399
R13352 VPWR.n700 VPWR.n699 4.06399
R13353 VPWR.n6090 VPWR.n6089 4.0132
R13354 VPWR.n1255 VPWR.n1254 4.0132
R13355 VPWR.n1881 VPWR.n1880 4.0132
R13356 VPWR.n2722 VPWR.n2721 4.0132
R13357 VPWR.n79 VPWR.n78 3.9624
R13358 VPWR.n3681 VPWR.n3642 3.9624
R13359 VPWR.n3619 VPWR 3.86082
R13360 VPWR.n6612 VPWR 3.81002
R13361 VPWR VPWR.n582 3.81002
R13362 VPWR VPWR.n1027 3.81002
R13363 VPWR.n1868 VPWR 3.81002
R13364 VPWR.n5401 VPWR 3.75923
R13365 VPWR.n902 VPWR 3.72662
R13366 VPWR.n5477 VPWR.n5476 3.53501
R13367 VPWR.n7669 VPWR.n7668 3.53475
R13368 VPWR.n6305 VPWR.n6278 3.50526
R13369 VPWR.n2602 VPWR.n2576 3.50526
R13370 VPWR.n5897 VPWR.n5896 3.50526
R13371 VPWR.n2425 VPWR.n2424 3.47425
R13372 VPWR.n5553 VPWR.n5552 3.47425
R13373 VPWR.n7114 VPWR.n7113 3.47425
R13374 VPWR.n7115 VPWR.n7114 3.47425
R13375 VPWR.n369 VPWR.n368 3.47425
R13376 VPWR.n4662 VPWR.n369 3.47425
R13377 VPWR.n393 VPWR.n392 3.47425
R13378 VPWR.n394 VPWR.n393 3.47425
R13379 VPWR.n2144 VPWR.n2143 3.47425
R13380 VPWR.n3677 VPWR.n3676 3.47425
R13381 VPWR.n2216 VPWR.n2215 3.47425
R13382 VPWR.n2217 VPWR.n2216 3.47425
R13383 VPWR.n3675 VPWR.n3673 3.43649
R13384 VPWR.n5676 VPWR.n5675 3.4105
R13385 VPWR.n7606 VPWR.n7605 3.4105
R13386 VPWR.n236 VPWR.n235 3.4105
R13387 VPWR.n6659 VPWR.n6658 3.4105
R13388 VPWR.n6665 VPWR.n6664 3.4105
R13389 VPWR.n6873 VPWR.n6872 3.4105
R13390 VPWR.n6901 VPWR.n6900 3.4105
R13391 VPWR.n6789 VPWR.n4931 3.4105
R13392 VPWR.n7475 VPWR.n7474 3.4105
R13393 VPWR.n5396 VPWR.n5393 3.4105
R13394 VPWR.n7210 VPWR.n7209 3.4105
R13395 VPWR.n7150 VPWR.n7149 3.4105
R13396 VPWR.n7165 VPWR.n7164 3.4105
R13397 VPWR VPWR.n7179 3.4105
R13398 VPWR.n7365 VPWR.n7364 3.4105
R13399 VPWR.n7315 VPWR.n7314 3.4105
R13400 VPWR.n7375 VPWR.n7374 3.4105
R13401 VPWR.n5328 VPWR.n5327 3.4105
R13402 VPWR.n5298 VPWR.n5297 3.4105
R13403 VPWR.n7023 VPWR.n7015 3.4105
R13404 VPWR.n563 VPWR.n562 3.4105
R13405 VPWR.n883 VPWR.n882 3.4105
R13406 VPWR.n832 VPWR.n831 3.4105
R13407 VPWR.n841 VPWR.n840 3.4105
R13408 VPWR.n4834 VPWR.n4833 3.4105
R13409 VPWR.n4761 VPWR.n318 3.4105
R13410 VPWR.n975 VPWR.n974 3.4105
R13411 VPWR.n722 VPWR.n721 3.4105
R13412 VPWR.n737 VPWR.n605 3.4105
R13413 VPWR.n4457 VPWR.n4456 3.4105
R13414 VPWR.n1296 VPWR.n1295 3.4105
R13415 VPWR.n4317 VPWR.n4316 3.4105
R13416 VPWR.n3786 VPWR.n3785 3.4105
R13417 VPWR.n1417 VPWR.n1416 3.4105
R13418 VPWR.n4129 VPWR.n4128 3.4105
R13419 VPWR.n1888 VPWR.n1885 3.4105
R13420 VPWR.n2029 VPWR.n2028 3.4105
R13421 VPWR.n4249 VPWR.n4248 3.4105
R13422 VPWR.n1820 VPWR.n1819 3.4105
R13423 VPWR.n2105 VPWR.n2104 3.4105
R13424 VPWR.n2781 VPWR.n2780 3.4105
R13425 VPWR.n2352 VPWR.n2351 3.4105
R13426 VPWR.n2995 VPWR.n2994 3.4105
R13427 VPWR.n7733 VPWR.n7732 3.4105
R13428 VPWR.n6427 VPWR.n6426 3.4105
R13429 VPWR.n3208 VPWR.n3207 3.4105
R13430 VPWR.n5991 VPWR.n5990 3.4105
R13431 VPWR.n7807 VPWR.n7806 3.4105
R13432 VPWR.n2550 VPWR.n2510 3.37141
R13433 VPWR.n1344 VPWR.n1342 3.37141
R13434 VPWR.n7086 VPWR.n7081 3.31258
R13435 VPWR.n51 VPWR 3.29747
R13436 VPWR.n181 VPWR 3.29747
R13437 VPWR.n7119 VPWR 3.29747
R13438 VPWR.n3313 VPWR.n3312 3.28365
R13439 VPWR.n3312 VPWR.n3302 3.273
R13440 VPWR.n7085 VPWR.n7082 3.23
R13441 VPWR.n7021 VPWR.n7020 3.20994
R13442 VPWR.n3309 VPWR.n3302 3.20311
R13443 VPWR.n7670 VPWR.n7669 3.2005
R13444 VPWR.n7085 VPWR.n7084 3.2005
R13445 VPWR.n6146 VPWR.n5827 3.16454
R13446 VPWR.n5305 VPWR.n5304 3.09667
R13447 VPWR.n859 VPWR.n822 3.06326
R13448 VPWR.n7598 VPWR.n7597 3.05891
R13449 VPWR.n2513 VPWR.n2511 3.01588
R13450 VPWR.n3227 VPWR.n3226 3.01588
R13451 VPWR.n3298 VPWR.n3297 3.01588
R13452 VPWR.n7722 VPWR.n7721 3.00117
R13453 VPWR.n7521 VPWR.n7520 3.00117
R13454 VPWR.n7407 VPWR.n277 3.00117
R13455 VPWR.n7075 VPWR.n4868 3.00117
R13456 VPWR.n354 VPWR.n337 3.00117
R13457 VPWR.n4488 VPWR.n4487 3.00117
R13458 VPWR.n1796 VPWR.n1733 3.00117
R13459 VPWR.n7626 VPWR.n7625 3.0005
R13460 VPWR.n6681 VPWR.n6680 3.0005
R13461 VPWR.n7489 VPWR.n7488 3.0005
R13462 VPWR.n5404 VPWR.n5403 3.0005
R13463 VPWR.n7178 VPWR.n7140 3.0005
R13464 VPWR.n7040 VPWR.n7039 3.0005
R13465 VPWR.n4848 VPWR.n4847 3.0005
R13466 VPWR.n856 VPWR.n855 3.0005
R13467 VPWR.n554 VPWR.n553 3.0005
R13468 VPWR.n711 VPWR.n710 3.0005
R13469 VPWR.n4592 VPWR.n4591 3.0005
R13470 VPWR.n1109 VPWR.n1108 3.0005
R13471 VPWR.n3789 VPWR.n3788 3.0005
R13472 VPWR.n4155 VPWR.n4154 3.0005
R13473 VPWR.n1924 VPWR.n1923 3.0005
R13474 VPWR.n2341 VPWR.n2340 3.0005
R13475 VPWR.n7770 VPWR.n7769 3.0005
R13476 VPWR.n6059 VPWR.n6058 2.99733
R13477 VPWR.n6691 VPWR.n6687 2.99733
R13478 VPWR.n3187 VPWR.n3186 2.98339
R13479 VPWR.n6407 VPWR.n6406 2.98339
R13480 VPWR.n5115 VPWR.n5114 2.98339
R13481 VPWR.n6343 VPWR.n6342 2.96248
R13482 VPWR.n2640 VPWR.n2639 2.96248
R13483 VPWR.n1332 VPWR.n1331 2.96248
R13484 VPWR.n3922 VPWR.n3921 2.94563
R13485 VPWR.n2328 VPWR.n2327 2.94563
R13486 VPWR.n6150 VPWR.n6149 2.76904
R13487 VPWR.n2544 VPWR.n2513 2.64665
R13488 VPWR.n3255 VPWR.n3254 2.64665
R13489 VPWR.n3298 VPWR.n3296 2.64665
R13490 VPWR.n6466 VPWR.n6465 2.64665
R13491 VPWR.n6491 VPWR.n6490 2.64665
R13492 VPWR.n6516 VPWR.n6515 2.64665
R13493 VPWR.n6543 VPWR.n6542 2.64665
R13494 VPWR.n4977 VPWR.n4976 2.64665
R13495 VPWR.n5151 VPWR.n5150 2.64665
R13496 VPWR.n5197 VPWR.n5196 2.64665
R13497 VPWR.n5568 VPWR.n5567 2.64665
R13498 VPWR.n1352 VPWR.n1351 2.64665
R13499 VPWR.n2308 VPWR.n2307 2.64665
R13500 VPWR.n3275 VPWR.n3274 2.50603
R13501 VPWR.n7229 VPWR.n7228 2.4386
R13502 VPWR.n3605 VPWR.n3604 2.4386
R13503 VPWR.n4511 VPWR.n4510 2.4268
R13504 VPWR.n5826 VPWR.n5824 2.37353
R13505 VPWR.n3321 VPWR 2.36572
R13506 VPWR.n4864 VPWR 2.36572
R13507 VPWR.n6252 VPWR.n5738 2.33701
R13508 VPWR.n6135 VPWR.n6134 2.33701
R13509 VPWR.n6117 VPWR.n6054 2.33701
R13510 VPWR.n2584 VPWR.n2583 2.33701
R13511 VPWR.n2585 VPWR.n2584 2.33701
R13512 VPWR.n47 VPWR.n46 2.33701
R13513 VPWR.n39 VPWR.n38 2.33701
R13514 VPWR.n35 VPWR.n34 2.33701
R13515 VPWR.n5021 VPWR.n5020 2.33701
R13516 VPWR.n7438 VPWR.n7437 2.33701
R13517 VPWR.n4924 VPWR.n4923 2.33701
R13518 VPWR.n6862 VPWR.n6861 2.33701
R13519 VPWR.n7336 VPWR.n7335 2.33701
R13520 VPWR.n5349 VPWR.n5348 2.33701
R13521 VPWR.n320 VPWR.n319 2.33701
R13522 VPWR.n904 VPWR.n903 2.33701
R13523 VPWR.n808 VPWR.n807 2.33701
R13524 VPWR.n509 VPWR.n508 2.33701
R13525 VPWR.n4500 VPWR.n4499 2.33701
R13526 VPWR.n3995 VPWR.n3994 2.33701
R13527 VPWR.n1643 VPWR.n1642 2.33701
R13528 VPWR.n1644 VPWR.n1643 2.33701
R13529 VPWR.n1955 VPWR.n1952 2.33701
R13530 VPWR.n1864 VPWR.n1863 2.33701
R13531 VPWR.n1870 VPWR.n1869 2.33701
R13532 VPWR.n1878 VPWR.n1877 2.33701
R13533 VPWR.n1602 VPWR.n1601 2.33701
R13534 VPWR.n2798 VPWR.n2797 2.33701
R13535 VPWR.n2707 VPWR.n2706 2.33701
R13536 VPWR.n5853 VPWR.n5852 2.33701
R13537 VPWR.n5738 VPWR.n5736 2.33701
R13538 VPWR.n6136 VPWR.n6135 2.33701
R13539 VPWR.n6054 VPWR.n6052 2.33701
R13540 VPWR.n7674 VPWR.n46 2.33701
R13541 VPWR.n7709 VPWR.n35 2.33701
R13542 VPWR.n5020 VPWR.n5019 2.33701
R13543 VPWR.n7464 VPWR.n7438 2.33701
R13544 VPWR.n6863 VPWR.n6862 2.33701
R13545 VPWR.n7337 VPWR.n7336 2.33701
R13546 VPWR.n903 VPWR.n902 2.33701
R13547 VPWR.n897 VPWR.n896 2.33701
R13548 VPWR.n896 VPWR.n895 2.33701
R13549 VPWR.n809 VPWR.n808 2.33701
R13550 VPWR.n4499 VPWR.n4498 2.33701
R13551 VPWR.n3996 VPWR.n3995 2.33701
R13552 VPWR.n1952 VPWR.n1951 2.33701
R13553 VPWR.n1863 VPWR.n1862 2.33701
R13554 VPWR.n1871 VPWR.n1870 2.33701
R13555 VPWR.n1877 VPWR.n1876 2.33701
R13556 VPWR.n1603 VPWR.n1602 2.33701
R13557 VPWR.n2893 VPWR.n2892 2.33701
R13558 VPWR.n5854 VPWR.n5853 2.33701
R13559 VPWR.n5379 VPWR.n5378 2.337
R13560 VPWR.n756 VPWR.n755 2.32777
R13561 VPWR.n755 VPWR.n754 2.32777
R13562 VPWR.n5164 VPWR.n5163 2.29662
R13563 VPWR.n5105 VPWR.n5104 2.29662
R13564 VPWR.n5106 VPWR.n5105 2.29662
R13565 VPWR.n5557 VPWR.n5466 2.29662
R13566 VPWR.n5498 VPWR.n5467 2.29662
R13567 VPWR.n3825 VPWR.n3778 2.29662
R13568 VPWR.n4084 VPWR.n1532 2.29662
R13569 VPWR.n4084 VPWR.n4083 2.29662
R13570 VPWR.n2126 VPWR.n1582 2.29662
R13571 VPWR.n2897 VPWR.n2896 2.29662
R13572 VPWR.n6478 VPWR.n6477 2.29662
R13573 VPWR.n3281 VPWR.n2384 2.29662
R13574 VPWR.n3264 VPWR.n3263 2.29662
R13575 VPWR.n3139 VPWR.n3138 2.29662
R13576 VPWR.n7525 VPWR.n160 2.29643
R13577 VPWR.n5317 VPWR.n5316 2.29643
R13578 VPWR.n7071 VPWR.n4870 2.29643
R13579 VPWR.n3827 VPWR.n3826 2.29643
R13580 VPWR.n4180 VPWR.n4179 2.29643
R13581 VPWR.n4097 VPWR.n1528 2.29643
R13582 VPWR.n1594 VPWR.n1583 2.29643
R13583 VPWR.n2561 VPWR.n2558 2.29643
R13584 VPWR.n5478 VPWR.n5477 2.28218
R13585 VPWR.n7036 VPWR.n4872 2.28218
R13586 VPWR.n4241 VPWR.n1461 2.28206
R13587 VPWR.n2842 VPWR.n2814 2.28206
R13588 VPWR.n7774 VPWR.n7773 2.28198
R13589 VPWR.n7299 VPWR.n289 2.28171
R13590 VPWR.n4066 VPWR.n4064 2.28171
R13591 VPWR.n569 VPWR.n470 2.28167
R13592 VPWR.n7669 VPWR.n103 2.28159
R13593 VPWR.n2415 VPWR.n2414 2.27488
R13594 VPWR.n5005 VPWR.n5004 2.27488
R13595 VPWR.n816 VPWR.n601 2.25932
R13596 VPWR.n1569 VPWR.n1568 2.23927
R13597 VPWR.n5047 VPWR.n5046 2.23542
R13598 VPWR.n6828 VPWR.n6827 2.23542
R13599 VPWR.n7228 VPWR.n7227 2.23542
R13600 VPWR.n3604 VPWR.n3603 2.23542
R13601 VPWR.n7668 VPWR.n7667 2.10848
R13602 VPWR.n5123 VPWR.n5122 1.93767
R13603 VPWR.n5621 VPWR.n5620 1.93767
R13604 VPWR.n5387 VPWR.n5386 1.93767
R13605 VPWR.n1054 VPWR.n1053 1.93767
R13606 VPWR.n1277 VPWR.n1276 1.93767
R13607 VPWR.n1897 VPWR.n1896 1.93767
R13608 VPWR.n1715 VPWR.n1714 1.93767
R13609 VPWR.n2745 VPWR.n2744 1.93767
R13610 VPWR.n6446 VPWR.n6445 1.93767
R13611 VPWR.n4724 VPWR.n4723 1.93767
R13612 VPWR.n4047 VPWR.n4046 1.93767
R13613 VPWR.n2361 VPWR.n2360 1.93767
R13614 VPWR VPWR.n2152 1.90463
R13615 VPWR.n6506 VPWR.n6505 1.88295
R13616 VPWR VPWR.n4459 1.88285
R13617 VPWR.n6481 VPWR.n6480 1.86464
R13618 VPWR.n5159 VPWR.n5145 1.86427
R13619 VPWR.n5555 VPWR.n5554 1.85065
R13620 VPWR.n3168 VPWR.n3167 1.85065
R13621 VPWR.n3882 VPWR.n3881 1.85065
R13622 VPWR.n2424 VPWR.n2423 1.81289
R13623 VPWR.n6919 VPWR.n4927 1.80429
R13624 VPWR.n7197 VPWR.n7196 1.80429
R13625 VPWR.n870 VPWR.n869 1.80429
R13626 VPWR.n4551 VPWR.n4550 1.80429
R13627 VPWR.n4325 VPWR.n1437 1.80429
R13628 VPWR.n4172 VPWR.n1486 1.80429
R13629 VPWR.n3163 VPWR.n3162 1.80429
R13630 VPWR.n7784 VPWR.n7783 1.80429
R13631 VPWR.n6747 VPWR.n4936 1.80429
R13632 VPWR.n3545 VPWR.n3544 1.80429
R13633 VPWR.n3488 VPWR.n3487 1.80429
R13634 VPWR.n6085 VPWR.n6084 1.80429
R13635 VPWR.n2075 VPWR.n2074 1.80353
R13636 VPWR.n6568 VPWR.n6567 1.80353
R13637 VPWR.n2852 VPWR.n2813 1.80353
R13638 VPWR.n6174 VPWR.n5820 1.80353
R13639 VPWR.n6992 VPWR.n6991 1.80347
R13640 VPWR.n4462 VPWR.n399 1.80347
R13641 VPWR.n4389 VPWR.n4388 1.80347
R13642 VPWR.n4232 VPWR.n1473 1.80347
R13643 VPWR.n3072 VPWR.n3071 1.80347
R13644 VPWR.n2555 VPWR 1.79885
R13645 VPWR.n5001 VPWR 1.79885
R13646 VPWR.n5165 VPWR 1.79885
R13647 VPWR.n5251 VPWR 1.79885
R13648 VPWR.n2146 VPWR.n2145 1.73737
R13649 VPWR.n2145 VPWR.n2144 1.73737
R13650 VPWR.n5378 VPWR.n5377 1.67669
R13651 VPWR.n2423 VPWR.n2422 1.66186
R13652 VPWR.n7105 VPWR.n7104 1.66186
R13653 VPWR.n3882 VPWR.n3876 1.66186
R13654 VPWR.n3675 VPWR.n3674 1.63881
R13655 VPWR.n3148 VPWR.n3147 1.6241
R13656 VPWR.n7593 VPWR.n7592 1.6241
R13657 VPWR.n5554 VPWR.n5553 1.6241
R13658 VPWR.n5541 VPWR.n5540 1.6241
R13659 VPWR.n7102 VPWR.n7101 1.6241
R13660 VPWR.n4512 VPWR.n4511 1.6241
R13661 VPWR.n4517 VPWR.n4516 1.6241
R13662 VPWR.n3667 VPWR.n3666 1.6241
R13663 VPWR.n6507 VPWR.n6506 1.62167
R13664 VPWR.n6483 VPWR.n6481 1.5112
R13665 VPWR.n5160 VPWR.n5159 1.51057
R13666 VPWR.n5095 VPWR.n5094 1.50646
R13667 VPWR.n5430 VPWR.n5429 1.50646
R13668 VPWR.n5353 VPWR.n5352 1.50646
R13669 VPWR.n480 VPWR.n479 1.50646
R13670 VPWR.n1022 VPWR.n1021 1.50646
R13671 VPWR.n1229 VPWR.n1228 1.50646
R13672 VPWR.n1849 VPWR.n1848 1.50646
R13673 VPWR.n1675 VPWR.n1674 1.50646
R13674 VPWR.n2694 VPWR.n2693 1.50646
R13675 VPWR.n6381 VPWR.n6380 1.50646
R13676 VPWR.n2582 VPWR.n2581 1.50646
R13677 VPWR.n7218 VPWR.n7217 1.50638
R13678 VPWR.n5187 VPWR.n5143 1.49961
R13679 VPWR.n6704 VPWR.n4941 1.49961
R13680 VPWR.n4197 VPWR.n4196 1.49961
R13681 VPWR.n1798 VPWR.n1731 1.49961
R13682 VPWR.n5004 VPWR.n5003 1.49961
R13683 VPWR.n2435 VPWR.n2434 1.49961
R13684 VPWR.n3121 VPWR.n2417 1.49961
R13685 VPWR.n3137 VPWR.n2415 1.49961
R13686 VPWR.n2944 VPWR.n2800 1.49956
R13687 VPWR.n5096 VPWR.n5093 1.49932
R13688 VPWR.n175 VPWR.n174 1.49932
R13689 VPWR.n6822 VPWR.n6820 1.49932
R13690 VPWR.n7445 VPWR.n7444 1.49932
R13691 VPWR.n5363 VPWR.n5347 1.49932
R13692 VPWR.n7272 VPWR.n7271 1.49932
R13693 VPWR.n7245 VPWR.n7233 1.49932
R13694 VPWR.n7329 VPWR.n7328 1.49932
R13695 VPWR.n677 VPWR.n639 1.49932
R13696 VPWR.n487 VPWR.n477 1.49932
R13697 VPWR.n892 VPWR.n583 1.49932
R13698 VPWR.n4801 VPWR.n4800 1.49932
R13699 VPWR.n1023 VPWR.n1020 1.49932
R13700 VPWR.n343 VPWR.n342 1.49932
R13701 VPWR.n4385 VPWR.n431 1.49932
R13702 VPWR.n3888 VPWR.n3887 1.49932
R13703 VPWR.n1961 VPWR.n1960 1.49932
R13704 VPWR.n3998 VPWR.n3997 1.49932
R13705 VPWR.n3588 VPWR.n1579 1.49932
R13706 VPWR.n3591 VPWR.n3590 1.49932
R13707 VPWR.n3641 VPWR.n1570 1.49932
R13708 VPWR.n3649 VPWR.n3648 1.49932
R13709 VPWR.n2696 VPWR.n2695 1.49932
R13710 VPWR.n2292 VPWR.n2291 1.49932
R13711 VPWR.n6383 VPWR.n6382 1.49932
R13712 VPWR.n61 VPWR.n50 1.49932
R13713 VPWR.n55 VPWR.n54 1.49932
R13714 VPWR.n3306 VPWR.n3305 1.49932
R13715 VPWR.n7086 VPWR.n7085 1.47352
R13716 VPWR.n497 VPWR.n496 1.41226
R13717 VPWR.n3881 VPWR.n3880 1.35979
R13718 VPWR.n7297 VPWR.n7296 1.35461
R13719 VPWR.n3951 VPWR.n3950 1.35461
R13720 VPWR.n3425 VPWR.n2269 1.35461
R13721 VPWR.n2649 VPWR.n2648 1.35461
R13722 VPWR.n7662 VPWR.n7661 1.35461
R13723 VPWR.n7519 VPWR.n7518 1.35461
R13724 VPWR.n3708 VPWR.n3707 1.35461
R13725 VPWR.n3364 VPWR.n3363 1.35461
R13726 VPWR.n6026 VPWR.n6025 1.35461
R13727 VPWR.n5662 VPWR.n5661 1.35459
R13728 VPWR.n5586 VPWR.n5585 1.35459
R13729 VPWR.n1308 VPWR.n444 1.35459
R13730 VPWR.n1944 VPWR.n1649 1.35459
R13731 VPWR.n1812 VPWR.n1811 1.35459
R13732 VPWR.n6458 VPWR.n6457 1.35459
R13733 VPWR.n6352 VPWR.n6351 1.35459
R13734 VPWR.n3279 VPWR.n3278 1.30773
R13735 VPWR.n3277 VPWR.n3276 1.30773
R13736 VPWR.n3167 VPWR.n3166 1.24652
R13737 VPWR.n3278 VPWR.n3277 1.1988
R13738 VPWR.n3276 VPWR.n3275 1.1988
R13739 VPWR.n6287 VPWR.n6286 1.16875
R13740 VPWR.n6306 VPWR.n6305 1.16875
R13741 VPWR.n6109 VPWR.n6059 1.16875
R13742 VPWR.n2603 VPWR.n2602 1.16875
R13743 VPWR.n5898 VPWR.n5897 1.16875
R13744 VPWR.n5931 VPWR.n5930 1.16875
R13745 VPWR.n7656 VPWR.n113 1.13896
R13746 VPWR.n7513 VPWR.n239 1.13896
R13747 VPWR.n6602 VPWR.n6601 1.13896
R13748 VPWR.n6996 VPWR.n6995 1.13896
R13749 VPWR.n7062 VPWR.n7061 1.13896
R13750 VPWR.n734 VPWR.n733 1.13896
R13751 VPWR.n4444 VPWR.n4443 1.13896
R13752 VPWR.n4393 VPWR.n4392 1.13896
R13753 VPWR.n1470 VPWR.n1453 1.13896
R13754 VPWR.n3716 VPWR.n1549 1.13896
R13755 VPWR.n2068 VPWR.n2067 1.13896
R13756 VPWR.n3540 VPWR.n3539 1.13896
R13757 VPWR.n1903 VPWR.n1902 1.13896
R13758 VPWR.n1283 VPWR.n1282 1.13896
R13759 VPWR.n1049 VPWR.n1008 1.13896
R13760 VPWR.n512 VPWR.n460 1.13896
R13761 VPWR.n5382 VPWR.n5211 1.13896
R13762 VPWR.n5627 VPWR.n5626 1.13896
R13763 VPWR.n5118 VPWR.n5073 1.13896
R13764 VPWR.n1710 VPWR.n1655 1.13896
R13765 VPWR.n6452 VPWR.n6451 1.13896
R13766 VPWR.n3372 VPWR.n2377 1.13896
R13767 VPWR.n7514 VPWR.n7513 1.13896
R13768 VPWR.n3716 VPWR.n3715 1.13896
R13769 VPWR.n7657 VPWR.n7656 1.13896
R13770 VPWR.n7610 VPWR.n131 1.13885
R13771 VPWR.n7433 VPWR.n256 1.13885
R13772 VPWR.n6877 VPWR.n6876 1.13885
R13773 VPWR.n7323 VPWR.n284 1.13885
R13774 VPWR.n7204 VPWR.n7203 1.13885
R13775 VPWR.n4793 VPWR.n301 1.13885
R13776 VPWR.n877 VPWR.n876 1.13885
R13777 VPWR.n4728 VPWR.n4727 1.13885
R13778 VPWR.n4570 VPWR.n4569 1.13885
R13779 VPWR.n3773 VPWR.n3772 1.13885
R13780 VPWR.n4298 VPWR.n4297 1.13885
R13781 VPWR.n4051 VPWR.n4050 1.13885
R13782 VPWR.n4133 VPWR.n4132 1.13885
R13783 VPWR.n4959 VPWR.n4958 1.13885
R13784 VPWR.n3068 VPWR.n3067 1.13885
R13785 VPWR.n5794 VPWR.n5793 1.13885
R13786 VPWR.n3202 VPWR.n3201 1.13885
R13787 VPWR.n7796 VPWR.n7795 1.13885
R13788 VPWR.n5716 VPWR.n5715 1.13885
R13789 VPWR.n2679 VPWR.n2652 1.13885
R13790 VPWR.n112 VPWR.n111 1.13717
R13791 VPWR.n238 VPWR.n237 1.13717
R13792 VPWR.n6766 VPWR.n6765 1.13717
R13793 VPWR.n5660 VPWR.n5659 1.13717
R13794 VPWR.n6599 VPWR.n6598 1.13717
R13795 VPWR.n7401 VPWR.n7400 1.13717
R13796 VPWR.n6777 VPWR.n6776 1.13717
R13797 VPWR.n5584 VPWR.n5583 1.13717
R13798 VPWR.n7006 VPWR.n7005 1.13717
R13799 VPWR.n7295 VPWR.n7294 1.13717
R13800 VPWR.n7201 VPWR.n7200 1.13717
R13801 VPWR.n5229 VPWR.n5228 1.13717
R13802 VPWR.n5296 VPWR.n5295 1.13717
R13803 VPWR.n4760 VPWR.n4759 1.13717
R13804 VPWR.n874 VPWR.n873 1.13717
R13805 VPWR.n977 VPWR.n976 1.13717
R13806 VPWR.n623 VPWR.n622 1.13717
R13807 VPWR.n4683 VPWR.n4682 1.13717
R13808 VPWR.n4555 VPWR.n4554 1.13717
R13809 VPWR.n1209 VPWR.n1208 1.13717
R13810 VPWR.n4432 VPWR.n4431 1.13717
R13811 VPWR.n3956 VPWR.n3955 1.13717
R13812 VPWR.n4283 VPWR.n4282 1.13717
R13813 VPWR.n1223 VPWR.n1222 1.13717
R13814 VPWR.n1415 VPWR.n1414 1.13717
R13815 VPWR.n4055 VPWR.n4054 1.13717
R13816 VPWR.n1501 VPWR.n1500 1.13717
R13817 VPWR.n1841 VPWR.n1840 1.13717
R13818 VPWR.n2034 VPWR.n2033 1.13717
R13819 VPWR.n1810 VPWR.n1809 1.13717
R13820 VPWR.n3537 VPWR.n3536 1.13717
R13821 VPWR.n2073 VPWR.n2072 1.13717
R13822 VPWR.n6570 VPWR.n6569 1.13717
R13823 VPWR.n2278 VPWR.n2277 1.13717
R13824 VPWR.n2997 VPWR.n2996 1.13717
R13825 VPWR.n2812 VPWR.n2811 1.13717
R13826 VPWR.n2470 VPWR.n2469 1.13717
R13827 VPWR.n5819 VPWR.n5818 1.13717
R13828 VPWR.n5760 VPWR.n5759 1.13717
R13829 VPWR.n5782 VPWR.n5781 1.13717
R13830 VPWR.n3070 VPWR.n3069 1.13717
R13831 VPWR.n3065 VPWR.n3062 1.13717
R13832 VPWR.n3016 VPWR.n3014 1.13717
R13833 VPWR.n3034 VPWR.n3033 1.13717
R13834 VPWR.n4966 VPWR.n4965 1.13717
R13835 VPWR.n5812 VPWR.n5811 1.13717
R13836 VPWR.n1472 VPWR.n1471 1.13717
R13837 VPWR.n4263 VPWR.n4262 1.13717
R13838 VPWR.n4269 VPWR.n4255 1.13717
R13839 VPWR.n4391 VPWR.n4390 1.13717
R13840 VPWR.n4413 VPWR.n4412 1.13717
R13841 VPWR.n4419 VPWR.n4405 1.13717
R13842 VPWR.n4442 VPWR.n4441 1.13717
R13843 VPWR.n4453 VPWR.n4452 1.13717
R13844 VPWR.n4446 VPWR.n416 1.13717
R13845 VPWR.n736 VPWR.n735 1.13717
R13846 VPWR.n725 VPWR.n724 1.13717
R13847 VPWR.n731 VPWR.n633 1.13717
R13848 VPWR.n7064 VPWR.n7063 1.13717
R13849 VPWR.n7053 VPWR.n7052 1.13717
R13850 VPWR.n7059 VPWR.n7045 1.13717
R13851 VPWR.n6994 VPWR.n6993 1.13717
R13852 VPWR.n4901 VPWR.n4900 1.13717
R13853 VPWR.n4907 VPWR.n4893 1.13717
R13854 VPWR.n6604 VPWR.n6603 1.13717
R13855 VPWR.n6668 VPWR.n6667 1.13717
R13856 VPWR.n6675 VPWR.n6674 1.13717
R13857 VPWR.n2047 VPWR.n2046 1.13717
R13858 VPWR.n2063 VPWR.n2062 1.13717
R13859 VPWR.n2066 VPWR.n1591 1.13717
R13860 VPWR.n4957 VPWR.n4955 1.13717
R13861 VPWR.n2482 VPWR.n2481 1.13717
R13862 VPWR.n3046 VPWR.n3045 1.13717
R13863 VPWR.n5792 VPWR.n5790 1.13717
R13864 VPWR.n3161 VPWR.n3160 1.13717
R13865 VPWR.n7803 VPWR.n7802 1.13717
R13866 VPWR.n3204 VPWR.n3203 1.13717
R13867 VPWR.n3199 VPWR.n3196 1.13717
R13868 VPWR.n3492 VPWR.n3491 1.13717
R13869 VPWR.n2181 VPWR.n2180 1.13717
R13870 VPWR.n2187 VPWR.n2173 1.13717
R13871 VPWR.n4149 VPWR.n4148 1.13717
R13872 VPWR.n4142 VPWR.n4141 1.13717
R13873 VPWR.n4131 VPWR.n4130 1.13717
R13874 VPWR.n4314 VPWR.n4313 1.13717
R13875 VPWR.n4307 VPWR.n4306 1.13717
R13876 VPWR.n4296 VPWR.n4295 1.13717
R13877 VPWR.n4586 VPWR.n4585 1.13717
R13878 VPWR.n4579 VPWR.n4578 1.13717
R13879 VPWR.n4568 VPWR.n4567 1.13717
R13880 VPWR.n850 VPWR.n849 1.13717
R13881 VPWR.n843 VPWR.n842 1.13717
R13882 VPWR.n879 VPWR.n878 1.13717
R13883 VPWR.n7174 VPWR.n7173 1.13717
R13884 VPWR.n7167 VPWR.n7166 1.13717
R13885 VPWR.n7206 VPWR.n7205 1.13717
R13886 VPWR.n6890 VPWR.n6889 1.13717
R13887 VPWR.n6897 VPWR.n6896 1.13717
R13888 VPWR.n6875 VPWR.n6874 1.13717
R13889 VPWR.n7631 VPWR.n7630 1.13717
R13890 VPWR.n141 VPWR.n140 1.13717
R13891 VPWR.n7612 VPWR.n7611 1.13717
R13892 VPWR.n3543 VPWR.n3542 1.13717
R13893 VPWR.n3502 VPWR.n3501 1.13717
R13894 VPWR.n2204 VPWR.n2203 1.13717
R13895 VPWR.n3520 VPWR.n3519 1.13717
R13896 VPWR.n2403 VPWR.n2402 1.13717
R13897 VPWR.n7734 VPWR.n24 1.13717
R13898 VPWR.n7756 VPWR.n7755 1.13717
R13899 VPWR.n7764 VPWR.n7763 1.13717
R13900 VPWR.n7794 VPWR.n7790 1.13717
R13901 VPWR.n6456 VPWR.n6455 1.13717
R13902 VPWR.n6354 VPWR.n6353 1.13717
R13903 VPWR.n2775 VPWR.n2774 1.13717
R13904 VPWR.n2737 VPWR.n2736 1.13717
R13905 VPWR.n6424 VPWR.n6423 1.13717
R13906 VPWR.n6376 VPWR.n6370 1.13717
R13907 VPWR.n1911 VPWR.n1910 1.13717
R13908 VPWR.n1918 VPWR.n1917 1.13717
R13909 VPWR.n1901 VPWR.n1899 1.13717
R13910 VPWR.n1292 VPWR.n1291 1.13717
R13911 VPWR.n1285 VPWR.n459 1.13717
R13912 VPWR.n1281 VPWR.n1279 1.13717
R13913 VPWR.n1000 VPWR.n999 1.13717
R13914 VPWR.n1006 VPWR.n993 1.13717
R13915 VPWR.n1052 VPWR.n1051 1.13717
R13916 VPWR.n541 VPWR.n474 1.13717
R13917 VPWR.n548 VPWR.n547 1.13717
R13918 VPWR.n515 VPWR.n514 1.13717
R13919 VPWR.n5415 VPWR.n5414 1.13717
R13920 VPWR.n5421 VPWR.n5408 1.13717
R13921 VPWR.n5385 VPWR.n5384 1.13717
R13922 VPWR.n5647 VPWR.n5646 1.13717
R13923 VPWR.n5653 VPWR.n5640 1.13717
R13924 VPWR.n5625 VPWR.n5623 1.13717
R13925 VPWR.n5678 VPWR.n5677 1.13717
R13926 VPWR.n5684 VPWR.n5086 1.13717
R13927 VPWR.n5121 VPWR.n5120 1.13717
R13928 VPWR.n1822 VPWR.n1821 1.13717
R13929 VPWR.n1828 VPWR.n1668 1.13717
R13930 VPWR.n1713 VPWR.n1712 1.13717
R13931 VPWR.n6450 VPWR.n6448 1.13717
R13932 VPWR.n2743 VPWR.n2742 1.13717
R13933 VPWR.n5722 VPWR.n5721 1.13717
R13934 VPWR.n5708 VPWR.n5707 1.13717
R13935 VPWR.n5714 VPWR.n5712 1.13717
R13936 VPWR.n2498 VPWR.n2495 1.13717
R13937 VPWR.n2659 VPWR.n2658 1.13717
R13938 VPWR.n2651 VPWR.n2650 1.13717
R13939 VPWR.n2676 VPWR.n2675 1.13717
R13940 VPWR.n3370 VPWR.n3369 1.13717
R13941 VPWR.n3411 VPWR.n3410 1.13717
R13942 VPWR.n2349 VPWR.n2287 1.13717
R13943 VPWR.n2363 VPWR.n2362 1.13717
R13944 VPWR.n3714 VPWR.n3712 1.13717
R13945 VPWR.n3985 VPWR.n3984 1.13717
R13946 VPWR.n3969 VPWR.n3968 1.13717
R13947 VPWR.n4049 VPWR.n4048 1.13717
R13948 VPWR.n3761 VPWR.n3760 1.13717
R13949 VPWR.n3745 VPWR.n3744 1.13717
R13950 VPWR.n3771 VPWR.n3770 1.13717
R13951 VPWR.n4753 VPWR.n4752 1.13717
R13952 VPWR.n4737 VPWR.n4736 1.13717
R13953 VPWR.n4726 VPWR.n4725 1.13717
R13954 VPWR.n4853 VPWR.n4852 1.13717
R13955 VPWR.n310 VPWR.n309 1.13717
R13956 VPWR.n4795 VPWR.n4794 1.13717
R13957 VPWR.n7394 VPWR.n7393 1.13717
R13958 VPWR.n7378 VPWR.n7377 1.13717
R13959 VPWR.n7325 VPWR.n7324 1.13717
R13960 VPWR.n7494 VPWR.n7493 1.13717
R13961 VPWR.n265 VPWR.n264 1.13717
R13962 VPWR.n7435 VPWR.n7434 1.13717
R13963 VPWR.n7511 VPWR.n7508 1.13717
R13964 VPWR.n254 VPWR.n250 1.13717
R13965 VPWR.n7517 VPWR.n7516 1.13717
R13966 VPWR.n1564 VPWR.n1563 1.13717
R13967 VPWR.n1548 VPWR.n1547 1.13717
R13968 VPWR.n3731 VPWR.n3730 1.13717
R13969 VPWR.n7654 VPWR.n7651 1.13717
R13970 VPWR.n126 VPWR.n125 1.13717
R13971 VPWR.n7660 VPWR.n7659 1.13717
R13972 VPWR.n2376 VPWR.n2375 1.13717
R13973 VPWR.n3398 VPWR.n3395 1.13717
R13974 VPWR.n3379 VPWR.n3378 1.13717
R13975 VPWR.n6005 VPWR.n6004 1.13717
R13976 VPWR.n5993 VPWR.n5992 1.13717
R13977 VPWR.n6019 VPWR.n6018 1.13717
R13978 VPWR.n6024 VPWR.n6023 1.13717
R13979 VPWR.n3066 VPWR.n3065 1.1368
R13980 VPWR.n4270 VPWR.n4269 1.1368
R13981 VPWR.n4420 VPWR.n4419 1.1368
R13982 VPWR.n4446 VPWR.n4445 1.1368
R13983 VPWR.n732 VPWR.n731 1.1368
R13984 VPWR.n7060 VPWR.n7059 1.1368
R13985 VPWR.n4908 VPWR.n4907 1.1368
R13986 VPWR.n6674 VPWR.n6575 1.1368
R13987 VPWR.n2064 VPWR.n2063 1.1368
R13988 VPWR.n5813 VPWR.n5812 1.1368
R13989 VPWR.n5783 VPWR.n5782 1.1368
R13990 VPWR.n3200 VPWR.n3199 1.1368
R13991 VPWR.n2188 VPWR.n2187 1.1368
R13992 VPWR.n6377 VPWR.n6376 1.1368
R13993 VPWR.n1917 VPWR.n1904 1.1368
R13994 VPWR.n1285 VPWR.n1284 1.1368
R13995 VPWR.n1007 VPWR.n1006 1.1368
R13996 VPWR.n547 VPWR.n540 1.1368
R13997 VPWR.n5422 VPWR.n5421 1.1368
R13998 VPWR.n5654 VPWR.n5653 1.1368
R13999 VPWR.n5685 VPWR.n5684 1.1368
R14000 VPWR.n1829 VPWR.n1828 1.1368
R14001 VPWR.n5709 VPWR.n5708 1.1368
R14002 VPWR.n7512 VPWR.n7511 1.1368
R14003 VPWR.n255 VPWR.n254 1.1368
R14004 VPWR.n127 VPWR.n126 1.1368
R14005 VPWR.n7655 VPWR.n7654 1.1368
R14006 VPWR.n3399 VPWR.n3398 1.1368
R14007 VPWR.n5993 VPWR.n5915 1.1368
R14008 VPWR.n2035 VPWR.n2034 1.13669
R14009 VPWR.n1414 VPWR.n419 1.13669
R14010 VPWR.n4433 VPWR.n4432 1.13669
R14011 VPWR.n624 VPWR.n623 1.13669
R14012 VPWR.n5295 VPWR.n4881 1.13669
R14013 VPWR.n7007 VPWR.n7006 1.13669
R14014 VPWR.n6600 VPWR.n6599 1.13669
R14015 VPWR.n2072 VPWR.n2070 1.13669
R14016 VPWR.n6571 VPWR.n6570 1.13669
R14017 VPWR.n2471 VPWR.n2470 1.13669
R14018 VPWR.n5818 VPWR.n5816 1.13669
R14019 VPWR.n3538 VPWR.n3537 1.13669
R14020 VPWR.n1502 VPWR.n1501 1.13669
R14021 VPWR.n4148 VPWR.n4134 1.13669
R14022 VPWR.n4284 VPWR.n4283 1.13669
R14023 VPWR.n4313 VPWR.n4299 1.13669
R14024 VPWR.n4556 VPWR.n4555 1.13669
R14025 VPWR.n4585 VPWR.n4571 1.13669
R14026 VPWR.n875 VPWR.n874 1.13669
R14027 VPWR.n849 VPWR.n597 1.13669
R14028 VPWR.n7202 VPWR.n7201 1.13669
R14029 VPWR.n7173 VPWR.n298 1.13669
R14030 VPWR.n6778 VPWR.n6777 1.13669
R14031 VPWR.n6890 VPWR.n6878 1.13669
R14032 VPWR.n6767 VPWR.n6766 1.13669
R14033 VPWR.n7632 VPWR.n7631 1.13669
R14034 VPWR.n3160 VPWR.n2392 1.13669
R14035 VPWR.n7802 VPWR.n7800 1.13669
R14036 VPWR.n7797 VPWR.n24 1.13669
R14037 VPWR.n7763 VPWR.n25 1.13669
R14038 VPWR.n6455 VPWR.n6453 1.13669
R14039 VPWR.n1842 VPWR.n1841 1.13669
R14040 VPWR.n1224 VPWR.n1223 1.13669
R14041 VPWR.n1210 VPWR.n1209 1.13669
R14042 VPWR.n978 VPWR.n977 1.13669
R14043 VPWR.n5228 VPWR.n5226 1.13669
R14044 VPWR.n5583 VPWR.n5425 1.13669
R14045 VPWR.n5659 VPWR.n5657 1.13669
R14046 VPWR.n1809 VPWR.n1807 1.13669
R14047 VPWR.n6355 VPWR.n6354 1.13669
R14048 VPWR.n2680 VPWR.n2498 1.13669
R14049 VPWR.n2678 VPWR.n2676 1.13669
R14050 VPWR.n4054 VPWR.n4052 1.13669
R14051 VPWR.n3986 VPWR.n3985 1.13669
R14052 VPWR.n3957 VPWR.n3956 1.13669
R14053 VPWR.n3762 VPWR.n3761 1.13669
R14054 VPWR.n4682 VPWR.n329 1.13669
R14055 VPWR.n4754 VPWR.n4753 1.13669
R14056 VPWR.n4759 VPWR.n4757 1.13669
R14057 VPWR.n4854 VPWR.n4853 1.13669
R14058 VPWR.n7294 VPWR.n7292 1.13669
R14059 VPWR.n7395 VPWR.n7394 1.13669
R14060 VPWR.n7400 VPWR.n7398 1.13669
R14061 VPWR.n7495 VPWR.n7494 1.13669
R14062 VPWR.n1565 VPWR.n1564 1.13669
R14063 VPWR.n3732 VPWR.n3731 1.13669
R14064 VPWR.n3371 VPWR.n3370 1.13669
R14065 VPWR.n822 VPWR.n821 1.12991
R14066 VPWR.n5162 VPWR.n5145 1.09272
R14067 VPWR.n5108 VPWR.n5107 1.09272
R14068 VPWR.n5240 VPWR.n5238 1.09272
R14069 VPWR.n7073 VPWR.n4869 1.09272
R14070 VPWR.n1251 VPWR.n1226 1.09272
R14071 VPWR.n6480 VPWR.n6479 1.09272
R14072 VPWR.n6400 VPWR.n6399 1.09272
R14073 VPWR.n2433 VPWR.n2432 1.09272
R14074 VPWR.n6850 VPWR.n6799 1.09216
R14075 VPWR.n648 VPWR.n646 1.09216
R14076 VPWR.n4486 VPWR.n397 1.09216
R14077 VPWR.n4625 VPWR.n375 1.09216
R14078 VPWR.n357 VPWR.n356 1.09216
R14079 VPWR.n7723 VPWR.n30 1.09216
R14080 VPWR.n664 VPWR.n643 1.09203
R14081 VPWR.n4506 VPWR.n4505 1.05773
R14082 VPWR.n3677 VPWR.n3643 1.05773
R14083 VPWR.n1478 VPWR.n1476 1.03351
R14084 VPWR.n6150 VPWR.n5826 0.935332
R14085 VPWR.n7128 VPWR.n7127 0.935332
R14086 VPWR.n6038 VPWR.n6037 0.935332
R14087 VPWR.n7162 VPWR 0.914786
R14088 VPWR.n1020 VPWR 0.899674
R14089 VPWR.n5467 VPWR 0.897835
R14090 VPWR.n1528 VPWR 0.896837
R14091 VPWR.n3307 VPWR 0.863992
R14092 VPWR.n904 VPWR 0.863992
R14093 VPWR.n894 VPWR 0.863992
R14094 VPWR.n1028 VPWR 0.863992
R14095 VPWR.n1865 VPWR 0.863992
R14096 VPWR.n3312 VPWR.n3311 0.842756
R14097 VPWR.n3616 VPWR 0.813198
R14098 VPWR.n3279 VPWR.n3272 0.802048
R14099 VPWR.n7667 VPWR.n7666 0.762405
R14100 VPWR.n1568 VPWR.n1567 0.762405
R14101 VPWR.n6907 VPWR.n6906 0.753441
R14102 VPWR.n495 VPWR.n494 0.753441
R14103 VPWR.n5594 VPWR.n5593 0.698804
R14104 VPWR VPWR.n5399 0.660817
R14105 VPWR.n6414 VPWR.n6413 0.656731
R14106 VPWR.n5670 VPWR.n5669 0.656731
R14107 VPWR.n5687 VPWR.n129 0.546928
R14108 VPWR.n538 VPWR.n300 0.546928
R14109 VPWR.n4273 VPWR.n1452 0.546928
R14110 VPWR.n6149 VPWR.n5827 0.539826
R14111 VPWR.n7133 VPWR.n7132 0.539826
R14112 VPWR.n6035 VPWR.n6034 0.539826
R14113 VPWR.n3921 VPWR.n3920 0.529114
R14114 VPWR.n2327 VPWR.n2326 0.529114
R14115 VPWR.n6058 VPWR.n6057 0.508436
R14116 VPWR.n6089 VPWR.n6088 0.508436
R14117 VPWR.n6690 VPWR.n6689 0.508436
R14118 VPWR.n7193 VPWR.n7192 0.508436
R14119 VPWR.n699 VPWR.n698 0.508436
R14120 VPWR.n6406 VPWR.n6405 0.491355
R14121 VPWR.n5114 VPWR.n5113 0.491355
R14122 VPWR.n7597 VPWR.n7596 0.415839
R14123 VPWR.n3017 VPWR.n2483 0.3805
R14124 VPWR.n3166 VPWR.n3165 0.378081
R14125 VPWR.n4217 VPWR.n1476 0.377983
R14126 VPWR.n7635 VPWR.n129 0.356928
R14127 VPWR.n7636 VPWR.n7635 0.356928
R14128 VPWR.n4858 VPWR.n300 0.356928
R14129 VPWR.n4858 VPWR.n4857 0.356928
R14130 VPWR.n4275 VPWR.n4273 0.356928
R14131 VPWR.n4275 VPWR.n4274 0.356928
R14132 VPWR.n696 VPWR.n695 0.356056
R14133 VPWR.n3002 VPWR.n3001 0.352216
R14134 VPWR.n2487 VPWR.n2206 0.347759
R14135 VPWR.n2369 VPWR.n2368 0.34507
R14136 VPWR.n3035 VPWR.n3034 0.342503
R14137 VPWR.n3017 VPWR.n3016 0.3424
R14138 VPWR.n3404 VPWR.n2287 0.3424
R14139 VPWR.n3017 VPWR.n2486 0.341811
R14140 VPWR.n3505 VPWR.n3494 0.341811
R14141 VPWR.n3505 VPWR.n3504 0.341811
R14142 VPWR.n2999 VPWR.n2998 0.341811
R14143 VPWR.n3404 VPWR.n2366 0.341811
R14144 VPWR.n2737 VPWR.n2491 0.31175
R14145 VPWR.n2205 VPWR.n2204 0.311379
R14146 VPWR.n3521 VPWR.n3520 0.311379
R14147 VPWR.n3410 VPWR.n3405 0.311379
R14148 VPWR.n2774 VPWR.n2684 0.311321
R14149 VPWR VPWR.n6611 0.305262
R14150 VPWR.n3879 VPWR.n3878 0.302565
R14151 VPWR.n3878 VPWR.n3877 0.302565
R14152 VPWR.n666 VPWR.n664 0.295115
R14153 VPWR.n5242 VPWR.n5240 0.294492
R14154 VPWR.n1253 VPWR.n1251 0.294492
R14155 VPWR.n650 VPWR.n648 0.294041
R14156 VPWR.n4627 VPWR.n4625 0.294041
R14157 VPWR.n356 VPWR.n355 0.294041
R14158 VPWR.n3311 VPWR 0.290856
R14159 VPWR VPWR.n5162 0.274365
R14160 VPWR.n6479 VPWR 0.274365
R14161 VPWR.n7020 VPWR.n7019 0.264807
R14162 VPWR.n3880 VPWR.n3879 0.264807
R14163 VPWR.n3311 VPWR 0.250033
R14164 VPWR.n5614 VPWR.n5613 0.246654
R14165 VPWR.n3827 VPWR.n3825 0.240185
R14166 VPWR.n7245 VPWR.n7244 0.23824
R14167 VPWR.n5107 VPWR 0.236604
R14168 VPWR.n5240 VPWR 0.236604
R14169 VPWR.n7073 VPWR 0.236604
R14170 VPWR.n1251 VPWR 0.236604
R14171 VPWR.n6399 VPWR 0.236604
R14172 VPWR VPWR.n2433 0.236604
R14173 VPWR.n664 VPWR 0.234963
R14174 VPWR VPWR.n6850 0.234145
R14175 VPWR.n648 VPWR 0.234145
R14176 VPWR VPWR.n397 0.234145
R14177 VPWR.n4625 VPWR 0.234145
R14178 VPWR.n356 VPWR 0.234145
R14179 VPWR.n30 VPWR 0.234145
R14180 VPWR.n7596 VPWR.n7595 0.227049
R14181 VPWR.n2291 VPWR 0.215749
R14182 VPWR.n4708 VPWR.n4707 0.21207
R14183 VPWR.n2336 VPWR.n2335 0.21207
R14184 VPWR.n1812 VPWR.n1798 0.205072
R14185 VPWR.n3707 VPWR.n3641 0.204272
R14186 VPWR.n5399 VPWR.n5345 0.203675
R14187 VPWR.n524 VPWR.n523 0.203675
R14188 VPWR.n1271 VPWR.n1270 0.203675
R14189 VPWR.n1891 VPWR.n1890 0.203675
R14190 VPWR.n2750 VPWR.n2749 0.203675
R14191 VPWR.n5162 VPWR 0.196835
R14192 VPWR.n5107 VPWR 0.196835
R14193 VPWR VPWR.n7073 0.196835
R14194 VPWR.n6479 VPWR 0.196835
R14195 VPWR.n6399 VPWR 0.196835
R14196 VPWR.n2433 VPWR 0.196835
R14197 VPWR.n6850 VPWR 0.196385
R14198 VPWR VPWR.n30 0.196385
R14199 VPWR.n397 VPWR 0.195082
R14200 VPWR.n4273 VPWR.n4272 0.1905
R14201 VPWR.n625 VPWR.n300 0.1905
R14202 VPWR.n6573 VPWR.n129 0.1905
R14203 VPWR.n4276 VPWR.n4275 0.1905
R14204 VPWR.n4859 VPWR.n4858 0.1905
R14205 VPWR.n7635 VPWR.n7634 0.1905
R14206 VPWR.n4857 VPWR.n4856 0.1905
R14207 VPWR.n7637 VPWR.n7636 0.1905
R14208 VPWR.n493 VPWR.n476 0.188735
R14209 VPWR.n497 VPWR.n495 0.188735
R14210 VPWR.n3336 VPWR.n3335 0.185115
R14211 VPWR.n7636 VPWR 0.183019
R14212 VPWR.n4857 VPWR 0.183019
R14213 VPWR.n4274 VPWR 0.183019
R14214 VPWR.n1047 VPWR.n1045 0.180551
R14215 VPWR.n4083 VPWR.n4082 0.180294
R14216 VPWR.n5318 VPWR.n5317 0.179926
R14217 VPWR.n5317 VPWR.n5315 0.179926
R14218 VPWR.n4182 VPWR.n4180 0.179926
R14219 VPWR.n4180 VPWR.n4178 0.179926
R14220 VPWR VPWR.n5187 0.179673
R14221 VPWR VPWR.n6704 0.179673
R14222 VPWR.n4196 VPWR 0.179673
R14223 VPWR.n5003 VPWR 0.179673
R14224 VPWR.n2434 VPWR 0.179673
R14225 VPWR.n3121 VPWR 0.179673
R14226 VPWR.n3137 VPWR 0.179673
R14227 VPWR.n2800 VPWR 0.179498
R14228 VPWR.n2371 VPWR 0.179389
R14229 VPWR.n7328 VPWR 0.178345
R14230 VPWR VPWR.n4801 0.178345
R14231 VPWR VPWR.n343 0.178345
R14232 VPWR.n3305 VPWR 0.178345
R14233 VPWR VPWR.n5093 0.177989
R14234 VPWR VPWR.n175 0.177989
R14235 VPWR.n6820 VPWR 0.177989
R14236 VPWR VPWR.n7445 0.177989
R14237 VPWR.n5363 VPWR 0.177989
R14238 VPWR.n7271 VPWR 0.177989
R14239 VPWR VPWR.n7245 0.177989
R14240 VPWR.n487 VPWR 0.177989
R14241 VPWR.n677 VPWR 0.177989
R14242 VPWR.n892 VPWR 0.177989
R14243 VPWR.n1023 VPWR 0.177989
R14244 VPWR VPWR.n4385 0.177989
R14245 VPWR.n3887 VPWR 0.177989
R14246 VPWR.n1960 VPWR 0.177989
R14247 VPWR.n3997 VPWR 0.177989
R14248 VPWR.n3588 VPWR 0.177989
R14249 VPWR.n3590 VPWR 0.177989
R14250 VPWR.n3641 VPWR 0.177989
R14251 VPWR VPWR.n3649 0.177989
R14252 VPWR.n2695 VPWR 0.177989
R14253 VPWR.n6382 VPWR 0.177989
R14254 VPWR VPWR.n61 0.177989
R14255 VPWR VPWR.n55 0.177989
R14256 VPWR.n5094 VPWR 0.171212
R14257 VPWR VPWR.n5430 0.171212
R14258 VPWR.n5352 VPWR 0.171212
R14259 VPWR VPWR.n480 0.171212
R14260 VPWR VPWR.n1022 0.171212
R14261 VPWR.n1228 VPWR 0.171212
R14262 VPWR VPWR.n1849 0.171212
R14263 VPWR.n1674 VPWR 0.171212
R14264 VPWR VPWR.n2694 0.171212
R14265 VPWR VPWR.n6381 0.171212
R14266 VPWR.n2581 VPWR 0.171212
R14267 VPWR.n5933 VPWR.n5932 0.160318
R14268 VPWR VPWR.n1594 0.15779
R14269 VPWR VPWR.n4097 0.156488
R14270 VPWR.n6288 VPWR.n6285 0.153014
R14271 VPWR.n86 VPWR.n85 0.152881
R14272 VPWR.n229 VPWR.n228 0.152881
R14273 VPWR.n7481 VPWR.n7480 0.152881
R14274 VPWR.n7192 VPWR.n7191 0.152881
R14275 VPWR.n3688 VPWR.n3687 0.152881
R14276 VPWR.n5984 VPWR.n5983 0.152881
R14277 VPWR.n6405 VPWR.n6404 0.151532
R14278 VPWR.n5113 VPWR.n5112 0.151532
R14279 VPWR.n5815 VPWR.n5814 0.151488
R14280 VPWR.n6589 VPWR.n6588 0.151488
R14281 VPWR.n7009 VPWR.n7008 0.151488
R14282 VPWR.n613 VPWR.n417 0.151488
R14283 VPWR.n4422 VPWR.n4421 0.151488
R14284 VPWR.n2037 VPWR.n2036 0.151488
R14285 VPWR.n7799 VPWR.n7798 0.151488
R14286 VPWR.n6769 VPWR.n6768 0.151488
R14287 VPWR.n6771 VPWR.n6770 0.151488
R14288 VPWR.n598 VPWR.n387 0.151488
R14289 VPWR.n1450 VPWR.n388 0.151488
R14290 VPWR.n2160 VPWR.n2159 0.151488
R14291 VPWR.n6357 VPWR.n6356 0.151488
R14292 VPWR.n5656 VPWR.n5655 0.151488
R14293 VPWR.n5424 VPWR.n5423 0.151488
R14294 VPWR.n980 VPWR.n979 0.151488
R14295 VPWR.n1212 VPWR.n1211 0.151488
R14296 VPWR.n1831 VPWR.n1830 0.151488
R14297 VPWR.n5912 VPWR.n5911 0.151488
R14298 VPWR.n7497 VPWR.n7496 0.151488
R14299 VPWR.n7397 VPWR.n7396 0.151488
R14300 VPWR.n4756 VPWR.n4755 0.151488
R14301 VPWR.n3736 VPWR.n3735 0.151488
R14302 VPWR.n3734 VPWR.n3733 0.151488
R14303 VPWR.n3524 VPWR.n3523 0.149872
R14304 VPWR.n7663 VPWR.n7662 0.145957
R14305 VPWR.n6146 VPWR.n6145 0.14432
R14306 VPWR.n7136 VPWR.n7135 0.14432
R14307 VPWR.n6030 VPWR.n6029 0.14432
R14308 VPWR.n3038 VPWR.n3037 0.143372
R14309 VPWR.n2395 VPWR.n2394 0.143372
R14310 VPWR.n2682 VPWR.n2681 0.143372
R14311 VPWR.n3401 VPWR.n3400 0.143372
R14312 VPWR VPWR.n2800 0.141026
R14313 VPWR.n5187 VPWR 0.140863
R14314 VPWR.n6704 VPWR 0.140863
R14315 VPWR.n4196 VPWR 0.140863
R14316 VPWR.n1798 VPWR 0.140863
R14317 VPWR.n5003 VPWR 0.140863
R14318 VPWR.n2434 VPWR 0.140863
R14319 VPWR VPWR.n3121 0.140863
R14320 VPWR VPWR.n3137 0.140863
R14321 VPWR.n5093 VPWR 0.140584
R14322 VPWR.n175 VPWR 0.140584
R14323 VPWR.n6820 VPWR 0.140584
R14324 VPWR.n7445 VPWR 0.140584
R14325 VPWR VPWR.n5363 0.140584
R14326 VPWR.n7271 VPWR 0.140584
R14327 VPWR VPWR.n487 0.140584
R14328 VPWR VPWR.n677 0.140584
R14329 VPWR VPWR.n1023 0.140584
R14330 VPWR.n4385 VPWR 0.140584
R14331 VPWR.n3887 VPWR 0.140584
R14332 VPWR.n1960 VPWR 0.140584
R14333 VPWR.n3997 VPWR 0.140584
R14334 VPWR VPWR.n3588 0.140584
R14335 VPWR.n3590 VPWR 0.140584
R14336 VPWR.n3649 VPWR 0.140584
R14337 VPWR.n2695 VPWR 0.140584
R14338 VPWR.n2291 VPWR 0.140584
R14339 VPWR.n6382 VPWR 0.140584
R14340 VPWR.n61 VPWR 0.140584
R14341 VPWR.n55 VPWR 0.140584
R14342 VPWR.n7328 VPWR 0.140228
R14343 VPWR.n4801 VPWR 0.140228
R14344 VPWR.n343 VPWR 0.140228
R14345 VPWR.n3305 VPWR 0.140228
R14346 VPWR VPWR.n892 0.139282
R14347 VPWR.n4272 VPWR.n4271 0.125931
R14348 VPWR.n4276 VPWR.n1451 0.125931
R14349 VPWR.n1654 VPWR.n1452 0.125931
R14350 VPWR.n3960 VPWR.n3959 0.125931
R14351 VPWR.n3345 VPWR.n3344 0.123577
R14352 VPWR.n5163 VPWR 0.120655
R14353 VPWR.n5104 VPWR 0.120655
R14354 VPWR.n5106 VPWR 0.120655
R14355 VPWR VPWR.n5557 0.120655
R14356 VPWR VPWR.n5498 0.120655
R14357 VPWR.n1532 VPWR 0.120655
R14358 VPWR.n4083 VPWR 0.120655
R14359 VPWR VPWR.n1582 0.120655
R14360 VPWR.n2896 VPWR 0.120655
R14361 VPWR.n6478 VPWR 0.120655
R14362 VPWR VPWR.n3281 0.120655
R14363 VPWR.n3263 VPWR 0.120655
R14364 VPWR.n3138 VPWR 0.120655
R14365 VPWR.n5104 VPWR 0.120399
R14366 VPWR VPWR.n1582 0.120399
R14367 VPWR.n5100 VPWR.n5098 0.120292
R14368 VPWR.n5102 VPWR.n5100 0.120292
R14369 VPWR.n5116 VPWR.n5111 0.120292
R14370 VPWR.n5203 VPWR.n5202 0.120292
R14371 VPWR.n5202 VPWR.n5200 0.120292
R14372 VPWR.n5200 VPWR.n5198 0.120292
R14373 VPWR.n5198 VPWR.n5195 0.120292
R14374 VPWR.n5195 VPWR.n5193 0.120292
R14375 VPWR.n5193 VPWR.n5191 0.120292
R14376 VPWR.n5182 VPWR.n5181 0.120292
R14377 VPWR.n5181 VPWR.n5179 0.120292
R14378 VPWR.n5175 VPWR.n5174 0.120292
R14379 VPWR.n5174 VPWR.n5172 0.120292
R14380 VPWR.n5169 VPWR.n5168 0.120292
R14381 VPWR.n5168 VPWR.n5166 0.120292
R14382 VPWR.n5161 VPWR.n5158 0.120292
R14383 VPWR.n5158 VPWR.n5156 0.120292
R14384 VPWR.n5156 VPWR.n5154 0.120292
R14385 VPWR.n5154 VPWR.n5152 0.120292
R14386 VPWR.n5152 VPWR.n5149 0.120292
R14387 VPWR.n5149 VPWR.n5147 0.120292
R14388 VPWR.n5147 VPWR.n5146 0.120292
R14389 VPWR.n6650 VPWR.n6649 0.120292
R14390 VPWR.n6649 VPWR.n6647 0.120292
R14391 VPWR.n6647 VPWR.n6645 0.120292
R14392 VPWR.n6645 VPWR.n6643 0.120292
R14393 VPWR.n6643 VPWR.n6640 0.120292
R14394 VPWR.n6640 VPWR.n6638 0.120292
R14395 VPWR.n6638 VPWR.n6636 0.120292
R14396 VPWR.n6636 VPWR.n6634 0.120292
R14397 VPWR.n6634 VPWR.n6632 0.120292
R14398 VPWR.n6632 VPWR.n6630 0.120292
R14399 VPWR.n6630 VPWR.n6628 0.120292
R14400 VPWR.n6625 VPWR.n6624 0.120292
R14401 VPWR.n6624 VPWR.n6623 0.120292
R14402 VPWR.n6623 VPWR.n6621 0.120292
R14403 VPWR.n6621 VPWR.n6619 0.120292
R14404 VPWR.n6619 VPWR.n6618 0.120292
R14405 VPWR.n6618 VPWR.n6617 0.120292
R14406 VPWR.n6713 VPWR.n6711 0.120292
R14407 VPWR.n6715 VPWR.n6713 0.120292
R14408 VPWR.n6717 VPWR.n6715 0.120292
R14409 VPWR.n6720 VPWR.n6717 0.120292
R14410 VPWR.n6722 VPWR.n6720 0.120292
R14411 VPWR.n6724 VPWR.n6722 0.120292
R14412 VPWR.n6726 VPWR.n6724 0.120292
R14413 VPWR.n6728 VPWR.n6726 0.120292
R14414 VPWR.n6730 VPWR.n6728 0.120292
R14415 VPWR.n6732 VPWR.n6730 0.120292
R14416 VPWR.n6733 VPWR.n6732 0.120292
R14417 VPWR.n6737 VPWR.n6736 0.120292
R14418 VPWR.n6742 VPWR.n6740 0.120292
R14419 VPWR.n6744 VPWR.n6742 0.120292
R14420 VPWR.n6746 VPWR.n6744 0.120292
R14421 VPWR.n7599 VPWR.n7594 0.120292
R14422 VPWR.n7594 VPWR.n7591 0.120292
R14423 VPWR.n7591 VPWR.n7589 0.120292
R14424 VPWR.n7589 VPWR.n7587 0.120292
R14425 VPWR.n7530 VPWR.n7528 0.120292
R14426 VPWR.n7531 VPWR.n7530 0.120292
R14427 VPWR.n7536 VPWR.n7534 0.120292
R14428 VPWR.n7538 VPWR.n7536 0.120292
R14429 VPWR.n7540 VPWR.n7538 0.120292
R14430 VPWR.n7543 VPWR.n7540 0.120292
R14431 VPWR.n7545 VPWR.n7543 0.120292
R14432 VPWR.n7547 VPWR.n7545 0.120292
R14433 VPWR.n7549 VPWR.n7547 0.120292
R14434 VPWR.n7551 VPWR.n7549 0.120292
R14435 VPWR.n7553 VPWR.n7551 0.120292
R14436 VPWR.n7555 VPWR.n7553 0.120292
R14437 VPWR.n7557 VPWR.n7555 0.120292
R14438 VPWR.n7561 VPWR.n7559 0.120292
R14439 VPWR.n7563 VPWR.n7561 0.120292
R14440 VPWR.n7565 VPWR.n7563 0.120292
R14441 VPWR.n7566 VPWR.n7565 0.120292
R14442 VPWR.n7571 VPWR.n7569 0.120292
R14443 VPWR.n7573 VPWR.n7571 0.120292
R14444 VPWR.n7575 VPWR.n7573 0.120292
R14445 VPWR.n7577 VPWR.n7575 0.120292
R14446 VPWR.n7579 VPWR.n7577 0.120292
R14447 VPWR.n7580 VPWR.n7579 0.120292
R14448 VPWR.n7523 VPWR.n7522 0.120292
R14449 VPWR.n203 VPWR.n201 0.120292
R14450 VPWR.n201 VPWR.n200 0.120292
R14451 VPWR.n200 VPWR.n198 0.120292
R14452 VPWR.n198 VPWR.n196 0.120292
R14453 VPWR.n196 VPWR.n194 0.120292
R14454 VPWR.n190 VPWR.n189 0.120292
R14455 VPWR.n189 VPWR.n188 0.120292
R14456 VPWR.n188 VPWR.n187 0.120292
R14457 VPWR.n187 VPWR.n185 0.120292
R14458 VPWR.n185 VPWR.n183 0.120292
R14459 VPWR.n178 VPWR.n176 0.120292
R14460 VPWR.n5437 VPWR.n5435 0.120292
R14461 VPWR.n5439 VPWR.n5437 0.120292
R14462 VPWR.n5441 VPWR.n5439 0.120292
R14463 VPWR.n5448 VPWR.n5446 0.120292
R14464 VPWR.n5450 VPWR.n5448 0.120292
R14465 VPWR.n5453 VPWR.n5450 0.120292
R14466 VPWR.n5455 VPWR.n5453 0.120292
R14467 VPWR.n5456 VPWR.n5455 0.120292
R14468 VPWR.n5462 VPWR.n5460 0.120292
R14469 VPWR.n5574 VPWR.n5573 0.120292
R14470 VPWR.n5573 VPWR.n5571 0.120292
R14471 VPWR.n5571 VPWR.n5569 0.120292
R14472 VPWR.n5569 VPWR.n5566 0.120292
R14473 VPWR.n5566 VPWR.n5564 0.120292
R14474 VPWR.n5564 VPWR.n5562 0.120292
R14475 VPWR.n5556 VPWR.n5546 0.120292
R14476 VPWR.n5546 VPWR.n5545 0.120292
R14477 VPWR.n5545 VPWR.n5544 0.120292
R14478 VPWR.n5544 VPWR.n5542 0.120292
R14479 VPWR.n5542 VPWR.n5539 0.120292
R14480 VPWR.n5537 VPWR.n5535 0.120292
R14481 VPWR.n5535 VPWR.n5533 0.120292
R14482 VPWR.n5533 VPWR.n5531 0.120292
R14483 VPWR.n5531 VPWR.n5529 0.120292
R14484 VPWR.n5529 VPWR.n5527 0.120292
R14485 VPWR.n5524 VPWR.n5523 0.120292
R14486 VPWR.n5523 VPWR.n5521 0.120292
R14487 VPWR.n5521 VPWR.n5519 0.120292
R14488 VPWR.n5519 VPWR.n5517 0.120292
R14489 VPWR.n5517 VPWR.n5514 0.120292
R14490 VPWR.n5514 VPWR.n5512 0.120292
R14491 VPWR.n5512 VPWR.n5510 0.120292
R14492 VPWR.n5510 VPWR.n5508 0.120292
R14493 VPWR.n5508 VPWR.n5506 0.120292
R14494 VPWR.n5506 VPWR.n5504 0.120292
R14495 VPWR.n5504 VPWR.n5502 0.120292
R14496 VPWR.n6990 VPWR.n6988 0.120292
R14497 VPWR.n6988 VPWR.n6986 0.120292
R14498 VPWR.n6986 VPWR.n6984 0.120292
R14499 VPWR.n6981 VPWR.n6980 0.120292
R14500 VPWR.n6980 VPWR.n6978 0.120292
R14501 VPWR.n6978 VPWR.n6976 0.120292
R14502 VPWR.n6976 VPWR.n6974 0.120292
R14503 VPWR.n6970 VPWR.n6969 0.120292
R14504 VPWR.n6969 VPWR.n6968 0.120292
R14505 VPWR.n6968 VPWR.n6967 0.120292
R14506 VPWR.n6967 VPWR.n6965 0.120292
R14507 VPWR.n6965 VPWR.n6963 0.120292
R14508 VPWR.n6959 VPWR.n6958 0.120292
R14509 VPWR.n6958 VPWR.n6956 0.120292
R14510 VPWR.n6950 VPWR.n6949 0.120292
R14511 VPWR.n6949 VPWR.n6948 0.120292
R14512 VPWR.n6948 VPWR.n6947 0.120292
R14513 VPWR.n6944 VPWR.n6943 0.120292
R14514 VPWR.n6943 VPWR.n6941 0.120292
R14515 VPWR.n6941 VPWR.n6939 0.120292
R14516 VPWR.n6939 VPWR.n6937 0.120292
R14517 VPWR.n6937 VPWR.n6934 0.120292
R14518 VPWR.n6934 VPWR.n6932 0.120292
R14519 VPWR.n6932 VPWR.n6930 0.120292
R14520 VPWR.n6930 VPWR.n6928 0.120292
R14521 VPWR.n6928 VPWR.n6926 0.120292
R14522 VPWR.n6864 VPWR.n6859 0.120292
R14523 VPWR.n6859 VPWR.n6858 0.120292
R14524 VPWR.n6858 VPWR.n6857 0.120292
R14525 VPWR.n6808 VPWR.n6806 0.120292
R14526 VPWR.n6810 VPWR.n6808 0.120292
R14527 VPWR.n6812 VPWR.n6810 0.120292
R14528 VPWR.n6814 VPWR.n6812 0.120292
R14529 VPWR.n6815 VPWR.n6814 0.120292
R14530 VPWR.n6819 VPWR.n6818 0.120292
R14531 VPWR.n6826 VPWR.n6824 0.120292
R14532 VPWR.n6829 VPWR.n6826 0.120292
R14533 VPWR.n6831 VPWR.n6829 0.120292
R14534 VPWR.n6833 VPWR.n6831 0.120292
R14535 VPWR.n6834 VPWR.n6833 0.120292
R14536 VPWR.n6835 VPWR.n6834 0.120292
R14537 VPWR.n6836 VPWR.n6835 0.120292
R14538 VPWR.n6842 VPWR.n6840 0.120292
R14539 VPWR.n6844 VPWR.n6842 0.120292
R14540 VPWR.n6846 VPWR.n6844 0.120292
R14541 VPWR.n6848 VPWR.n6846 0.120292
R14542 VPWR.n6849 VPWR.n6848 0.120292
R14543 VPWR.n7472 VPWR.n7470 0.120292
R14544 VPWR.n7470 VPWR.n7468 0.120292
R14545 VPWR.n7468 VPWR.n7466 0.120292
R14546 VPWR.n7463 VPWR.n7462 0.120292
R14547 VPWR.n7462 VPWR.n7461 0.120292
R14548 VPWR.n7461 VPWR.n7460 0.120292
R14549 VPWR.n7456 VPWR.n7455 0.120292
R14550 VPWR.n7454 VPWR.n7452 0.120292
R14551 VPWR.n7448 VPWR.n7447 0.120292
R14552 VPWR.n7447 VPWR.n7446 0.120292
R14553 VPWR.n5356 VPWR.n5355 0.120292
R14554 VPWR.n5357 VPWR.n5356 0.120292
R14555 VPWR.n5358 VPWR.n5357 0.120292
R14556 VPWR.n5369 VPWR.n5367 0.120292
R14557 VPWR.n5371 VPWR.n5369 0.120292
R14558 VPWR.n5373 VPWR.n5371 0.120292
R14559 VPWR.n5374 VPWR.n5373 0.120292
R14560 VPWR.n5323 VPWR.n5322 0.120292
R14561 VPWR.n5322 VPWR.n5320 0.120292
R14562 VPWR.n5320 VPWR.n5318 0.120292
R14563 VPWR.n5244 VPWR.n5242 0.120292
R14564 VPWR.n5246 VPWR.n5244 0.120292
R14565 VPWR.n5247 VPWR.n5246 0.120292
R14566 VPWR.n5252 VPWR.n5250 0.120292
R14567 VPWR.n5259 VPWR.n5256 0.120292
R14568 VPWR.n5261 VPWR.n5259 0.120292
R14569 VPWR.n5263 VPWR.n5261 0.120292
R14570 VPWR.n5265 VPWR.n5263 0.120292
R14571 VPWR.n5267 VPWR.n5265 0.120292
R14572 VPWR.n5269 VPWR.n5267 0.120292
R14573 VPWR.n5271 VPWR.n5269 0.120292
R14574 VPWR.n5273 VPWR.n5271 0.120292
R14575 VPWR.n5279 VPWR.n5278 0.120292
R14576 VPWR.n5284 VPWR.n5283 0.120292
R14577 VPWR.n5307 VPWR.n5306 0.120292
R14578 VPWR.n7078 VPWR.n7077 0.120292
R14579 VPWR.n7088 VPWR.n7087 0.120292
R14580 VPWR.n7089 VPWR.n7088 0.120292
R14581 VPWR.n7091 VPWR.n7089 0.120292
R14582 VPWR.n7093 VPWR.n7091 0.120292
R14583 VPWR.n7103 VPWR.n7100 0.120292
R14584 VPWR.n7106 VPWR.n7103 0.120292
R14585 VPWR.n7108 VPWR.n7106 0.120292
R14586 VPWR.n7110 VPWR.n7108 0.120292
R14587 VPWR.n7111 VPWR.n7110 0.120292
R14588 VPWR.n7112 VPWR.n7111 0.120292
R14589 VPWR.n7116 VPWR.n7112 0.120292
R14590 VPWR.n7129 VPWR.n7126 0.120292
R14591 VPWR.n7134 VPWR.n7129 0.120292
R14592 VPWR.n7137 VPWR.n7134 0.120292
R14593 VPWR.n7139 VPWR.n7137 0.120292
R14594 VPWR.n7220 VPWR.n7219 0.120292
R14595 VPWR.n7222 VPWR.n7220 0.120292
R14596 VPWR.n7224 VPWR.n7222 0.120292
R14597 VPWR.n7270 VPWR.n7269 0.120292
R14598 VPWR.n7269 VPWR.n7268 0.120292
R14599 VPWR.n7268 VPWR.n7267 0.120292
R14600 VPWR.n7267 VPWR.n7265 0.120292
R14601 VPWR.n7265 VPWR.n7263 0.120292
R14602 VPWR.n7263 VPWR.n7261 0.120292
R14603 VPWR.n7261 VPWR.n7259 0.120292
R14604 VPWR.n7256 VPWR.n7255 0.120292
R14605 VPWR.n7255 VPWR.n7253 0.120292
R14606 VPWR.n7253 VPWR.n7251 0.120292
R14607 VPWR.n7251 VPWR.n7249 0.120292
R14608 VPWR.n7244 VPWR.n7242 0.120292
R14609 VPWR.n7242 VPWR.n7241 0.120292
R14610 VPWR.n7241 VPWR.n7240 0.120292
R14611 VPWR.n7237 VPWR.n7236 0.120292
R14612 VPWR.n7284 VPWR.n7282 0.120292
R14613 VPWR.n7286 VPWR.n7284 0.120292
R14614 VPWR.n7362 VPWR.n7360 0.120292
R14615 VPWR.n7360 VPWR.n7358 0.120292
R14616 VPWR.n7358 VPWR.n7356 0.120292
R14617 VPWR.n7356 VPWR.n7354 0.120292
R14618 VPWR.n7354 VPWR.n7352 0.120292
R14619 VPWR.n7348 VPWR.n7347 0.120292
R14620 VPWR.n7344 VPWR.n7343 0.120292
R14621 VPWR.n7338 VPWR.n7333 0.120292
R14622 VPWR.n7333 VPWR.n7332 0.120292
R14623 VPWR.n7332 VPWR.n7331 0.120292
R14624 VPWR.n486 VPWR.n484 0.120292
R14625 VPWR.n500 VPWR.n498 0.120292
R14626 VPWR.n502 VPWR.n500 0.120292
R14627 VPWR.n503 VPWR.n502 0.120292
R14628 VPWR.n510 VPWR.n507 0.120292
R14629 VPWR.n969 VPWR.n968 0.120292
R14630 VPWR.n968 VPWR.n967 0.120292
R14631 VPWR.n967 VPWR.n965 0.120292
R14632 VPWR.n965 VPWR.n963 0.120292
R14633 VPWR.n963 VPWR.n961 0.120292
R14634 VPWR.n961 VPWR.n959 0.120292
R14635 VPWR.n652 VPWR.n650 0.120292
R14636 VPWR.n654 VPWR.n652 0.120292
R14637 VPWR.n655 VPWR.n654 0.120292
R14638 VPWR.n660 VPWR.n659 0.120292
R14639 VPWR.n667 VPWR.n666 0.120292
R14640 VPWR.n668 VPWR.n667 0.120292
R14641 VPWR.n669 VPWR.n668 0.120292
R14642 VPWR.n674 VPWR.n672 0.120292
R14643 VPWR.n676 VPWR.n674 0.120292
R14644 VPWR.n747 VPWR.n745 0.120292
R14645 VPWR.n749 VPWR.n747 0.120292
R14646 VPWR.n750 VPWR.n749 0.120292
R14647 VPWR.n758 VPWR.n757 0.120292
R14648 VPWR.n759 VPWR.n758 0.120292
R14649 VPWR.n760 VPWR.n759 0.120292
R14650 VPWR.n764 VPWR.n763 0.120292
R14651 VPWR.n765 VPWR.n764 0.120292
R14652 VPWR.n770 VPWR.n768 0.120292
R14653 VPWR.n772 VPWR.n770 0.120292
R14654 VPWR.n774 VPWR.n772 0.120292
R14655 VPWR.n776 VPWR.n774 0.120292
R14656 VPWR.n778 VPWR.n776 0.120292
R14657 VPWR.n780 VPWR.n778 0.120292
R14658 VPWR.n782 VPWR.n780 0.120292
R14659 VPWR.n787 VPWR.n785 0.120292
R14660 VPWR.n789 VPWR.n787 0.120292
R14661 VPWR.n791 VPWR.n789 0.120292
R14662 VPWR.n793 VPWR.n791 0.120292
R14663 VPWR.n795 VPWR.n793 0.120292
R14664 VPWR.n797 VPWR.n795 0.120292
R14665 VPWR.n799 VPWR.n797 0.120292
R14666 VPWR.n801 VPWR.n799 0.120292
R14667 VPWR.n803 VPWR.n801 0.120292
R14668 VPWR.n804 VPWR.n803 0.120292
R14669 VPWR.n811 VPWR.n810 0.120292
R14670 VPWR.n812 VPWR.n811 0.120292
R14671 VPWR.n814 VPWR.n812 0.120292
R14672 VPWR.n820 VPWR.n818 0.120292
R14673 VPWR.n891 VPWR.n889 0.120292
R14674 VPWR.n899 VPWR.n898 0.120292
R14675 VPWR.n900 VPWR.n899 0.120292
R14676 VPWR.n907 VPWR.n906 0.120292
R14677 VPWR.n913 VPWR.n911 0.120292
R14678 VPWR.n915 VPWR.n913 0.120292
R14679 VPWR.n917 VPWR.n915 0.120292
R14680 VPWR.n919 VPWR.n917 0.120292
R14681 VPWR.n921 VPWR.n919 0.120292
R14682 VPWR.n923 VPWR.n921 0.120292
R14683 VPWR.n925 VPWR.n923 0.120292
R14684 VPWR.n927 VPWR.n925 0.120292
R14685 VPWR.n929 VPWR.n927 0.120292
R14686 VPWR.n931 VPWR.n929 0.120292
R14687 VPWR.n933 VPWR.n931 0.120292
R14688 VPWR.n935 VPWR.n933 0.120292
R14689 VPWR.n937 VPWR.n935 0.120292
R14690 VPWR.n939 VPWR.n937 0.120292
R14691 VPWR.n941 VPWR.n939 0.120292
R14692 VPWR.n943 VPWR.n941 0.120292
R14693 VPWR.n944 VPWR.n943 0.120292
R14694 VPWR.n945 VPWR.n944 0.120292
R14695 VPWR.n948 VPWR.n946 0.120292
R14696 VPWR.n946 VPWR.n322 0.120292
R14697 VPWR.n4765 VPWR.n322 0.120292
R14698 VPWR.n4828 VPWR.n4827 0.120292
R14699 VPWR.n4827 VPWR.n4825 0.120292
R14700 VPWR.n4825 VPWR.n4824 0.120292
R14701 VPWR.n4824 VPWR.n4822 0.120292
R14702 VPWR.n4819 VPWR.n4818 0.120292
R14703 VPWR.n4818 VPWR.n4816 0.120292
R14704 VPWR.n4816 VPWR.n4814 0.120292
R14705 VPWR.n4811 VPWR.n4810 0.120292
R14706 VPWR.n4810 VPWR.n4808 0.120292
R14707 VPWR.n4804 VPWR.n4803 0.120292
R14708 VPWR.n4803 VPWR.n4802 0.120292
R14709 VPWR.n1024 VPWR.n1019 0.120292
R14710 VPWR.n1029 VPWR.n1019 0.120292
R14711 VPWR.n1031 VPWR.n1030 0.120292
R14712 VPWR.n1032 VPWR.n1031 0.120292
R14713 VPWR.n1037 VPWR.n1035 0.120292
R14714 VPWR.n1039 VPWR.n1037 0.120292
R14715 VPWR.n1041 VPWR.n1039 0.120292
R14716 VPWR.n1202 VPWR.n1200 0.120292
R14717 VPWR.n1200 VPWR.n1198 0.120292
R14718 VPWR.n1198 VPWR.n1196 0.120292
R14719 VPWR.n1196 VPWR.n1194 0.120292
R14720 VPWR.n1194 VPWR.n1191 0.120292
R14721 VPWR.n1187 VPWR.n1186 0.120292
R14722 VPWR.n1183 VPWR.n1182 0.120292
R14723 VPWR.n1182 VPWR.n1180 0.120292
R14724 VPWR.n1177 VPWR.n1176 0.120292
R14725 VPWR.n1176 VPWR.n1174 0.120292
R14726 VPWR.n1174 VPWR.n1172 0.120292
R14727 VPWR.n1172 VPWR.n1170 0.120292
R14728 VPWR.n1170 VPWR.n1167 0.120292
R14729 VPWR.n1167 VPWR.n1165 0.120292
R14730 VPWR.n1165 VPWR.n1163 0.120292
R14731 VPWR.n1163 VPWR.n1161 0.120292
R14732 VPWR.n1161 VPWR.n1159 0.120292
R14733 VPWR.n1159 VPWR.n1157 0.120292
R14734 VPWR.n1157 VPWR.n1155 0.120292
R14735 VPWR.n1152 VPWR.n1151 0.120292
R14736 VPWR.n1151 VPWR.n1149 0.120292
R14737 VPWR.n1149 VPWR.n1148 0.120292
R14738 VPWR.n1148 VPWR.n1147 0.120292
R14739 VPWR.n1143 VPWR.n1141 0.120292
R14740 VPWR.n1137 VPWR.n1136 0.120292
R14741 VPWR.n1132 VPWR.n1131 0.120292
R14742 VPWR.n4466 VPWR.n4464 0.120292
R14743 VPWR.n4468 VPWR.n4466 0.120292
R14744 VPWR.n4469 VPWR.n4468 0.120292
R14745 VPWR.n4474 VPWR.n4472 0.120292
R14746 VPWR.n4476 VPWR.n4474 0.120292
R14747 VPWR.n4478 VPWR.n4476 0.120292
R14748 VPWR.n4480 VPWR.n4478 0.120292
R14749 VPWR.n4482 VPWR.n4480 0.120292
R14750 VPWR.n4483 VPWR.n4482 0.120292
R14751 VPWR.n4490 VPWR.n4489 0.120292
R14752 VPWR.n4497 VPWR.n4496 0.120292
R14753 VPWR.n4504 VPWR.n4503 0.120292
R14754 VPWR.n4509 VPWR.n4507 0.120292
R14755 VPWR.n4513 VPWR.n4509 0.120292
R14756 VPWR.n4515 VPWR.n4513 0.120292
R14757 VPWR.n4518 VPWR.n4515 0.120292
R14758 VPWR.n4519 VPWR.n4518 0.120292
R14759 VPWR.n4520 VPWR.n4519 0.120292
R14760 VPWR.n4521 VPWR.n4520 0.120292
R14761 VPWR.n4527 VPWR.n4525 0.120292
R14762 VPWR.n4615 VPWR.n4613 0.120292
R14763 VPWR.n4617 VPWR.n4615 0.120292
R14764 VPWR.n4619 VPWR.n4617 0.120292
R14765 VPWR.n4620 VPWR.n4619 0.120292
R14766 VPWR.n4629 VPWR.n4627 0.120292
R14767 VPWR.n4631 VPWR.n4629 0.120292
R14768 VPWR.n4632 VPWR.n4631 0.120292
R14769 VPWR.n373 VPWR.n372 0.120292
R14770 VPWR.n4640 VPWR.n4639 0.120292
R14771 VPWR.n4645 VPWR.n4643 0.120292
R14772 VPWR.n4646 VPWR.n4645 0.120292
R14773 VPWR.n4652 VPWR.n4651 0.120292
R14774 VPWR.n4658 VPWR.n4656 0.120292
R14775 VPWR.n4659 VPWR.n4658 0.120292
R14776 VPWR.n4660 VPWR.n4659 0.120292
R14777 VPWR.n4661 VPWR.n4660 0.120292
R14778 VPWR.n4672 VPWR.n4669 0.120292
R14779 VPWR.n4674 VPWR.n4672 0.120292
R14780 VPWR.n4676 VPWR.n4674 0.120292
R14781 VPWR.n366 VPWR.n364 0.120292
R14782 VPWR.n360 VPWR.n359 0.120292
R14783 VPWR.n355 VPWR.n338 0.120292
R14784 VPWR.n351 VPWR.n338 0.120292
R14785 VPWR.n351 VPWR.n350 0.120292
R14786 VPWR.n346 VPWR.n345 0.120292
R14787 VPWR.n345 VPWR.n344 0.120292
R14788 VPWR.n1232 VPWR.n1231 0.120292
R14789 VPWR.n1237 VPWR.n1235 0.120292
R14790 VPWR.n1239 VPWR.n1237 0.120292
R14791 VPWR.n1240 VPWR.n1239 0.120292
R14792 VPWR.n1245 VPWR.n1244 0.120292
R14793 VPWR.n1250 VPWR.n1248 0.120292
R14794 VPWR.n1256 VPWR.n1253 0.120292
R14795 VPWR.n1312 VPWR.n1310 0.120292
R14796 VPWR.n1314 VPWR.n1312 0.120292
R14797 VPWR.n1317 VPWR.n1314 0.120292
R14798 VPWR.n1319 VPWR.n1317 0.120292
R14799 VPWR.n1321 VPWR.n1319 0.120292
R14800 VPWR.n1322 VPWR.n1321 0.120292
R14801 VPWR.n1328 VPWR.n1326 0.120292
R14802 VPWR.n1329 VPWR.n1328 0.120292
R14803 VPWR.n1335 VPWR.n1333 0.120292
R14804 VPWR.n1339 VPWR.n1335 0.120292
R14805 VPWR.n1340 VPWR.n1339 0.120292
R14806 VPWR.n1346 VPWR.n1345 0.120292
R14807 VPWR.n1348 VPWR.n1346 0.120292
R14808 VPWR.n1350 VPWR.n1348 0.120292
R14809 VPWR.n1353 VPWR.n1350 0.120292
R14810 VPWR.n1355 VPWR.n1353 0.120292
R14811 VPWR.n1357 VPWR.n1355 0.120292
R14812 VPWR.n1358 VPWR.n1357 0.120292
R14813 VPWR.n1363 VPWR.n1361 0.120292
R14814 VPWR.n1364 VPWR.n1363 0.120292
R14815 VPWR.n1368 VPWR.n441 0.120292
R14816 VPWR.n440 VPWR.n439 0.120292
R14817 VPWR.n1377 VPWR.n439 0.120292
R14818 VPWR.n1379 VPWR.n1378 0.120292
R14819 VPWR.n1426 VPWR.n1424 0.120292
R14820 VPWR.n4387 VPWR.n4386 0.120292
R14821 VPWR.n4381 VPWR.n4380 0.120292
R14822 VPWR.n4377 VPWR.n4376 0.120292
R14823 VPWR.n4376 VPWR.n4374 0.120292
R14824 VPWR.n4374 VPWR.n4372 0.120292
R14825 VPWR.n4372 VPWR.n4371 0.120292
R14826 VPWR.n4371 VPWR.n4370 0.120292
R14827 VPWR.n4370 VPWR.n4368 0.120292
R14828 VPWR.n4368 VPWR.n4367 0.120292
R14829 VPWR.n4363 VPWR.n4362 0.120292
R14830 VPWR.n4357 VPWR.n4356 0.120292
R14831 VPWR.n4356 VPWR.n4355 0.120292
R14832 VPWR.n4351 VPWR.n4350 0.120292
R14833 VPWR.n4345 VPWR.n4344 0.120292
R14834 VPWR.n4344 VPWR.n4342 0.120292
R14835 VPWR.n4342 VPWR.n4340 0.120292
R14836 VPWR.n4340 VPWR.n4338 0.120292
R14837 VPWR.n4338 VPWR.n4335 0.120292
R14838 VPWR.n4335 VPWR.n4333 0.120292
R14839 VPWR.n4333 VPWR.n4331 0.120292
R14840 VPWR.n4331 VPWR.n4329 0.120292
R14841 VPWR.n4329 VPWR.n4327 0.120292
R14842 VPWR.n3810 VPWR.n3808 0.120292
R14843 VPWR.n3811 VPWR.n3810 0.120292
R14844 VPWR.n3863 VPWR.n3862 0.120292
R14845 VPWR.n3862 VPWR.n3860 0.120292
R14846 VPWR.n3849 VPWR.n3848 0.120292
R14847 VPWR.n3848 VPWR.n3846 0.120292
R14848 VPWR.n3846 VPWR.n3844 0.120292
R14849 VPWR.n3844 VPWR.n3842 0.120292
R14850 VPWR.n3842 VPWR.n3841 0.120292
R14851 VPWR.n3841 VPWR.n3839 0.120292
R14852 VPWR.n3835 VPWR.n3834 0.120292
R14853 VPWR.n3834 VPWR.n3832 0.120292
R14854 VPWR.n3832 VPWR.n3831 0.120292
R14855 VPWR.n3831 VPWR.n3830 0.120292
R14856 VPWR.n3830 VPWR.n3829 0.120292
R14857 VPWR.n3875 VPWR.n3873 0.120292
R14858 VPWR.n3883 VPWR.n3875 0.120292
R14859 VPWR.n3923 VPWR.n3918 0.120292
R14860 VPWR.n3915 VPWR.n3914 0.120292
R14861 VPWR.n3914 VPWR.n3912 0.120292
R14862 VPWR.n3904 VPWR.n3903 0.120292
R14863 VPWR.n3898 VPWR.n3896 0.120292
R14864 VPWR.n3896 VPWR.n3894 0.120292
R14865 VPWR.n3894 VPWR.n3892 0.120292
R14866 VPWR.n3892 VPWR.n3890 0.120292
R14867 VPWR.n1855 VPWR.n1854 0.120292
R14868 VPWR.n1861 VPWR.n1844 0.120292
R14869 VPWR.n1866 VPWR.n1844 0.120292
R14870 VPWR.n1874 VPWR.n1873 0.120292
R14871 VPWR.n1882 VPWR.n1879 0.120292
R14872 VPWR.n1949 VPWR.n1948 0.120292
R14873 VPWR.n1957 VPWR.n1956 0.120292
R14874 VPWR.n1958 VPWR.n1957 0.120292
R14875 VPWR.n1965 VPWR.n1963 0.120292
R14876 VPWR.n1967 VPWR.n1965 0.120292
R14877 VPWR.n1969 VPWR.n1967 0.120292
R14878 VPWR.n1972 VPWR.n1969 0.120292
R14879 VPWR.n1974 VPWR.n1972 0.120292
R14880 VPWR.n1976 VPWR.n1974 0.120292
R14881 VPWR.n1978 VPWR.n1976 0.120292
R14882 VPWR.n1980 VPWR.n1978 0.120292
R14883 VPWR.n1982 VPWR.n1980 0.120292
R14884 VPWR.n1984 VPWR.n1982 0.120292
R14885 VPWR.n1985 VPWR.n1984 0.120292
R14886 VPWR.n1990 VPWR.n1988 0.120292
R14887 VPWR.n1992 VPWR.n1990 0.120292
R14888 VPWR.n1994 VPWR.n1992 0.120292
R14889 VPWR.n1996 VPWR.n1994 0.120292
R14890 VPWR.n1998 VPWR.n1996 0.120292
R14891 VPWR.n2003 VPWR.n2002 0.120292
R14892 VPWR.n2004 VPWR.n2003 0.120292
R14893 VPWR.n2005 VPWR.n2004 0.120292
R14894 VPWR.n2014 VPWR.n2013 0.120292
R14895 VPWR.n4231 VPWR.n4229 0.120292
R14896 VPWR.n4229 VPWR.n4228 0.120292
R14897 VPWR.n4225 VPWR.n4224 0.120292
R14898 VPWR.n4224 VPWR.n4222 0.120292
R14899 VPWR.n4222 VPWR.n4220 0.120292
R14900 VPWR.n4220 VPWR.n4219 0.120292
R14901 VPWR.n4214 VPWR.n4210 0.120292
R14902 VPWR.n4210 VPWR.n4209 0.120292
R14903 VPWR.n4209 VPWR.n4208 0.120292
R14904 VPWR.n4208 VPWR.n4206 0.120292
R14905 VPWR.n4203 VPWR.n4202 0.120292
R14906 VPWR.n4193 VPWR.n4192 0.120292
R14907 VPWR.n4192 VPWR.n4190 0.120292
R14908 VPWR.n4190 VPWR.n4188 0.120292
R14909 VPWR.n4185 VPWR.n4184 0.120292
R14910 VPWR.n4184 VPWR.n4182 0.120292
R14911 VPWR.n4117 VPWR.n4116 0.120292
R14912 VPWR.n4116 VPWR.n4114 0.120292
R14913 VPWR.n4104 VPWR.n4103 0.120292
R14914 VPWR.n4103 VPWR.n4102 0.120292
R14915 VPWR.n4102 VPWR.n4101 0.120292
R14916 VPWR.n4101 VPWR.n4100 0.120292
R14917 VPWR.n4100 VPWR.n4099 0.120292
R14918 VPWR.n4096 VPWR.n4094 0.120292
R14919 VPWR.n4094 VPWR.n4092 0.120292
R14920 VPWR.n4092 VPWR.n4090 0.120292
R14921 VPWR.n4090 VPWR.n4089 0.120292
R14922 VPWR.n4089 VPWR.n4087 0.120292
R14923 VPWR.n4082 VPWR.n4080 0.120292
R14924 VPWR.n4080 VPWR.n4079 0.120292
R14925 VPWR.n4079 VPWR.n4078 0.120292
R14926 VPWR.n4071 VPWR.n1537 0.120292
R14927 VPWR.n4069 VPWR.n4068 0.120292
R14928 VPWR.n4028 VPWR.n4027 0.120292
R14929 VPWR.n4027 VPWR.n4025 0.120292
R14930 VPWR.n4025 VPWR.n4023 0.120292
R14931 VPWR.n4023 VPWR.n4021 0.120292
R14932 VPWR.n4018 VPWR.n4017 0.120292
R14933 VPWR.n4017 VPWR.n4015 0.120292
R14934 VPWR.n4015 VPWR.n4013 0.120292
R14935 VPWR.n4013 VPWR.n4011 0.120292
R14936 VPWR.n4011 VPWR.n4009 0.120292
R14937 VPWR.n4009 VPWR.n4007 0.120292
R14938 VPWR.n4003 VPWR.n4002 0.120292
R14939 VPWR.n4002 VPWR.n4001 0.120292
R14940 VPWR.n4001 VPWR.n4000 0.120292
R14941 VPWR.n1679 VPWR.n1677 0.120292
R14942 VPWR.n1680 VPWR.n1679 0.120292
R14943 VPWR.n1685 VPWR.n1683 0.120292
R14944 VPWR.n1686 VPWR.n1685 0.120292
R14945 VPWR.n1691 VPWR.n1689 0.120292
R14946 VPWR.n1693 VPWR.n1691 0.120292
R14947 VPWR.n1695 VPWR.n1693 0.120292
R14948 VPWR.n1697 VPWR.n1695 0.120292
R14949 VPWR.n1699 VPWR.n1698 0.120292
R14950 VPWR.n1704 VPWR.n1702 0.120292
R14951 VPWR.n1706 VPWR.n1704 0.120292
R14952 VPWR.n1708 VPWR.n1706 0.120292
R14953 VPWR.n1797 VPWR.n1732 0.120292
R14954 VPWR.n1736 VPWR.n1732 0.120292
R14955 VPWR.n1790 VPWR.n1788 0.120292
R14956 VPWR.n1785 VPWR.n1784 0.120292
R14957 VPWR.n1784 VPWR.n1782 0.120292
R14958 VPWR.n1782 VPWR.n1780 0.120292
R14959 VPWR.n1780 VPWR.n1778 0.120292
R14960 VPWR.n1778 VPWR.n1775 0.120292
R14961 VPWR.n1775 VPWR.n1773 0.120292
R14962 VPWR.n1773 VPWR.n1771 0.120292
R14963 VPWR.n1771 VPWR.n1769 0.120292
R14964 VPWR.n1769 VPWR.n1767 0.120292
R14965 VPWR.n1767 VPWR.n1765 0.120292
R14966 VPWR.n1765 VPWR.n1763 0.120292
R14967 VPWR.n1760 VPWR.n1759 0.120292
R14968 VPWR.n1759 VPWR.n1758 0.120292
R14969 VPWR.n1758 VPWR.n1757 0.120292
R14970 VPWR.n1756 VPWR.n1755 0.120292
R14971 VPWR.n1755 VPWR.n1754 0.120292
R14972 VPWR.n1751 VPWR.n1750 0.120292
R14973 VPWR.n2118 VPWR.n2117 0.120292
R14974 VPWR.n2117 VPWR.n2116 0.120292
R14975 VPWR.n1629 VPWR.n1627 0.120292
R14976 VPWR.n1627 VPWR.n1625 0.120292
R14977 VPWR.n1625 VPWR.n1623 0.120292
R14978 VPWR.n1623 VPWR.n1621 0.120292
R14979 VPWR.n1621 VPWR.n1619 0.120292
R14980 VPWR.n1619 VPWR.n1617 0.120292
R14981 VPWR.n1617 VPWR.n1615 0.120292
R14982 VPWR.n1615 VPWR.n1613 0.120292
R14983 VPWR.n1613 VPWR.n1611 0.120292
R14984 VPWR.n1611 VPWR.n1609 0.120292
R14985 VPWR.n1609 VPWR.n1607 0.120292
R14986 VPWR.n1607 VPWR.n1605 0.120292
R14987 VPWR.n1604 VPWR.n1599 0.120292
R14988 VPWR.n1599 VPWR.n1598 0.120292
R14989 VPWR.n1598 VPWR.n1597 0.120292
R14990 VPWR.n2130 VPWR.n2128 0.120292
R14991 VPWR.n2132 VPWR.n2130 0.120292
R14992 VPWR.n2134 VPWR.n2132 0.120292
R14993 VPWR.n2137 VPWR.n2134 0.120292
R14994 VPWR.n2139 VPWR.n2137 0.120292
R14995 VPWR.n2140 VPWR.n2139 0.120292
R14996 VPWR.n2148 VPWR.n2147 0.120292
R14997 VPWR.n2149 VPWR.n2148 0.120292
R14998 VPWR.n2150 VPWR.n2149 0.120292
R14999 VPWR.n2156 VPWR.n2154 0.120292
R15000 VPWR.n3587 VPWR.n3585 0.120292
R15001 VPWR.n3595 VPWR.n3594 0.120292
R15002 VPWR.n3597 VPWR.n3595 0.120292
R15003 VPWR.n3599 VPWR.n3597 0.120292
R15004 VPWR.n3608 VPWR.n3607 0.120292
R15005 VPWR.n3609 VPWR.n3608 0.120292
R15006 VPWR.n3611 VPWR.n3609 0.120292
R15007 VPWR.n3613 VPWR.n3611 0.120292
R15008 VPWR.n3615 VPWR.n3613 0.120292
R15009 VPWR.n3617 VPWR.n3615 0.120292
R15010 VPWR.n3622 VPWR.n1576 0.120292
R15011 VPWR.n3623 VPWR.n3622 0.120292
R15012 VPWR.n3624 VPWR.n3623 0.120292
R15013 VPWR.n3629 VPWR.n3627 0.120292
R15014 VPWR.n3631 VPWR.n3629 0.120292
R15015 VPWR.n3632 VPWR.n3631 0.120292
R15016 VPWR.n3633 VPWR.n3632 0.120292
R15017 VPWR.n3634 VPWR.n3633 0.120292
R15018 VPWR.n3640 VPWR.n3638 0.120292
R15019 VPWR.n3678 VPWR.n3672 0.120292
R15020 VPWR.n3672 VPWR.n3671 0.120292
R15021 VPWR.n3671 VPWR.n3670 0.120292
R15022 VPWR.n3670 VPWR.n3668 0.120292
R15023 VPWR.n3668 VPWR.n3665 0.120292
R15024 VPWR.n3661 VPWR.n3660 0.120292
R15025 VPWR.n3656 VPWR.n3655 0.120292
R15026 VPWR.n3652 VPWR.n3651 0.120292
R15027 VPWR.n3651 VPWR.n3650 0.120292
R15028 VPWR.n2699 VPWR.n2698 0.120292
R15029 VPWR.n2700 VPWR.n2699 0.120292
R15030 VPWR.n2704 VPWR.n2703 0.120292
R15031 VPWR.n2705 VPWR.n2704 0.120292
R15032 VPWR.n2710 VPWR.n2705 0.120292
R15033 VPWR.n2723 VPWR.n2720 0.120292
R15034 VPWR.n2985 VPWR.n2984 0.120292
R15035 VPWR.n2980 VPWR.n2979 0.120292
R15036 VPWR.n2975 VPWR.n2973 0.120292
R15037 VPWR.n2973 VPWR.n2972 0.120292
R15038 VPWR.n2972 VPWR.n2971 0.120292
R15039 VPWR.n2968 VPWR.n2967 0.120292
R15040 VPWR.n2967 VPWR.n2965 0.120292
R15041 VPWR.n2965 VPWR.n2963 0.120292
R15042 VPWR.n2963 VPWR.n2961 0.120292
R15043 VPWR.n2961 VPWR.n2958 0.120292
R15044 VPWR.n2958 VPWR.n2956 0.120292
R15045 VPWR.n2956 VPWR.n2954 0.120292
R15046 VPWR.n2954 VPWR.n2952 0.120292
R15047 VPWR.n2952 VPWR.n2950 0.120292
R15048 VPWR.n2950 VPWR.n2948 0.120292
R15049 VPWR.n2948 VPWR.n2946 0.120292
R15050 VPWR.n2941 VPWR.n2940 0.120292
R15051 VPWR.n2940 VPWR.n2938 0.120292
R15052 VPWR.n2938 VPWR.n2937 0.120292
R15053 VPWR.n2937 VPWR.n2935 0.120292
R15054 VPWR.n2935 VPWR.n2933 0.120292
R15055 VPWR.n2819 VPWR.n2817 0.120292
R15056 VPWR.n2855 VPWR.n2854 0.120292
R15057 VPWR.n2861 VPWR.n2860 0.120292
R15058 VPWR.n2862 VPWR.n2861 0.120292
R15059 VPWR.n2864 VPWR.n2862 0.120292
R15060 VPWR.n2866 VPWR.n2864 0.120292
R15061 VPWR.n2867 VPWR.n2866 0.120292
R15062 VPWR.n2872 VPWR.n2870 0.120292
R15063 VPWR.n2874 VPWR.n2872 0.120292
R15064 VPWR.n2876 VPWR.n2874 0.120292
R15065 VPWR.n2879 VPWR.n2876 0.120292
R15066 VPWR.n2880 VPWR.n2879 0.120292
R15067 VPWR.n2886 VPWR.n2884 0.120292
R15068 VPWR.n2888 VPWR.n2886 0.120292
R15069 VPWR.n2890 VPWR.n2888 0.120292
R15070 VPWR.n2891 VPWR.n2890 0.120292
R15071 VPWR.n2923 VPWR.n2922 0.120292
R15072 VPWR.n2922 VPWR.n2921 0.120292
R15073 VPWR.n2921 VPWR.n2920 0.120292
R15074 VPWR.n2917 VPWR.n2916 0.120292
R15075 VPWR.n2916 VPWR.n2914 0.120292
R15076 VPWR.n2914 VPWR.n2912 0.120292
R15077 VPWR.n2912 VPWR.n2910 0.120292
R15078 VPWR.n2910 VPWR.n2907 0.120292
R15079 VPWR.n2907 VPWR.n2905 0.120292
R15080 VPWR.n2905 VPWR.n2903 0.120292
R15081 VPWR.n2900 VPWR.n2899 0.120292
R15082 VPWR.n3450 VPWR.n3448 0.120292
R15083 VPWR.n3448 VPWR.n3446 0.120292
R15084 VPWR.n3446 VPWR.n3444 0.120292
R15085 VPWR.n3444 VPWR.n3442 0.120292
R15086 VPWR.n2219 VPWR.n2218 0.120292
R15087 VPWR.n2224 VPWR.n2222 0.120292
R15088 VPWR.n2226 VPWR.n2224 0.120292
R15089 VPWR.n2228 VPWR.n2226 0.120292
R15090 VPWR.n2231 VPWR.n2228 0.120292
R15091 VPWR.n2233 VPWR.n2231 0.120292
R15092 VPWR.n2236 VPWR.n2233 0.120292
R15093 VPWR.n2239 VPWR.n2237 0.120292
R15094 VPWR.n2240 VPWR.n2239 0.120292
R15095 VPWR.n2241 VPWR.n2240 0.120292
R15096 VPWR.n2242 VPWR.n2241 0.120292
R15097 VPWR.n2248 VPWR.n2246 0.120292
R15098 VPWR.n2250 VPWR.n2248 0.120292
R15099 VPWR.n2252 VPWR.n2250 0.120292
R15100 VPWR.n2255 VPWR.n2252 0.120292
R15101 VPWR.n2257 VPWR.n2255 0.120292
R15102 VPWR.n2259 VPWR.n2257 0.120292
R15103 VPWR.n2261 VPWR.n2259 0.120292
R15104 VPWR.n2263 VPWR.n2261 0.120292
R15105 VPWR.n2265 VPWR.n2263 0.120292
R15106 VPWR.n2267 VPWR.n2265 0.120292
R15107 VPWR.n2268 VPWR.n2267 0.120292
R15108 VPWR.n3434 VPWR.n3432 0.120292
R15109 VPWR.n3432 VPWR.n3430 0.120292
R15110 VPWR.n3430 VPWR.n3428 0.120292
R15111 VPWR.n2329 VPWR.n2324 0.120292
R15112 VPWR.n2324 VPWR.n2322 0.120292
R15113 VPWR.n2322 VPWR.n2320 0.120292
R15114 VPWR.n2320 VPWR.n2318 0.120292
R15115 VPWR.n2315 VPWR.n2314 0.120292
R15116 VPWR.n2314 VPWR.n2313 0.120292
R15117 VPWR.n2313 VPWR.n2311 0.120292
R15118 VPWR.n2311 VPWR.n2309 0.120292
R15119 VPWR.n2309 VPWR.n2306 0.120292
R15120 VPWR.n2306 VPWR.n2304 0.120292
R15121 VPWR.n2304 VPWR.n2302 0.120292
R15122 VPWR.n2302 VPWR.n2300 0.120292
R15123 VPWR.n2300 VPWR.n2298 0.120292
R15124 VPWR.n2298 VPWR.n2296 0.120292
R15125 VPWR.n2296 VPWR.n2294 0.120292
R15126 VPWR.n6387 VPWR.n6385 0.120292
R15127 VPWR.n6388 VPWR.n6387 0.120292
R15128 VPWR.n6394 VPWR.n6393 0.120292
R15129 VPWR.n6398 VPWR.n6397 0.120292
R15130 VPWR.n6408 VPWR.n6403 0.120292
R15131 VPWR.n6462 VPWR.n6460 0.120292
R15132 VPWR.n6464 VPWR.n6462 0.120292
R15133 VPWR.n6467 VPWR.n6464 0.120292
R15134 VPWR.n6469 VPWR.n6467 0.120292
R15135 VPWR.n6471 VPWR.n6469 0.120292
R15136 VPWR.n6473 VPWR.n6471 0.120292
R15137 VPWR.n6485 VPWR.n6484 0.120292
R15138 VPWR.n6487 VPWR.n6485 0.120292
R15139 VPWR.n6489 VPWR.n6487 0.120292
R15140 VPWR.n6492 VPWR.n6489 0.120292
R15141 VPWR.n6494 VPWR.n6492 0.120292
R15142 VPWR.n6495 VPWR.n6494 0.120292
R15143 VPWR.n6496 VPWR.n6495 0.120292
R15144 VPWR.n6502 VPWR.n6500 0.120292
R15145 VPWR.n6503 VPWR.n6502 0.120292
R15146 VPWR.n6504 VPWR.n6503 0.120292
R15147 VPWR.n6510 VPWR.n6508 0.120292
R15148 VPWR.n6512 VPWR.n6510 0.120292
R15149 VPWR.n6514 VPWR.n6512 0.120292
R15150 VPWR.n6517 VPWR.n6514 0.120292
R15151 VPWR.n6519 VPWR.n6517 0.120292
R15152 VPWR.n6520 VPWR.n6519 0.120292
R15153 VPWR.n6521 VPWR.n6520 0.120292
R15154 VPWR.n6526 VPWR.n6525 0.120292
R15155 VPWR.n6527 VPWR.n6526 0.120292
R15156 VPWR.n4983 VPWR.n4978 0.120292
R15157 VPWR.n4985 VPWR.n4983 0.120292
R15158 VPWR.n4987 VPWR.n4985 0.120292
R15159 VPWR.n4988 VPWR.n4987 0.120292
R15160 VPWR.n4993 VPWR.n4992 0.120292
R15161 VPWR.n4994 VPWR.n4993 0.120292
R15162 VPWR.n5000 VPWR.n4998 0.120292
R15163 VPWR.n5002 VPWR.n5000 0.120292
R15164 VPWR.n5009 VPWR.n5007 0.120292
R15165 VPWR.n5010 VPWR.n5009 0.120292
R15166 VPWR.n5015 VPWR.n5013 0.120292
R15167 VPWR.n5052 VPWR.n5050 0.120292
R15168 VPWR.n5050 VPWR.n5048 0.120292
R15169 VPWR.n5048 VPWR.n5045 0.120292
R15170 VPWR.n5045 VPWR.n5043 0.120292
R15171 VPWR.n5043 VPWR.n5041 0.120292
R15172 VPWR.n5041 VPWR.n5040 0.120292
R15173 VPWR.n5040 VPWR.n5039 0.120292
R15174 VPWR.n5036 VPWR.n5035 0.120292
R15175 VPWR.n5035 VPWR.n5033 0.120292
R15176 VPWR.n5029 VPWR.n5028 0.120292
R15177 VPWR.n5028 VPWR.n5027 0.120292
R15178 VPWR.n7718 VPWR.n32 0.120292
R15179 VPWR.n7714 VPWR.n7713 0.120292
R15180 VPWR.n7713 VPWR.n7711 0.120292
R15181 VPWR.n7708 VPWR.n7707 0.120292
R15182 VPWR.n7707 VPWR.n7706 0.120292
R15183 VPWR.n7706 VPWR.n7705 0.120292
R15184 VPWR.n7702 VPWR.n7701 0.120292
R15185 VPWR.n7701 VPWR.n7699 0.120292
R15186 VPWR.n7695 VPWR.n7694 0.120292
R15187 VPWR.n7694 VPWR.n7693 0.120292
R15188 VPWR.n7693 VPWR.n7692 0.120292
R15189 VPWR.n7689 VPWR.n7688 0.120292
R15190 VPWR.n7688 VPWR.n7687 0.120292
R15191 VPWR.n7682 VPWR.n7680 0.120292
R15192 VPWR.n7680 VPWR.n7678 0.120292
R15193 VPWR.n7678 VPWR.n7677 0.120292
R15194 VPWR.n7677 VPWR.n7676 0.120292
R15195 VPWR.n7672 VPWR.n7671 0.120292
R15196 VPWR.n80 VPWR.n77 0.120292
R15197 VPWR.n74 VPWR.n73 0.120292
R15198 VPWR.n73 VPWR.n71 0.120292
R15199 VPWR.n71 VPWR.n69 0.120292
R15200 VPWR.n64 VPWR.n62 0.120292
R15201 VPWR.n58 VPWR.n56 0.120292
R15202 VPWR.n2586 VPWR.n2580 0.120292
R15203 VPWR.n2587 VPWR.n2586 0.120292
R15204 VPWR.n2588 VPWR.n2587 0.120292
R15205 VPWR.n2578 VPWR.n2577 0.120292
R15206 VPWR.n2599 VPWR.n2597 0.120292
R15207 VPWR.n2601 VPWR.n2599 0.120292
R15208 VPWR.n2605 VPWR.n2601 0.120292
R15209 VPWR.n2607 VPWR.n2606 0.120292
R15210 VPWR.n2608 VPWR.n2607 0.120292
R15211 VPWR.n2613 VPWR.n2611 0.120292
R15212 VPWR.n2575 VPWR.n2573 0.120292
R15213 VPWR.n2573 VPWR.n2571 0.120292
R15214 VPWR.n2571 VPWR.n2569 0.120292
R15215 VPWR.n2569 VPWR.n2567 0.120292
R15216 VPWR.n2567 VPWR.n2565 0.120292
R15217 VPWR.n2565 VPWR.n2563 0.120292
R15218 VPWR.n2557 VPWR.n2556 0.120292
R15219 VPWR.n2553 VPWR.n2552 0.120292
R15220 VPWR.n2551 VPWR.n2509 0.120292
R15221 VPWR.n2547 VPWR.n2509 0.120292
R15222 VPWR.n2547 VPWR.n2546 0.120292
R15223 VPWR.n2546 VPWR.n2545 0.120292
R15224 VPWR.n2545 VPWR.n2512 0.120292
R15225 VPWR.n2541 VPWR.n2512 0.120292
R15226 VPWR.n2541 VPWR.n2540 0.120292
R15227 VPWR.n2539 VPWR.n2515 0.120292
R15228 VPWR.n2535 VPWR.n2515 0.120292
R15229 VPWR.n2535 VPWR.n2534 0.120292
R15230 VPWR.n2532 VPWR.n2518 0.120292
R15231 VPWR.n2527 VPWR.n2525 0.120292
R15232 VPWR.n2525 VPWR.n2523 0.120292
R15233 VPWR.n2522 VPWR.n2521 0.120292
R15234 VPWR.n2449 VPWR.n2448 0.120292
R15235 VPWR.n2448 VPWR.n2447 0.120292
R15236 VPWR.n2447 VPWR.n2446 0.120292
R15237 VPWR.n2446 VPWR.n2444 0.120292
R15238 VPWR.n2441 VPWR.n2440 0.120292
R15239 VPWR.n2440 VPWR.n2439 0.120292
R15240 VPWR.n3127 VPWR.n3125 0.120292
R15241 VPWR.n3129 VPWR.n3127 0.120292
R15242 VPWR.n3132 VPWR.n3129 0.120292
R15243 VPWR.n3134 VPWR.n3132 0.120292
R15244 VPWR.n3136 VPWR.n3134 0.120292
R15245 VPWR.n3149 VPWR.n3143 0.120292
R15246 VPWR.n3151 VPWR.n3149 0.120292
R15247 VPWR.n3220 VPWR.n3218 0.120292
R15248 VPWR.n3222 VPWR.n3220 0.120292
R15249 VPWR.n3224 VPWR.n3222 0.120292
R15250 VPWR.n3225 VPWR.n3224 0.120292
R15251 VPWR.n3280 VPWR.n3271 0.120292
R15252 VPWR.n3271 VPWR.n3270 0.120292
R15253 VPWR.n3270 VPWR.n3269 0.120292
R15254 VPWR.n3269 VPWR.n3268 0.120292
R15255 VPWR.n3268 VPWR.n3266 0.120292
R15256 VPWR.n3262 VPWR.n3261 0.120292
R15257 VPWR.n3261 VPWR.n3260 0.120292
R15258 VPWR.n3260 VPWR.n3258 0.120292
R15259 VPWR.n3258 VPWR.n3256 0.120292
R15260 VPWR.n3256 VPWR.n3253 0.120292
R15261 VPWR.n3253 VPWR.n3251 0.120292
R15262 VPWR.n3251 VPWR.n3249 0.120292
R15263 VPWR.n3249 VPWR.n3247 0.120292
R15264 VPWR.n3247 VPWR.n3245 0.120292
R15265 VPWR.n3242 VPWR.n3241 0.120292
R15266 VPWR.n3233 VPWR.n3232 0.120292
R15267 VPWR.n3293 VPWR.n3291 0.120292
R15268 VPWR.n3295 VPWR.n3293 0.120292
R15269 VPWR.n3299 VPWR.n3295 0.120292
R15270 VPWR.n3329 VPWR.n3327 0.120292
R15271 VPWR.n3327 VPWR.n3325 0.120292
R15272 VPWR.n3325 VPWR.n3323 0.120292
R15273 VPWR.n3318 VPWR.n3316 0.120292
R15274 VPWR.n3310 VPWR.n3303 0.120292
R15275 VPWR.n3304 VPWR.n3303 0.120292
R15276 VPWR.n6290 VPWR.n6289 0.120292
R15277 VPWR.n6290 VPWR.n6283 0.120292
R15278 VPWR.n6294 VPWR.n6283 0.120292
R15279 VPWR.n6295 VPWR.n6294 0.120292
R15280 VPWR.n6296 VPWR.n6295 0.120292
R15281 VPWR.n6300 VPWR.n6281 0.120292
R15282 VPWR.n6302 VPWR.n6301 0.120292
R15283 VPWR.n6302 VPWR.n6279 0.120292
R15284 VPWR.n6308 VPWR.n6279 0.120292
R15285 VPWR.n6310 VPWR.n6309 0.120292
R15286 VPWR.n6311 VPWR.n6310 0.120292
R15287 VPWR.n6316 VPWR.n6314 0.120292
R15288 VPWR.n6277 VPWR.n6276 0.120292
R15289 VPWR.n6276 VPWR.n6274 0.120292
R15290 VPWR.n6274 VPWR.n6272 0.120292
R15291 VPWR.n6272 VPWR.n6270 0.120292
R15292 VPWR.n6270 VPWR.n6268 0.120292
R15293 VPWR.n6268 VPWR.n6266 0.120292
R15294 VPWR.n6262 VPWR.n6261 0.120292
R15295 VPWR.n6261 VPWR.n6259 0.120292
R15296 VPWR.n6259 VPWR.n6258 0.120292
R15297 VPWR.n6254 VPWR.n6253 0.120292
R15298 VPWR.n6253 VPWR.n5737 0.120292
R15299 VPWR.n6249 VPWR.n5737 0.120292
R15300 VPWR.n6248 VPWR.n6247 0.120292
R15301 VPWR.n6247 VPWR.n5740 0.120292
R15302 VPWR.n6243 VPWR.n5740 0.120292
R15303 VPWR.n6243 VPWR.n6242 0.120292
R15304 VPWR.n6242 VPWR.n5742 0.120292
R15305 VPWR.n6238 VPWR.n5742 0.120292
R15306 VPWR.n6238 VPWR.n6237 0.120292
R15307 VPWR.n6237 VPWR.n6236 0.120292
R15308 VPWR.n6236 VPWR.n5744 0.120292
R15309 VPWR.n6232 VPWR.n5744 0.120292
R15310 VPWR.n6232 VPWR.n6231 0.120292
R15311 VPWR.n6227 VPWR.n6226 0.120292
R15312 VPWR.n6226 VPWR.n6224 0.120292
R15313 VPWR.n6223 VPWR.n6221 0.120292
R15314 VPWR.n6217 VPWR.n6216 0.120292
R15315 VPWR.n6173 VPWR.n6172 0.120292
R15316 VPWR.n6172 VPWR.n6170 0.120292
R15317 VPWR.n6170 VPWR.n6168 0.120292
R15318 VPWR.n6168 VPWR.n6166 0.120292
R15319 VPWR.n6166 VPWR.n6164 0.120292
R15320 VPWR.n6164 VPWR.n6162 0.120292
R15321 VPWR.n6158 VPWR.n6157 0.120292
R15322 VPWR.n6157 VPWR.n5823 0.120292
R15323 VPWR.n6152 VPWR.n6151 0.120292
R15324 VPWR.n6151 VPWR.n5825 0.120292
R15325 VPWR.n6144 VPWR.n5825 0.120292
R15326 VPWR.n6144 VPWR.n6143 0.120292
R15327 VPWR.n6143 VPWR.n6142 0.120292
R15328 VPWR.n6142 VPWR.n5829 0.120292
R15329 VPWR VPWR.n5829 0.120292
R15330 VPWR.n6137 VPWR.n6047 0.120292
R15331 VPWR.n6132 VPWR.n6047 0.120292
R15332 VPWR.n6132 VPWR.n6131 0.120292
R15333 VPWR.n6130 VPWR.n6129 0.120292
R15334 VPWR.n6129 VPWR.n6050 0.120292
R15335 VPWR.n6125 VPWR.n6050 0.120292
R15336 VPWR.n6125 VPWR.n6124 0.120292
R15337 VPWR.n6124 VPWR.n6123 0.120292
R15338 VPWR.n6119 VPWR.n6118 0.120292
R15339 VPWR.n6118 VPWR.n6053 0.120292
R15340 VPWR.n6114 VPWR.n6053 0.120292
R15341 VPWR.n6113 VPWR.n6112 0.120292
R15342 VPWR.n6112 VPWR.n6111 0.120292
R15343 VPWR.n5841 VPWR.n5839 0.120292
R15344 VPWR.n5843 VPWR.n5841 0.120292
R15345 VPWR.n5845 VPWR.n5843 0.120292
R15346 VPWR.n5847 VPWR.n5845 0.120292
R15347 VPWR.n5856 VPWR.n5855 0.120292
R15348 VPWR.n5857 VPWR.n5856 0.120292
R15349 VPWR.n5858 VPWR.n5857 0.120292
R15350 VPWR.n5863 VPWR.n5861 0.120292
R15351 VPWR.n5865 VPWR.n5863 0.120292
R15352 VPWR.n5867 VPWR.n5865 0.120292
R15353 VPWR.n5870 VPWR.n5867 0.120292
R15354 VPWR.n5872 VPWR.n5870 0.120292
R15355 VPWR.n5874 VPWR.n5872 0.120292
R15356 VPWR.n5876 VPWR.n5874 0.120292
R15357 VPWR.n5878 VPWR.n5876 0.120292
R15358 VPWR.n5880 VPWR.n5878 0.120292
R15359 VPWR.n5882 VPWR.n5880 0.120292
R15360 VPWR.n5883 VPWR.n5882 0.120292
R15361 VPWR.n5888 VPWR.n5886 0.120292
R15362 VPWR.n5889 VPWR.n5888 0.120292
R15363 VPWR.n5895 VPWR.n5893 0.120292
R15364 VPWR.n5900 VPWR.n5895 0.120292
R15365 VPWR.n5902 VPWR.n5901 0.120292
R15366 VPWR.n5903 VPWR.n5902 0.120292
R15367 VPWR.n6040 VPWR.n6039 0.120292
R15368 VPWR.n6039 VPWR.n6036 0.120292
R15369 VPWR.n6036 VPWR.n6031 0.120292
R15370 VPWR.n6031 VPWR.n6028 0.120292
R15371 VPWR.n5954 VPWR.n5921 0.120292
R15372 VPWR.n5954 VPWR.n5953 0.120292
R15373 VPWR.n5948 VPWR.n5923 0.120292
R15374 VPWR.n5948 VPWR.n5947 0.120292
R15375 VPWR.n5947 VPWR.n5946 0.120292
R15376 VPWR.n5946 VPWR.n5925 0.120292
R15377 VPWR.n5940 VPWR.n5939 0.120292
R15378 VPWR.n5939 VPWR.n5928 0.120292
R15379 VPWR.n5935 VPWR.n5928 0.120292
R15380 VPWR.n5935 VPWR.n5934 0.120292
R15381 VPWR VPWR.n7525 0.12003
R15382 VPWR.n7525 VPWR 0.12003
R15383 VPWR VPWR.n4870 0.12003
R15384 VPWR.n4870 VPWR 0.12003
R15385 VPWR VPWR.n3827 0.12003
R15386 VPWR VPWR.n7663 0.12003
R15387 VPWR VPWR.n2558 0.12003
R15388 VPWR.n1054 VPWR.n1047 0.116104
R15389 VPWR.n3165 VPWR.n3164 0.113774
R15390 VPWR.n3920 VPWR.n3919 0.113774
R15391 VPWR.n2326 VPWR.n2325 0.113774
R15392 VPWR.n6747 VPWR.n6746 0.109682
R15393 VPWR.n6921 VPWR.n6919 0.109682
R15394 VPWR.n7196 VPWR.n7139 0.109682
R15395 VPWR.n869 VPWR.n820 0.109682
R15396 VPWR.n4550 VPWR.n4532 0.109682
R15397 VPWR.n4327 VPWR.n4325 0.109682
R15398 VPWR.n4173 VPWR.n4172 0.109682
R15399 VPWR.n3545 VPWR.n2156 0.109682
R15400 VPWR.n3487 VPWR.n2208 0.109682
R15401 VPWR.n3163 VPWR.n3151 0.109682
R15402 VPWR.n2075 VPWR.n1629 0.109342
R15403 VPWR.n2854 VPWR.n2852 0.109342
R15404 VPWR.n6567 VPWR.n4978 0.109342
R15405 VPWR.n6174 VPWR.n6173 0.109342
R15406 VPWR.n6991 VPWR.n6990 0.108642
R15407 VPWR.n4464 VPWR.n4462 0.108642
R15408 VPWR.n4388 VPWR.n4387 0.108642
R15409 VPWR.n4232 VPWR.n4231 0.108642
R15410 VPWR.n3072 VPWR.n2453 0.108642
R15411 VPWR.n5306 VPWR.n5303 0.107271
R15412 VPWR.n685 VPWR.n684 0.107271
R15413 VPWR.n1130 VPWR.n1128 0.107271
R15414 VPWR.n1424 VPWR.n1423 0.107271
R15415 VPWR.n2116 VPWR.n2114 0.107271
R15416 VPWR.n2821 VPWR.n2819 0.107271
R15417 VPWR.n6213 VPWR.n6212 0.107271
R15418 VPWR.n6332 VPWR.n6331 0.106285
R15419 VPWR.n2629 VPWR.n2628 0.106285
R15420 VPWR.n1069 VPWR.n1068 0.106285
R15421 VPWR.n7600 VPWR.n7599 0.105969
R15422 VPWR.n6866 VPWR.n6865 0.105969
R15423 VPWR.n4613 VPWR.n4611 0.105969
R15424 VPWR.n3808 VPWR.n3806 0.105969
R15425 VPWR.n3585 VPWR.n3583 0.105969
R15426 VPWR.n3452 VPWR.n3450 0.105969
R15427 VPWR.n3218 VPWR.n3216 0.105969
R15428 VPWR.n5839 VPWR.n5837 0.105969
R15429 VPWR.n626 VPWR.n625 0.105956
R15430 VPWR.n4859 VPWR.n299 0.105956
R15431 VPWR.n539 VPWR.n538 0.105956
R15432 VPWR.n4856 VPWR.n4855 0.105956
R15433 VPWR.n5094 VPWR 0.104136
R15434 VPWR.n5430 VPWR 0.104136
R15435 VPWR.n5352 VPWR 0.104136
R15436 VPWR.n480 VPWR 0.104136
R15437 VPWR.n1022 VPWR 0.104136
R15438 VPWR.n1228 VPWR 0.104136
R15439 VPWR.n1849 VPWR 0.104136
R15440 VPWR.n1674 VPWR 0.104136
R15441 VPWR.n2694 VPWR 0.104136
R15442 VPWR.n6381 VPWR 0.104136
R15443 VPWR.n2581 VPWR 0.104136
R15444 VPWR.n5932 VPWR 0.102383
R15445 VPWR.n7666 VPWR.n7665 0.102087
R15446 VPWR.n220 VPWR.n219 0.102087
R15447 VPWR.n6689 VPWR.n6688 0.102087
R15448 VPWR.n7425 VPWR.n7424 0.102087
R15449 VPWR.n698 VPWR.n697 0.102087
R15450 VPWR.n1567 VPWR.n1566 0.102087
R15451 VPWR.n5975 VPWR.n5974 0.102087
R15452 VPWR.n484 VPWR 0.0994583
R15453 VPWR.n4381 VPWR 0.0994583
R15454 VPWR.n5188 VPWR 0.0981562
R15455 VPWR VPWR.n5186 0.0981562
R15456 VPWR.n6705 VPWR 0.0981562
R15457 VPWR.n6625 VPWR 0.0981562
R15458 VPWR.n7534 VPWR 0.0981562
R15459 VPWR.n7559 VPWR 0.0981562
R15460 VPWR VPWR.n179 0.0981562
R15461 VPWR.n5435 VPWR 0.0981562
R15462 VPWR.n5446 VPWR 0.0981562
R15463 VPWR.n5559 VPWR 0.0981562
R15464 VPWR VPWR.n5556 0.0981562
R15465 VPWR.n5524 VPWR 0.0981562
R15466 VPWR.n5499 VPWR 0.0981562
R15467 VPWR VPWR.n6921 0.0981562
R15468 VPWR.n6806 VPWR 0.0981562
R15469 VPWR.n6840 VPWR 0.0981562
R15470 VPWR.n7448 VPWR 0.0981562
R15471 VPWR.n5362 VPWR 0.0981562
R15472 VPWR.n5278 VPWR 0.0981562
R15473 VPWR VPWR.n4871 0.0981562
R15474 VPWR.n7077 VPWR 0.0981562
R15475 VPWR.n7118 VPWR 0.0981562
R15476 VPWR.n7121 VPWR 0.0981562
R15477 VPWR.n7219 VPWR 0.0981562
R15478 VPWR VPWR.n7339 0.0981562
R15479 VPWR.n491 VPWR 0.0981562
R15480 VPWR.n498 VPWR 0.0981562
R15481 VPWR.n659 VPWR 0.0981562
R15482 VPWR.n906 VPWR 0.0981562
R15483 VPWR.n911 VPWR 0.0981562
R15484 VPWR.n4828 VPWR 0.0981562
R15485 VPWR.n4804 VPWR 0.0981562
R15486 VPWR.n1045 VPWR 0.0981562
R15487 VPWR VPWR.n1202 0.0981562
R15488 VPWR.n1177 VPWR 0.0981562
R15489 VPWR.n1152 VPWR 0.0981562
R15490 VPWR.n4494 VPWR 0.0981562
R15491 VPWR.n4525 VPWR 0.0981562
R15492 VPWR.n4529 VPWR 0.0981562
R15493 VPWR.n4621 VPWR 0.0981562
R15494 VPWR.n4664 VPWR 0.0981562
R15495 VPWR.n4669 VPWR 0.0981562
R15496 VPWR.n361 VPWR 0.0981562
R15497 VPWR VPWR.n360 0.0981562
R15498 VPWR.n346 VPWR 0.0981562
R15499 VPWR.n1361 VPWR 0.0981562
R15500 VPWR.n1369 VPWR 0.0981562
R15501 VPWR VPWR.n1368 0.0981562
R15502 VPWR VPWR.n3849 0.0981562
R15503 VPWR VPWR.n3835 0.0981562
R15504 VPWR.n3909 VPWR 0.0981562
R15505 VPWR VPWR.n3898 0.0981562
R15506 VPWR.n1854 VPWR 0.0981562
R15507 VPWR.n1859 VPWR 0.0981562
R15508 VPWR.n1873 VPWR 0.0981562
R15509 VPWR.n1956 VPWR 0.0981562
R15510 VPWR.n1988 VPWR 0.0981562
R15511 VPWR.n4118 VPWR 0.0981562
R15512 VPWR.n4104 VPWR 0.0981562
R15513 VPWR VPWR.n4069 0.0981562
R15514 VPWR.n1760 VPWR 0.0981562
R15515 VPWR VPWR.n1746 0.0981562
R15516 VPWR VPWR.n3661 0.0981562
R15517 VPWR VPWR.n3656 0.0981562
R15518 VPWR.n3652 VPWR 0.0981562
R15519 VPWR.n2715 VPWR 0.0981562
R15520 VPWR VPWR.n2985 0.0981562
R15521 VPWR VPWR.n2941 0.0981562
R15522 VPWR.n2884 VPWR 0.0981562
R15523 VPWR.n2927 VPWR 0.0981562
R15524 VPWR VPWR.n2208 0.0981562
R15525 VPWR.n2211 VPWR 0.0981562
R15526 VPWR.n2243 VPWR 0.0981562
R15527 VPWR.n3436 VPWR 0.0981562
R15528 VPWR.n6393 VPWR 0.0981562
R15529 VPWR.n6403 VPWR 0.0981562
R15530 VPWR.n6474 VPWR 0.0981562
R15531 VPWR.n6500 VPWR 0.0981562
R15532 VPWR.n6508 VPWR 0.0981562
R15533 VPWR.n6522 VPWR 0.0981562
R15534 VPWR.n4992 VPWR 0.0981562
R15535 VPWR.n4998 VPWR 0.0981562
R15536 VPWR.n5013 VPWR 0.0981562
R15537 VPWR VPWR.n59 0.0981562
R15538 VPWR VPWR.n2539 0.0981562
R15539 VPWR VPWR.n2533 0.0981562
R15540 VPWR VPWR.n2527 0.0981562
R15541 VPWR VPWR.n3113 0.0981562
R15542 VPWR.n2441 VPWR 0.0981562
R15543 VPWR.n3143 VPWR 0.0981562
R15544 VPWR.n3242 VPWR 0.0981562
R15545 VPWR.n3229 VPWR 0.0981562
R15546 VPWR.n3237 VPWR 0.0981562
R15547 VPWR.n3320 VPWR 0.0981562
R15548 VPWR VPWR.n3319 0.0981562
R15549 VPWR VPWR.n3318 0.0981562
R15550 VPWR.n6263 VPWR 0.0981562
R15551 VPWR VPWR.n6230 0.0981562
R15552 VPWR.n6227 VPWR 0.0981562
R15553 VPWR.n6159 VPWR 0.0981562
R15554 VPWR VPWR.n6158 0.0981562
R15555 VPWR.n5886 VPWR 0.0981562
R15556 VPWR.n5893 VPWR 0.0981562
R15557 VPWR.n5921 VPWR 0.0981562
R15558 VPWR.n5923 VPWR 0.0981562
R15559 VPWR VPWR.n5940 0.0981562
R15560 VPWR VPWR.n7456 0.0968542
R15561 VPWR VPWR.n7348 0.0968542
R15562 VPWR.n818 VPWR 0.0968542
R15563 VPWR.n4532 VPWR 0.0968542
R15564 VPWR.n4651 VPWR 0.0968542
R15565 VPWR VPWR.n1426 0.0968542
R15566 VPWR VPWR.n4351 0.0968542
R15567 VPWR VPWR.n3853 0.0968542
R15568 VPWR.n3904 VPWR 0.0968542
R15569 VPWR VPWR.n4173 0.0968542
R15570 VPWR.n2154 VPWR 0.0968542
R15571 VPWR VPWR.n64 0.0968542
R15572 VPWR.n3017 VPWR.n3002 0.0942472
R15573 VPWR.n3505 VPWR.n2206 0.0942472
R15574 VPWR.n3404 VPWR.n2371 0.0940635
R15575 VPWR VPWR.n5106 0.0930549
R15576 VPWR.n3281 VPWR 0.0930549
R15577 VPWR.n7783 VPWR 0.0875462
R15578 VPWR.n7522 VPWR.n7519 0.0863232
R15579 VPWR.n7297 VPWR.n7286 0.0863232
R15580 VPWR.n3950 VPWR.n3883 0.0863232
R15581 VPWR.n3428 VPWR.n3425 0.0863232
R15582 VPWR.n3363 VPWR.n3299 0.0863232
R15583 VPWR.n6028 VPWR.n6026 0.0863232
R15584 VPWR.n6574 VPWR.n6573 0.0859812
R15585 VPWR.n7634 VPWR.n7633 0.0859812
R15586 VPWR.n5687 VPWR.n5686 0.0859812
R15587 VPWR.n7637 VPWR.n128 0.0859812
R15588 VPWR.n5662 VPWR.n5203 0.0857946
R15589 VPWR.n5586 VPWR.n5574 0.0857946
R15590 VPWR.n1310 VPWR.n1308 0.0857946
R15591 VPWR.n1945 VPWR.n1944 0.0857946
R15592 VPWR.n6460 VPWR.n6458 0.0857946
R15593 VPWR.n6351 VPWR.n6277 0.0857946
R15594 VPWR VPWR.n6703 0.0851354
R15595 VPWR.n6530 VPWR 0.0851354
R15596 VPWR.n2648 VPWR.n2575 0.0850212
R15597 VPWR.n2457 VPWR 0.0830437
R15598 VPWR.n2391 VPWR 0.0830437
R15599 VPWR.n2677 VPWR 0.0830437
R15600 VPWR.n2378 VPWR 0.0830437
R15601 VPWR.n5163 VPWR 0.0826382
R15602 VPWR.n5557 VPWR 0.0826382
R15603 VPWR.n5498 VPWR 0.0826382
R15604 VPWR.n3825 VPWR 0.0826382
R15605 VPWR.n2896 VPWR 0.0826382
R15606 VPWR VPWR.n6478 0.0826382
R15607 VPWR.n3138 VPWR 0.0826382
R15608 VPWR.n3263 VPWR 0.0826382
R15609 VPWR.n4097 VPWR 0.0822696
R15610 VPWR.n1594 VPWR 0.0822696
R15611 VPWR.n2558 VPWR 0.0822696
R15612 VPWR VPWR.n1532 0.0813361
R15613 VPWR.n3936 VPWR.n3935 0.0760162
R15614 VPWR.n6573 VPWR.n6572 0.0660062
R15615 VPWR.n7634 VPWR.n130 0.0660062
R15616 VPWR.n5688 VPWR.n5687 0.0660062
R15617 VPWR.n7638 VPWR.n7637 0.0660062
R15618 VPWR.n6285 VPWR 0.0657573
R15619 VPWR.n5605 VPWR.n5604 0.0620385
R15620 VPWR.n5098 VPWR 0.0603958
R15621 VPWR.n5103 VPWR 0.0603958
R15622 VPWR.n5111 VPWR 0.0603958
R15623 VPWR.n5182 VPWR 0.0603958
R15624 VPWR.n5175 VPWR 0.0603958
R15625 VPWR.n5169 VPWR 0.0603958
R15626 VPWR VPWR.n5161 0.0603958
R15627 VPWR VPWR.n6653 0.0603958
R15628 VPWR.n6650 VPWR 0.0603958
R15629 VPWR VPWR.n4938 0.0603958
R15630 VPWR.n6711 VPWR 0.0603958
R15631 VPWR.n6736 VPWR 0.0603958
R15632 VPWR.n6740 VPWR 0.0603958
R15633 VPWR.n158 VPWR 0.0603958
R15634 VPWR.n7528 VPWR 0.0603958
R15635 VPWR.n7569 VPWR 0.0603958
R15636 VPWR VPWR.n7526 0.0603958
R15637 VPWR VPWR.n7524 0.0603958
R15638 VPWR VPWR.n7523 0.0603958
R15639 VPWR.n191 VPWR 0.0603958
R15640 VPWR VPWR.n190 0.0603958
R15641 VPWR.n180 VPWR 0.0603958
R15642 VPWR VPWR.n178 0.0603958
R15643 VPWR.n5431 VPWR 0.0603958
R15644 VPWR.n5432 VPWR 0.0603958
R15645 VPWR.n5442 VPWR 0.0603958
R15646 VPWR.n5443 VPWR 0.0603958
R15647 VPWR VPWR.n5456 0.0603958
R15648 VPWR.n5457 VPWR 0.0603958
R15649 VPWR.n5460 VPWR 0.0603958
R15650 VPWR VPWR.n5558 0.0603958
R15651 VPWR VPWR.n5537 0.0603958
R15652 VPWR VPWR.n5497 0.0603958
R15653 VPWR.n6981 VPWR 0.0603958
R15654 VPWR.n6971 VPWR 0.0603958
R15655 VPWR VPWR.n6970 0.0603958
R15656 VPWR.n6960 VPWR 0.0603958
R15657 VPWR VPWR.n6959 0.0603958
R15658 VPWR VPWR.n6954 0.0603958
R15659 VPWR.n6951 VPWR 0.0603958
R15660 VPWR VPWR.n6950 0.0603958
R15661 VPWR.n6944 VPWR 0.0603958
R15662 VPWR.n6923 VPWR 0.0603958
R15663 VPWR VPWR.n6922 0.0603958
R15664 VPWR.n6865 VPWR 0.0603958
R15665 VPWR VPWR.n6864 0.0603958
R15666 VPWR.n6797 VPWR 0.0603958
R15667 VPWR.n6804 VPWR 0.0603958
R15668 VPWR.n6815 VPWR 0.0603958
R15669 VPWR.n6818 VPWR 0.0603958
R15670 VPWR.n6824 VPWR 0.0603958
R15671 VPWR.n6837 VPWR 0.0603958
R15672 VPWR.n6851 VPWR 0.0603958
R15673 VPWR.n7406 VPWR 0.0603958
R15674 VPWR.n7463 VPWR 0.0603958
R15675 VPWR.n7457 VPWR 0.0603958
R15676 VPWR.n7455 VPWR 0.0603958
R15677 VPWR VPWR.n7454 0.0603958
R15678 VPWR VPWR.n7451 0.0603958
R15679 VPWR.n5355 VPWR 0.0603958
R15680 VPWR.n5359 VPWR 0.0603958
R15681 VPWR.n5364 VPWR 0.0603958
R15682 VPWR.n5367 VPWR 0.0603958
R15683 VPWR.n5375 VPWR 0.0603958
R15684 VPWR.n5380 VPWR 0.0603958
R15685 VPWR.n5234 VPWR 0.0603958
R15686 VPWR.n5239 VPWR 0.0603958
R15687 VPWR.n5250 VPWR 0.0603958
R15688 VPWR.n5253 VPWR 0.0603958
R15689 VPWR.n5256 VPWR 0.0603958
R15690 VPWR.n5274 VPWR 0.0603958
R15691 VPWR.n5275 VPWR 0.0603958
R15692 VPWR.n5279 VPWR 0.0603958
R15693 VPWR.n5283 VPWR 0.0603958
R15694 VPWR.n5285 VPWR 0.0603958
R15695 VPWR.n5308 VPWR 0.0603958
R15696 VPWR VPWR.n5307 0.0603958
R15697 VPWR.n7072 VPWR 0.0603958
R15698 VPWR.n7074 VPWR 0.0603958
R15699 VPWR VPWR.n7078 0.0603958
R15700 VPWR.n7079 VPWR 0.0603958
R15701 VPWR.n7087 VPWR 0.0603958
R15702 VPWR.n7095 VPWR 0.0603958
R15703 VPWR.n7096 VPWR 0.0603958
R15704 VPWR.n7097 VPWR 0.0603958
R15705 VPWR.n7100 VPWR 0.0603958
R15706 VPWR.n7117 VPWR 0.0603958
R15707 VPWR VPWR.n7121 0.0603958
R15708 VPWR.n7122 VPWR 0.0603958
R15709 VPWR VPWR.n7122 0.0603958
R15710 VPWR.n7123 VPWR 0.0603958
R15711 VPWR.n7126 VPWR 0.0603958
R15712 VPWR VPWR.n7224 0.0603958
R15713 VPWR.n7225 VPWR 0.0603958
R15714 VPWR VPWR.n7225 0.0603958
R15715 VPWR.n7226 VPWR 0.0603958
R15716 VPWR VPWR.n7270 0.0603958
R15717 VPWR.n7256 VPWR 0.0603958
R15718 VPWR VPWR.n7247 0.0603958
R15719 VPWR VPWR.n7246 0.0603958
R15720 VPWR.n7237 VPWR 0.0603958
R15721 VPWR.n7277 VPWR 0.0603958
R15722 VPWR.n7278 VPWR 0.0603958
R15723 VPWR.n7279 VPWR 0.0603958
R15724 VPWR.n7282 VPWR 0.0603958
R15725 VPWR.n7349 VPWR 0.0603958
R15726 VPWR.n7347 VPWR 0.0603958
R15727 VPWR.n7344 VPWR 0.0603958
R15728 VPWR.n7340 VPWR 0.0603958
R15729 VPWR VPWR.n7338 0.0603958
R15730 VPWR.n481 VPWR 0.0603958
R15731 VPWR VPWR.n486 0.0603958
R15732 VPWR.n488 VPWR 0.0603958
R15733 VPWR.n492 VPWR 0.0603958
R15734 VPWR VPWR.n503 0.0603958
R15735 VPWR.n504 VPWR 0.0603958
R15736 VPWR.n507 VPWR 0.0603958
R15737 VPWR.n574 VPWR 0.0603958
R15738 VPWR.n647 VPWR 0.0603958
R15739 VPWR.n656 VPWR 0.0603958
R15740 VPWR.n663 VPWR 0.0603958
R15741 VPWR.n672 VPWR 0.0603958
R15742 VPWR.n678 VPWR 0.0603958
R15743 VPWR.n679 VPWR 0.0603958
R15744 VPWR VPWR.n679 0.0603958
R15745 VPWR.n680 VPWR 0.0603958
R15746 VPWR.n684 VPWR 0.0603958
R15747 VPWR.n745 VPWR 0.0603958
R15748 VPWR.n750 VPWR 0.0603958
R15749 VPWR VPWR.n603 0.0603958
R15750 VPWR.n757 VPWR 0.0603958
R15751 VPWR.n763 VPWR 0.0603958
R15752 VPWR.n768 VPWR 0.0603958
R15753 VPWR.n783 VPWR 0.0603958
R15754 VPWR.n785 VPWR 0.0603958
R15755 VPWR.n810 VPWR 0.0603958
R15756 VPWR.n815 VPWR 0.0603958
R15757 VPWR.n889 VPWR 0.0603958
R15758 VPWR VPWR.n891 0.0603958
R15759 VPWR.n893 VPWR 0.0603958
R15760 VPWR.n898 VPWR 0.0603958
R15761 VPWR.n901 VPWR 0.0603958
R15762 VPWR.n905 VPWR 0.0603958
R15763 VPWR VPWR.n581 0.0603958
R15764 VPWR.n950 VPWR 0.0603958
R15765 VPWR VPWR.n949 0.0603958
R15766 VPWR VPWR.n948 0.0603958
R15767 VPWR.n4822 VPWR 0.0603958
R15768 VPWR.n4819 VPWR 0.0603958
R15769 VPWR.n4811 VPWR 0.0603958
R15770 VPWR VPWR.n4807 0.0603958
R15771 VPWR.n1024 VPWR 0.0603958
R15772 VPWR.n1030 VPWR 0.0603958
R15773 VPWR.n1035 VPWR 0.0603958
R15774 VPWR.n1042 VPWR 0.0603958
R15775 VPWR.n1188 VPWR 0.0603958
R15776 VPWR VPWR.n1187 0.0603958
R15777 VPWR.n1183 VPWR 0.0603958
R15778 VPWR.n1144 VPWR 0.0603958
R15779 VPWR VPWR.n1143 0.0603958
R15780 VPWR.n1137 VPWR 0.0603958
R15781 VPWR.n1133 VPWR 0.0603958
R15782 VPWR VPWR.n1132 0.0603958
R15783 VPWR VPWR.n1130 0.0603958
R15784 VPWR.n4472 VPWR 0.0603958
R15785 VPWR.n4484 VPWR 0.0603958
R15786 VPWR.n4489 VPWR 0.0603958
R15787 VPWR.n4491 VPWR 0.0603958
R15788 VPWR.n4495 VPWR 0.0603958
R15789 VPWR.n4497 VPWR 0.0603958
R15790 VPWR.n4496 VPWR 0.0603958
R15791 VPWR.n4503 VPWR 0.0603958
R15792 VPWR.n4507 VPWR 0.0603958
R15793 VPWR.n4522 VPWR 0.0603958
R15794 VPWR VPWR.n4527 0.0603958
R15795 VPWR.n4528 VPWR 0.0603958
R15796 VPWR.n4624 VPWR 0.0603958
R15797 VPWR VPWR.n373 0.0603958
R15798 VPWR.n4637 VPWR 0.0603958
R15799 VPWR.n4639 VPWR 0.0603958
R15800 VPWR.n4643 VPWR 0.0603958
R15801 VPWR.n4647 VPWR 0.0603958
R15802 VPWR VPWR.n4652 0.0603958
R15803 VPWR.n4653 VPWR 0.0603958
R15804 VPWR.n4656 VPWR 0.0603958
R15805 VPWR.n4665 VPWR 0.0603958
R15806 VPWR.n4666 VPWR 0.0603958
R15807 VPWR.n359 VPWR 0.0603958
R15808 VPWR VPWR.n349 0.0603958
R15809 VPWR.n1231 VPWR 0.0603958
R15810 VPWR.n1235 VPWR 0.0603958
R15811 VPWR VPWR.n1227 0.0603958
R15812 VPWR.n1244 VPWR 0.0603958
R15813 VPWR.n1245 VPWR 0.0603958
R15814 VPWR.n1248 VPWR 0.0603958
R15815 VPWR.n1323 VPWR 0.0603958
R15816 VPWR.n1326 VPWR 0.0603958
R15817 VPWR.n1333 VPWR 0.0603958
R15818 VPWR.n1345 VPWR 0.0603958
R15819 VPWR.n1367 VPWR 0.0603958
R15820 VPWR.n441 VPWR 0.0603958
R15821 VPWR VPWR.n440 0.0603958
R15822 VPWR.n1378 VPWR 0.0603958
R15823 VPWR.n1428 VPWR 0.0603958
R15824 VPWR VPWR.n1427 0.0603958
R15825 VPWR VPWR.n4384 0.0603958
R15826 VPWR.n4380 VPWR 0.0603958
R15827 VPWR.n4377 VPWR 0.0603958
R15828 VPWR.n4364 VPWR 0.0603958
R15829 VPWR VPWR.n4363 0.0603958
R15830 VPWR VPWR.n4361 0.0603958
R15831 VPWR.n4358 VPWR 0.0603958
R15832 VPWR VPWR.n4357 0.0603958
R15833 VPWR.n4352 VPWR 0.0603958
R15834 VPWR.n4350 VPWR 0.0603958
R15835 VPWR VPWR.n4349 0.0603958
R15836 VPWR VPWR.n4348 0.0603958
R15837 VPWR.n4345 VPWR 0.0603958
R15838 VPWR.n3814 VPWR 0.0603958
R15839 VPWR.n3815 VPWR 0.0603958
R15840 VPWR.n3864 VPWR 0.0603958
R15841 VPWR VPWR.n3863 0.0603958
R15842 VPWR.n3857 VPWR 0.0603958
R15843 VPWR VPWR.n3856 0.0603958
R15844 VPWR VPWR.n3855 0.0603958
R15845 VPWR.n3853 VPWR 0.0603958
R15846 VPWR.n3850 VPWR 0.0603958
R15847 VPWR.n3839 VPWR 0.0603958
R15848 VPWR.n3836 VPWR 0.0603958
R15849 VPWR.n3829 VPWR 0.0603958
R15850 VPWR VPWR.n3828 0.0603958
R15851 VPWR VPWR.n3779 0.0603958
R15852 VPWR.n3869 VPWR 0.0603958
R15853 VPWR.n3870 VPWR 0.0603958
R15854 VPWR.n3873 VPWR 0.0603958
R15855 VPWR.n3915 VPWR 0.0603958
R15856 VPWR VPWR.n3908 0.0603958
R15857 VPWR VPWR.n3907 0.0603958
R15858 VPWR.n3903 VPWR 0.0603958
R15859 VPWR.n3900 VPWR 0.0603958
R15860 VPWR VPWR.n3899 0.0603958
R15861 VPWR.n1850 VPWR 0.0603958
R15862 VPWR.n1851 VPWR 0.0603958
R15863 VPWR VPWR.n1855 0.0603958
R15864 VPWR.n1856 VPWR 0.0603958
R15865 VPWR VPWR.n1859 0.0603958
R15866 VPWR.n1860 VPWR 0.0603958
R15867 VPWR.n1861 VPWR 0.0603958
R15868 VPWR.n1867 VPWR 0.0603958
R15869 VPWR.n1872 VPWR 0.0603958
R15870 VPWR VPWR.n1874 0.0603958
R15871 VPWR.n1875 VPWR 0.0603958
R15872 VPWR.n1879 VPWR 0.0603958
R15873 VPWR.n1948 VPWR 0.0603958
R15874 VPWR.n1950 VPWR 0.0603958
R15875 VPWR.n1959 VPWR 0.0603958
R15876 VPWR.n1963 VPWR 0.0603958
R15877 VPWR.n1999 VPWR 0.0603958
R15878 VPWR.n2002 VPWR 0.0603958
R15879 VPWR.n2008 VPWR 0.0603958
R15880 VPWR.n2009 VPWR 0.0603958
R15881 VPWR.n2010 VPWR 0.0603958
R15882 VPWR.n2013 VPWR 0.0603958
R15883 VPWR.n4225 VPWR 0.0603958
R15884 VPWR.n1477 VPWR 0.0603958
R15885 VPWR VPWR.n1477 0.0603958
R15886 VPWR.n4216 VPWR 0.0603958
R15887 VPWR VPWR.n4215 0.0603958
R15888 VPWR VPWR.n4214 0.0603958
R15889 VPWR.n4203 VPWR 0.0603958
R15890 VPWR.n4199 VPWR 0.0603958
R15891 VPWR VPWR.n4198 0.0603958
R15892 VPWR VPWR.n4195 0.0603958
R15893 VPWR VPWR.n4194 0.0603958
R15894 VPWR VPWR.n4193 0.0603958
R15895 VPWR.n4185 VPWR 0.0603958
R15896 VPWR.n4175 VPWR 0.0603958
R15897 VPWR VPWR.n4174 0.0603958
R15898 VPWR VPWR.n4117 0.0603958
R15899 VPWR.n4111 VPWR 0.0603958
R15900 VPWR.n4111 VPWR 0.0603958
R15901 VPWR VPWR.n4110 0.0603958
R15902 VPWR VPWR.n4109 0.0603958
R15903 VPWR VPWR.n4107 0.0603958
R15904 VPWR.n4099 VPWR 0.0603958
R15905 VPWR VPWR.n4098 0.0603958
R15906 VPWR VPWR.n4096 0.0603958
R15907 VPWR.n4087 VPWR 0.0603958
R15908 VPWR VPWR.n4086 0.0603958
R15909 VPWR.n1535 VPWR 0.0603958
R15910 VPWR.n1537 VPWR 0.0603958
R15911 VPWR VPWR.n4070 0.0603958
R15912 VPWR.n4018 VPWR 0.0603958
R15913 VPWR.n4004 VPWR 0.0603958
R15914 VPWR VPWR.n4003 0.0603958
R15915 VPWR.n1677 VPWR 0.0603958
R15916 VPWR.n1683 VPWR 0.0603958
R15917 VPWR.n1689 VPWR 0.0603958
R15918 VPWR.n1698 VPWR 0.0603958
R15919 VPWR.n1702 VPWR 0.0603958
R15920 VPWR VPWR.n1797 0.0603958
R15921 VPWR.n1792 VPWR 0.0603958
R15922 VPWR VPWR.n1791 0.0603958
R15923 VPWR VPWR.n1790 0.0603958
R15924 VPWR.n1785 VPWR 0.0603958
R15925 VPWR VPWR.n1756 0.0603958
R15926 VPWR.n1751 VPWR 0.0603958
R15927 VPWR.n1747 VPWR 0.0603958
R15928 VPWR VPWR.n1745 0.0603958
R15929 VPWR.n1745 VPWR 0.0603958
R15930 VPWR VPWR.n1743 0.0603958
R15931 VPWR.n2119 VPWR 0.0603958
R15932 VPWR VPWR.n2118 0.0603958
R15933 VPWR VPWR.n1604 0.0603958
R15934 VPWR VPWR.n1595 0.0603958
R15935 VPWR VPWR.n1584 0.0603958
R15936 VPWR.n2125 VPWR 0.0603958
R15937 VPWR.n2128 VPWR 0.0603958
R15938 VPWR VPWR.n2140 0.0603958
R15939 VPWR.n2141 VPWR 0.0603958
R15940 VPWR.n2147 VPWR 0.0603958
R15941 VPWR.n2151 VPWR 0.0603958
R15942 VPWR VPWR.n3587 0.0603958
R15943 VPWR.n3589 VPWR 0.0603958
R15944 VPWR.n3594 VPWR 0.0603958
R15945 VPWR.n3600 VPWR 0.0603958
R15946 VPWR.n3601 VPWR 0.0603958
R15947 VPWR.n3607 VPWR 0.0603958
R15948 VPWR.n3618 VPWR 0.0603958
R15949 VPWR VPWR.n1576 0.0603958
R15950 VPWR.n3627 VPWR 0.0603958
R15951 VPWR.n3635 VPWR 0.0603958
R15952 VPWR.n3638 VPWR 0.0603958
R15953 VPWR.n3679 VPWR 0.0603958
R15954 VPWR VPWR.n3678 0.0603958
R15955 VPWR.n3662 VPWR 0.0603958
R15956 VPWR.n3660 VPWR 0.0603958
R15957 VPWR.n3657 VPWR 0.0603958
R15958 VPWR.n2698 VPWR 0.0603958
R15959 VPWR.n2703 VPWR 0.0603958
R15960 VPWR.n2711 VPWR 0.0603958
R15961 VPWR.n2712 VPWR 0.0603958
R15962 VPWR.n2716 VPWR 0.0603958
R15963 VPWR VPWR.n2716 0.0603958
R15964 VPWR.n2717 VPWR 0.0603958
R15965 VPWR.n2720 VPWR 0.0603958
R15966 VPWR.n2986 VPWR 0.0603958
R15967 VPWR.n2984 VPWR 0.0603958
R15968 VPWR.n2981 VPWR 0.0603958
R15969 VPWR VPWR.n2980 0.0603958
R15970 VPWR VPWR.n2978 0.0603958
R15971 VPWR VPWR.n2977 0.0603958
R15972 VPWR VPWR.n2975 0.0603958
R15973 VPWR.n2968 VPWR 0.0603958
R15974 VPWR.n2942 VPWR 0.0603958
R15975 VPWR.n2933 VPWR 0.0603958
R15976 VPWR.n2803 VPWR 0.0603958
R15977 VPWR.n2815 VPWR 0.0603958
R15978 VPWR.n2817 VPWR 0.0603958
R15979 VPWR.n2860 VPWR 0.0603958
R15980 VPWR.n2870 VPWR 0.0603958
R15981 VPWR.n2881 VPWR 0.0603958
R15982 VPWR VPWR.n2926 0.0603958
R15983 VPWR.n2923 VPWR 0.0603958
R15984 VPWR.n2917 VPWR 0.0603958
R15985 VPWR.n2903 VPWR 0.0603958
R15986 VPWR.n2900 VPWR 0.0603958
R15987 VPWR.n2218 VPWR 0.0603958
R15988 VPWR.n2222 VPWR 0.0603958
R15989 VPWR.n2237 VPWR 0.0603958
R15990 VPWR.n2246 VPWR 0.0603958
R15991 VPWR VPWR.n3435 0.0603958
R15992 VPWR VPWR.n3434 0.0603958
R15993 VPWR.n2315 VPWR 0.0603958
R15994 VPWR.n6385 VPWR 0.0603958
R15995 VPWR.n6389 VPWR 0.0603958
R15996 VPWR.n6394 VPWR 0.0603958
R15997 VPWR.n6397 VPWR 0.0603958
R15998 VPWR.n6475 VPWR 0.0603958
R15999 VPWR.n6484 VPWR 0.0603958
R16000 VPWR.n6525 VPWR 0.0603958
R16001 VPWR.n5007 VPWR 0.0603958
R16002 VPWR.n5016 VPWR 0.0603958
R16003 VPWR.n5054 VPWR 0.0603958
R16004 VPWR VPWR.n5053 0.0603958
R16005 VPWR VPWR.n5052 0.0603958
R16006 VPWR.n5036 VPWR 0.0603958
R16007 VPWR.n5030 VPWR 0.0603958
R16008 VPWR VPWR.n5029 0.0603958
R16009 VPWR.n5024 VPWR 0.0603958
R16010 VPWR VPWR.n5023 0.0603958
R16011 VPWR.n7720 VPWR 0.0603958
R16012 VPWR VPWR.n7719 0.0603958
R16013 VPWR VPWR.n7718 0.0603958
R16014 VPWR.n7714 VPWR 0.0603958
R16015 VPWR.n7708 VPWR 0.0603958
R16016 VPWR.n7702 VPWR 0.0603958
R16017 VPWR.n7696 VPWR 0.0603958
R16018 VPWR VPWR.n7695 0.0603958
R16019 VPWR.n7689 VPWR 0.0603958
R16020 VPWR.n7684 VPWR 0.0603958
R16021 VPWR VPWR.n7683 0.0603958
R16022 VPWR VPWR.n7682 0.0603958
R16023 VPWR.n7673 VPWR 0.0603958
R16024 VPWR VPWR.n7672 0.0603958
R16025 VPWR.n7664 VPWR 0.0603958
R16026 VPWR.n74 VPWR 0.0603958
R16027 VPWR.n66 VPWR 0.0603958
R16028 VPWR VPWR.n65 0.0603958
R16029 VPWR.n62 VPWR 0.0603958
R16030 VPWR VPWR.n60 0.0603958
R16031 VPWR VPWR.n58 0.0603958
R16032 VPWR VPWR.n2580 0.0603958
R16033 VPWR VPWR.n2578 0.0603958
R16034 VPWR.n2593 VPWR 0.0603958
R16035 VPWR.n2594 VPWR 0.0603958
R16036 VPWR.n2597 VPWR 0.0603958
R16037 VPWR.n2606 VPWR 0.0603958
R16038 VPWR.n2611 VPWR 0.0603958
R16039 VPWR.n2559 VPWR 0.0603958
R16040 VPWR VPWR.n2557 0.0603958
R16041 VPWR.n2553 VPWR 0.0603958
R16042 VPWR VPWR.n2551 0.0603958
R16043 VPWR VPWR.n2532 0.0603958
R16044 VPWR.n2528 VPWR 0.0603958
R16045 VPWR.n2523 VPWR 0.0603958
R16046 VPWR VPWR.n2522 0.0603958
R16047 VPWR.n3115 VPWR 0.0603958
R16048 VPWR VPWR.n3114 0.0603958
R16049 VPWR VPWR.n3112 0.0603958
R16050 VPWR.n3112 VPWR 0.0603958
R16051 VPWR.n2450 VPWR 0.0603958
R16052 VPWR VPWR.n2449 0.0603958
R16053 VPWR VPWR.n2438 0.0603958
R16054 VPWR VPWR.n2437 0.0603958
R16055 VPWR.n2429 VPWR 0.0603958
R16056 VPWR VPWR.n2429 0.0603958
R16057 VPWR.n3120 VPWR 0.0603958
R16058 VPWR.n3122 VPWR 0.0603958
R16059 VPWR.n3125 VPWR 0.0603958
R16060 VPWR.n3282 VPWR 0.0603958
R16061 VPWR VPWR.n3280 0.0603958
R16062 VPWR VPWR.n3262 0.0603958
R16063 VPWR VPWR.n3236 0.0603958
R16064 VPWR.n3236 VPWR 0.0603958
R16065 VPWR.n3233 VPWR 0.0603958
R16066 VPWR.n3287 VPWR 0.0603958
R16067 VPWR.n3288 VPWR 0.0603958
R16068 VPWR.n3291 VPWR 0.0603958
R16069 VPWR.n3316 VPWR 0.0603958
R16070 VPWR VPWR.n3315 0.0603958
R16071 VPWR VPWR.n3310 0.0603958
R16072 VPWR VPWR.n6288 0.0603958
R16073 VPWR.n6289 VPWR 0.0603958
R16074 VPWR VPWR.n6281 0.0603958
R16075 VPWR.n6301 VPWR 0.0603958
R16076 VPWR.n6309 VPWR 0.0603958
R16077 VPWR.n6314 VPWR 0.0603958
R16078 VPWR VPWR.n6262 0.0603958
R16079 VPWR.n6255 VPWR 0.0603958
R16080 VPWR VPWR.n6254 0.0603958
R16081 VPWR VPWR.n6248 0.0603958
R16082 VPWR.n6224 VPWR 0.0603958
R16083 VPWR VPWR.n6223 0.0603958
R16084 VPWR.n6218 VPWR 0.0603958
R16085 VPWR VPWR.n6217 0.0603958
R16086 VPWR.n6213 VPWR 0.0603958
R16087 VPWR VPWR.n5823 0.0603958
R16088 VPWR.n6153 VPWR 0.0603958
R16089 VPWR VPWR.n6152 0.0603958
R16090 VPWR VPWR.n6138 0.0603958
R16091 VPWR VPWR.n6137 0.0603958
R16092 VPWR VPWR.n6130 0.0603958
R16093 VPWR.n6120 VPWR 0.0603958
R16094 VPWR VPWR.n6119 0.0603958
R16095 VPWR VPWR.n6113 0.0603958
R16096 VPWR.n5848 VPWR 0.0603958
R16097 VPWR.n5849 VPWR 0.0603958
R16098 VPWR.n5855 VPWR 0.0603958
R16099 VPWR.n5861 VPWR 0.0603958
R16100 VPWR.n5890 VPWR 0.0603958
R16101 VPWR VPWR.n5900 0.0603958
R16102 VPWR.n5901 VPWR 0.0603958
R16103 VPWR.n5904 VPWR 0.0603958
R16104 VPWR.n6040 VPWR 0.0603958
R16105 VPWR.n5953 VPWR 0.0603958
R16106 VPWR VPWR.n5952 0.0603958
R16107 VPWR VPWR.n5925 0.0603958
R16108 VPWR.n5942 VPWR 0.0603958
R16109 VPWR VPWR.n5941 0.0603958
R16110 VPWR.n5934 VPWR 0.0603958
R16111 VPWR VPWR.n5933 0.0603958
R16112 VPWR.n4046 VPWR.n4045 0.059272
R16113 VPWR.n4687 VPWR.n4676 0.0590938
R16114 VPWR.n1717 VPWR.n1715 0.0586222
R16115 VPWR.n5324 VPWR.n5323 0.0577917
R16116 VPWR.n971 VPWR.n969 0.0577917
R16117 VPWR.n1204 VPWR.n1203 0.0577917
R16118 VPWR.n2991 VPWR.n2989 0.0577917
R16119 VPWR.n5123 VPWR.n5116 0.0561015
R16120 VPWR.n5620 VPWR.n5462 0.0561015
R16121 VPWR.n5387 VPWR.n5380 0.0561015
R16122 VPWR.n1276 VPWR.n1256 0.0561015
R16123 VPWR.n1896 VPWR.n1882 0.0561015
R16124 VPWR.n1715 VPWR.n1708 0.0561015
R16125 VPWR.n2745 VPWR.n2723 0.0561015
R16126 VPWR.n2614 VPWR.n2613 0.0561015
R16127 VPWR.n6317 VPWR.n6316 0.0561015
R16128 VPWR.n6445 VPWR.n6408 0.0561015
R16129 VPWR.n3001 VPWR.n2999 0.0548679
R16130 VPWR.n81 VPWR.n80 0.0547995
R16131 VPWR.n4723 VPWR.n366 0.0547995
R16132 VPWR.n3924 VPWR.n3923 0.0547995
R16133 VPWR.n4046 VPWR.n4028 0.0547995
R16134 VPWR.n3683 VPWR.n3682 0.0547995
R16135 VPWR.n2360 VPWR.n2329 0.0547995
R16136 VPWR.n3330 VPWR.n3329 0.0547995
R16137 VPWR.n5401 VPWR.n5400 0.0512937
R16138 VPWR.n556 VPWR.n555 0.0512937
R16139 VPWR.n1262 VPWR.n1261 0.0512937
R16140 VPWR.n2759 VPWR.n2758 0.0512937
R16141 VPWR.n6085 VPWR 0.0497858
R16142 VPWR.n5124 VPWR.n5123 0.0496664
R16143 VPWR.n5620 VPWR.n5619 0.0496664
R16144 VPWR.n5388 VPWR.n5387 0.0496664
R16145 VPWR.n1056 VPWR.n1054 0.0496664
R16146 VPWR.n4723 VPWR.n4722 0.0496664
R16147 VPWR.n1276 VPWR.n1275 0.0496664
R16148 VPWR.n3925 VPWR.n3924 0.0496664
R16149 VPWR.n1896 VPWR.n1895 0.0496664
R16150 VPWR.n3684 VPWR.n3683 0.0496664
R16151 VPWR.n2746 VPWR.n2745 0.0496664
R16152 VPWR.n2360 VPWR.n2359 0.0496664
R16153 VPWR.n6445 VPWR.n6444 0.0496664
R16154 VPWR.n82 VPWR.n81 0.0496664
R16155 VPWR.n2616 VPWR.n2614 0.0496664
R16156 VPWR.n3332 VPWR.n3330 0.0496664
R16157 VPWR.n6319 VPWR.n6317 0.0496664
R16158 VPWR VPWR.n5496 0.047375
R16159 VPWR.n2017 VPWR 0.047375
R16160 VPWR.n3109 VPWR 0.047375
R16161 VPWR.n6696 VPWR.n6695 0.0460729
R16162 VPWR.n5490 VPWR.n5489 0.0460729
R16163 VPWR.n6795 VPWR.n6794 0.0460729
R16164 VPWR.n692 VPWR.n691 0.0460729
R16165 VPWR.n589 VPWR.n588 0.0460729
R16166 VPWR.n1119 VPWR.n1118 0.0460729
R16167 VPWR.n4602 VPWR.n4601 0.0460729
R16168 VPWR.n3799 VPWR.n3798 0.0460729
R16169 VPWR.n3574 VPWR.n3573 0.0460729
R16170 VPWR.n2830 VPWR.n2829 0.0460729
R16171 VPWR.n3461 VPWR.n3460 0.0460729
R16172 VPWR.n6539 VPWR.n6538 0.0460729
R16173 VPWR.n3101 VPWR.n3100 0.0460729
R16174 VPWR.n6203 VPWR.n6202 0.0460729
R16175 VPWR.n4860 VPWR.n4859 0.0460313
R16176 VPWR.n517 VPWR.n510 0.0446272
R16177 VPWR.n5959 VPWR.n5958 0.0433251
R16178 VPWR.n204 VPWR.n203 0.0433251
R16179 VPWR.n7473 VPWR.n7472 0.0433251
R16180 VPWR.n7363 VPWR.n7362 0.0433251
R16181 VPWR.n4832 VPWR.n4831 0.0433251
R16182 VPWR.n5131 VPWR.n5130 0.0421667
R16183 VPWR.n225 VPWR.n224 0.0421667
R16184 VPWR.n5610 VPWR.n5609 0.0421667
R16185 VPWR.n7486 VPWR.n7485 0.0421667
R16186 VPWR.n529 VPWR.n528 0.0421667
R16187 VPWR.n4845 VPWR.n4844 0.0421667
R16188 VPWR.n1065 VPWR.n1064 0.0421667
R16189 VPWR.n4713 VPWR.n4712 0.0421667
R16190 VPWR.n1267 VPWR.n1266 0.0421667
R16191 VPWR.n3932 VPWR.n3931 0.0421667
R16192 VPWR.n4040 VPWR.n4039 0.0421667
R16193 VPWR.n1723 VPWR.n1722 0.0421667
R16194 VPWR.n3693 VPWR.n3692 0.0421667
R16195 VPWR.n2755 VPWR.n2754 0.0421667
R16196 VPWR.n6438 VPWR.n6437 0.0421667
R16197 VPWR.n91 VPWR.n90 0.0421667
R16198 VPWR.n2625 VPWR.n2624 0.0421667
R16199 VPWR.n3341 VPWR.n3340 0.0421667
R16200 VPWR.n6328 VPWR.n6327 0.0421667
R16201 VPWR.n5980 VPWR.n5979 0.0421667
R16202 VPWR.n520 VPWR.n518 0.0408646
R16203 VPWR.n2495 VPWR.n2494 0.0393514
R16204 VPWR.n111 VPWR.n109 0.0393514
R16205 VPWR.n237 VPWR.n167 0.0393514
R16206 VPWR.n5121 VPWR.n5117 0.0393514
R16207 VPWR.n7435 VPWR.n7429 0.0393514
R16208 VPWR.n5623 VPWR.n5622 0.0393514
R16209 VPWR.n7325 VPWR.n7319 0.0393514
R16210 VPWR.n5385 VPWR.n5381 0.0393514
R16211 VPWR.n4795 VPWR.n4789 0.0393514
R16212 VPWR.n515 VPWR.n511 0.0393514
R16213 VPWR.n4725 VPWR.n335 0.0393514
R16214 VPWR.n1052 VPWR.n1048 0.0393514
R16215 VPWR.n3770 VPWR.n3768 0.0393514
R16216 VPWR.n1279 VPWR.n1278 0.0393514
R16217 VPWR.n4048 VPWR.n3992 0.0393514
R16218 VPWR.n1899 VPWR.n1898 0.0393514
R16219 VPWR.n1713 VPWR.n1709 0.0393514
R16220 VPWR.n1547 VPWR.n1545 0.0393514
R16221 VPWR.n2362 VPWR.n2289 0.0393514
R16222 VPWR.n6448 VPWR.n6447 0.0393514
R16223 VPWR.n5712 VPWR.n5711 0.0393514
R16224 VPWR.n2375 VPWR.n2373 0.0393514
R16225 VPWR.n5992 VPWR.n5920 0.0393514
R16226 VPWR.n6433 VPWR.n6432 0.0382581
R16227 VPWR.n5135 VPWR.n5134 0.0382581
R16228 VPWR.n3676 VPWR.n3675 0.0382581
R16229 VPWR.n235 VPWR 0.0369583
R16230 VPWR VPWR.n7475 0.0369583
R16231 VPWR VPWR.n4764 0.0369583
R16232 VPWR.n4059 VPWR 0.0369583
R16233 VPWR.n5990 VPWR 0.0369583
R16234 VPWR.n6656 VPWR.n6655 0.035973
R16235 VPWR.n5471 VPWR.n5470 0.0356562
R16236 VPWR.n6916 VPWR.n6915 0.0356562
R16237 VPWR.n7031 VPWR.n7030 0.0356562
R16238 VPWR.n7189 VPWR.n7188 0.0356562
R16239 VPWR.n865 VPWR.n864 0.0356562
R16240 VPWR.n1384 VPWR.n1383 0.0356562
R16241 VPWR.n4236 VPWR.n4235 0.0356562
R16242 VPWR.n2080 VPWR.n2079 0.0356562
R16243 VPWR.n3551 VPWR.n3550 0.0356562
R16244 VPWR.n2848 VPWR.n2847 0.0356562
R16245 VPWR.n3484 VPWR.n3483 0.0356562
R16246 VPWR.n6563 VPWR.n6562 0.0356562
R16247 VPWR.n3078 VPWR.n3077 0.0356562
R16248 VPWR.n3172 VPWR.n3171 0.0356562
R16249 VPWR.n6180 VPWR.n6179 0.0356562
R16250 VPWR.n6106 VPWR.n6105 0.0356562
R16251 VPWR VPWR.n6660 0.0343542
R16252 VPWR.n216 VPWR.n214 0.0343542
R16253 VPWR.n7421 VPWR.n7419 0.0343542
R16254 VPWR.n5342 VPWR.n5340 0.0343542
R16255 VPWR.n7306 VPWR.n7304 0.0343542
R16256 VPWR VPWR.n717 0.0343542
R16257 VPWR.n4782 VPWR.n4781 0.0343542
R16258 VPWR.n1075 VPWR.n1074 0.0343542
R16259 VPWR VPWR.n403 0.0343542
R16260 VPWR.n4704 VPWR.n4702 0.0343542
R16261 VPWR.n3942 VPWR.n3941 0.0343542
R16262 VPWR.n4033 VPWR.n4032 0.0343542
R16263 VPWR.n3700 VPWR.n3699 0.0343542
R16264 VPWR.n2332 VPWR.n2330 0.0343542
R16265 VPWR.n98 VPWR.n97 0.0343542
R16266 VPWR.n2635 VPWR.n2634 0.0343542
R16267 VPWR.n3351 VPWR.n3350 0.0343542
R16268 VPWR.n6338 VPWR.n6337 0.0343542
R16269 VPWR.n5971 VPWR.n5969 0.0343542
R16270 VPWR.n7736 VPWR.n7735 0.0342838
R16271 VPWR.n7614 VPWR.n7613 0.0342838
R16272 VPWR.n6597 VPWR.n6596 0.0342838
R16273 VPWR.n6785 VPWR.n6784 0.0342838
R16274 VPWR.n7004 VPWR.n7003 0.0342838
R16275 VPWR.n7157 VPWR.n294 0.0342838
R16276 VPWR.n5292 VPWR.n5291 0.0342838
R16277 VPWR.n593 VPWR.n592 0.0342838
R16278 VPWR.n621 VPWR.n620 0.0342838
R16279 VPWR.n4563 VPWR.n4562 0.0342838
R16280 VPWR.n4430 VPWR.n4429 0.0342838
R16281 VPWR.n4291 VPWR.n4290 0.0342838
R16282 VPWR.n1411 VPWR.n1410 0.0342838
R16283 VPWR.n1517 VPWR.n1506 0.0342838
R16284 VPWR.n2032 VPWR.n2031 0.0342838
R16285 VPWR.n3532 VPWR.n3531 0.0342838
R16286 VPWR.n1590 VPWR.n1589 0.0342838
R16287 VPWR.n4954 VPWR.n4953 0.0342838
R16288 VPWR.n3497 VPWR.n3496 0.0342838
R16289 VPWR.n2480 VPWR.n2479 0.0342838
R16290 VPWR.n2468 VPWR.n2467 0.0342838
R16291 VPWR.n5789 VPWR.n5788 0.0342838
R16292 VPWR.n2389 VPWR.n2388 0.0342838
R16293 VPWR.n6060 VPWR.n2 0.0342838
R16294 VPWR.n5675 VPWR 0.0330521
R16295 VPWR.n6737 VPWR 0.0330521
R16296 VPWR.n6763 VPWR 0.0330521
R16297 VPWR.n176 VPWR 0.0330521
R16298 VPWR VPWR.n5599 0.0330521
R16299 VPWR.n7452 VPWR 0.0330521
R16300 VPWR VPWR.n5284 0.0330521
R16301 VPWR.n7236 VPWR 0.0330521
R16302 VPWR.n7279 VPWR 0.0330521
R16303 VPWR.n7343 VPWR 0.0330521
R16304 VPWR.n562 VPWR 0.0330521
R16305 VPWR.n680 VPWR 0.0330521
R16306 VPWR.n1186 VPWR 0.0330521
R16307 VPWR.n1131 VPWR 0.0330521
R16308 VPWR VPWR.n4490 0.0330521
R16309 VPWR.n4545 VPWR 0.0330521
R16310 VPWR.n4640 VPWR 0.0330521
R16311 VPWR.n1232 VPWR 0.0330521
R16312 VPWR VPWR.n1250 0.0330521
R16313 VPWR.n1296 VPWR 0.0330521
R16314 VPWR VPWR.n1379 0.0330521
R16315 VPWR.n4362 VPWR 0.0330521
R16316 VPWR.n4321 VPWR 0.0330521
R16317 VPWR.n1932 VPWR 0.0330521
R16318 VPWR VPWR.n1949 0.0330521
R16319 VPWR.n4202 VPWR 0.0330521
R16320 VPWR.n4169 VPWR 0.0330521
R16321 VPWR.n4118 VPWR 0.0330521
R16322 VPWR.n4071 VPWR 0.0330521
R16323 VPWR.n1699 VPWR 0.0330521
R16324 VPWR.n1819 VPWR 0.0330521
R16325 VPWR.n1788 VPWR 0.0330521
R16326 VPWR.n1750 VPWR 0.0330521
R16327 VPWR.n1743 VPWR 0.0330521
R16328 VPWR VPWR.n3640 0.0330521
R16329 VPWR.n2781 VPWR 0.0330521
R16330 VPWR.n2979 VPWR 0.0330521
R16331 VPWR.n2899 VPWR 0.0330521
R16332 VPWR.n2219 VPWR 0.0330521
R16333 VPWR VPWR.n6398 0.0330521
R16334 VPWR VPWR.n6427 0.0330521
R16335 VPWR.n7780 VPWR 0.0330521
R16336 VPWR.n7683 VPWR 0.0330521
R16337 VPWR.n7671 VPWR 0.0330521
R16338 VPWR.n56 VPWR 0.0330521
R16339 VPWR.n2552 VPWR 0.0330521
R16340 VPWR.n3113 VPWR 0.0330521
R16341 VPWR VPWR.n6300 0.0330521
R16342 VPWR.n6221 VPWR 0.0330521
R16343 VPWR.n6216 VPWR 0.0330521
R16344 VPWR.n7627 VPWR.n7626 0.0325946
R16345 VPWR.n6886 VPWR.n6885 0.0325946
R16346 VPWR.n7179 VPWR.n7178 0.0325946
R16347 VPWR.n855 VPWR.n853 0.0325946
R16348 VPWR.n4591 VPWR.n4589 0.0325946
R16349 VPWR.n3788 VPWR.n3786 0.0325946
R16350 VPWR.n4154 VPWR.n4152 0.0325946
R16351 VPWR.n2170 VPWR.n2169 0.0325946
R16352 VPWR.n3054 VPWR.n3053 0.0325946
R16353 VPWR.n6072 VPWR.n6071 0.0325946
R16354 VPWR.n5188 VPWR 0.03175
R16355 VPWR.n6705 VPWR 0.03175
R16356 VPWR.n4938 VPWR 0.03175
R16357 VPWR VPWR.n158 0.03175
R16358 VPWR.n7524 VPWR 0.03175
R16359 VPWR.n191 VPWR 0.03175
R16360 VPWR VPWR.n5431 0.03175
R16361 VPWR VPWR.n5442 0.03175
R16362 VPWR.n5457 VPWR 0.03175
R16363 VPWR.n5559 VPWR 0.03175
R16364 VPWR.n5558 VPWR 0.03175
R16365 VPWR.n5499 VPWR 0.03175
R16366 VPWR.n6971 VPWR 0.03175
R16367 VPWR.n6954 VPWR 0.03175
R16368 VPWR.n6951 VPWR 0.03175
R16369 VPWR.n6923 VPWR 0.03175
R16370 VPWR VPWR.n6797 0.03175
R16371 VPWR.n6851 VPWR 0.03175
R16372 VPWR.n7406 VPWR 0.03175
R16373 VPWR.n5364 VPWR 0.03175
R16374 VPWR.n5375 VPWR 0.03175
R16375 VPWR VPWR.n5234 0.03175
R16376 VPWR VPWR.n5239 0.03175
R16377 VPWR.n5253 VPWR 0.03175
R16378 VPWR VPWR.n5274 0.03175
R16379 VPWR VPWR.n5285 0.03175
R16380 VPWR.n5308 VPWR 0.03175
R16381 VPWR VPWR.n7096 0.03175
R16382 VPWR.n7097 VPWR 0.03175
R16383 VPWR.n7123 VPWR 0.03175
R16384 VPWR VPWR.n7226 0.03175
R16385 VPWR.n7247 VPWR 0.03175
R16386 VPWR VPWR.n7277 0.03175
R16387 VPWR.n504 VPWR 0.03175
R16388 VPWR VPWR.n574 0.03175
R16389 VPWR VPWR.n647 0.03175
R16390 VPWR VPWR.n663 0.03175
R16391 VPWR VPWR.n678 0.03175
R16392 VPWR.n603 VPWR 0.03175
R16393 VPWR VPWR.n783 0.03175
R16394 VPWR VPWR.n893 0.03175
R16395 VPWR.n950 VPWR 0.03175
R16396 VPWR.n949 VPWR 0.03175
R16397 VPWR.n1188 VPWR 0.03175
R16398 VPWR.n1144 VPWR 0.03175
R16399 VPWR.n1133 VPWR 0.03175
R16400 VPWR.n4484 VPWR 0.03175
R16401 VPWR VPWR.n4495 0.03175
R16402 VPWR.n4621 VPWR 0.03175
R16403 VPWR VPWR.n4624 0.03175
R16404 VPWR.n4653 VPWR 0.03175
R16405 VPWR VPWR.n4665 0.03175
R16406 VPWR.n1323 VPWR 0.03175
R16407 VPWR.n4358 VPWR 0.03175
R16408 VPWR.n4349 VPWR 0.03175
R16409 VPWR VPWR.n3815 0.03175
R16410 VPWR.n3864 VPWR 0.03175
R16411 VPWR.n3857 VPWR 0.03175
R16412 VPWR.n3828 VPWR 0.03175
R16413 VPWR.n3779 VPWR 0.03175
R16414 VPWR VPWR.n3869 0.03175
R16415 VPWR.n3908 VPWR 0.03175
R16416 VPWR.n3900 VPWR 0.03175
R16417 VPWR VPWR.n1860 0.03175
R16418 VPWR VPWR.n1959 0.03175
R16419 VPWR VPWR.n2009 0.03175
R16420 VPWR.n2010 VPWR 0.03175
R16421 VPWR.n4216 VPWR 0.03175
R16422 VPWR.n4198 VPWR 0.03175
R16423 VPWR.n4194 VPWR 0.03175
R16424 VPWR.n4175 VPWR 0.03175
R16425 VPWR.n4110 VPWR 0.03175
R16426 VPWR.n4086 VPWR 0.03175
R16427 VPWR VPWR.n1535 0.03175
R16428 VPWR.n4004 VPWR 0.03175
R16429 VPWR.n1791 VPWR 0.03175
R16430 VPWR.n2119 VPWR 0.03175
R16431 VPWR.n1584 VPWR 0.03175
R16432 VPWR.n2141 VPWR 0.03175
R16433 VPWR VPWR.n3589 0.03175
R16434 VPWR.n3601 VPWR 0.03175
R16435 VPWR.n3635 VPWR 0.03175
R16436 VPWR.n2717 VPWR 0.03175
R16437 VPWR.n2978 VPWR 0.03175
R16438 VPWR.n2977 VPWR 0.03175
R16439 VPWR VPWR.n2803 0.03175
R16440 VPWR VPWR.n2815 0.03175
R16441 VPWR.n2927 VPWR 0.03175
R16442 VPWR.n2926 VPWR 0.03175
R16443 VPWR VPWR.n2211 0.03175
R16444 VPWR.n3436 VPWR 0.03175
R16445 VPWR.n3435 VPWR 0.03175
R16446 VPWR VPWR.n6474 0.03175
R16447 VPWR.n6475 VPWR 0.03175
R16448 VPWR.n6522 VPWR 0.03175
R16449 VPWR VPWR.n5016 0.03175
R16450 VPWR.n5054 VPWR 0.03175
R16451 VPWR.n5053 VPWR 0.03175
R16452 VPWR.n5030 VPWR 0.03175
R16453 VPWR.n7720 VPWR 0.03175
R16454 VPWR.n7719 VPWR 0.03175
R16455 VPWR.n7696 VPWR 0.03175
R16456 VPWR.n7673 VPWR 0.03175
R16457 VPWR.n66 VPWR 0.03175
R16458 VPWR.n2594 VPWR 0.03175
R16459 VPWR.n2559 VPWR 0.03175
R16460 VPWR.n3115 VPWR 0.03175
R16461 VPWR.n2450 VPWR 0.03175
R16462 VPWR.n2437 VPWR 0.03175
R16463 VPWR VPWR.n3120 0.03175
R16464 VPWR.n3282 VPWR 0.03175
R16465 VPWR VPWR.n3287 0.03175
R16466 VPWR.n3315 VPWR 0.03175
R16467 VPWR.n6263 VPWR 0.03175
R16468 VPWR.n6255 VPWR 0.03175
R16469 VPWR.n6218 VPWR 0.03175
R16470 VPWR.n6153 VPWR 0.03175
R16471 VPWR.n6138 VPWR 0.03175
R16472 VPWR.n6120 VPWR 0.03175
R16473 VPWR VPWR.n5848 0.03175
R16474 VPWR.n5849 VPWR 0.03175
R16475 VPWR VPWR.n5904 0.03175
R16476 VPWR.n5942 VPWR 0.03175
R16477 VPWR.n7788 VPWR.n7787 0.0309054
R16478 VPWR.n6583 VPWR.n6582 0.0309054
R16479 VPWR.n7429 VPWR.n7428 0.0309054
R16480 VPWR.n4914 VPWR.n4913 0.0309054
R16481 VPWR.n7319 VPWR.n7318 0.0309054
R16482 VPWR.n4875 VPWR.n4874 0.0309054
R16483 VPWR.n4789 VPWR.n4788 0.0309054
R16484 VPWR.n608 VPWR.n607 0.0309054
R16485 VPWR.n335 VPWR.n334 0.0309054
R16486 VPWR.n4439 VPWR.n4438 0.0309054
R16487 VPWR.n3768 VPWR.n3767 0.0309054
R16488 VPWR.n425 VPWR.n424 0.0309054
R16489 VPWR.n3992 VPWR.n3991 0.0309054
R16490 VPWR.n1465 VPWR.n1464 0.0309054
R16491 VPWR.n1632 VPWR.n1631 0.0309054
R16492 VPWR.n4974 VPWR.n4973 0.0309054
R16493 VPWR.n2728 VPWR.n2727 0.0309054
R16494 VPWR.n5752 VPWR.n5751 0.0309054
R16495 VPWR.n3154 VPWR.n3153 0.0309054
R16496 VPWR.n6081 VPWR.n6080 0.0309054
R16497 VPWR.n5920 VPWR.n5919 0.0309054
R16498 VPWR VPWR.n7068 0.0296459
R16499 VPWR.n740 VPWR 0.0296459
R16500 VPWR VPWR.n1405 0.0291458
R16501 VPWR VPWR.n2026 0.0291458
R16502 VPWR VPWR.n2102 0.0291458
R16503 VPWR.n5664 VPWR.n5662 0.0284688
R16504 VPWR.n5588 VPWR.n5586 0.0284688
R16505 VPWR.n1308 VPWR.n1307 0.0284688
R16506 VPWR.n1944 VPWR.n1943 0.0284688
R16507 VPWR.n1813 VPWR.n1812 0.0284688
R16508 VPWR.n6458 VPWR.n5066 0.0284688
R16509 VPWR.n6351 VPWR.n6350 0.0284688
R16510 VPWR.n7519 VPWR.n162 0.0282455
R16511 VPWR.n7298 VPWR.n7297 0.0282455
R16512 VPWR.n3950 VPWR.n3949 0.0282455
R16513 VPWR.n3707 VPWR.n3706 0.0282455
R16514 VPWR.n3425 VPWR.n3424 0.0282455
R16515 VPWR.n7662 VPWR.n104 0.0282455
R16516 VPWR.n2648 VPWR.n2647 0.0282455
R16517 VPWR.n6026 VPWR.n5906 0.0282455
R16518 VPWR.n3363 VPWR.n3362 0.0282455
R16519 VPWR.n6606 VPWR.n6605 0.0278438
R16520 VPWR.n6654 VPWR 0.0278438
R16521 VPWR.n7616 VPWR 0.0278438
R16522 VPWR VPWR.n7405 0.0278438
R16523 VPWR.n7159 VPWR 0.0278438
R16524 VPWR VPWR.n7365 0.0278438
R16525 VPWR.n3190 VPWR 0.0278438
R16526 VPWR VPWR.n0 0.0278438
R16527 VPWR.n2672 VPWR.n2671 0.027527
R16528 VPWR.n7643 VPWR.n7642 0.027527
R16529 VPWR.n5083 VPWR.n5082 0.027527
R16530 VPWR.n7489 VPWR.n275 0.027527
R16531 VPWR.n5637 VPWR.n5636 0.027527
R16532 VPWR.n7389 VPWR.n7388 0.027527
R16533 VPWR.n5405 VPWR.n5404 0.027527
R16534 VPWR.n4848 VPWR.n317 0.027527
R16535 VPWR.n553 VPWR.n551 0.027527
R16536 VPWR.n4748 VPWR.n4747 0.027527
R16537 VPWR.n990 VPWR.n989 0.027527
R16538 VPWR.n3756 VPWR.n3755 0.027527
R16539 VPWR.n456 VPWR.n455 0.027527
R16540 VPWR.n3980 VPWR.n3979 0.027527
R16541 VPWR.n1923 VPWR.n1921 0.027527
R16542 VPWR.n1665 VPWR.n1664 0.027527
R16543 VPWR.n6367 VPWR.n6366 0.027527
R16544 VPWR.n5704 VPWR.n5703 0.027527
R16545 VPWR.n3387 VPWR.n3386 0.027527
R16546 VPWR.n5999 VPWR.n5998 0.027527
R16547 VPWR.n6684 VPWR.n6683 0.0265417
R16548 VPWR.n7623 VPWR.n7622 0.0265417
R16549 VPWR.n5484 VPWR.n5483 0.0265417
R16550 VPWR.n7025 VPWR.n7024 0.0265417
R16551 VPWR.n704 VPWR.n703 0.0265417
R16552 VPWR VPWR.n4834 0.0265417
R16553 VPWR.n1112 VPWR.n1111 0.0265417
R16554 VPWR.n4595 VPWR.n4594 0.0265417
R16555 VPWR.n1400 VPWR.n1399 0.0265417
R16556 VPWR.n3792 VPWR.n3791 0.0265417
R16557 VPWR.n4247 VPWR.n4246 0.0265417
R16558 VPWR.n1510 VPWR.n1509 0.0265417
R16559 VPWR.n2096 VPWR.n2095 0.0265417
R16560 VPWR.n3567 VPWR.n3566 0.0265417
R16561 VPWR.n2837 VPWR.n2836 0.0265417
R16562 VPWR.n3468 VPWR.n3467 0.0265417
R16563 VPWR.n6547 VPWR.n6546 0.0265417
R16564 VPWR.n7744 VPWR.n7743 0.0265417
R16565 VPWR.n3094 VPWR.n3093 0.0265417
R16566 VPWR.n3184 VPWR.n3183 0.0265417
R16567 VPWR.n6196 VPWR.n6195 0.0265417
R16568 VPWR.n6094 VPWR.n6093 0.0265417
R16569 VPWR.n4277 VPWR.n4276 0.0260562
R16570 VPWR.n3959 VPWR.n3958 0.0260562
R16571 VPWR.n2503 VPWR.n2502 0.0258378
R16572 VPWR.n119 VPWR.n118 0.0258378
R16573 VPWR.n7768 VPWR.n7767 0.0258378
R16574 VPWR.n7747 VPWR.n7746 0.0258378
R16575 VPWR.n7737 VPWR.n7736 0.0258378
R16576 VPWR.n28 VPWR.n27 0.0258378
R16577 VPWR.n243 VPWR.n242 0.0258378
R16578 VPWR.n7615 VPWR.n7614 0.0258378
R16579 VPWR.n156 VPWR.n155 0.0258378
R16580 VPWR.n6593 VPWR.n6592 0.0258378
R16581 VPWR.n6596 VPWR.n6595 0.0258378
R16582 VPWR.n4944 VPWR.n4943 0.0258378
R16583 VPWR.n6679 VPWR.n6678 0.0258378
R16584 VPWR.n272 VPWR.n271 0.0258378
R16585 VPWR.n6784 VPWR.n6783 0.0258378
R16586 VPWR.n6787 VPWR.n6786 0.0258378
R16587 VPWR.n7000 VPWR.n6999 0.0258378
R16588 VPWR.n7003 VPWR.n7002 0.0258378
R16589 VPWR.n4885 VPWR.n4884 0.0258378
R16590 VPWR.n4890 VPWR.n4889 0.0258378
R16591 VPWR.n7385 VPWR.n7384 0.0258378
R16592 VPWR.n7158 VPWR.n7157 0.0258378
R16593 VPWR.n7208 VPWR.n7207 0.0258378
R16594 VPWR.n5289 VPWR.n5288 0.0258378
R16595 VPWR.n5291 VPWR.n5290 0.0258378
R16596 VPWR.n7013 VPWR.n7012 0.0258378
R16597 VPWR.n7042 VPWR.n7041 0.0258378
R16598 VPWR.n4778 VPWR.n4776 0.0258378
R16599 VPWR.n592 VPWR.n591 0.0258378
R16600 VPWR.n881 VPWR.n880 0.0258378
R16601 VPWR.n617 VPWR.n616 0.0258378
R16602 VPWR.n620 VPWR.n619 0.0258378
R16603 VPWR.n630 VPWR.n629 0.0258378
R16604 VPWR.n709 VPWR.n708 0.0258378
R16605 VPWR.n4744 VPWR.n4743 0.0258378
R16606 VPWR.n4562 VPWR.n4561 0.0258378
R16607 VPWR.n4565 VPWR.n4564 0.0258378
R16608 VPWR.n4426 VPWR.n4425 0.0258378
R16609 VPWR.n4429 VPWR.n4428 0.0258378
R16610 VPWR.n413 VPWR.n412 0.0258378
R16611 VPWR.n1107 VPWR.n1106 0.0258378
R16612 VPWR.n3752 VPWR.n3751 0.0258378
R16613 VPWR.n4290 VPWR.n4289 0.0258378
R16614 VPWR.n4293 VPWR.n4292 0.0258378
R16615 VPWR.n1408 VPWR.n1407 0.0258378
R16616 VPWR.n1410 VPWR.n1409 0.0258378
R16617 VPWR.n4397 VPWR.n4396 0.0258378
R16618 VPWR.n4402 VPWR.n4401 0.0258378
R16619 VPWR.n3976 VPWR.n3975 0.0258378
R16620 VPWR.n1518 VPWR.n1517 0.0258378
R16621 VPWR.n1508 VPWR.n1507 0.0258378
R16622 VPWR.n1640 VPWR.n1639 0.0258378
R16623 VPWR.n2031 VPWR.n2030 0.0258378
R16624 VPWR.n1457 VPWR.n1456 0.0258378
R16625 VPWR.n4252 VPWR.n4251 0.0258378
R16626 VPWR.n3531 VPWR.n3530 0.0258378
R16627 VPWR.n3534 VPWR.n3533 0.0258378
R16628 VPWR.n3723 VPWR.n3722 0.0258378
R16629 VPWR.n2107 VPWR.n2106 0.0258378
R16630 VPWR.n1589 VPWR.n1588 0.0258378
R16631 VPWR.n2054 VPWR.n2053 0.0258378
R16632 VPWR.n2059 VPWR.n2058 0.0258378
R16633 VPWR.n4950 VPWR.n4949 0.0258378
R16634 VPWR.n4953 VPWR.n4952 0.0258378
R16635 VPWR.n5803 VPWR.n5802 0.0258378
R16636 VPWR.n5808 VPWR.n5807 0.0258378
R16637 VPWR.n3414 VPWR.n2272 0.0258378
R16638 VPWR.n2778 VPWR.n2777 0.0258378
R16639 VPWR.n2195 VPWR.n2194 0.0258378
R16640 VPWR.n2200 VPWR.n2199 0.0258378
R16641 VPWR.n3499 VPWR.n3498 0.0258378
R16642 VPWR.n2477 VPWR.n2476 0.0258378
R16643 VPWR.n3025 VPWR.n3024 0.0258378
R16644 VPWR.n3030 VPWR.n3029 0.0258378
R16645 VPWR.n2463 VPWR.n2462 0.0258378
R16646 VPWR.n2467 VPWR.n2466 0.0258378
R16647 VPWR.n5785 VPWR.n5784 0.0258378
R16648 VPWR.n5788 VPWR.n5787 0.0258378
R16649 VPWR.n5773 VPWR.n5772 0.0258378
R16650 VPWR.n5778 VPWR.n5777 0.0258378
R16651 VPWR.n2411 VPWR.n2410 0.0258378
R16652 VPWR.n3193 VPWR.n3192 0.0258378
R16653 VPWR.n2388 VPWR.n2387 0.0258378
R16654 VPWR.n3206 VPWR.n3205 0.0258378
R16655 VPWR.n6070 VPWR.n6069 0.0258378
R16656 VPWR.n6063 VPWR.n6062 0.0258378
R16657 VPWR.n6061 VPWR.n6060 0.0258378
R16658 VPWR.n7805 VPWR.n7804 0.0258378
R16659 VPWR.n5068 VPWR.n5067 0.0258378
R16660 VPWR.n5728 VPWR.n5727 0.0258378
R16661 VPWR.n6013 VPWR.n6012 0.0258378
R16662 VPWR.n6681 VPWR.n4942 0.0252396
R16663 VPWR.n6660 VPWR.n6659 0.0252396
R16664 VPWR.n7625 VPWR.n153 0.0252396
R16665 VPWR.n5481 VPWR.n5480 0.0252396
R16666 VPWR.n5470 VPWR.n5469 0.0252396
R16667 VPWR.n6917 VPWR.n6916 0.0252396
R16668 VPWR.n6904 VPWR.n6903 0.0252396
R16669 VPWR.n7039 VPWR.n7038 0.0252396
R16670 VPWR.n7030 VPWR.n7029 0.0252396
R16671 VPWR.n7190 VPWR.n7189 0.0252396
R16672 VPWR VPWR.n7140 0.0252396
R16673 VPWR.n712 VPWR.n711 0.0252396
R16674 VPWR.n717 VPWR.n605 0.0252396
R16675 VPWR.n866 VPWR.n865 0.0252396
R16676 VPWR.n1109 VPWR.n1103 0.0252396
R16677 VPWR.n403 VPWR.n400 0.0252396
R16678 VPWR.n4546 VPWR.n4545 0.0252396
R16679 VPWR.n4592 VPWR.n379 0.0252396
R16680 VPWR.n1397 VPWR.n1396 0.0252396
R16681 VPWR.n1383 VPWR.n1382 0.0252396
R16682 VPWR.n4322 VPWR.n4321 0.0252396
R16683 VPWR.n4244 VPWR.n4243 0.0252396
R16684 VPWR.n4235 VPWR.n4234 0.0252396
R16685 VPWR.n4170 VPWR.n4169 0.0252396
R16686 VPWR.n4156 VPWR.n4155 0.0252396
R16687 VPWR.n2093 VPWR.n2092 0.0252396
R16688 VPWR.n2079 VPWR.n2078 0.0252396
R16689 VPWR.n3550 VPWR.n3549 0.0252396
R16690 VPWR.n3564 VPWR.n3563 0.0252396
R16691 VPWR.n2840 VPWR.n2839 0.0252396
R16692 VPWR.n2849 VPWR.n2848 0.0252396
R16693 VPWR.n3485 VPWR.n3484 0.0252396
R16694 VPWR.n3471 VPWR.n3470 0.0252396
R16695 VPWR.n6550 VPWR.n6549 0.0252396
R16696 VPWR.n6564 VPWR.n6563 0.0252396
R16697 VPWR.n7781 VPWR.n7780 0.0252396
R16698 VPWR.n7771 VPWR.n7770 0.0252396
R16699 VPWR.n3091 VPWR.n3090 0.0252396
R16700 VPWR.n3077 VPWR.n3076 0.0252396
R16701 VPWR.n3171 VPWR.n3170 0.0252396
R16702 VPWR.n3181 VPWR.n3180 0.0252396
R16703 VPWR.n6193 VPWR.n6192 0.0252396
R16704 VPWR.n6179 VPWR.n6178 0.0252396
R16705 VPWR.n6107 VPWR.n6106 0.0252396
R16706 VPWR.n6097 VPWR.n6096 0.0252396
R16707 VPWR.n2506 VPWR.n2505 0.0241486
R16708 VPWR.n107 VPWR.n106 0.0241486
R16709 VPWR.n7790 VPWR.n7789 0.0241486
R16710 VPWR.n165 VPWR.n164 0.0241486
R16711 VPWR.n6765 VPWR.n6764 0.0241486
R16712 VPWR.n5207 VPWR.n5206 0.0241486
R16713 VPWR.n6604 VPWR.n6584 0.0241486
R16714 VPWR.n282 VPWR.n281 0.0241486
R16715 VPWR.n6776 VPWR.n6775 0.0241486
R16716 VPWR.n5578 VPWR.n5577 0.0241486
R16717 VPWR.n6993 VPWR.n4915 0.0241486
R16718 VPWR.n7289 VPWR.n7288 0.0241486
R16719 VPWR.n7200 VPWR.n7199 0.0241486
R16720 VPWR.n5221 VPWR.n5220 0.0241486
R16721 VPWR.n7064 VPWR.n4876 0.0241486
R16722 VPWR.n327 VPWR.n326 0.0241486
R16723 VPWR.n873 VPWR.n872 0.0241486
R16724 VPWR.n468 VPWR.n467 0.0241486
R16725 VPWR.n736 VPWR.n609 0.0241486
R16726 VPWR.n4679 VPWR.n4678 0.0241486
R16727 VPWR.n4554 VPWR.n4553 0.0241486
R16728 VPWR.n1016 VPWR.n1015 0.0241486
R16729 VPWR.n4441 VPWR.n4440 0.0241486
R16730 VPWR.n3954 VPWR.n3953 0.0241486
R16731 VPWR.n4282 VPWR.n4281 0.0241486
R16732 VPWR.n1221 VPWR.n1220 0.0241486
R16733 VPWR.n4390 VPWR.n426 0.0241486
R16734 VPWR.n1542 VPWR.n1541 0.0241486
R16735 VPWR.n1500 VPWR.n1499 0.0241486
R16736 VPWR.n1839 VPWR.n1838 0.0241486
R16737 VPWR.n1472 VPWR.n1466 0.0241486
R16738 VPWR.n1802 VPWR.n1801 0.0241486
R16739 VPWR.n3543 VPWR.n2158 0.0241486
R16740 VPWR.n3711 VPWR.n3710 0.0241486
R16741 VPWR.n2073 VPWR.n1633 0.0241486
R16742 VPWR.n6569 VPWR.n4975 0.0241486
R16743 VPWR.n2276 VPWR.n2275 0.0241486
R16744 VPWR.n2688 VPWR.n2687 0.0241486
R16745 VPWR.n3491 VPWR.n3490 0.0241486
R16746 VPWR.n2812 VPWR.n2809 0.0241486
R16747 VPWR.n3070 VPWR.n2455 0.0241486
R16748 VPWR.n5819 VPWR.n5753 0.0241486
R16749 VPWR.n3161 VPWR.n3155 0.0241486
R16750 VPWR.n6083 VPWR.n6082 0.0241486
R16751 VPWR.n5071 VPWR.n5070 0.0241486
R16752 VPWR.n5731 VPWR.n5730 0.0241486
R16753 VPWR.n3368 VPWR.n3367 0.0241486
R16754 VPWR.n5908 VPWR.n5907 0.0241486
R16755 VPWR.n7457 VPWR 0.0239375
R16756 VPWR.n7349 VPWR 0.0239375
R16757 VPWR VPWR.n676 0.0239375
R16758 VPWR.n765 VPWR 0.0239375
R16759 VPWR.n815 VPWR 0.0239375
R16760 VPWR VPWR.n856 0.0239375
R16761 VPWR.n4529 VPWR 0.0239375
R16762 VPWR.n4647 VPWR 0.0239375
R16763 VPWR.n4361 VPWR 0.0239375
R16764 VPWR.n4352 VPWR 0.0239375
R16765 VPWR.n3789 VPWR 0.0239375
R16766 VPWR.n3855 VPWR 0.0239375
R16767 VPWR.n3907 VPWR 0.0239375
R16768 VPWR.n4199 VPWR 0.0239375
R16769 VPWR.n4174 VPWR 0.0239375
R16770 VPWR.n4098 VPWR 0.0239375
R16771 VPWR.n2151 VPWR 0.0239375
R16772 VPWR.n65 VPWR 0.0239375
R16773 VPWR VPWR.n5102 0.0226354
R16774 VPWR VPWR.n5103 0.0226354
R16775 VPWR.n5191 VPWR 0.0226354
R16776 VPWR.n5186 VPWR 0.0226354
R16777 VPWR.n5179 VPWR 0.0226354
R16778 VPWR.n5172 VPWR 0.0226354
R16779 VPWR.n5166 VPWR 0.0226354
R16780 VPWR.n5146 VPWR 0.0226354
R16781 VPWR.n6653 VPWR 0.0226354
R16782 VPWR.n6628 VPWR 0.0226354
R16783 VPWR.n6617 VPWR 0.0226354
R16784 VPWR.n6733 VPWR 0.0226354
R16785 VPWR.n7587 VPWR 0.0226354
R16786 VPWR.n7531 VPWR 0.0226354
R16787 VPWR VPWR.n7557 0.0226354
R16788 VPWR.n7566 VPWR 0.0226354
R16789 VPWR.n7580 VPWR 0.0226354
R16790 VPWR.n7526 VPWR 0.0226354
R16791 VPWR.n194 VPWR 0.0226354
R16792 VPWR.n183 VPWR 0.0226354
R16793 VPWR.n180 VPWR 0.0226354
R16794 VPWR.n179 VPWR 0.0226354
R16795 VPWR.n5432 VPWR 0.0226354
R16796 VPWR VPWR.n5441 0.0226354
R16797 VPWR.n5443 VPWR 0.0226354
R16798 VPWR.n5562 VPWR 0.0226354
R16799 VPWR.n5539 VPWR 0.0226354
R16800 VPWR.n5527 VPWR 0.0226354
R16801 VPWR.n5502 VPWR 0.0226354
R16802 VPWR.n5497 VPWR 0.0226354
R16803 VPWR.n6984 VPWR 0.0226354
R16804 VPWR.n6974 VPWR 0.0226354
R16805 VPWR.n6963 VPWR 0.0226354
R16806 VPWR.n6960 VPWR 0.0226354
R16807 VPWR.n6956 VPWR 0.0226354
R16808 VPWR.n6947 VPWR 0.0226354
R16809 VPWR.n6926 VPWR 0.0226354
R16810 VPWR.n6922 VPWR 0.0226354
R16811 VPWR.n6857 VPWR 0.0226354
R16812 VPWR VPWR.n6804 0.0226354
R16813 VPWR VPWR.n6819 0.0226354
R16814 VPWR VPWR.n6836 0.0226354
R16815 VPWR.n6837 VPWR 0.0226354
R16816 VPWR VPWR.n6849 0.0226354
R16817 VPWR.n7466 VPWR 0.0226354
R16818 VPWR.n7460 VPWR 0.0226354
R16819 VPWR.n7451 VPWR 0.0226354
R16820 VPWR.n7446 VPWR 0.0226354
R16821 VPWR VPWR.n5358 0.0226354
R16822 VPWR.n5359 VPWR 0.0226354
R16823 VPWR VPWR.n5362 0.0226354
R16824 VPWR VPWR.n5374 0.0226354
R16825 VPWR.n5315 VPWR 0.0226354
R16826 VPWR.n5247 VPWR 0.0226354
R16827 VPWR VPWR.n5252 0.0226354
R16828 VPWR.n5275 VPWR 0.0226354
R16829 VPWR VPWR.n7072 0.0226354
R16830 VPWR.n7074 VPWR 0.0226354
R16831 VPWR.n7079 VPWR 0.0226354
R16832 VPWR VPWR.n7093 0.0226354
R16833 VPWR VPWR.n7095 0.0226354
R16834 VPWR VPWR.n7116 0.0226354
R16835 VPWR VPWR.n7117 0.0226354
R16836 VPWR.n7118 VPWR 0.0226354
R16837 VPWR.n7259 VPWR 0.0226354
R16838 VPWR.n7249 VPWR 0.0226354
R16839 VPWR.n7246 VPWR 0.0226354
R16840 VPWR.n7240 VPWR 0.0226354
R16841 VPWR VPWR.n7278 0.0226354
R16842 VPWR.n7316 VPWR 0.0226354
R16843 VPWR.n7352 VPWR 0.0226354
R16844 VPWR.n7340 VPWR 0.0226354
R16845 VPWR.n7339 VPWR 0.0226354
R16846 VPWR.n7331 VPWR 0.0226354
R16847 VPWR.n488 VPWR 0.0226354
R16848 VPWR VPWR.n491 0.0226354
R16849 VPWR.n492 VPWR 0.0226354
R16850 VPWR.n959 VPWR 0.0226354
R16851 VPWR VPWR.n655 0.0226354
R16852 VPWR.n656 VPWR 0.0226354
R16853 VPWR.n660 VPWR 0.0226354
R16854 VPWR.n669 VPWR 0.0226354
R16855 VPWR.n760 VPWR 0.0226354
R16856 VPWR VPWR.n782 0.0226354
R16857 VPWR.n804 VPWR 0.0226354
R16858 VPWR VPWR.n814 0.0226354
R16859 VPWR VPWR.n900 0.0226354
R16860 VPWR.n901 VPWR 0.0226354
R16861 VPWR VPWR.n905 0.0226354
R16862 VPWR.n907 VPWR 0.0226354
R16863 VPWR.n581 VPWR 0.0226354
R16864 VPWR VPWR.n945 0.0226354
R16865 VPWR.n4765 VPWR 0.0226354
R16866 VPWR.n4831 VPWR 0.0226354
R16867 VPWR.n4814 VPWR 0.0226354
R16868 VPWR.n4807 VPWR 0.0226354
R16869 VPWR.n4802 VPWR 0.0226354
R16870 VPWR VPWR.n1029 0.0226354
R16871 VPWR.n1032 VPWR 0.0226354
R16872 VPWR.n1042 VPWR 0.0226354
R16873 VPWR.n1203 VPWR 0.0226354
R16874 VPWR.n1191 VPWR 0.0226354
R16875 VPWR.n1180 VPWR 0.0226354
R16876 VPWR.n1155 VPWR 0.0226354
R16877 VPWR.n1147 VPWR 0.0226354
R16878 VPWR.n1141 VPWR 0.0226354
R16879 VPWR.n1136 VPWR 0.0226354
R16880 VPWR.n4491 VPWR 0.0226354
R16881 VPWR VPWR.n4494 0.0226354
R16882 VPWR VPWR.n4504 0.0226354
R16883 VPWR VPWR.n4521 0.0226354
R16884 VPWR.n4522 VPWR 0.0226354
R16885 VPWR VPWR.n4528 0.0226354
R16886 VPWR VPWR.n4620 0.0226354
R16887 VPWR.n4632 VPWR 0.0226354
R16888 VPWR.n372 VPWR 0.0226354
R16889 VPWR VPWR.n4637 0.0226354
R16890 VPWR VPWR.n4646 0.0226354
R16891 VPWR.n4661 VPWR 0.0226354
R16892 VPWR VPWR.n4664 0.0226354
R16893 VPWR.n4666 VPWR 0.0226354
R16894 VPWR.n364 VPWR 0.0226354
R16895 VPWR.n361 VPWR 0.0226354
R16896 VPWR.n350 VPWR 0.0226354
R16897 VPWR.n349 VPWR 0.0226354
R16898 VPWR.n344 VPWR 0.0226354
R16899 VPWR.n1240 VPWR 0.0226354
R16900 VPWR.n1227 VPWR 0.0226354
R16901 VPWR VPWR.n1322 0.0226354
R16902 VPWR.n1329 VPWR 0.0226354
R16903 VPWR.n1340 VPWR 0.0226354
R16904 VPWR.n1358 VPWR 0.0226354
R16905 VPWR VPWR.n1367 0.0226354
R16906 VPWR.n1369 VPWR 0.0226354
R16907 VPWR VPWR.n1377 0.0226354
R16908 VPWR.n1428 VPWR 0.0226354
R16909 VPWR.n1427 VPWR 0.0226354
R16910 VPWR.n4364 VPWR 0.0226354
R16911 VPWR.n4355 VPWR 0.0226354
R16912 VPWR.n4348 VPWR 0.0226354
R16913 VPWR VPWR.n3814 0.0226354
R16914 VPWR.n3860 VPWR 0.0226354
R16915 VPWR.n3856 VPWR 0.0226354
R16916 VPWR.n3850 VPWR 0.0226354
R16917 VPWR.n3836 VPWR 0.0226354
R16918 VPWR.n3870 VPWR 0.0226354
R16919 VPWR.n3918 VPWR 0.0226354
R16920 VPWR.n3912 VPWR 0.0226354
R16921 VPWR.n3909 VPWR 0.0226354
R16922 VPWR.n3899 VPWR 0.0226354
R16923 VPWR.n3890 VPWR 0.0226354
R16924 VPWR VPWR.n1850 0.0226354
R16925 VPWR.n1851 VPWR 0.0226354
R16926 VPWR.n1856 VPWR 0.0226354
R16927 VPWR VPWR.n1866 0.0226354
R16928 VPWR.n1867 VPWR 0.0226354
R16929 VPWR VPWR.n1872 0.0226354
R16930 VPWR.n1875 VPWR 0.0226354
R16931 VPWR.n1945 VPWR 0.0226354
R16932 VPWR.n1950 VPWR 0.0226354
R16933 VPWR VPWR.n1958 0.0226354
R16934 VPWR.n1985 VPWR 0.0226354
R16935 VPWR VPWR.n1998 0.0226354
R16936 VPWR.n1999 VPWR 0.0226354
R16937 VPWR.n2005 VPWR 0.0226354
R16938 VPWR VPWR.n2008 0.0226354
R16939 VPWR.n2014 VPWR 0.0226354
R16940 VPWR.n4219 VPWR 0.0226354
R16941 VPWR.n4215 VPWR 0.0226354
R16942 VPWR.n4195 VPWR 0.0226354
R16943 VPWR.n4188 VPWR 0.0226354
R16944 VPWR.n4178 VPWR 0.0226354
R16945 VPWR.n4107 VPWR 0.0226354
R16946 VPWR.n4078 VPWR 0.0226354
R16947 VPWR.n4070 VPWR 0.0226354
R16948 VPWR.n4068 VPWR 0.0226354
R16949 VPWR.n4021 VPWR 0.0226354
R16950 VPWR.n4007 VPWR 0.0226354
R16951 VPWR.n4000 VPWR 0.0226354
R16952 VPWR.n1680 VPWR 0.0226354
R16953 VPWR.n1686 VPWR 0.0226354
R16954 VPWR VPWR.n1697 0.0226354
R16955 VPWR VPWR.n1736 0.0226354
R16956 VPWR.n1792 VPWR 0.0226354
R16957 VPWR.n1763 VPWR 0.0226354
R16958 VPWR.n1757 VPWR 0.0226354
R16959 VPWR.n1754 VPWR 0.0226354
R16960 VPWR.n1747 VPWR 0.0226354
R16961 VPWR.n1746 VPWR 0.0226354
R16962 VPWR.n1605 VPWR 0.0226354
R16963 VPWR.n1597 VPWR 0.0226354
R16964 VPWR.n1595 VPWR 0.0226354
R16965 VPWR.n2125 VPWR 0.0226354
R16966 VPWR VPWR.n2150 0.0226354
R16967 VPWR VPWR.n3599 0.0226354
R16968 VPWR VPWR.n3600 0.0226354
R16969 VPWR.n3618 VPWR 0.0226354
R16970 VPWR.n3624 VPWR 0.0226354
R16971 VPWR VPWR.n3634 0.0226354
R16972 VPWR.n3682 VPWR 0.0226354
R16973 VPWR.n3679 VPWR 0.0226354
R16974 VPWR.n3665 VPWR 0.0226354
R16975 VPWR.n3662 VPWR 0.0226354
R16976 VPWR.n3657 VPWR 0.0226354
R16977 VPWR.n3655 VPWR 0.0226354
R16978 VPWR.n3650 VPWR 0.0226354
R16979 VPWR.n2700 VPWR 0.0226354
R16980 VPWR VPWR.n2710 0.0226354
R16981 VPWR VPWR.n2711 0.0226354
R16982 VPWR.n2712 VPWR 0.0226354
R16983 VPWR VPWR.n2715 0.0226354
R16984 VPWR.n2989 VPWR 0.0226354
R16985 VPWR.n2986 VPWR 0.0226354
R16986 VPWR.n2981 VPWR 0.0226354
R16987 VPWR.n2971 VPWR 0.0226354
R16988 VPWR.n2946 VPWR 0.0226354
R16989 VPWR.n2942 VPWR 0.0226354
R16990 VPWR.n2855 VPWR 0.0226354
R16991 VPWR.n2867 VPWR 0.0226354
R16992 VPWR VPWR.n2880 0.0226354
R16993 VPWR.n2881 VPWR 0.0226354
R16994 VPWR VPWR.n2891 0.0226354
R16995 VPWR.n2920 VPWR 0.0226354
R16996 VPWR.n3442 VPWR 0.0226354
R16997 VPWR VPWR.n2236 0.0226354
R16998 VPWR VPWR.n2242 0.0226354
R16999 VPWR.n2243 VPWR 0.0226354
R17000 VPWR VPWR.n2268 0.0226354
R17001 VPWR.n2353 VPWR 0.0226354
R17002 VPWR.n2318 VPWR 0.0226354
R17003 VPWR.n2294 VPWR 0.0226354
R17004 VPWR VPWR.n6388 0.0226354
R17005 VPWR.n6389 VPWR 0.0226354
R17006 VPWR VPWR.n6473 0.0226354
R17007 VPWR VPWR.n6496 0.0226354
R17008 VPWR.n6504 VPWR 0.0226354
R17009 VPWR VPWR.n6521 0.0226354
R17010 VPWR.n6527 VPWR 0.0226354
R17011 VPWR.n4988 VPWR 0.0226354
R17012 VPWR.n4994 VPWR 0.0226354
R17013 VPWR VPWR.n5002 0.0226354
R17014 VPWR.n5010 VPWR 0.0226354
R17015 VPWR VPWR.n5015 0.0226354
R17016 VPWR.n5039 VPWR 0.0226354
R17017 VPWR.n5033 VPWR 0.0226354
R17018 VPWR.n5027 VPWR 0.0226354
R17019 VPWR.n5024 VPWR 0.0226354
R17020 VPWR.n5023 VPWR 0.0226354
R17021 VPWR VPWR.n32 0.0226354
R17022 VPWR.n7711 VPWR 0.0226354
R17023 VPWR.n7705 VPWR 0.0226354
R17024 VPWR.n7699 VPWR 0.0226354
R17025 VPWR.n7692 VPWR 0.0226354
R17026 VPWR.n7687 VPWR 0.0226354
R17027 VPWR.n7684 VPWR 0.0226354
R17028 VPWR.n7676 VPWR 0.0226354
R17029 VPWR.n7664 VPWR 0.0226354
R17030 VPWR.n77 VPWR 0.0226354
R17031 VPWR.n69 VPWR 0.0226354
R17032 VPWR.n60 VPWR 0.0226354
R17033 VPWR.n59 VPWR 0.0226354
R17034 VPWR.n2588 VPWR 0.0226354
R17035 VPWR.n2577 VPWR 0.0226354
R17036 VPWR VPWR.n2593 0.0226354
R17037 VPWR VPWR.n2605 0.0226354
R17038 VPWR.n2608 VPWR 0.0226354
R17039 VPWR.n2563 VPWR 0.0226354
R17040 VPWR.n2556 VPWR 0.0226354
R17041 VPWR.n2540 VPWR 0.0226354
R17042 VPWR.n2534 VPWR 0.0226354
R17043 VPWR.n2533 VPWR 0.0226354
R17044 VPWR VPWR.n2518 0.0226354
R17045 VPWR.n2528 VPWR 0.0226354
R17046 VPWR.n2521 VPWR 0.0226354
R17047 VPWR.n3114 VPWR 0.0226354
R17048 VPWR.n2453 VPWR 0.0226354
R17049 VPWR.n2444 VPWR 0.0226354
R17050 VPWR.n2439 VPWR 0.0226354
R17051 VPWR.n2438 VPWR 0.0226354
R17052 VPWR.n3122 VPWR 0.0226354
R17053 VPWR VPWR.n3136 0.0226354
R17054 VPWR VPWR.n3225 0.0226354
R17055 VPWR.n3266 VPWR 0.0226354
R17056 VPWR.n3245 VPWR 0.0226354
R17057 VPWR.n3241 VPWR 0.0226354
R17058 VPWR VPWR.n3229 0.0226354
R17059 VPWR.n3237 VPWR 0.0226354
R17060 VPWR.n3232 VPWR 0.0226354
R17061 VPWR.n3288 VPWR 0.0226354
R17062 VPWR.n3323 VPWR 0.0226354
R17063 VPWR.n3320 VPWR 0.0226354
R17064 VPWR.n3319 VPWR 0.0226354
R17065 VPWR VPWR.n3304 0.0226354
R17066 VPWR.n6296 VPWR 0.0226354
R17067 VPWR VPWR.n6308 0.0226354
R17068 VPWR.n6311 VPWR 0.0226354
R17069 VPWR.n6266 VPWR 0.0226354
R17070 VPWR.n6258 VPWR 0.0226354
R17071 VPWR.n6249 VPWR 0.0226354
R17072 VPWR.n6231 VPWR 0.0226354
R17073 VPWR.n6230 VPWR 0.0226354
R17074 VPWR.n6162 VPWR 0.0226354
R17075 VPWR.n6159 VPWR 0.0226354
R17076 VPWR.n6131 VPWR 0.0226354
R17077 VPWR.n6123 VPWR 0.0226354
R17078 VPWR.n6114 VPWR 0.0226354
R17079 VPWR.n6111 VPWR 0.0226354
R17080 VPWR VPWR.n5847 0.0226354
R17081 VPWR.n5858 VPWR 0.0226354
R17082 VPWR.n5883 VPWR 0.0226354
R17083 VPWR.n5890 VPWR 0.0226354
R17084 VPWR VPWR.n5903 0.0226354
R17085 VPWR.n5958 VPWR 0.0226354
R17086 VPWR.n5952 VPWR 0.0226354
R17087 VPWR.n5941 VPWR 0.0226354
R17088 VPWR.n2667 VPWR.n2666 0.0224595
R17089 VPWR.n2674 VPWR.n2673 0.0224595
R17090 VPWR.n2655 VPWR.n2654 0.0224595
R17091 VPWR.n2658 VPWR.n2657 0.0224595
R17092 VPWR.n125 VPWR.n121 0.0224595
R17093 VPWR.n124 VPWR.n123 0.0224595
R17094 VPWR.n7645 VPWR.n7644 0.0224595
R17095 VPWR.n7648 VPWR.n7647 0.0224595
R17096 VPWR.n7767 VPWR.n7766 0.0224595
R17097 VPWR.n7764 VPWR.n7749 0.0224595
R17098 VPWR.n250 VPWR.n245 0.0224595
R17099 VPWR.n249 VPWR.n248 0.0224595
R17100 VPWR.n7502 VPWR.n7501 0.0224595
R17101 VPWR.n7505 VPWR.n7504 0.0224595
R17102 VPWR.n135 VPWR.n134 0.0224595
R17103 VPWR.n140 VPWR.n139 0.0224595
R17104 VPWR.n5078 VPWR.n5077 0.0224595
R17105 VPWR.n5085 VPWR.n5084 0.0224595
R17106 VPWR.n5088 VPWR.n5087 0.0224595
R17107 VPWR.n5677 VPWR.n5676 0.0224595
R17108 VPWR.n6675 VPWR.n4946 0.0224595
R17109 VPWR.n6678 VPWR.n6677 0.0224595
R17110 VPWR.n7493 VPWR.n274 0.0224595
R17111 VPWR.n7492 VPWR.n7491 0.0224595
R17112 VPWR.n260 VPWR.n259 0.0224595
R17113 VPWR.n6900 VPWR.n6899 0.0224595
R17114 VPWR.n6897 VPWR.n4931 0.0224595
R17115 VPWR.n5632 VPWR.n5631 0.0224595
R17116 VPWR.n5639 VPWR.n5638 0.0224595
R17117 VPWR.n5642 VPWR.n5641 0.0224595
R17118 VPWR.n5646 VPWR.n5645 0.0224595
R17119 VPWR.n4893 VPWR.n4887 0.0224595
R17120 VPWR.n4891 VPWR.n4890 0.0224595
R17121 VPWR.n7393 VPWR.n7387 0.0224595
R17122 VPWR.n7392 VPWR.n7391 0.0224595
R17123 VPWR.n7314 VPWR.n287 0.0224595
R17124 VPWR.n7151 VPWR.n7150 0.0224595
R17125 VPWR.n7166 VPWR.n7165 0.0224595
R17126 VPWR.n5397 VPWR.n5395 0.0224595
R17127 VPWR.n5407 VPWR.n5406 0.0224595
R17128 VPWR.n5410 VPWR.n5409 0.0224595
R17129 VPWR.n5414 VPWR.n5413 0.0224595
R17130 VPWR.n7045 VPWR.n7015 0.0224595
R17131 VPWR.n7043 VPWR.n7042 0.0224595
R17132 VPWR.n4852 VPWR.n316 0.0224595
R17133 VPWR.n4851 VPWR.n4850 0.0224595
R17134 VPWR.n305 VPWR.n304 0.0224595
R17135 VPWR.n833 VPWR.n832 0.0224595
R17136 VPWR.n842 VPWR.n841 0.0224595
R17137 VPWR.n533 VPWR.n532 0.0224595
R17138 VPWR.n550 VPWR.n549 0.0224595
R17139 VPWR.n473 VPWR.n472 0.0224595
R17140 VPWR.n563 VPWR.n474 0.0224595
R17141 VPWR.n633 VPWR.n632 0.0224595
R17142 VPWR.n708 VPWR.n707 0.0224595
R17143 VPWR.n4752 VPWR.n4746 0.0224595
R17144 VPWR.n4751 VPWR.n4750 0.0224595
R17145 VPWR.n4732 VPWR.n4731 0.0224595
R17146 VPWR.n4573 VPWR.n4572 0.0224595
R17147 VPWR.n4578 VPWR.n4577 0.0224595
R17148 VPWR.n985 VPWR.n984 0.0224595
R17149 VPWR.n992 VPWR.n991 0.0224595
R17150 VPWR.n995 VPWR.n994 0.0224595
R17151 VPWR.n999 VPWR.n998 0.0224595
R17152 VPWR.n416 VPWR.n415 0.0224595
R17153 VPWR.n1106 VPWR.n1105 0.0224595
R17154 VPWR.n3760 VPWR.n3754 0.0224595
R17155 VPWR.n3759 VPWR.n3758 0.0224595
R17156 VPWR.n3740 VPWR.n3739 0.0224595
R17157 VPWR.n4301 VPWR.n4300 0.0224595
R17158 VPWR.n4306 VPWR.n4305 0.0224595
R17159 VPWR.n451 VPWR.n450 0.0224595
R17160 VPWR.n458 VPWR.n457 0.0224595
R17161 VPWR.n446 VPWR.n445 0.0224595
R17162 VPWR.n1295 VPWR.n1292 0.0224595
R17163 VPWR.n4405 VPWR.n4399 0.0224595
R17164 VPWR.n4403 VPWR.n4402 0.0224595
R17165 VPWR.n3984 VPWR.n3978 0.0224595
R17166 VPWR.n3983 VPWR.n3982 0.0224595
R17167 VPWR.n3964 VPWR.n3963 0.0224595
R17168 VPWR.n4136 VPWR.n4135 0.0224595
R17169 VPWR.n4141 VPWR.n4140 0.0224595
R17170 VPWR.n1889 VPWR.n1887 0.0224595
R17171 VPWR.n1920 VPWR.n1919 0.0224595
R17172 VPWR.n1906 VPWR.n1905 0.0224595
R17173 VPWR.n1910 VPWR.n1909 0.0224595
R17174 VPWR.n4255 VPWR.n4249 0.0224595
R17175 VPWR.n4253 VPWR.n4252 0.0224595
R17176 VPWR.n1660 VPWR.n1659 0.0224595
R17177 VPWR.n1667 VPWR.n1666 0.0224595
R17178 VPWR.n1670 VPWR.n1669 0.0224595
R17179 VPWR.n1821 VPWR.n1820 0.0224595
R17180 VPWR.n2175 VPWR.n2174 0.0224595
R17181 VPWR.n2180 VPWR.n2179 0.0224595
R17182 VPWR.n3730 VPWR.n3725 0.0224595
R17183 VPWR.n3729 VPWR.n3728 0.0224595
R17184 VPWR.n1557 VPWR.n1556 0.0224595
R17185 VPWR.n1560 VPWR.n1559 0.0224595
R17186 VPWR.n2062 VPWR.n2056 0.0224595
R17187 VPWR.n2060 VPWR.n2059 0.0224595
R17188 VPWR.n5811 VPWR.n5805 0.0224595
R17189 VPWR.n5809 VPWR.n5808 0.0224595
R17190 VPWR.n3412 VPWR.n3411 0.0224595
R17191 VPWR.n2338 VPWR.n2273 0.0224595
R17192 VPWR.n2351 VPWR.n2350 0.0224595
R17193 VPWR.n2346 VPWR.n2345 0.0224595
R17194 VPWR.n2730 VPWR.n2729 0.0224595
R17195 VPWR.n2735 VPWR.n2734 0.0224595
R17196 VPWR.n2768 VPWR.n2767 0.0224595
R17197 VPWR.n2780 VPWR.n2775 0.0224595
R17198 VPWR.n2196 VPWR.n2195 0.0224595
R17199 VPWR.n2203 VPWR.n2202 0.0224595
R17200 VPWR.n3033 VPWR.n3027 0.0224595
R17201 VPWR.n3031 VPWR.n3030 0.0224595
R17202 VPWR.n3045 VPWR.n3041 0.0224595
R17203 VPWR.n3043 VPWR.n3042 0.0224595
R17204 VPWR.n5781 VPWR.n5775 0.0224595
R17205 VPWR.n5779 VPWR.n5778 0.0224595
R17206 VPWR.n2412 VPWR.n2411 0.0224595
R17207 VPWR.n3196 VPWR.n3195 0.0224595
R17208 VPWR.n6069 VPWR.n6068 0.0224595
R17209 VPWR.n6066 VPWR.n6065 0.0224595
R17210 VPWR.n6362 VPWR.n6361 0.0224595
R17211 VPWR.n6369 VPWR.n6368 0.0224595
R17212 VPWR.n6420 VPWR.n6419 0.0224595
R17213 VPWR.n6426 VPWR.n6424 0.0224595
R17214 VPWR.n5699 VPWR.n5698 0.0224595
R17215 VPWR.n5706 VPWR.n5705 0.0224595
R17216 VPWR.n5718 VPWR.n5717 0.0224595
R17217 VPWR.n5721 VPWR.n5720 0.0224595
R17218 VPWR.n3378 VPWR.n3375 0.0224595
R17219 VPWR.n3377 VPWR.n3376 0.0224595
R17220 VPWR.n3389 VPWR.n3388 0.0224595
R17221 VPWR.n3392 VPWR.n3391 0.0224595
R17222 VPWR.n6018 VPWR.n6015 0.0224595
R17223 VPWR.n6017 VPWR.n6016 0.0224595
R17224 VPWR.n6001 VPWR.n6000 0.0224595
R17225 VPWR.n5918 VPWR.n5917 0.0224595
R17226 VPWR.n860 VPWR.n859 0.0217384
R17227 VPWR.n5133 VPWR.n5132 0.0213333
R17228 VPWR.n223 VPWR.n222 0.0213333
R17229 VPWR.n5608 VPWR.n5607 0.0213333
R17230 VPWR.n7488 VPWR.n7487 0.0213333
R17231 VPWR.n5392 VPWR 0.0213333
R17232 VPWR VPWR.n5391 0.0213333
R17233 VPWR.n5403 VPWR.n5216 0.0213333
R17234 VPWR VPWR.n5273 0.0213333
R17235 VPWR.n4871 VPWR 0.0213333
R17236 VPWR.n481 VPWR 0.0213333
R17237 VPWR.n554 VPWR.n530 0.0213333
R17238 VPWR.n4847 VPWR.n4846 0.0213333
R17239 VPWR.n4808 VPWR 0.0213333
R17240 VPWR VPWR.n1041 0.0213333
R17241 VPWR.n1067 VPWR.n1066 0.0213333
R17242 VPWR.n4469 VPWR 0.0213333
R17243 VPWR VPWR.n4483 0.0213333
R17244 VPWR.n4711 VPWR.n4710 0.0213333
R17245 VPWR.n1265 VPWR.n1264 0.0213333
R17246 VPWR.n1364 VPWR 0.0213333
R17247 VPWR.n4386 VPWR 0.0213333
R17248 VPWR.n4384 VPWR 0.0213333
R17249 VPWR.n4367 VPWR 0.0213333
R17250 VPWR.n3811 VPWR 0.0213333
R17251 VPWR.n3934 VPWR.n3933 0.0213333
R17252 VPWR.n1884 VPWR 0.0213333
R17253 VPWR VPWR.n1883 0.0213333
R17254 VPWR.n1924 VPWR.n1650 0.0213333
R17255 VPWR.n4228 VPWR 0.0213333
R17256 VPWR.n4206 VPWR 0.0213333
R17257 VPWR.n4114 VPWR 0.0213333
R17258 VPWR.n4109 VPWR 0.0213333
R17259 VPWR.n4038 VPWR.n4037 0.0213333
R17260 VPWR.n1725 VPWR.n1724 0.0213333
R17261 VPWR VPWR.n3617 0.0213333
R17262 VPWR.n3695 VPWR.n3694 0.0213333
R17263 VPWR.n2757 VPWR.n2756 0.0213333
R17264 VPWR.n6436 VPWR.n6435 0.0213333
R17265 VPWR.n93 VPWR.n92 0.0213333
R17266 VPWR.n2627 VPWR.n2626 0.0213333
R17267 VPWR.n3343 VPWR.n3342 0.0213333
R17268 VPWR.n6330 VPWR.n6329 0.0213333
R17269 VPWR VPWR.n5889 0.0213333
R17270 VPWR.n5978 VPWR.n5977 0.0213333
R17271 VPWR.n115 VPWR.n114 0.0202124
R17272 VPWR.n7653 VPWR.n7652 0.0202124
R17273 VPWR.n241 VPWR.n240 0.0202124
R17274 VPWR.n7510 VPWR.n7509 0.0202124
R17275 VPWR.n133 VPWR.n132 0.0202124
R17276 VPWR.n7608 VPWR.n7607 0.0202124
R17277 VPWR.n5075 VPWR.n5074 0.0202124
R17278 VPWR.n5209 VPWR.n5208 0.0202124
R17279 VPWR.n4948 VPWR.n4947 0.0202124
R17280 VPWR.n6586 VPWR.n6585 0.0202124
R17281 VPWR.n258 VPWR.n257 0.0202124
R17282 VPWR.n7431 VPWR.n7430 0.0202124
R17283 VPWR.n4933 VPWR.n4932 0.0202124
R17284 VPWR.n6780 VPWR.n6779 0.0202124
R17285 VPWR.n5629 VPWR.n5628 0.0202124
R17286 VPWR.n5580 VPWR.n5579 0.0202124
R17287 VPWR.n4883 VPWR.n4882 0.0202124
R17288 VPWR.n4910 VPWR.n4909 0.0202124
R17289 VPWR.n286 VPWR.n285 0.0202124
R17290 VPWR.n7321 VPWR.n7320 0.0202124
R17291 VPWR.n7147 VPWR.n7146 0.0202124
R17292 VPWR.n296 VPWR.n295 0.0202124
R17293 VPWR.n5213 VPWR.n5212 0.0202124
R17294 VPWR.n5223 VPWR.n5222 0.0202124
R17295 VPWR.n7011 VPWR.n7010 0.0202124
R17296 VPWR.n4878 VPWR.n4877 0.0202124
R17297 VPWR.n303 VPWR.n302 0.0202124
R17298 VPWR.n4791 VPWR.n4790 0.0202124
R17299 VPWR.n830 VPWR.n829 0.0202124
R17300 VPWR.n595 VPWR.n594 0.0202124
R17301 VPWR.n537 VPWR.n536 0.0202124
R17302 VPWR.n462 VPWR.n461 0.0202124
R17303 VPWR.n628 VPWR.n627 0.0202124
R17304 VPWR.n611 VPWR.n610 0.0202124
R17305 VPWR.n4730 VPWR.n4729 0.0202124
R17306 VPWR.n331 VPWR.n330 0.0202124
R17307 VPWR.n386 VPWR.n385 0.0202124
R17308 VPWR.n4558 VPWR.n4557 0.0202124
R17309 VPWR.n982 VPWR.n981 0.0202124
R17310 VPWR.n1010 VPWR.n1009 0.0202124
R17311 VPWR.n411 VPWR.n410 0.0202124
R17312 VPWR.n4435 VPWR.n4434 0.0202124
R17313 VPWR.n3738 VPWR.n3737 0.0202124
R17314 VPWR.n3764 VPWR.n3763 0.0202124
R17315 VPWR.n1449 VPWR.n1448 0.0202124
R17316 VPWR.n4286 VPWR.n4285 0.0202124
R17317 VPWR.n448 VPWR.n447 0.0202124
R17318 VPWR.n1215 VPWR.n1214 0.0202124
R17319 VPWR.n4395 VPWR.n4394 0.0202124
R17320 VPWR.n421 VPWR.n420 0.0202124
R17321 VPWR.n3962 VPWR.n3961 0.0202124
R17322 VPWR.n3988 VPWR.n3987 0.0202124
R17323 VPWR.n1495 VPWR.n1494 0.0202124
R17324 VPWR.n1504 VPWR.n1503 0.0202124
R17325 VPWR.n1653 VPWR.n1652 0.0202124
R17326 VPWR.n1833 VPWR.n1832 0.0202124
R17327 VPWR.n1455 VPWR.n1454 0.0202124
R17328 VPWR.n1468 VPWR.n1467 0.0202124
R17329 VPWR.n1657 VPWR.n1656 0.0202124
R17330 VPWR.n1804 VPWR.n1803 0.0202124
R17331 VPWR.n2162 VPWR.n2161 0.0202124
R17332 VPWR.n3526 VPWR.n3525 0.0202124
R17333 VPWR.n3718 VPWR.n3717 0.0202124
R17334 VPWR.n1554 VPWR.n1553 0.0202124
R17335 VPWR.n2039 VPWR.n2038 0.0202124
R17336 VPWR.n1635 VPWR.n1634 0.0202124
R17337 VPWR.n5796 VPWR.n5795 0.0202124
R17338 VPWR.n4968 VPWR.n4967 0.0202124
R17339 VPWR.n2282 VPWR.n2281 0.0202124
R17340 VPWR.n2739 VPWR.n2738 0.0202124
R17341 VPWR.n2773 VPWR.n2772 0.0202124
R17342 VPWR.n3507 VPWR.n3506 0.0202124
R17343 VPWR.n2192 VPWR.n2191 0.0202124
R17344 VPWR.n3020 VPWR.n3019 0.0202124
R17345 VPWR.n2460 VPWR.n2459 0.0202124
R17346 VPWR.n3064 VPWR.n3063 0.0202124
R17347 VPWR.n5766 VPWR.n5765 0.0202124
R17348 VPWR.n5762 VPWR.n5761 0.0202124
R17349 VPWR.n3158 VPWR.n3157 0.0202124
R17350 VPWR.n3198 VPWR.n3197 0.0202124
R17351 VPWR.n7 VPWR.n6 0.0202124
R17352 VPWR.n16 VPWR.n15 0.0202124
R17353 VPWR.n7792 VPWR.n7791 0.0202124
R17354 VPWR.n6359 VPWR.n6358 0.0202124
R17355 VPWR.n6422 VPWR.n6421 0.0202124
R17356 VPWR.n5691 VPWR.n5690 0.0202124
R17357 VPWR.n5724 VPWR.n5723 0.0202124
R17358 VPWR.n2500 VPWR.n2499 0.0202124
R17359 VPWR.n2381 VPWR.n2380 0.0202124
R17360 VPWR.n3397 VPWR.n3396 0.0202124
R17361 VPWR.n6021 VPWR.n6020 0.0202124
R17362 VPWR.n5996 VPWR.n5995 0.0202124
R17363 VPWR.n5673 VPWR.n5672 0.0200312
R17364 VPWR.n6699 VPWR.n6698 0.0200312
R17365 VPWR.n6694 VPWR.n6693 0.0200312
R17366 VPWR.n6683 VPWR.n6682 0.0200312
R17367 VPWR VPWR.n6750 0.0200312
R17368 VPWR.n7624 VPWR.n7623 0.0200312
R17369 VPWR.n7604 VPWR.n7603 0.0200312
R17370 VPWR.n212 VPWR.n211 0.0200312
R17371 VPWR.n5597 VPWR.n5596 0.0200312
R17372 VPWR.n5493 VPWR.n5492 0.0200312
R17373 VPWR.n5488 VPWR.n5487 0.0200312
R17374 VPWR.n5483 VPWR.n5482 0.0200312
R17375 VPWR.n6871 VPWR.n6870 0.0200312
R17376 VPWR.n7417 VPWR.n7416 0.0200312
R17377 VPWR.n5338 VPWR.n5337 0.0200312
R17378 VPWR.n5300 VPWR.n5299 0.0200312
R17379 VPWR.n7018 VPWR.n7017 0.0200312
R17380 VPWR.n7026 VPWR.n7025 0.0200312
R17381 VPWR.n7027 VPWR 0.0200312
R17382 VPWR.n7212 VPWR.n7211 0.0200312
R17383 VPWR.n7302 VPWR.n7301 0.0200312
R17384 VPWR VPWR.n7315 0.0200312
R17385 VPWR.n567 VPWR.n566 0.0200312
R17386 VPWR.n689 VPWR.n688 0.0200312
R17387 VPWR.n694 VPWR.n693 0.0200312
R17388 VPWR.n705 VPWR.n704 0.0200312
R17389 VPWR.n741 VPWR 0.0200312
R17390 VPWR.n587 VPWR.n586 0.0200312
R17391 VPWR.n885 VPWR.n884 0.0200312
R17392 VPWR.n4779 VPWR.n4775 0.0200312
R17393 VPWR.n1078 VPWR.n1077 0.0200312
R17394 VPWR.n1123 VPWR.n1121 0.0200312
R17395 VPWR.n1117 VPWR.n1116 0.0200312
R17396 VPWR.n1111 VPWR.n1110 0.0200312
R17397 VPWR.n4594 VPWR.n4593 0.0200312
R17398 VPWR.n4600 VPWR.n4599 0.0200312
R17399 VPWR.n4606 VPWR.n4604 0.0200312
R17400 VPWR.n4700 VPWR.n4699 0.0200312
R17401 VPWR.n1299 VPWR.n1298 0.0200312
R17402 VPWR.n1419 VPWR.n1418 0.0200312
R17403 VPWR.n1404 VPWR.n1403 0.0200312
R17404 VPWR.n1399 VPWR.n1398 0.0200312
R17405 VPWR.n3791 VPWR.n3790 0.0200312
R17406 VPWR.n3797 VPWR.n3796 0.0200312
R17407 VPWR.n3802 VPWR.n3801 0.0200312
R17408 VPWR.n3945 VPWR.n3944 0.0200312
R17409 VPWR.n1935 VPWR.n1934 0.0200312
R17410 VPWR.n2023 VPWR.n2022 0.0200312
R17411 VPWR.n2025 VPWR.n2024 0.0200312
R17412 VPWR.n4246 VPWR.n4245 0.0200312
R17413 VPWR.n1509 VPWR.n1488 0.0200312
R17414 VPWR.n1515 VPWR.n1514 0.0200312
R17415 VPWR.n4127 VPWR.n4126 0.0200312
R17416 VPWR.n4030 VPWR.n4029 0.0200312
R17417 VPWR.n1817 VPWR.n1816 0.0200312
R17418 VPWR.n2101 VPWR.n2100 0.0200312
R17419 VPWR.n2095 VPWR.n2094 0.0200312
R17420 VPWR.n3566 VPWR.n3565 0.0200312
R17421 VPWR.n3572 VPWR.n3571 0.0200312
R17422 VPWR.n3578 VPWR.n3576 0.0200312
R17423 VPWR.n3703 VPWR.n3702 0.0200312
R17424 VPWR.n2784 VPWR.n2783 0.0200312
R17425 VPWR.n2827 VPWR.n2826 0.0200312
R17426 VPWR.n2832 VPWR.n2831 0.0200312
R17427 VPWR.n2838 VPWR.n2837 0.0200312
R17428 VPWR.n3469 VPWR.n3468 0.0200312
R17429 VPWR.n3463 VPWR.n3462 0.0200312
R17430 VPWR.n3458 VPWR.n3457 0.0200312
R17431 VPWR.n3416 VPWR.n3415 0.0200312
R17432 VPWR VPWR.n2352 0.0200312
R17433 VPWR.n6417 VPWR.n6416 0.0200312
R17434 VPWR.n6536 VPWR.n6535 0.0200312
R17435 VPWR.n6541 VPWR.n6540 0.0200312
R17436 VPWR.n6548 VPWR.n6547 0.0200312
R17437 VPWR.n7745 VPWR.n7744 0.0200312
R17438 VPWR.n7739 VPWR.n7738 0.0200312
R17439 VPWR.n7731 VPWR.n7730 0.0200312
R17440 VPWR.n101 VPWR.n100 0.0200312
R17441 VPWR.n2638 VPWR.n2637 0.0200312
R17442 VPWR.n3105 VPWR.n3103 0.0200312
R17443 VPWR.n3099 VPWR.n3098 0.0200312
R17444 VPWR.n3093 VPWR.n3092 0.0200312
R17445 VPWR.n3183 VPWR.n3182 0.0200312
R17446 VPWR.n3211 VPWR.n3209 0.0200312
R17447 VPWR.n3354 VPWR.n3353 0.0200312
R17448 VPWR.n6341 VPWR.n6340 0.0200312
R17449 VPWR.n6207 VPWR.n6205 0.0200312
R17450 VPWR.n6201 VPWR.n6200 0.0200312
R17451 VPWR.n6195 VPWR.n6194 0.0200312
R17452 VPWR.n6095 VPWR.n6094 0.0200312
R17453 VPWR.n5833 VPWR.n1 0.0200312
R17454 VPWR.n5967 VPWR.n5966 0.0200312
R17455 VPWR.n2668 VPWR.n2667 0.0190811
R17456 VPWR.n2675 VPWR.n2669 0.0190811
R17457 VPWR.n7651 VPWR.n7650 0.0190811
R17458 VPWR.n7649 VPWR.n7648 0.0190811
R17459 VPWR.n7508 VPWR.n7507 0.0190811
R17460 VPWR.n7506 VPWR.n7505 0.0190811
R17461 VPWR.n150 VPWR.n149 0.0190811
R17462 VPWR.n5079 VPWR.n5078 0.0190811
R17463 VPWR.n5086 VPWR.n5080 0.0190811
R17464 VPWR.n6665 VPWR.n6579 0.0190811
R17465 VPWR.n264 VPWR.n263 0.0190811
R17466 VPWR.n262 VPWR.n261 0.0190811
R17467 VPWR.n6882 VPWR.n6881 0.0190811
R17468 VPWR.n5633 VPWR.n5632 0.0190811
R17469 VPWR.n5640 VPWR.n5634 0.0190811
R17470 VPWR.n4898 VPWR.n4897 0.0190811
R17471 VPWR.n7377 VPWR.n7376 0.0190811
R17472 VPWR.n7375 VPWR.n288 0.0190811
R17473 VPWR.n7144 VPWR.n7143 0.0190811
R17474 VPWR.n5397 VPWR.n5396 0.0190811
R17475 VPWR.n5408 VPWR.n5214 0.0190811
R17476 VPWR.n7050 VPWR.n7049 0.0190811
R17477 VPWR.n309 VPWR.n308 0.0190811
R17478 VPWR.n307 VPWR.n306 0.0190811
R17479 VPWR.n827 VPWR.n826 0.0190811
R17480 VPWR.n534 VPWR.n533 0.0190811
R17481 VPWR.n548 VPWR.n535 0.0190811
R17482 VPWR.n722 VPWR.n637 0.0190811
R17483 VPWR.n4736 VPWR.n4735 0.0190811
R17484 VPWR.n4734 VPWR.n4733 0.0190811
R17485 VPWR.n383 VPWR.n382 0.0190811
R17486 VPWR.n986 VPWR.n985 0.0190811
R17487 VPWR.n993 VPWR.n987 0.0190811
R17488 VPWR.n4456 VPWR.n4455 0.0190811
R17489 VPWR.n3744 VPWR.n3743 0.0190811
R17490 VPWR.n3742 VPWR.n3741 0.0190811
R17491 VPWR.n4316 VPWR.n1446 0.0190811
R17492 VPWR.n452 VPWR.n451 0.0190811
R17493 VPWR.n459 VPWR.n453 0.0190811
R17494 VPWR.n4410 VPWR.n4409 0.0190811
R17495 VPWR.n3968 VPWR.n3967 0.0190811
R17496 VPWR.n3966 VPWR.n3965 0.0190811
R17497 VPWR.n1492 VPWR.n1491 0.0190811
R17498 VPWR.n1889 VPWR.n1888 0.0190811
R17499 VPWR.n1918 VPWR.n1651 0.0190811
R17500 VPWR.n4260 VPWR.n4259 0.0190811
R17501 VPWR.n1661 VPWR.n1660 0.0190811
R17502 VPWR.n1668 VPWR.n1662 0.0190811
R17503 VPWR.n2166 VPWR.n2165 0.0190811
R17504 VPWR.n1563 VPWR.n1562 0.0190811
R17505 VPWR.n1561 VPWR.n1560 0.0190811
R17506 VPWR.n2044 VPWR.n2043 0.0190811
R17507 VPWR.n2349 VPWR.n2348 0.0190811
R17508 VPWR.n2347 VPWR.n2346 0.0190811
R17509 VPWR.n2731 VPWR.n2730 0.0190811
R17510 VPWR.n2736 VPWR.n2732 0.0190811
R17511 VPWR.n3514 VPWR.n3513 0.0190811
R17512 VPWR.n3012 VPWR.n3011 0.0190811
R17513 VPWR.n3060 VPWR.n3059 0.0190811
R17514 VPWR.n2397 VPWR.n2396 0.0190811
R17515 VPWR.n6078 VPWR.n6077 0.0190811
R17516 VPWR.n6363 VPWR.n6362 0.0190811
R17517 VPWR.n6370 VPWR.n6364 0.0190811
R17518 VPWR.n5700 VPWR.n5699 0.0190811
R17519 VPWR.n5707 VPWR.n5701 0.0190811
R17520 VPWR.n3395 VPWR.n3394 0.0190811
R17521 VPWR.n3393 VPWR.n3392 0.0190811
R17522 VPWR.n6004 VPWR.n6003 0.0190811
R17523 VPWR.n6685 VPWR.n6684 0.0187292
R17524 VPWR.n7622 VPWR.n7621 0.0187292
R17525 VPWR.n157 VPWR 0.0187292
R17526 VPWR.n234 VPWR.n232 0.0187292
R17527 VPWR.n5485 VPWR.n5484 0.0187292
R17528 VPWR.n6789 VPWR.n6788 0.0187292
R17529 VPWR.n7409 VPWR.n276 0.0187292
R17530 VPWR.n7478 VPWR.n7477 0.0187292
R17531 VPWR.n7164 VPWR.n7155 0.0187292
R17532 VPWR VPWR.n293 0.0187292
R17533 VPWR.n7369 VPWR.n7367 0.0187292
R17534 VPWR.n703 VPWR.n702 0.0187292
R17535 VPWR.n840 VPWR.n837 0.0187292
R17536 VPWR.n584 VPWR 0.0187292
R17537 VPWR.n4768 VPWR.n318 0.0187292
R17538 VPWR.n4838 VPWR.n4836 0.0187292
R17539 VPWR.n1087 VPWR.n1086 0.0187292
R17540 VPWR.n1113 VPWR.n1112 0.0187292
R17541 VPWR.n4596 VPWR.n4595 0.0187292
R17542 VPWR.n4692 VPWR.n4690 0.0187292
R17543 VPWR.n4722 VPWR.n4720 0.0187292
R17544 VPWR.n1401 VPWR.n1400 0.0187292
R17545 VPWR.n3793 VPWR.n3792 0.0187292
R17546 VPWR.n3926 VPWR.n3925 0.0187292
R17547 VPWR.n1511 VPWR.n1510 0.0187292
R17548 VPWR.n1519 VPWR 0.0187292
R17549 VPWR.n4063 VPWR.n4062 0.0187292
R17550 VPWR.n2097 VPWR.n2096 0.0187292
R17551 VPWR.n3568 VPWR.n3567 0.0187292
R17552 VPWR.n3685 VPWR.n3684 0.0187292
R17553 VPWR.n2994 VPWR.n2792 0.0187292
R17554 VPWR.n2836 VPWR.n2835 0.0187292
R17555 VPWR.n3467 VPWR.n3466 0.0187292
R17556 VPWR.n2359 VPWR.n2358 0.0187292
R17557 VPWR.n6546 VPWR.n6545 0.0187292
R17558 VPWR.n7743 VPWR.n7742 0.0187292
R17559 VPWR.n29 VPWR 0.0187292
R17560 VPWR.n83 VPWR.n82 0.0187292
R17561 VPWR.n3095 VPWR.n3094 0.0187292
R17562 VPWR.n3185 VPWR.n3184 0.0187292
R17563 VPWR VPWR.n2386 0.0187292
R17564 VPWR.n3333 VPWR.n3332 0.0187292
R17565 VPWR.n6197 VPWR.n6196 0.0187292
R17566 VPWR.n6093 VPWR.n6092 0.0187292
R17567 VPWR VPWR.n7808 0.0187292
R17568 VPWR.n5989 VPWR.n5987 0.0187292
R17569 VPWR VPWR.n5959 0.0185211
R17570 VPWR VPWR.n204 0.0185211
R17571 VPWR.n7473 VPWR 0.0185211
R17572 VPWR.n7363 VPWR 0.0185211
R17573 VPWR.n4832 VPWR 0.0185211
R17574 VPWR.n5125 VPWR.n5124 0.0174271
R17575 VPWR.n5128 VPWR.n5127 0.0174271
R17576 VPWR.n230 VPWR.n227 0.0174271
R17577 VPWR.n5619 VPWR.n5617 0.0174271
R17578 VPWR.n5615 VPWR.n5612 0.0174271
R17579 VPWR VPWR.n279 0.0174271
R17580 VPWR.n7483 VPWR.n7482 0.0174271
R17581 VPWR.n5389 VPWR.n5388 0.0174271
R17582 VPWR.n5398 VPWR 0.0174271
R17583 VPWR.n7373 VPWR.n7372 0.0174271
R17584 VPWR.n521 VPWR.n520 0.0174271
R17585 VPWR.n526 VPWR.n525 0.0174271
R17586 VPWR VPWR.n324 0.0174271
R17587 VPWR.n4842 VPWR.n4841 0.0174271
R17588 VPWR.n1058 VPWR.n1056 0.0174271
R17589 VPWR.n1062 VPWR.n1061 0.0174271
R17590 VPWR.n4688 VPWR 0.0174271
R17591 VPWR.n4717 VPWR.n4715 0.0174271
R17592 VPWR.n1275 VPWR.n1274 0.0174271
R17593 VPWR.n1272 VPWR.n1269 0.0174271
R17594 VPWR.n1406 VPWR 0.0174271
R17595 VPWR.n3929 VPWR.n3928 0.0174271
R17596 VPWR.n1895 VPWR.n1894 0.0174271
R17597 VPWR.n1892 VPWR 0.0174271
R17598 VPWR.n2027 VPWR 0.0174271
R17599 VPWR.n4248 VPWR 0.0174271
R17600 VPWR.n4060 VPWR 0.0174271
R17601 VPWR.n4043 VPWR.n4042 0.0174271
R17602 VPWR.n1720 VPWR.n1719 0.0174271
R17603 VPWR.n2103 VPWR 0.0174271
R17604 VPWR.n3690 VPWR.n3689 0.0174271
R17605 VPWR.n2747 VPWR.n2746 0.0174271
R17606 VPWR.n2752 VPWR.n2751 0.0174271
R17607 VPWR.n2356 VPWR.n2355 0.0174271
R17608 VPWR.n6444 VPWR.n6443 0.0174271
R17609 VPWR.n6441 VPWR.n6440 0.0174271
R17610 VPWR.n7725 VPWR 0.0174271
R17611 VPWR.n88 VPWR.n87 0.0174271
R17612 VPWR.n2618 VPWR.n2616 0.0174271
R17613 VPWR.n2622 VPWR.n2621 0.0174271
R17614 VPWR.n3338 VPWR.n3337 0.0174271
R17615 VPWR.n6321 VPWR.n6319 0.0174271
R17616 VPWR.n6325 VPWR.n6324 0.0174271
R17617 VPWR.n5985 VPWR.n5982 0.0174271
R17618 VPWR.n5478 VPWR.n5475 0.0173937
R17619 VPWR.n7036 VPWR.n7035 0.0173937
R17620 VPWR.n2671 VPWR.n2670 0.0173919
R17621 VPWR.n7754 VPWR.n7753 0.0173919
R17622 VPWR.n247 VPWR.n246 0.0173919
R17623 VPWR.n7629 VPWR.n7628 0.0173919
R17624 VPWR.n5082 VPWR.n5081 0.0173919
R17625 VPWR.n6578 VPWR.n6577 0.0173919
R17626 VPWR.n7490 VPWR.n7489 0.0173919
R17627 VPWR.n6888 VPWR.n6887 0.0173919
R17628 VPWR.n5636 VPWR.n5635 0.0173919
R17629 VPWR.n4896 VPWR.n4895 0.0173919
R17630 VPWR.n7390 VPWR.n7389 0.0173919
R17631 VPWR.n7176 VPWR.n7175 0.0173919
R17632 VPWR.n5404 VPWR.n5215 0.0173919
R17633 VPWR.n7048 VPWR.n7047 0.0173919
R17634 VPWR.n4849 VPWR.n4848 0.0173919
R17635 VPWR.n852 VPWR.n851 0.0173919
R17636 VPWR.n553 VPWR.n552 0.0173919
R17637 VPWR.n636 VPWR.n635 0.0173919
R17638 VPWR.n4749 VPWR.n4748 0.0173919
R17639 VPWR.n4588 VPWR.n4587 0.0173919
R17640 VPWR.n989 VPWR.n988 0.0173919
R17641 VPWR.n409 VPWR.n408 0.0173919
R17642 VPWR.n3757 VPWR.n3756 0.0173919
R17643 VPWR.n3782 VPWR.n1447 0.0173919
R17644 VPWR.n455 VPWR.n454 0.0173919
R17645 VPWR.n4408 VPWR.n4407 0.0173919
R17646 VPWR.n3981 VPWR.n3980 0.0173919
R17647 VPWR.n4151 VPWR.n4150 0.0173919
R17648 VPWR.n1923 VPWR.n1922 0.0173919
R17649 VPWR.n4258 VPWR.n4257 0.0173919
R17650 VPWR.n1664 VPWR.n1663 0.0173919
R17651 VPWR.n2172 VPWR.n2171 0.0173919
R17652 VPWR.n3727 VPWR.n3726 0.0173919
R17653 VPWR.n2042 VPWR.n2041 0.0173919
R17654 VPWR.n4962 VPWR.n4961 0.0173919
R17655 VPWR.n2340 VPWR.n2339 0.0173919
R17656 VPWR.n2766 VPWR.n2765 0.0173919
R17657 VPWR.n3518 VPWR.n3517 0.0173919
R17658 VPWR.n3008 VPWR.n3007 0.0173919
R17659 VPWR.n3056 VPWR.n3055 0.0173919
R17660 VPWR.n5756 VPWR.n5755 0.0173919
R17661 VPWR.n2401 VPWR.n2400 0.0173919
R17662 VPWR.n6074 VPWR.n6073 0.0173919
R17663 VPWR.n6366 VPWR.n6365 0.0173919
R17664 VPWR.n5703 VPWR.n5702 0.0173919
R17665 VPWR.n3386 VPWR.n3385 0.0173919
R17666 VPWR.n5998 VPWR.n5997 0.0173919
R17667 VPWR.n4241 VPWR.n4240 0.0172664
R17668 VPWR.n2843 VPWR.n2842 0.0172664
R17669 VPWR.n3705 VPWR.n3704 0.0172634
R17670 VPWR.n103 VPWR.n102 0.0172634
R17671 VPWR VPWR.n517 0.017219
R17672 VPWR.n7300 VPWR.n7299 0.017135
R17673 VPWR.n4064 VPWR.n1539 0.017135
R17674 VPWR.n7775 VPWR.n7774 0.0169468
R17675 VPWR.n7774 VPWR.n7772 0.0169468
R17676 VPWR.n1814 VPWR.n1813 0.0169447
R17677 VPWR.n1815 VPWR.n1814 0.0169447
R17678 VPWR.n569 VPWR.n568 0.0169447
R17679 VPWR.n570 VPWR.n569 0.0169447
R17680 VPWR.n7659 VPWR.n7658 0.0168788
R17681 VPWR.n112 VPWR.n108 0.0168788
R17682 VPWR.n7516 VPWR.n7515 0.0168788
R17683 VPWR.n238 VPWR.n166 0.0168788
R17684 VPWR.n6766 VPWR.n4935 0.0168788
R17685 VPWR.n7611 VPWR.n7609 0.0168788
R17686 VPWR.n5120 VPWR.n5119 0.0168788
R17687 VPWR.n5659 VPWR.n5210 0.0168788
R17688 VPWR.n6599 VPWR.n6591 0.0168788
R17689 VPWR.n6603 VPWR.n6587 0.0168788
R17690 VPWR.n7400 VPWR.n7399 0.0168788
R17691 VPWR.n7434 VPWR.n7432 0.0168788
R17692 VPWR.n6777 VPWR.n6773 0.0168788
R17693 VPWR.n6875 VPWR.n6781 0.0168788
R17694 VPWR.n5625 VPWR.n5624 0.0168788
R17695 VPWR.n5583 VPWR.n5581 0.0168788
R17696 VPWR.n7006 VPWR.n6998 0.0168788
R17697 VPWR.n6994 VPWR.n4911 0.0168788
R17698 VPWR.n7294 VPWR.n7293 0.0168788
R17699 VPWR.n7324 VPWR.n7322 0.0168788
R17700 VPWR.n7201 VPWR.n4862 0.0168788
R17701 VPWR.n7205 VPWR.n297 0.0168788
R17702 VPWR.n5384 VPWR.n5383 0.0168788
R17703 VPWR.n5228 VPWR.n5224 0.0168788
R17704 VPWR.n5295 VPWR.n5294 0.0168788
R17705 VPWR.n7063 VPWR.n4879 0.0168788
R17706 VPWR.n4759 VPWR.n4758 0.0168788
R17707 VPWR.n4794 VPWR.n4792 0.0168788
R17708 VPWR.n874 VPWR.n600 0.0168788
R17709 VPWR.n878 VPWR.n596 0.0168788
R17710 VPWR.n514 VPWR.n513 0.0168788
R17711 VPWR.n977 VPWR.n463 0.0168788
R17712 VPWR.n623 VPWR.n615 0.0168788
R17713 VPWR.n735 VPWR.n612 0.0168788
R17714 VPWR.n4682 VPWR.n4681 0.0168788
R17715 VPWR.n4726 VPWR.n332 0.0168788
R17716 VPWR.n4555 VPWR.n390 0.0168788
R17717 VPWR.n4568 VPWR.n4559 0.0168788
R17718 VPWR.n1051 VPWR.n1050 0.0168788
R17719 VPWR.n1209 VPWR.n1011 0.0168788
R17720 VPWR.n4432 VPWR.n4424 0.0168788
R17721 VPWR.n4442 VPWR.n4436 0.0168788
R17722 VPWR.n3956 VPWR.n3775 0.0168788
R17723 VPWR.n3771 VPWR.n3765 0.0168788
R17724 VPWR.n4283 VPWR.n4279 0.0168788
R17725 VPWR.n4296 VPWR.n4287 0.0168788
R17726 VPWR.n1281 VPWR.n1280 0.0168788
R17727 VPWR.n1223 VPWR.n1216 0.0168788
R17728 VPWR.n1414 VPWR.n1413 0.0168788
R17729 VPWR.n4391 VPWR.n422 0.0168788
R17730 VPWR.n4054 VPWR.n4053 0.0168788
R17731 VPWR.n4049 VPWR.n3989 0.0168788
R17732 VPWR.n1501 VPWR.n1497 0.0168788
R17733 VPWR.n4131 VPWR.n1505 0.0168788
R17734 VPWR.n1901 VPWR.n1900 0.0168788
R17735 VPWR.n1841 VPWR.n1834 0.0168788
R17736 VPWR.n2034 VPWR.n1638 0.0168788
R17737 VPWR.n1471 VPWR.n1469 0.0168788
R17738 VPWR.n1712 VPWR.n1711 0.0168788
R17739 VPWR.n1809 VPWR.n1805 0.0168788
R17740 VPWR.n3542 VPWR.n3541 0.0168788
R17741 VPWR.n3537 VPWR.n3527 0.0168788
R17742 VPWR.n3714 VPWR.n3713 0.0168788
R17743 VPWR.n1548 VPWR.n1544 0.0168788
R17744 VPWR.n2066 VPWR.n2065 0.0168788
R17745 VPWR.n2072 VPWR.n1636 0.0168788
R17746 VPWR.n4957 VPWR.n4956 0.0168788
R17747 VPWR.n6570 VPWR.n4969 0.0168788
R17748 VPWR.n2470 VPWR.n2461 0.0168788
R17749 VPWR.n3069 VPWR.n2456 0.0168788
R17750 VPWR.n5792 VPWR.n5791 0.0168788
R17751 VPWR.n5818 VPWR.n5763 0.0168788
R17752 VPWR.n3160 VPWR.n3159 0.0168788
R17753 VPWR.n3203 VPWR.n2390 0.0168788
R17754 VPWR.n5 VPWR.n4 0.0168788
R17755 VPWR.n7802 VPWR.n17 0.0168788
R17756 VPWR.n7794 VPWR.n7793 0.0168788
R17757 VPWR.n24 VPWR.n22 0.0168788
R17758 VPWR.n6450 VPWR.n6449 0.0168788
R17759 VPWR.n6455 VPWR.n5072 0.0168788
R17760 VPWR.n5714 VPWR.n5713 0.0168788
R17761 VPWR.n6354 VPWR.n5725 0.0168788
R17762 VPWR.n2498 VPWR.n2497 0.0168788
R17763 VPWR.n2651 VPWR.n2501 0.0168788
R17764 VPWR.n3370 VPWR.n2382 0.0168788
R17765 VPWR.n2376 VPWR.n2372 0.0168788
R17766 VPWR.n6023 VPWR.n6022 0.0168788
R17767 VPWR.n5994 VPWR.n5993 0.0168788
R17768 VPWR.n7299 VPWR.n7298 0.0167522
R17769 VPWR.n4064 VPWR.n4063 0.0167522
R17770 VPWR.n4242 VPWR.n4241 0.0166276
R17771 VPWR.n2842 VPWR.n2841 0.0166276
R17772 VPWR.n3706 VPWR.n3705 0.0166244
R17773 VPWR.n104 VPWR.n103 0.0166244
R17774 VPWR.n5479 VPWR.n5478 0.016499
R17775 VPWR.n7037 VPWR.n7036 0.016499
R17776 VPWR VPWR.n5230 0.016125
R17777 VPWR VPWR.n7023 0.016125
R17778 VPWR.n972 VPWR 0.016125
R17779 VPWR VPWR.n1089 0.016125
R17780 VPWR.n2992 VPWR 0.016125
R17781 VPWR VPWR.n2341 0.016125
R17782 VPWR.n2657 VPWR.n2656 0.0157027
R17783 VPWR.n2504 VPWR.n2503 0.0157027
R17784 VPWR.n2505 VPWR.n2504 0.0157027
R17785 VPWR.n2650 VPWR.n2506 0.0157027
R17786 VPWR.n7660 VPWR.n107 0.0157027
R17787 VPWR.n106 VPWR.n105 0.0157027
R17788 VPWR.n121 VPWR.n120 0.0157027
R17789 VPWR.n123 VPWR.n122 0.0157027
R17790 VPWR.n7789 VPWR.n7788 0.0157027
R17791 VPWR.n7517 VPWR.n165 0.0157027
R17792 VPWR.n164 VPWR.n163 0.0157027
R17793 VPWR.n245 VPWR.n244 0.0157027
R17794 VPWR.n248 VPWR.n247 0.0157027
R17795 VPWR.n6764 VPWR.n4937 0.0157027
R17796 VPWR.n5676 VPWR.n5090 0.0157027
R17797 VPWR.n5205 VPWR.n5204 0.0157027
R17798 VPWR.n5206 VPWR.n5205 0.0157027
R17799 VPWR.n5660 VPWR.n5207 0.0157027
R17800 VPWR.n6584 VPWR.n6583 0.0157027
R17801 VPWR.n7404 VPWR.n7403 0.0157027
R17802 VPWR.n7401 VPWR.n282 0.0157027
R17803 VPWR.n281 VPWR.n280 0.0157027
R17804 VPWR.n274 VPWR.n273 0.0157027
R17805 VPWR.n7491 VPWR.n7490 0.0157027
R17806 VPWR.n6775 VPWR.n6774 0.0157027
R17807 VPWR.n5645 VPWR.n5644 0.0157027
R17808 VPWR.n5576 VPWR.n5575 0.0157027
R17809 VPWR.n5577 VPWR.n5576 0.0157027
R17810 VPWR.n5584 VPWR.n5578 0.0157027
R17811 VPWR.n4915 VPWR.n4914 0.0157027
R17812 VPWR.n7295 VPWR.n7289 0.0157027
R17813 VPWR.n7288 VPWR.n7287 0.0157027
R17814 VPWR.n7387 VPWR.n7386 0.0157027
R17815 VPWR.n7391 VPWR.n7390 0.0157027
R17816 VPWR.n7199 VPWR.n7198 0.0157027
R17817 VPWR.n5413 VPWR.n5412 0.0157027
R17818 VPWR.n5219 VPWR.n5218 0.0157027
R17819 VPWR.n5220 VPWR.n5219 0.0157027
R17820 VPWR.n5229 VPWR.n5221 0.0157027
R17821 VPWR.n5326 VPWR.n5325 0.0157027
R17822 VPWR.n4876 VPWR.n4875 0.0157027
R17823 VPWR.n4763 VPWR.n4762 0.0157027
R17824 VPWR.n4760 VPWR.n327 0.0157027
R17825 VPWR.n326 VPWR.n325 0.0157027
R17826 VPWR.n4777 VPWR.n316 0.0157027
R17827 VPWR.n4850 VPWR.n4849 0.0157027
R17828 VPWR.n872 VPWR.n871 0.0157027
R17829 VPWR.n564 VPWR.n563 0.0157027
R17830 VPWR.n466 VPWR.n465 0.0157027
R17831 VPWR.n467 VPWR.n466 0.0157027
R17832 VPWR.n976 VPWR.n468 0.0157027
R17833 VPWR.n970 VPWR.n469 0.0157027
R17834 VPWR.n609 VPWR.n608 0.0157027
R17835 VPWR.n4686 VPWR.n4685 0.0157027
R17836 VPWR.n4683 VPWR.n4679 0.0157027
R17837 VPWR.n4678 VPWR.n4677 0.0157027
R17838 VPWR.n4746 VPWR.n4745 0.0157027
R17839 VPWR.n4750 VPWR.n4749 0.0157027
R17840 VPWR.n4553 VPWR.n4552 0.0157027
R17841 VPWR.n998 VPWR.n997 0.0157027
R17842 VPWR.n1014 VPWR.n1013 0.0157027
R17843 VPWR.n1015 VPWR.n1014 0.0157027
R17844 VPWR.n1208 VPWR.n1016 0.0157027
R17845 VPWR.n1206 VPWR.n1205 0.0157027
R17846 VPWR.n4440 VPWR.n4439 0.0157027
R17847 VPWR.n3955 VPWR.n3954 0.0157027
R17848 VPWR.n3953 VPWR.n3952 0.0157027
R17849 VPWR.n3754 VPWR.n3753 0.0157027
R17850 VPWR.n3758 VPWR.n3757 0.0157027
R17851 VPWR.n4281 VPWR.n4280 0.0157027
R17852 VPWR.n1295 VPWR.n1294 0.0157027
R17853 VPWR.n1219 VPWR.n1218 0.0157027
R17854 VPWR.n1220 VPWR.n1219 0.0157027
R17855 VPWR.n1222 VPWR.n1221 0.0157027
R17856 VPWR.n426 VPWR.n425 0.0157027
R17857 VPWR.n4058 VPWR.n4057 0.0157027
R17858 VPWR.n4055 VPWR.n1542 0.0157027
R17859 VPWR.n1541 VPWR.n1540 0.0157027
R17860 VPWR.n3978 VPWR.n3977 0.0157027
R17861 VPWR.n3982 VPWR.n3981 0.0157027
R17862 VPWR.n1499 VPWR.n1498 0.0157027
R17863 VPWR.n1909 VPWR.n1908 0.0157027
R17864 VPWR.n1837 VPWR.n1836 0.0157027
R17865 VPWR.n1838 VPWR.n1837 0.0157027
R17866 VPWR.n1840 VPWR.n1839 0.0157027
R17867 VPWR.n1466 VPWR.n1465 0.0157027
R17868 VPWR.n1820 VPWR.n1672 0.0157027
R17869 VPWR.n1800 VPWR.n1799 0.0157027
R17870 VPWR.n1801 VPWR.n1800 0.0157027
R17871 VPWR.n1810 VPWR.n1802 0.0157027
R17872 VPWR.n2158 VPWR.n2157 0.0157027
R17873 VPWR.n3712 VPWR.n3711 0.0157027
R17874 VPWR.n3710 VPWR.n3709 0.0157027
R17875 VPWR.n3725 VPWR.n3724 0.0157027
R17876 VPWR.n3728 VPWR.n3727 0.0157027
R17877 VPWR.n1633 VPWR.n1632 0.0157027
R17878 VPWR.n4975 VPWR.n4974 0.0157027
R17879 VPWR.n2277 VPWR.n2276 0.0157027
R17880 VPWR.n2272 VPWR.n2271 0.0157027
R17881 VPWR.n3413 VPWR.n3412 0.0157027
R17882 VPWR.n2339 VPWR.n2338 0.0157027
R17883 VPWR.n2767 VPWR.n2766 0.0157027
R17884 VPWR.n2780 VPWR.n2779 0.0157027
R17885 VPWR.n2777 VPWR.n2776 0.0157027
R17886 VPWR.n2996 VPWR.n2688 0.0157027
R17887 VPWR.n2990 VPWR.n2689 0.0157027
R17888 VPWR.n3490 VPWR.n3489 0.0157027
R17889 VPWR.n2809 VPWR.n2808 0.0157027
R17890 VPWR.n2455 VPWR.n2454 0.0157027
R17891 VPWR.n5753 VPWR.n5752 0.0157027
R17892 VPWR.n3155 VPWR.n3154 0.0157027
R17893 VPWR.n6082 VPWR.n6081 0.0157027
R17894 VPWR.n6426 VPWR.n6425 0.0157027
R17895 VPWR.n5069 VPWR.n5068 0.0157027
R17896 VPWR.n5070 VPWR.n5069 0.0157027
R17897 VPWR.n6456 VPWR.n5071 0.0157027
R17898 VPWR.n5720 VPWR.n5719 0.0157027
R17899 VPWR.n5729 VPWR.n5728 0.0157027
R17900 VPWR.n5730 VPWR.n5729 0.0157027
R17901 VPWR.n6353 VPWR.n5731 0.0157027
R17902 VPWR.n3369 VPWR.n3368 0.0157027
R17903 VPWR.n3367 VPWR.n3366 0.0157027
R17904 VPWR.n3366 VPWR.n3365 0.0157027
R17905 VPWR.n3375 VPWR.n3374 0.0157027
R17906 VPWR.n6024 VPWR.n5908 0.0157027
R17907 VPWR.n6012 VPWR.n6011 0.0157027
R17908 VPWR.n6015 VPWR.n6014 0.0157027
R17909 VPWR.n2077 VPWR.n2075 0.0153255
R17910 VPWR.n2852 VPWR.n2851 0.0153255
R17911 VPWR.n6567 VPWR.n6566 0.0153255
R17912 VPWR.n6177 VPWR.n6174 0.0153255
R17913 VPWR.n6991 VPWR.n4916 0.0150286
R17914 VPWR.n4462 VPWR.n4461 0.0150286
R17915 VPWR.n4388 VPWR.n428 0.0150286
R17916 VPWR.n4233 VPWR.n4232 0.0150286
R17917 VPWR.n3075 VPWR.n3072 0.0150286
R17918 VPWR.n5129 VPWR.n5128 0.0148229
R17919 VPWR.n6610 VPWR.n6609 0.0148229
R17920 VPWR.n6664 VPWR.n6663 0.0148229
R17921 VPWR.n6760 VPWR.n6759 0.0148229
R17922 VPWR.n227 VPWR.n226 0.0148229
R17923 VPWR.n5612 VPWR.n5611 0.0148229
R17924 VPWR.n5474 VPWR.n5473 0.0148229
R17925 VPWR.n6913 VPWR.n6912 0.0148229
R17926 VPWR VPWR.n6792 0.0148229
R17927 VPWR.n7484 VPWR.n7483 0.0148229
R17928 VPWR VPWR.n5393 0.0148229
R17929 VPWR.n7034 VPWR.n7033 0.0148229
R17930 VPWR.n7186 VPWR.n7185 0.0148229
R17931 VPWR.n7313 VPWR 0.0148229
R17932 VPWR.n7374 VPWR.n7373 0.0148229
R17933 VPWR.n527 VPWR.n526 0.0148229
R17934 VPWR.n716 VPWR.n715 0.0148229
R17935 VPWR.n721 VPWR.n720 0.0148229
R17936 VPWR.n862 VPWR.n861 0.0148229
R17937 VPWR.n4843 VPWR.n4842 0.0148229
R17938 VPWR.n4836 VPWR 0.0148229
R17939 VPWR.n1063 VPWR.n1062 0.0148229
R17940 VPWR.n4458 VPWR.n402 0.0148229
R17941 VPWR.n4457 VPWR.n406 0.0148229
R17942 VPWR.n4542 VPWR.n4541 0.0148229
R17943 VPWR.n4715 VPWR.n4714 0.0148229
R17944 VPWR.n1269 VPWR.n1268 0.0148229
R17945 VPWR.n1391 VPWR.n1389 0.0148229
R17946 VPWR.n1387 VPWR.n1386 0.0148229
R17947 VPWR.n4318 VPWR.n4317 0.0148229
R17948 VPWR.n3930 VPWR.n3929 0.0148229
R17949 VPWR VPWR.n1885 0.0148229
R17950 VPWR.n4239 VPWR.n4238 0.0148229
R17951 VPWR.n4166 VPWR.n4165 0.0148229
R17952 VPWR.n4042 VPWR.n4041 0.0148229
R17953 VPWR.n1721 VPWR.n1720 0.0148229
R17954 VPWR.n2087 VPWR.n2085 0.0148229
R17955 VPWR.n2083 VPWR.n2082 0.0148229
R17956 VPWR.n3554 VPWR.n3553 0.0148229
R17957 VPWR.n3691 VPWR.n3690 0.0148229
R17958 VPWR.n2753 VPWR.n2752 0.0148229
R17959 VPWR.n2845 VPWR.n2844 0.0148229
R17960 VPWR.n3481 VPWR.n3480 0.0148229
R17961 VPWR.n2355 VPWR.n2354 0.0148229
R17962 VPWR.n6440 VPWR.n6439 0.0148229
R17963 VPWR.n6558 VPWR.n6556 0.0148229
R17964 VPWR.n6560 VPWR.n6559 0.0148229
R17965 VPWR.n7777 VPWR.n7776 0.0148229
R17966 VPWR.n89 VPWR.n88 0.0148229
R17967 VPWR.n2623 VPWR.n2622 0.0148229
R17968 VPWR.n3085 VPWR.n3083 0.0148229
R17969 VPWR.n3081 VPWR.n3080 0.0148229
R17970 VPWR.n3175 VPWR.n3174 0.0148229
R17971 VPWR.n3339 VPWR.n3338 0.0148229
R17972 VPWR.n6326 VPWR.n6325 0.0148229
R17973 VPWR.n6187 VPWR.n6185 0.0148229
R17974 VPWR.n6183 VPWR.n6182 0.0148229
R17975 VPWR.n6103 VPWR.n6102 0.0148229
R17976 VPWR.n5982 VPWR.n5981 0.0148229
R17977 VPWR.n7640 VPWR.n7639 0.0145155
R17978 VPWR.n252 VPWR.n251 0.0145155
R17979 VPWR.n145 VPWR.n144 0.0145155
R17980 VPWR.n144 VPWR.n143 0.0145155
R17981 VPWR.n5682 VPWR.n5681 0.0145155
R17982 VPWR.n5681 VPWR.n5680 0.0145155
R17983 VPWR.n6672 VPWR.n6671 0.0145155
R17984 VPWR.n6671 VPWR.n6670 0.0145155
R17985 VPWR.n269 VPWR.n268 0.0145155
R17986 VPWR.n268 VPWR.n267 0.0145155
R17987 VPWR.n6893 VPWR.n6892 0.0145155
R17988 VPWR.n6894 VPWR.n6893 0.0145155
R17989 VPWR.n5651 VPWR.n5650 0.0145155
R17990 VPWR.n5650 VPWR.n5649 0.0145155
R17991 VPWR.n4905 VPWR.n4904 0.0145155
R17992 VPWR.n4904 VPWR.n4903 0.0145155
R17993 VPWR.n7382 VPWR.n7381 0.0145155
R17994 VPWR.n7381 VPWR.n7380 0.0145155
R17995 VPWR.n7171 VPWR.n7170 0.0145155
R17996 VPWR.n7170 VPWR.n7169 0.0145155
R17997 VPWR.n5419 VPWR.n5418 0.0145155
R17998 VPWR.n5418 VPWR.n5417 0.0145155
R17999 VPWR.n7057 VPWR.n7056 0.0145155
R18000 VPWR.n7056 VPWR.n7055 0.0145155
R18001 VPWR.n314 VPWR.n313 0.0145155
R18002 VPWR.n313 VPWR.n312 0.0145155
R18003 VPWR.n847 VPWR.n846 0.0145155
R18004 VPWR.n846 VPWR.n845 0.0145155
R18005 VPWR.n545 VPWR.n544 0.0145155
R18006 VPWR.n544 VPWR.n543 0.0145155
R18007 VPWR.n729 VPWR.n728 0.0145155
R18008 VPWR.n728 VPWR.n727 0.0145155
R18009 VPWR.n4741 VPWR.n4740 0.0145155
R18010 VPWR.n4740 VPWR.n4739 0.0145155
R18011 VPWR.n4583 VPWR.n4582 0.0145155
R18012 VPWR.n4582 VPWR.n4581 0.0145155
R18013 VPWR.n1004 VPWR.n1003 0.0145155
R18014 VPWR.n1003 VPWR.n1002 0.0145155
R18015 VPWR.n4449 VPWR.n4448 0.0145155
R18016 VPWR.n4450 VPWR.n4449 0.0145155
R18017 VPWR.n3749 VPWR.n3748 0.0145155
R18018 VPWR.n3748 VPWR.n3747 0.0145155
R18019 VPWR.n4311 VPWR.n4310 0.0145155
R18020 VPWR.n4310 VPWR.n4309 0.0145155
R18021 VPWR.n1288 VPWR.n1287 0.0145155
R18022 VPWR.n1289 VPWR.n1288 0.0145155
R18023 VPWR.n4417 VPWR.n4416 0.0145155
R18024 VPWR.n4416 VPWR.n4415 0.0145155
R18025 VPWR.n3973 VPWR.n3972 0.0145155
R18026 VPWR.n3972 VPWR.n3971 0.0145155
R18027 VPWR.n4146 VPWR.n4145 0.0145155
R18028 VPWR.n4145 VPWR.n4144 0.0145155
R18029 VPWR.n1915 VPWR.n1914 0.0145155
R18030 VPWR.n1914 VPWR.n1913 0.0145155
R18031 VPWR.n4267 VPWR.n4266 0.0145155
R18032 VPWR.n4266 VPWR.n4265 0.0145155
R18033 VPWR.n1826 VPWR.n1825 0.0145155
R18034 VPWR.n1825 VPWR.n1824 0.0145155
R18035 VPWR.n2185 VPWR.n2184 0.0145155
R18036 VPWR.n2184 VPWR.n2183 0.0145155
R18037 VPWR.n3720 VPWR.n3719 0.0145155
R18038 VPWR.n2051 VPWR.n2050 0.0145155
R18039 VPWR.n2050 VPWR.n2049 0.0145155
R18040 VPWR.n5800 VPWR.n5799 0.0145155
R18041 VPWR.n5799 VPWR.n5798 0.0145155
R18042 VPWR.n3408 VPWR.n3407 0.0145155
R18043 VPWR.n3407 VPWR.n3406 0.0145155
R18044 VPWR.n2770 VPWR.n2769 0.0145155
R18045 VPWR.n3509 VPWR.n3508 0.0145155
R18046 VPWR.n3004 VPWR.n3003 0.0145155
R18047 VPWR.n3049 VPWR.n3048 0.0145155
R18048 VPWR.n3050 VPWR.n3049 0.0145155
R18049 VPWR.n5770 VPWR.n5769 0.0145155
R18050 VPWR.n5769 VPWR.n5768 0.0145155
R18051 VPWR.n2406 VPWR.n2405 0.0145155
R18052 VPWR.n2407 VPWR.n2406 0.0145155
R18053 VPWR.n11 VPWR.n10 0.0145155
R18054 VPWR.n12 VPWR.n11 0.0145155
R18055 VPWR.n7759 VPWR.n7758 0.0145155
R18056 VPWR.n7760 VPWR.n7759 0.0145155
R18057 VPWR.n6374 VPWR.n6373 0.0145155
R18058 VPWR.n6373 VPWR.n6372 0.0145155
R18059 VPWR.n5695 VPWR.n5694 0.0145155
R18060 VPWR.n5694 VPWR.n5693 0.0145155
R18061 VPWR.n2663 VPWR.n2662 0.0145155
R18062 VPWR.n2662 VPWR.n2661 0.0145155
R18063 VPWR.n3382 VPWR.n3381 0.0145155
R18064 VPWR.n3383 VPWR.n3382 0.0145155
R18065 VPWR.n6009 VPWR.n6008 0.0145155
R18066 VPWR.n6008 VPWR.n6007 0.0145155
R18067 VPWR.n2675 VPWR.n2674 0.0140135
R18068 VPWR.n2658 VPWR.n2655 0.0140135
R18069 VPWR.n125 VPWR.n124 0.0140135
R18070 VPWR.n7651 VPWR.n7645 0.0140135
R18071 VPWR.n7787 VPWR.n7786 0.0140135
R18072 VPWR.n7751 VPWR.n7750 0.0140135
R18073 VPWR.n7755 VPWR.n7754 0.0140135
R18074 VPWR.n250 VPWR.n249 0.0140135
R18075 VPWR.n7508 VPWR.n7502 0.0140135
R18076 VPWR.n148 VPWR.n147 0.0140135
R18077 VPWR.n151 VPWR.n150 0.0140135
R18078 VPWR.n7630 VPWR.n7629 0.0140135
R18079 VPWR.n5086 VPWR.n5085 0.0140135
R18080 VPWR.n5677 VPWR.n5088 0.0140135
R18081 VPWR.n6667 VPWR.n6578 0.0140135
R18082 VPWR.n6666 VPWR.n6665 0.0140135
R18083 VPWR.n6582 VPWR.n6581 0.0140135
R18084 VPWR.n7493 VPWR.n7492 0.0140135
R18085 VPWR.n264 VPWR.n260 0.0140135
R18086 VPWR.n6880 VPWR.n6879 0.0140135
R18087 VPWR.n6883 VPWR.n6882 0.0140135
R18088 VPWR.n6889 VPWR.n6888 0.0140135
R18089 VPWR.n5640 VPWR.n5639 0.0140135
R18090 VPWR.n5646 VPWR.n5642 0.0140135
R18091 VPWR.n4900 VPWR.n4896 0.0140135
R18092 VPWR.n4899 VPWR.n4898 0.0140135
R18093 VPWR.n4913 VPWR.n4912 0.0140135
R18094 VPWR.n7393 VPWR.n7392 0.0140135
R18095 VPWR.n7377 VPWR.n287 0.0140135
R18096 VPWR.n7142 VPWR.n7141 0.0140135
R18097 VPWR.n7145 VPWR.n7144 0.0140135
R18098 VPWR.n7175 VPWR.n7174 0.0140135
R18099 VPWR.n5408 VPWR.n5407 0.0140135
R18100 VPWR.n5414 VPWR.n5410 0.0140135
R18101 VPWR.n7052 VPWR.n7048 0.0140135
R18102 VPWR.n7051 VPWR.n7050 0.0140135
R18103 VPWR.n4874 VPWR.n4873 0.0140135
R18104 VPWR.n4852 VPWR.n4851 0.0140135
R18105 VPWR.n309 VPWR.n305 0.0140135
R18106 VPWR.n825 VPWR.n824 0.0140135
R18107 VPWR.n828 VPWR.n827 0.0140135
R18108 VPWR.n851 VPWR.n850 0.0140135
R18109 VPWR.n549 VPWR.n548 0.0140135
R18110 VPWR.n474 VPWR.n473 0.0140135
R18111 VPWR.n724 VPWR.n636 0.0140135
R18112 VPWR.n723 VPWR.n722 0.0140135
R18113 VPWR.n607 VPWR.n606 0.0140135
R18114 VPWR.n4752 VPWR.n4751 0.0140135
R18115 VPWR.n4736 VPWR.n4732 0.0140135
R18116 VPWR.n381 VPWR.n380 0.0140135
R18117 VPWR.n384 VPWR.n383 0.0140135
R18118 VPWR.n4587 VPWR.n4586 0.0140135
R18119 VPWR.n993 VPWR.n992 0.0140135
R18120 VPWR.n999 VPWR.n995 0.0140135
R18121 VPWR.n4453 VPWR.n409 0.0140135
R18122 VPWR.n4456 VPWR.n4454 0.0140135
R18123 VPWR.n4438 VPWR.n4437 0.0140135
R18124 VPWR.n3760 VPWR.n3759 0.0140135
R18125 VPWR.n3744 VPWR.n3740 0.0140135
R18126 VPWR.n1445 VPWR.n1444 0.0140135
R18127 VPWR.n4316 VPWR.n4315 0.0140135
R18128 VPWR.n4314 VPWR.n1447 0.0140135
R18129 VPWR.n459 VPWR.n458 0.0140135
R18130 VPWR.n1292 VPWR.n446 0.0140135
R18131 VPWR.n4412 VPWR.n4408 0.0140135
R18132 VPWR.n4411 VPWR.n4410 0.0140135
R18133 VPWR.n424 VPWR.n423 0.0140135
R18134 VPWR.n3984 VPWR.n3983 0.0140135
R18135 VPWR.n3968 VPWR.n3964 0.0140135
R18136 VPWR.n1490 VPWR.n1489 0.0140135
R18137 VPWR.n1493 VPWR.n1492 0.0140135
R18138 VPWR.n4150 VPWR.n4149 0.0140135
R18139 VPWR.n1919 VPWR.n1918 0.0140135
R18140 VPWR.n1910 VPWR.n1906 0.0140135
R18141 VPWR.n4262 VPWR.n4258 0.0140135
R18142 VPWR.n4261 VPWR.n4260 0.0140135
R18143 VPWR.n1464 VPWR.n1463 0.0140135
R18144 VPWR.n1668 VPWR.n1667 0.0140135
R18145 VPWR.n1821 VPWR.n1670 0.0140135
R18146 VPWR.n2164 VPWR.n2163 0.0140135
R18147 VPWR.n2167 VPWR.n2166 0.0140135
R18148 VPWR.n2173 VPWR.n2172 0.0140135
R18149 VPWR.n3730 VPWR.n3729 0.0140135
R18150 VPWR.n1563 VPWR.n1557 0.0140135
R18151 VPWR.n2046 VPWR.n2042 0.0140135
R18152 VPWR.n2045 VPWR.n2044 0.0140135
R18153 VPWR.n1631 VPWR.n1630 0.0140135
R18154 VPWR.n4965 VPWR.n4962 0.0140135
R18155 VPWR.n4964 VPWR.n4963 0.0140135
R18156 VPWR.n4973 VPWR.n4972 0.0140135
R18157 VPWR.n3411 VPWR.n2273 0.0140135
R18158 VPWR.n2350 VPWR.n2349 0.0140135
R18159 VPWR.n2736 VPWR.n2735 0.0140135
R18160 VPWR.n2775 VPWR.n2768 0.0140135
R18161 VPWR.n3512 VPWR.n3511 0.0140135
R18162 VPWR.n3515 VPWR.n3514 0.0140135
R18163 VPWR.n3519 VPWR.n3518 0.0140135
R18164 VPWR.n3014 VPWR.n3008 0.0140135
R18165 VPWR.n3013 VPWR.n3012 0.0140135
R18166 VPWR.n3010 VPWR.n3009 0.0140135
R18167 VPWR.n3062 VPWR.n3056 0.0140135
R18168 VPWR.n3061 VPWR.n3060 0.0140135
R18169 VPWR.n3058 VPWR.n3057 0.0140135
R18170 VPWR.n5759 VPWR.n5756 0.0140135
R18171 VPWR.n5758 VPWR.n5757 0.0140135
R18172 VPWR.n5751 VPWR.n5750 0.0140135
R18173 VPWR.n3153 VPWR.n3152 0.0140135
R18174 VPWR.n2398 VPWR.n2397 0.0140135
R18175 VPWR.n2402 VPWR.n2401 0.0140135
R18176 VPWR.n6080 VPWR.n6079 0.0140135
R18177 VPWR.n6077 VPWR.n6076 0.0140135
R18178 VPWR.n6075 VPWR.n6074 0.0140135
R18179 VPWR.n6370 VPWR.n6369 0.0140135
R18180 VPWR.n6424 VPWR.n6420 0.0140135
R18181 VPWR.n5707 VPWR.n5706 0.0140135
R18182 VPWR.n5721 VPWR.n5718 0.0140135
R18183 VPWR.n3378 VPWR.n3377 0.0140135
R18184 VPWR.n3395 VPWR.n3389 0.0140135
R18185 VPWR.n6018 VPWR.n6017 0.0140135
R18186 VPWR.n6004 VPWR.n6001 0.0140135
R18187 VPWR.n6919 VPWR.n6918 0.0139925
R18188 VPWR.n7196 VPWR.n7195 0.0139925
R18189 VPWR.n869 VPWR.n868 0.0139925
R18190 VPWR.n4550 VPWR.n4549 0.0139925
R18191 VPWR.n4325 VPWR.n4324 0.0139925
R18192 VPWR.n4172 VPWR.n4171 0.0139925
R18193 VPWR.n3169 VPWR.n3163 0.0139925
R18194 VPWR.n6749 VPWR.n6747 0.0139925
R18195 VPWR.n3548 VPWR.n3545 0.0139925
R18196 VPWR.n3487 VPWR.n3486 0.0139925
R18197 VPWR.n7783 VPWR.n7782 0.0139925
R18198 VPWR.n6108 VPWR.n6085 0.0139925
R18199 VPWR.n5136 VPWR.n5133 0.0135208
R18200 VPWR.n6608 VPWR.n6607 0.0135208
R18201 VPWR.n6758 VPWR.n6756 0.0135208
R18202 VPWR.n6754 VPWR.n6752 0.0135208
R18203 VPWR.n7618 VPWR 0.0135208
R18204 VPWR.n222 VPWR.n221 0.0135208
R18205 VPWR.n5607 VPWR.n5606 0.0135208
R18206 VPWR.n6911 VPWR.n6909 0.0135208
R18207 VPWR.n7488 VPWR.n7426 0.0135208
R18208 VPWR.n5403 VPWR.n5402 0.0135208
R18209 VPWR.n7184 VPWR.n7183 0.0135208
R18210 VPWR.n7182 VPWR.n7181 0.0135208
R18211 VPWR.n7161 VPWR 0.0135208
R18212 VPWR.n7312 VPWR.n7311 0.0135208
R18213 VPWR.n7367 VPWR 0.0135208
R18214 VPWR.n557 VPWR.n554 0.0135208
R18215 VPWR VPWR.n570 0.0135208
R18216 VPWR.n714 VPWR.n713 0.0135208
R18217 VPWR.n4847 VPWR.n4786 0.0135208
R18218 VPWR.n1070 VPWR.n1067 0.0135208
R18219 VPWR.n1102 VPWR.n1100 0.0135208
R18220 VPWR.n4540 VPWR.n4538 0.0135208
R18221 VPWR.n4536 VPWR.n4534 0.0135208
R18222 VPWR.n4710 VPWR.n4709 0.0135208
R18223 VPWR.n1264 VPWR.n1263 0.0135208
R18224 VPWR.n1395 VPWR.n1393 0.0135208
R18225 VPWR.n1443 VPWR.n1441 0.0135208
R18226 VPWR.n3937 VPWR.n3934 0.0135208
R18227 VPWR.n1926 VPWR.n1924 0.0135208
R18228 VPWR.n4164 VPWR.n4162 0.0135208
R18229 VPWR.n4160 VPWR.n4158 0.0135208
R18230 VPWR.n4037 VPWR.n4036 0.0135208
R18231 VPWR.n1726 VPWR.n1725 0.0135208
R18232 VPWR.n2109 VPWR 0.0135208
R18233 VPWR.n2091 VPWR.n2089 0.0135208
R18234 VPWR.n3558 VPWR.n3556 0.0135208
R18235 VPWR.n3562 VPWR.n3560 0.0135208
R18236 VPWR.n3696 VPWR.n3695 0.0135208
R18237 VPWR.n2760 VPWR.n2757 0.0135208
R18238 VPWR.n3479 VPWR.n3477 0.0135208
R18239 VPWR.n3475 VPWR.n3473 0.0135208
R18240 VPWR.n2341 VPWR.n2337 0.0135208
R18241 VPWR.n6435 VPWR.n6434 0.0135208
R18242 VPWR.n6554 VPWR.n6552 0.0135208
R18243 VPWR.n94 VPWR.n93 0.0135208
R18244 VPWR.n2630 VPWR.n2627 0.0135208
R18245 VPWR.n3089 VPWR.n3087 0.0135208
R18246 VPWR.n3177 VPWR.n3176 0.0135208
R18247 VPWR.n3179 VPWR.n3178 0.0135208
R18248 VPWR VPWR.n3189 0.0135208
R18249 VPWR.n3346 VPWR.n3343 0.0135208
R18250 VPWR.n6333 VPWR.n6330 0.0135208
R18251 VPWR.n6191 VPWR.n6189 0.0135208
R18252 VPWR.n6101 VPWR.n6100 0.0135208
R18253 VPWR.n6099 VPWR.n6098 0.0135208
R18254 VPWR.n6087 VPWR 0.0135208
R18255 VPWR.n5977 VPWR.n5976 0.0135208
R18256 VPWR.n7609 VPWR.n7608 0.0130912
R18257 VPWR.n5210 VPWR.n5209 0.0130912
R18258 VPWR.n6587 VPWR.n6586 0.0130912
R18259 VPWR.n7432 VPWR.n7431 0.0130912
R18260 VPWR.n6781 VPWR.n6780 0.0130912
R18261 VPWR.n5581 VPWR.n5580 0.0130912
R18262 VPWR.n4911 VPWR.n4910 0.0130912
R18263 VPWR.n7322 VPWR.n7321 0.0130912
R18264 VPWR.n297 VPWR.n296 0.0130912
R18265 VPWR.n5224 VPWR.n5223 0.0130912
R18266 VPWR.n4879 VPWR.n4878 0.0130912
R18267 VPWR.n4792 VPWR.n4791 0.0130912
R18268 VPWR.n596 VPWR.n595 0.0130912
R18269 VPWR.n463 VPWR.n462 0.0130912
R18270 VPWR.n612 VPWR.n611 0.0130912
R18271 VPWR.n332 VPWR.n331 0.0130912
R18272 VPWR.n4559 VPWR.n4558 0.0130912
R18273 VPWR.n1011 VPWR.n1010 0.0130912
R18274 VPWR.n4436 VPWR.n4435 0.0130912
R18275 VPWR.n3765 VPWR.n3764 0.0130912
R18276 VPWR.n4287 VPWR.n4286 0.0130912
R18277 VPWR.n1216 VPWR.n1215 0.0130912
R18278 VPWR.n422 VPWR.n421 0.0130912
R18279 VPWR.n3989 VPWR.n3988 0.0130912
R18280 VPWR.n1505 VPWR.n1504 0.0130912
R18281 VPWR.n1834 VPWR.n1833 0.0130912
R18282 VPWR.n1469 VPWR.n1468 0.0130912
R18283 VPWR.n1805 VPWR.n1804 0.0130912
R18284 VPWR.n3527 VPWR.n3526 0.0130912
R18285 VPWR.n1636 VPWR.n1635 0.0130912
R18286 VPWR.n4969 VPWR.n4968 0.0130912
R18287 VPWR.n2281 VPWR.n2280 0.0130912
R18288 VPWR.n2365 VPWR.n2364 0.0130912
R18289 VPWR.n2740 VPWR.n2739 0.0130912
R18290 VPWR.n3019 VPWR.n3018 0.0130912
R18291 VPWR.n2485 VPWR.n2484 0.0130912
R18292 VPWR.n2461 VPWR.n2460 0.0130912
R18293 VPWR.n5763 VPWR.n5762 0.0130912
R18294 VPWR.n3159 VPWR.n3158 0.0130912
R18295 VPWR.n6 VPWR.n5 0.0130912
R18296 VPWR.n17 VPWR.n16 0.0130912
R18297 VPWR.n7793 VPWR.n7792 0.0130912
R18298 VPWR.n22 VPWR.n21 0.0130912
R18299 VPWR.n6421 VPWR.n5072 0.0130912
R18300 VPWR.n5725 VPWR.n5724 0.0130912
R18301 VPWR.n2497 VPWR.n2496 0.0130912
R18302 VPWR.n2501 VPWR.n2500 0.0130912
R18303 VPWR.n2382 VPWR.n2381 0.0130912
R18304 VPWR.n6022 VPWR.n6021 0.0130912
R18305 VPWR.n5995 VPWR.n5994 0.0130912
R18306 VPWR.n2279 VPWR.n2278 0.0126061
R18307 VPWR.n2742 VPWR.n2741 0.0126061
R18308 VPWR.n2483 VPWR.n2482 0.0126061
R18309 VPWR.n7786 VPWR.n7785 0.0123243
R18310 VPWR.n7766 VPWR.n7765 0.0123243
R18311 VPWR.n7748 VPWR.n7747 0.0123243
R18312 VPWR.n149 VPWR.n148 0.0123243
R18313 VPWR.n136 VPWR.n135 0.0123243
R18314 VPWR.n138 VPWR.n137 0.0123243
R18315 VPWR.n6677 VPWR.n6676 0.0123243
R18316 VPWR.n6881 VPWR.n6880 0.0123243
R18317 VPWR.n6899 VPWR.n6898 0.0123243
R18318 VPWR.n4930 VPWR.n4929 0.0123243
R18319 VPWR.n4892 VPWR.n4891 0.0123243
R18320 VPWR.n7143 VPWR.n7142 0.0123243
R18321 VPWR.n7152 VPWR.n7151 0.0123243
R18322 VPWR.n7154 VPWR.n7153 0.0123243
R18323 VPWR.n7044 VPWR.n7043 0.0123243
R18324 VPWR.n826 VPWR.n825 0.0123243
R18325 VPWR.n834 VPWR.n833 0.0123243
R18326 VPWR.n836 VPWR.n835 0.0123243
R18327 VPWR.n707 VPWR.n706 0.0123243
R18328 VPWR.n382 VPWR.n381 0.0123243
R18329 VPWR.n4574 VPWR.n4573 0.0123243
R18330 VPWR.n4576 VPWR.n4575 0.0123243
R18331 VPWR.n1105 VPWR.n1104 0.0123243
R18332 VPWR.n1446 VPWR.n1445 0.0123243
R18333 VPWR.n4302 VPWR.n4301 0.0123243
R18334 VPWR.n4304 VPWR.n4303 0.0123243
R18335 VPWR.n4404 VPWR.n4403 0.0123243
R18336 VPWR.n1491 VPWR.n1490 0.0123243
R18337 VPWR.n4137 VPWR.n4136 0.0123243
R18338 VPWR.n4139 VPWR.n4138 0.0123243
R18339 VPWR.n4254 VPWR.n4253 0.0123243
R18340 VPWR.n2165 VPWR.n2164 0.0123243
R18341 VPWR.n2176 VPWR.n2175 0.0123243
R18342 VPWR.n2178 VPWR.n2177 0.0123243
R18343 VPWR.n2061 VPWR.n2060 0.0123243
R18344 VPWR.n5810 VPWR.n5809 0.0123243
R18345 VPWR.n4972 VPWR.n4971 0.0123243
R18346 VPWR.n3513 VPWR.n3512 0.0123243
R18347 VPWR.n2197 VPWR.n2196 0.0123243
R18348 VPWR.n2201 VPWR.n2200 0.0123243
R18349 VPWR.n3032 VPWR.n3031 0.0123243
R18350 VPWR.n3011 VPWR.n3010 0.0123243
R18351 VPWR.n3044 VPWR.n3043 0.0123243
R18352 VPWR.n3059 VPWR.n3058 0.0123243
R18353 VPWR.n5780 VPWR.n5779 0.0123243
R18354 VPWR.n5750 VPWR.n5749 0.0123243
R18355 VPWR.n2413 VPWR.n2412 0.0123243
R18356 VPWR.n3194 VPWR.n3193 0.0123243
R18357 VPWR.n6079 VPWR.n6078 0.0123243
R18358 VPWR.n6068 VPWR.n6067 0.0123243
R18359 VPWR.n6064 VPWR.n6063 0.0123243
R18360 VPWR.n5672 VPWR.n5671 0.0122188
R18361 VPWR.n6703 VPWR.n6702 0.0122188
R18362 VPWR.n7601 VPWR.n7600 0.0122188
R18363 VPWR.n211 VPWR.n210 0.0122188
R18364 VPWR.n214 VPWR.n213 0.0122188
R18365 VPWR.n5599 VPWR.n5598 0.0122188
R18366 VPWR.n5596 VPWR.n5595 0.0122188
R18367 VPWR.n5496 VPWR.n5495 0.0122188
R18368 VPWR.n6867 VPWR.n6866 0.0122188
R18369 VPWR.n279 VPWR.n278 0.0122188
R18370 VPWR.n7416 VPWR.n7415 0.0122188
R18371 VPWR.n7419 VPWR.n7418 0.0122188
R18372 VPWR.n5340 VPWR.n5339 0.0122188
R18373 VPWR.n5337 VPWR.n5336 0.0122188
R18374 VPWR.n5330 VPWR 0.0122188
R18375 VPWR.n5230 VPWR.n5217 0.0122188
R18376 VPWR.n5303 VPWR.n5302 0.0122188
R18377 VPWR.n7214 VPWR.n7213 0.0122188
R18378 VPWR.n7301 VPWR.n7300 0.0122188
R18379 VPWR.n7304 VPWR.n7303 0.0122188
R18380 VPWR.n568 VPWR.n567 0.0122188
R18381 VPWR.n973 VPWR.n972 0.0122188
R18382 VPWR.n686 VPWR.n685 0.0122188
R18383 VPWR.n585 VPWR.n584 0.0122188
R18384 VPWR.n324 VPWR.n323 0.0122188
R18385 VPWR.n1076 VPWR.n1075 0.0122188
R18386 VPWR.n1080 VPWR.n1078 0.0122188
R18387 VPWR.n1089 VPWR.n1088 0.0122188
R18388 VPWR.n1128 VPWR.n1126 0.0122188
R18389 VPWR.n4611 VPWR.n4609 0.0122188
R18390 VPWR.n4689 VPWR.n4688 0.0122188
R18391 VPWR.n4699 VPWR.n4698 0.0122188
R18392 VPWR.n4702 VPWR.n4701 0.0122188
R18393 VPWR.n1301 VPWR.n1299 0.0122188
R18394 VPWR.n1423 VPWR.n1422 0.0122188
R18395 VPWR.n3806 VPWR.n3805 0.0122188
R18396 VPWR.n3946 VPWR.n3945 0.0122188
R18397 VPWR.n3943 VPWR.n3942 0.0122188
R18398 VPWR.n1933 VPWR.n1932 0.0122188
R18399 VPWR.n1937 VPWR.n1935 0.0122188
R18400 VPWR.n2018 VPWR.n2017 0.0122188
R18401 VPWR.n4122 VPWR.n4121 0.0122188
R18402 VPWR.n4061 VPWR.n4060 0.0122188
R18403 VPWR.n4029 VPWR.n1539 0.0122188
R18404 VPWR.n4032 VPWR.n4031 0.0122188
R18405 VPWR.n1816 VPWR.n1815 0.0122188
R18406 VPWR.n2114 VPWR.n2112 0.0122188
R18407 VPWR.n3583 VPWR.n3581 0.0122188
R18408 VPWR.n3704 VPWR.n3703 0.0122188
R18409 VPWR.n3701 VPWR.n3700 0.0122188
R18410 VPWR.n2786 VPWR.n2784 0.0122188
R18411 VPWR.n2993 VPWR.n2992 0.0122188
R18412 VPWR.n2822 VPWR.n2821 0.0122188
R18413 VPWR.n3453 VPWR.n3452 0.0122188
R18414 VPWR.n6416 VPWR.n6415 0.0122188
R18415 VPWR.n6531 VPWR.n6530 0.0122188
R18416 VPWR.n7726 VPWR.n7725 0.0122188
R18417 VPWR.n102 VPWR.n101 0.0122188
R18418 VPWR.n99 VPWR.n98 0.0122188
R18419 VPWR.n2636 VPWR.n2635 0.0122188
R18420 VPWR.n2641 VPWR.n2638 0.0122188
R18421 VPWR.n3109 VPWR.n3108 0.0122188
R18422 VPWR.n3216 VPWR.n3214 0.0122188
R18423 VPWR.n3356 VPWR.n3354 0.0122188
R18424 VPWR.n3352 VPWR.n3351 0.0122188
R18425 VPWR.n6339 VPWR.n6338 0.0122188
R18426 VPWR.n6344 VPWR.n6341 0.0122188
R18427 VPWR.n6212 VPWR.n6210 0.0122188
R18428 VPWR.n5837 VPWR.n5836 0.0122188
R18429 VPWR.n5966 VPWR.n5965 0.0122188
R18430 VPWR.n5969 VPWR.n5968 0.0122188
R18431 VPWR.n1729 VPWR.n1728 0.0120783
R18432 VPWR.n1718 VPWR.n1717 0.01206
R18433 VPWR.n2998 VPWR.n2997 0.0118576
R18434 VPWR.n2811 VPWR.n2486 0.0118576
R18435 VPWR.n3494 VPWR.n3492 0.0118576
R18436 VPWR.n3504 VPWR.n3502 0.0118576
R18437 VPWR.n2366 VPWR.n2363 0.0118576
R18438 VPWR.n3141 VPWR.n3140 0.0117355
R18439 VPWR.n5548 VPWR.n5547 0.0117355
R18440 VPWR.n6909 VPWR.n6908 0.0115187
R18441 VPWR.n4785 VPWR.n4783 0.0114378
R18442 VPWR.n4035 VPWR.n4034 0.0114378
R18443 VPWR.n4045 VPWR.n4044 0.0114077
R18444 VPWR.n859 VPWR.n858 0.0111911
R18445 VPWR.n5138 VPWR.n5137 0.0109167
R18446 VPWR.n5140 VPWR.n5138 0.0109167
R18447 VPWR.n5671 VPWR.n5668 0.0109167
R18448 VPWR.n5666 VPWR.n5664 0.0109167
R18449 VPWR.n6697 VPWR.n6696 0.0109167
R18450 VPWR.n6662 VPWR.n6661 0.0109167
R18451 VPWR.n6762 VPWR.n6761 0.0109167
R18452 VPWR.n6759 VPWR.n6758 0.0109167
R18453 VPWR.n7605 VPWR.n157 0.0109167
R18454 VPWR.n208 VPWR.n206 0.0109167
R18455 VPWR.n210 VPWR.n208 0.0109167
R18456 VPWR.n217 VPWR.n216 0.0109167
R18457 VPWR.n5603 VPWR.n5602 0.0109167
R18458 VPWR.n5602 VPWR.n5601 0.0109167
R18459 VPWR.n5595 VPWR.n5592 0.0109167
R18460 VPWR.n5590 VPWR.n5588 0.0109167
R18461 VPWR.n5491 VPWR.n5490 0.0109167
R18462 VPWR.n5475 VPWR.n5474 0.0109167
R18463 VPWR.n5472 VPWR.n5471 0.0109167
R18464 VPWR.n6915 VPWR.n6914 0.0109167
R18465 VPWR.n6912 VPWR.n6911 0.0109167
R18466 VPWR VPWR.n6901 0.0109167
R18467 VPWR.n6872 VPWR.n6795 0.0109167
R18468 VPWR.n7413 VPWR.n7411 0.0109167
R18469 VPWR.n7415 VPWR.n7413 0.0109167
R18470 VPWR.n7422 VPWR.n7421 0.0109167
R18471 VPWR.n5344 VPWR.n5343 0.0109167
R18472 VPWR.n5343 VPWR.n5342 0.0109167
R18473 VPWR.n5336 VPWR.n5334 0.0109167
R18474 VPWR.n5332 VPWR.n5330 0.0109167
R18475 VPWR.n5298 VPWR.n5287 0.0109167
R18476 VPWR.n7035 VPWR.n7034 0.0109167
R18477 VPWR.n7032 VPWR.n7031 0.0109167
R18478 VPWR.n7188 VPWR.n7187 0.0109167
R18479 VPWR.n7185 VPWR.n7184 0.0109167
R18480 VPWR.n7149 VPWR 0.0109167
R18481 VPWR.n7210 VPWR.n293 0.0109167
R18482 VPWR.n7307 VPWR.n7306 0.0109167
R18483 VPWR.n559 VPWR.n558 0.0109167
R18484 VPWR.n561 VPWR.n559 0.0109167
R18485 VPWR.n691 VPWR.n690 0.0109167
R18486 VPWR.n719 VPWR.n718 0.0109167
R18487 VPWR.n864 VPWR.n863 0.0109167
R18488 VPWR.n861 VPWR.n860 0.0109167
R18489 VPWR.n831 VPWR 0.0109167
R18490 VPWR.n883 VPWR.n589 0.0109167
R18491 VPWR.n4772 VPWR.n4770 0.0109167
R18492 VPWR.n4774 VPWR.n4772 0.0109167
R18493 VPWR.n4775 VPWR 0.0109167
R18494 VPWR.n4783 VPWR.n4782 0.0109167
R18495 VPWR.n1072 VPWR.n1071 0.0109167
R18496 VPWR.n1074 VPWR.n1072 0.0109167
R18497 VPWR.n1082 VPWR.n1080 0.0109167
R18498 VPWR.n1086 VPWR.n1084 0.0109167
R18499 VPWR.n1120 VPWR.n1119 0.0109167
R18500 VPWR.n405 VPWR.n404 0.0109167
R18501 VPWR.n4544 VPWR.n4543 0.0109167
R18502 VPWR.n4541 VPWR.n4540 0.0109167
R18503 VPWR.n4603 VPWR.n4602 0.0109167
R18504 VPWR.n4696 VPWR.n4694 0.0109167
R18505 VPWR.n4698 VPWR.n4696 0.0109167
R18506 VPWR.n4705 VPWR.n4704 0.0109167
R18507 VPWR.n1260 VPWR.n1259 0.0109167
R18508 VPWR.n1259 VPWR.n1258 0.0109167
R18509 VPWR.n1303 VPWR.n1301 0.0109167
R18510 VPWR.n1307 VPWR.n1305 0.0109167
R18511 VPWR.n1417 VPWR.n1406 0.0109167
R18512 VPWR.n1389 VPWR.n1387 0.0109167
R18513 VPWR.n1385 VPWR.n1384 0.0109167
R18514 VPWR.n4320 VPWR.n4319 0.0109167
R18515 VPWR.n4317 VPWR.n1443 0.0109167
R18516 VPWR.n3800 VPWR.n3799 0.0109167
R18517 VPWR.n3948 VPWR.n3947 0.0109167
R18518 VPWR.n3947 VPWR.n3946 0.0109167
R18519 VPWR.n3941 VPWR.n3939 0.0109167
R18520 VPWR.n1929 VPWR.n1928 0.0109167
R18521 VPWR.n1931 VPWR.n1929 0.0109167
R18522 VPWR.n1939 VPWR.n1937 0.0109167
R18523 VPWR.n1943 VPWR.n1941 0.0109167
R18524 VPWR.n2028 VPWR.n2027 0.0109167
R18525 VPWR.n4240 VPWR.n4239 0.0109167
R18526 VPWR.n4237 VPWR.n4236 0.0109167
R18527 VPWR.n4168 VPWR.n4167 0.0109167
R18528 VPWR.n4165 VPWR.n4164 0.0109167
R18529 VPWR.n4128 VPWR.n1519 0.0109167
R18530 VPWR.n4034 VPWR.n4033 0.0109167
R18531 VPWR.n1730 VPWR.n1729 0.0109167
R18532 VPWR.n2104 VPWR.n2103 0.0109167
R18533 VPWR.n2085 VPWR.n2083 0.0109167
R18534 VPWR.n2081 VPWR.n2080 0.0109167
R18535 VPWR.n3552 VPWR.n3551 0.0109167
R18536 VPWR.n3556 VPWR.n3554 0.0109167
R18537 VPWR.n3575 VPWR.n3574 0.0109167
R18538 VPWR.n3699 VPWR.n3698 0.0109167
R18539 VPWR.n2762 VPWR.n2761 0.0109167
R18540 VPWR.n2764 VPWR.n2762 0.0109167
R18541 VPWR.n2788 VPWR.n2786 0.0109167
R18542 VPWR.n2792 VPWR.n2790 0.0109167
R18543 VPWR.n2829 VPWR.n2828 0.0109167
R18544 VPWR.n2844 VPWR.n2843 0.0109167
R18545 VPWR.n2847 VPWR.n2846 0.0109167
R18546 VPWR.n3483 VPWR.n3482 0.0109167
R18547 VPWR.n3480 VPWR.n3479 0.0109167
R18548 VPWR.n3460 VPWR.n3459 0.0109167
R18549 VPWR.n3422 VPWR.n3420 0.0109167
R18550 VPWR.n3420 VPWR.n3418 0.0109167
R18551 VPWR VPWR.n3416 0.0109167
R18552 VPWR.n2333 VPWR.n2332 0.0109167
R18553 VPWR.n6431 VPWR.n6430 0.0109167
R18554 VPWR.n6430 VPWR.n6429 0.0109167
R18555 VPWR.n6415 VPWR.n6412 0.0109167
R18556 VPWR.n6410 VPWR.n5066 0.0109167
R18557 VPWR.n6538 VPWR.n6537 0.0109167
R18558 VPWR.n6559 VPWR.n6558 0.0109167
R18559 VPWR.n6562 VPWR.n6561 0.0109167
R18560 VPWR.n7779 VPWR.n7778 0.0109167
R18561 VPWR.n7776 VPWR.n7775 0.0109167
R18562 VPWR.n7732 VPWR.n29 0.0109167
R18563 VPWR.n97 VPWR.n96 0.0109167
R18564 VPWR.n2632 VPWR.n2631 0.0109167
R18565 VPWR.n2634 VPWR.n2632 0.0109167
R18566 VPWR.n2643 VPWR.n2641 0.0109167
R18567 VPWR.n2647 VPWR.n2645 0.0109167
R18568 VPWR.n3102 VPWR.n3101 0.0109167
R18569 VPWR.n3083 VPWR.n3081 0.0109167
R18570 VPWR.n3079 VPWR.n3078 0.0109167
R18571 VPWR.n3173 VPWR.n3172 0.0109167
R18572 VPWR.n3176 VPWR.n3175 0.0109167
R18573 VPWR.n3208 VPWR.n2386 0.0109167
R18574 VPWR.n3360 VPWR.n3358 0.0109167
R18575 VPWR.n3358 VPWR.n3356 0.0109167
R18576 VPWR.n3350 VPWR.n3348 0.0109167
R18577 VPWR.n6335 VPWR.n6334 0.0109167
R18578 VPWR.n6337 VPWR.n6335 0.0109167
R18579 VPWR.n6346 VPWR.n6344 0.0109167
R18580 VPWR.n6350 VPWR.n6348 0.0109167
R18581 VPWR.n6204 VPWR.n6203 0.0109167
R18582 VPWR.n6185 VPWR.n6183 0.0109167
R18583 VPWR.n6181 VPWR.n6180 0.0109167
R18584 VPWR.n6105 VPWR.n6104 0.0109167
R18585 VPWR.n6102 VPWR.n6101 0.0109167
R18586 VPWR.n7808 VPWR.n7807 0.0109167
R18587 VPWR.n5963 VPWR.n5961 0.0109167
R18588 VPWR.n5965 VPWR.n5963 0.0109167
R18589 VPWR.n5972 VPWR.n5971 0.0109167
R18590 VPWR.n4945 VPWR.n4944 0.0106351
R18591 VPWR.n4886 VPWR.n4885 0.0106351
R18592 VPWR.n7014 VPWR.n7013 0.0106351
R18593 VPWR.n631 VPWR.n630 0.0106351
R18594 VPWR.n414 VPWR.n413 0.0106351
R18595 VPWR.n4398 VPWR.n4397 0.0106351
R18596 VPWR.n1458 VPWR.n1457 0.0106351
R18597 VPWR.n2055 VPWR.n2054 0.0106351
R18598 VPWR.n5804 VPWR.n5803 0.0106351
R18599 VPWR.n3026 VPWR.n3025 0.0106351
R18600 VPWR.n3040 VPWR.n3039 0.0106351
R18601 VPWR.n5774 VPWR.n5773 0.0106351
R18602 VPWR.n7068 VPWR 0.0101142
R18603 VPWR VPWR.n740 0.0101142
R18604 VPWR.n126 VPWR.n115 0.00975758
R18605 VPWR.n117 VPWR.n116 0.00975758
R18606 VPWR.n7641 VPWR.n7640 0.00975758
R18607 VPWR.n7654 VPWR.n7653 0.00975758
R18608 VPWR.n254 VPWR.n241 0.00975758
R18609 VPWR.n253 VPWR.n252 0.00975758
R18610 VPWR.n7499 VPWR.n7498 0.00975758
R18611 VPWR.n7511 VPWR.n7510 0.00975758
R18612 VPWR.n7631 VPWR.n133 0.00975758
R18613 VPWR.n146 VPWR.n145 0.00975758
R18614 VPWR.n143 VPWR.n142 0.00975758
R18615 VPWR.n5684 VPWR.n5075 0.00975758
R18616 VPWR.n5683 VPWR.n5682 0.00975758
R18617 VPWR.n5680 VPWR.n5679 0.00975758
R18618 VPWR.n6674 VPWR.n4948 0.00975758
R18619 VPWR.n6673 VPWR.n6672 0.00975758
R18620 VPWR.n6670 VPWR.n6669 0.00975758
R18621 VPWR.n7494 VPWR.n258 0.00975758
R18622 VPWR.n270 VPWR.n269 0.00975758
R18623 VPWR.n267 VPWR.n266 0.00975758
R18624 VPWR.n6890 VPWR.n4933 0.00975758
R18625 VPWR.n6892 VPWR.n6891 0.00975758
R18626 VPWR.n6895 VPWR.n6894 0.00975758
R18627 VPWR.n5653 VPWR.n5629 0.00975758
R18628 VPWR.n5652 VPWR.n5651 0.00975758
R18629 VPWR.n5649 VPWR.n5648 0.00975758
R18630 VPWR.n4907 VPWR.n4883 0.00975758
R18631 VPWR.n4906 VPWR.n4905 0.00975758
R18632 VPWR.n4903 VPWR.n4902 0.00975758
R18633 VPWR.n7394 VPWR.n286 0.00975758
R18634 VPWR.n7383 VPWR.n7382 0.00975758
R18635 VPWR.n7380 VPWR.n7379 0.00975758
R18636 VPWR.n7173 VPWR.n7147 0.00975758
R18637 VPWR.n7172 VPWR.n7171 0.00975758
R18638 VPWR.n7169 VPWR.n7168 0.00975758
R18639 VPWR.n5421 VPWR.n5213 0.00975758
R18640 VPWR.n5420 VPWR.n5419 0.00975758
R18641 VPWR.n5417 VPWR.n5416 0.00975758
R18642 VPWR.n7059 VPWR.n7011 0.00975758
R18643 VPWR.n7058 VPWR.n7057 0.00975758
R18644 VPWR.n7055 VPWR.n7054 0.00975758
R18645 VPWR.n4853 VPWR.n303 0.00975758
R18646 VPWR.n315 VPWR.n314 0.00975758
R18647 VPWR.n312 VPWR.n311 0.00975758
R18648 VPWR.n849 VPWR.n830 0.00975758
R18649 VPWR.n848 VPWR.n847 0.00975758
R18650 VPWR.n845 VPWR.n844 0.00975758
R18651 VPWR.n547 VPWR.n537 0.00975758
R18652 VPWR.n546 VPWR.n545 0.00975758
R18653 VPWR.n543 VPWR.n542 0.00975758
R18654 VPWR.n731 VPWR.n628 0.00975758
R18655 VPWR.n730 VPWR.n729 0.00975758
R18656 VPWR.n727 VPWR.n726 0.00975758
R18657 VPWR.n4753 VPWR.n4730 0.00975758
R18658 VPWR.n4742 VPWR.n4741 0.00975758
R18659 VPWR.n4739 VPWR.n4738 0.00975758
R18660 VPWR.n4585 VPWR.n386 0.00975758
R18661 VPWR.n4584 VPWR.n4583 0.00975758
R18662 VPWR.n4581 VPWR.n4580 0.00975758
R18663 VPWR.n1006 VPWR.n982 0.00975758
R18664 VPWR.n1005 VPWR.n1004 0.00975758
R18665 VPWR.n1002 VPWR.n1001 0.00975758
R18666 VPWR.n4446 VPWR.n411 0.00975758
R18667 VPWR.n4448 VPWR.n4447 0.00975758
R18668 VPWR.n4451 VPWR.n4450 0.00975758
R18669 VPWR.n3761 VPWR.n3738 0.00975758
R18670 VPWR.n3750 VPWR.n3749 0.00975758
R18671 VPWR.n3747 VPWR.n3746 0.00975758
R18672 VPWR.n4313 VPWR.n1449 0.00975758
R18673 VPWR.n4312 VPWR.n4311 0.00975758
R18674 VPWR.n4309 VPWR.n4308 0.00975758
R18675 VPWR.n1285 VPWR.n448 0.00975758
R18676 VPWR.n1287 VPWR.n1286 0.00975758
R18677 VPWR.n1290 VPWR.n1289 0.00975758
R18678 VPWR.n4419 VPWR.n4395 0.00975758
R18679 VPWR.n4418 VPWR.n4417 0.00975758
R18680 VPWR.n4415 VPWR.n4414 0.00975758
R18681 VPWR.n3985 VPWR.n3962 0.00975758
R18682 VPWR.n3974 VPWR.n3973 0.00975758
R18683 VPWR.n3971 VPWR.n3970 0.00975758
R18684 VPWR.n4148 VPWR.n1495 0.00975758
R18685 VPWR.n4147 VPWR.n4146 0.00975758
R18686 VPWR.n4144 VPWR.n4143 0.00975758
R18687 VPWR.n1917 VPWR.n1653 0.00975758
R18688 VPWR.n1916 VPWR.n1915 0.00975758
R18689 VPWR.n1913 VPWR.n1912 0.00975758
R18690 VPWR.n4269 VPWR.n1455 0.00975758
R18691 VPWR.n4268 VPWR.n4267 0.00975758
R18692 VPWR.n4265 VPWR.n4264 0.00975758
R18693 VPWR.n1828 VPWR.n1657 0.00975758
R18694 VPWR.n1827 VPWR.n1826 0.00975758
R18695 VPWR.n1824 VPWR.n1823 0.00975758
R18696 VPWR.n2187 VPWR.n2162 0.00975758
R18697 VPWR.n2186 VPWR.n2185 0.00975758
R18698 VPWR.n2183 VPWR.n2182 0.00975758
R18699 VPWR.n3731 VPWR.n3718 0.00975758
R18700 VPWR.n3721 VPWR.n3720 0.00975758
R18701 VPWR.n1552 VPWR.n1551 0.00975758
R18702 VPWR.n1564 VPWR.n1554 0.00975758
R18703 VPWR.n2063 VPWR.n2039 0.00975758
R18704 VPWR.n2052 VPWR.n2051 0.00975758
R18705 VPWR.n2049 VPWR.n2048 0.00975758
R18706 VPWR.n5812 VPWR.n5796 0.00975758
R18707 VPWR.n5801 VPWR.n5800 0.00975758
R18708 VPWR.n5798 VPWR.n5797 0.00975758
R18709 VPWR.n4967 VPWR.n4966 0.00975758
R18710 VPWR.n3410 VPWR.n2282 0.00975758
R18711 VPWR.n3409 VPWR.n3408 0.00975758
R18712 VPWR.n2287 VPWR.n2286 0.00975758
R18713 VPWR.n2738 VPWR.n2737 0.00975758
R18714 VPWR.n2726 VPWR.n2725 0.00975758
R18715 VPWR.n2771 VPWR.n2770 0.00975758
R18716 VPWR.n2774 VPWR.n2773 0.00975758
R18717 VPWR.n3520 VPWR.n3507 0.00975758
R18718 VPWR.n3510 VPWR.n3509 0.00975758
R18719 VPWR.n2190 VPWR.n2189 0.00975758
R18720 VPWR.n2204 VPWR.n2192 0.00975758
R18721 VPWR.n3034 VPWR.n3020 0.00975758
R18722 VPWR.n3022 VPWR.n3021 0.00975758
R18723 VPWR.n3005 VPWR.n3004 0.00975758
R18724 VPWR.n3016 VPWR.n3015 0.00975758
R18725 VPWR.n3048 VPWR.n3047 0.00975758
R18726 VPWR.n3051 VPWR.n3050 0.00975758
R18727 VPWR.n3065 VPWR.n3064 0.00975758
R18728 VPWR.n5782 VPWR.n5766 0.00975758
R18729 VPWR.n5771 VPWR.n5770 0.00975758
R18730 VPWR.n5768 VPWR.n5767 0.00975758
R18731 VPWR.n5761 VPWR.n5760 0.00975758
R18732 VPWR.n2405 VPWR.n2404 0.00975758
R18733 VPWR.n2408 VPWR.n2407 0.00975758
R18734 VPWR.n3199 VPWR.n3198 0.00975758
R18735 VPWR.n8 VPWR.n7 0.00975758
R18736 VPWR.n10 VPWR.n9 0.00975758
R18737 VPWR.n13 VPWR.n12 0.00975758
R18738 VPWR.n15 VPWR.n14 0.00975758
R18739 VPWR.n7758 VPWR.n7757 0.00975758
R18740 VPWR.n7761 VPWR.n7760 0.00975758
R18741 VPWR.n7763 VPWR.n7762 0.00975758
R18742 VPWR.n6376 VPWR.n6359 0.00975758
R18743 VPWR.n6375 VPWR.n6374 0.00975758
R18744 VPWR.n6372 VPWR.n6371 0.00975758
R18745 VPWR.n6423 VPWR.n6422 0.00975758
R18746 VPWR.n5708 VPWR.n5691 0.00975758
R18747 VPWR.n5696 VPWR.n5695 0.00975758
R18748 VPWR.n5693 VPWR.n5692 0.00975758
R18749 VPWR.n5723 VPWR.n5722 0.00975758
R18750 VPWR.n2676 VPWR.n2653 0.00975758
R18751 VPWR.n2664 VPWR.n2663 0.00975758
R18752 VPWR.n2661 VPWR.n2660 0.00975758
R18753 VPWR.n3381 VPWR.n3380 0.00975758
R18754 VPWR.n3384 VPWR.n3383 0.00975758
R18755 VPWR.n3398 VPWR.n3397 0.00975758
R18756 VPWR.n6020 VPWR.n6019 0.00975758
R18757 VPWR.n6010 VPWR.n6009 0.00975758
R18758 VPWR.n6007 VPWR.n6006 0.00975758
R18759 VPWR.n6005 VPWR.n5996 0.00975758
R18760 VPWR.n5668 VPWR.n5666 0.00961458
R18761 VPWR.n6663 VPWR.n6662 0.00961458
R18762 VPWR.n6761 VPWR.n6760 0.00961458
R18763 VPWR.n7620 VPWR.n7618 0.00961458
R18764 VPWR.n206 VPWR.n162 0.00961458
R18765 VPWR.n218 VPWR.n217 0.00961458
R18766 VPWR.n5592 VPWR.n5590 0.00961458
R18767 VPWR.n5473 VPWR.n5472 0.00961458
R18768 VPWR.n6914 VPWR.n6913 0.00961458
R18769 VPWR.n6902 VPWR 0.00961458
R18770 VPWR.n6792 VPWR.n6791 0.00961458
R18771 VPWR.n7411 VPWR.n7409 0.00961458
R18772 VPWR.n7423 VPWR.n7422 0.00961458
R18773 VPWR.n5334 VPWR.n5332 0.00961458
R18774 VPWR.n5301 VPWR.n5300 0.00961458
R18775 VPWR.n7033 VPWR.n7032 0.00961458
R18776 VPWR.n7187 VPWR.n7186 0.00961458
R18777 VPWR VPWR.n7148 0.00961458
R18778 VPWR.n7163 VPWR.n7161 0.00961458
R18779 VPWR.n7309 VPWR.n7307 0.00961458
R18780 VPWR.n688 VPWR.n687 0.00961458
R18781 VPWR.n720 VPWR.n719 0.00961458
R18782 VPWR.n863 VPWR.n862 0.00961458
R18783 VPWR VPWR.n823 0.00961458
R18784 VPWR.n4770 VPWR.n4768 0.00961458
R18785 VPWR.n1084 VPWR.n1082 0.00961458
R18786 VPWR.n1125 VPWR.n1123 0.00961458
R18787 VPWR.n406 VPWR.n405 0.00961458
R18788 VPWR.n4543 VPWR.n4542 0.00961458
R18789 VPWR.n4599 VPWR.n4598 0.00961458
R18790 VPWR.n4694 VPWR.n4692 0.00961458
R18791 VPWR.n4706 VPWR.n4705 0.00961458
R18792 VPWR.n1305 VPWR.n1303 0.00961458
R18793 VPWR.n1386 VPWR.n1385 0.00961458
R18794 VPWR.n4319 VPWR.n4318 0.00961458
R18795 VPWR.n3796 VPWR.n3795 0.00961458
R18796 VPWR.n3949 VPWR.n3948 0.00961458
R18797 VPWR.n3939 VPWR.n3938 0.00961458
R18798 VPWR.n1941 VPWR.n1939 0.00961458
R18799 VPWR.n2022 VPWR.n2020 0.00961458
R18800 VPWR.n4238 VPWR.n4237 0.00961458
R18801 VPWR.n4167 VPWR.n4166 0.00961458
R18802 VPWR.n1514 VPWR.n1513 0.00961458
R18803 VPWR.n2111 VPWR.n2109 0.00961458
R18804 VPWR.n2082 VPWR.n2081 0.00961458
R18805 VPWR.n3553 VPWR.n3552 0.00961458
R18806 VPWR.n3571 VPWR.n3570 0.00961458
R18807 VPWR.n3698 VPWR.n3697 0.00961458
R18808 VPWR.n2790 VPWR.n2788 0.00961458
R18809 VPWR.n2826 VPWR.n2824 0.00961458
R18810 VPWR.n2846 VPWR.n2845 0.00961458
R18811 VPWR.n3482 VPWR.n3481 0.00961458
R18812 VPWR.n3465 VPWR.n3463 0.00961458
R18813 VPWR.n3424 VPWR.n3422 0.00961458
R18814 VPWR.n2334 VPWR.n2333 0.00961458
R18815 VPWR.n6412 VPWR.n6410 0.00961458
R18816 VPWR.n6535 VPWR.n6533 0.00961458
R18817 VPWR.n6561 VPWR.n6560 0.00961458
R18818 VPWR.n7778 VPWR.n7777 0.00961458
R18819 VPWR.n7741 VPWR.n7739 0.00961458
R18820 VPWR.n96 VPWR.n95 0.00961458
R18821 VPWR.n2645 VPWR.n2643 0.00961458
R18822 VPWR.n3107 VPWR.n3105 0.00961458
R18823 VPWR.n3080 VPWR.n3079 0.00961458
R18824 VPWR.n3174 VPWR.n3173 0.00961458
R18825 VPWR.n3189 VPWR.n3188 0.00961458
R18826 VPWR.n3362 VPWR.n3360 0.00961458
R18827 VPWR.n3348 VPWR.n3347 0.00961458
R18828 VPWR.n6348 VPWR.n6346 0.00961458
R18829 VPWR.n6209 VPWR.n6207 0.00961458
R18830 VPWR.n6182 VPWR.n6181 0.00961458
R18831 VPWR.n6104 VPWR.n6103 0.00961458
R18832 VPWR.n6091 VPWR.n6087 0.00961458
R18833 VPWR.n5961 VPWR.n5906 0.00961458
R18834 VPWR.n5973 VPWR.n5972 0.00961458
R18835 VPWR.n3037 VPWR.n3036 0.00956852
R18836 VPWR.n2394 VPWR.n2393 0.00956852
R18837 VPWR.n2683 VPWR.n2682 0.00956852
R18838 VPWR.n3402 VPWR.n3401 0.00956852
R18839 VPWR.n2495 VPWR.n2493 0.00894595
R18840 VPWR.n2650 VPWR.n2649 0.00894595
R18841 VPWR.n7661 VPWR.n7660 0.00894595
R18842 VPWR.n111 VPWR.n110 0.00894595
R18843 VPWR.n7790 VPWR.n7784 0.00894595
R18844 VPWR.n7755 VPWR.n7751 0.00894595
R18845 VPWR.n7734 VPWR.n7733 0.00894595
R18846 VPWR.n7518 VPWR.n7517 0.00894595
R18847 VPWR.n237 VPWR.n236 0.00894595
R18848 VPWR.n6765 VPWR.n4936 0.00894595
R18849 VPWR.n7630 VPWR.n151 0.00894595
R18850 VPWR.n7612 VPWR.n7606 0.00894595
R18851 VPWR.n5122 VPWR.n5121 0.00894595
R18852 VPWR.n5661 VPWR.n5660 0.00894595
R18853 VPWR.n6598 VPWR.n6594 0.00894595
R18854 VPWR.n4946 VPWR.n4945 0.00894595
R18855 VPWR.n6667 VPWR.n6666 0.00894595
R18856 VPWR.n6658 VPWR.n6604 0.00894595
R18857 VPWR.n7402 VPWR.n7401 0.00894595
R18858 VPWR.n7474 VPWR.n7435 0.00894595
R18859 VPWR.n6776 VPWR.n4927 0.00894595
R18860 VPWR.n6889 VPWR.n6883 0.00894595
R18861 VPWR.n6874 VPWR.n6873 0.00894595
R18862 VPWR.n5623 VPWR.n5621 0.00894595
R18863 VPWR.n5585 VPWR.n5584 0.00894595
R18864 VPWR.n7005 VPWR.n7001 0.00894595
R18865 VPWR.n4887 VPWR.n4886 0.00894595
R18866 VPWR.n4900 VPWR.n4899 0.00894595
R18867 VPWR.n6993 VPWR.n6992 0.00894595
R18868 VPWR.n7296 VPWR.n7295 0.00894595
R18869 VPWR.n7364 VPWR.n7325 0.00894595
R18870 VPWR.n7200 VPWR.n7197 0.00894595
R18871 VPWR.n7174 VPWR.n7145 0.00894595
R18872 VPWR.n7209 VPWR.n7206 0.00894595
R18873 VPWR.n5386 VPWR.n5385 0.00894595
R18874 VPWR.n5327 VPWR.n5229 0.00894595
R18875 VPWR.n5297 VPWR.n5296 0.00894595
R18876 VPWR.n7015 VPWR.n7014 0.00894595
R18877 VPWR.n7052 VPWR.n7051 0.00894595
R18878 VPWR.n7065 VPWR.n7064 0.00894595
R18879 VPWR.n4761 VPWR.n4760 0.00894595
R18880 VPWR.n4833 VPWR.n4795 0.00894595
R18881 VPWR.n873 VPWR.n870 0.00894595
R18882 VPWR.n850 VPWR.n828 0.00894595
R18883 VPWR.n882 VPWR.n879 0.00894595
R18884 VPWR.n516 VPWR.n515 0.00894595
R18885 VPWR.n976 VPWR.n975 0.00894595
R18886 VPWR.n622 VPWR.n618 0.00894595
R18887 VPWR.n632 VPWR.n631 0.00894595
R18888 VPWR.n724 VPWR.n723 0.00894595
R18889 VPWR.n737 VPWR.n736 0.00894595
R18890 VPWR.n4684 VPWR.n4683 0.00894595
R18891 VPWR.n4725 VPWR.n4724 0.00894595
R18892 VPWR.n4554 VPWR.n4551 0.00894595
R18893 VPWR.n4586 VPWR.n384 0.00894595
R18894 VPWR.n4567 VPWR.n4566 0.00894595
R18895 VPWR.n1053 VPWR.n1052 0.00894595
R18896 VPWR.n1208 VPWR.n1207 0.00894595
R18897 VPWR.n4431 VPWR.n4427 0.00894595
R18898 VPWR.n415 VPWR.n414 0.00894595
R18899 VPWR.n4454 VPWR.n4453 0.00894595
R18900 VPWR.n4441 VPWR.n399 0.00894595
R18901 VPWR.n3955 VPWR.n3951 0.00894595
R18902 VPWR.n3770 VPWR.n3769 0.00894595
R18903 VPWR.n4282 VPWR.n1437 0.00894595
R18904 VPWR.n4315 VPWR.n4314 0.00894595
R18905 VPWR.n4295 VPWR.n4294 0.00894595
R18906 VPWR.n1279 VPWR.n1277 0.00894595
R18907 VPWR.n1222 VPWR.n444 0.00894595
R18908 VPWR.n1416 VPWR.n1415 0.00894595
R18909 VPWR.n4399 VPWR.n4398 0.00894595
R18910 VPWR.n4412 VPWR.n4411 0.00894595
R18911 VPWR.n4390 VPWR.n4389 0.00894595
R18912 VPWR.n4056 VPWR.n4055 0.00894595
R18913 VPWR.n4048 VPWR.n4047 0.00894595
R18914 VPWR.n1500 VPWR.n1486 0.00894595
R18915 VPWR.n4149 VPWR.n1493 0.00894595
R18916 VPWR.n4130 VPWR.n4129 0.00894595
R18917 VPWR.n1899 VPWR.n1897 0.00894595
R18918 VPWR.n1840 VPWR.n1649 0.00894595
R18919 VPWR.n2033 VPWR.n2029 0.00894595
R18920 VPWR.n4249 VPWR.n1458 0.00894595
R18921 VPWR.n4262 VPWR.n4261 0.00894595
R18922 VPWR.n1473 VPWR.n1472 0.00894595
R18923 VPWR.n1714 VPWR.n1713 0.00894595
R18924 VPWR.n1811 VPWR.n1810 0.00894595
R18925 VPWR.n3544 VPWR.n3543 0.00894595
R18926 VPWR.n2173 VPWR.n2167 0.00894595
R18927 VPWR.n3536 VPWR.n3535 0.00894595
R18928 VPWR.n3712 VPWR.n3708 0.00894595
R18929 VPWR.n1547 VPWR.n1546 0.00894595
R18930 VPWR.n2105 VPWR.n1591 0.00894595
R18931 VPWR.n2056 VPWR.n2055 0.00894595
R18932 VPWR.n2046 VPWR.n2045 0.00894595
R18933 VPWR.n2074 VPWR.n2073 0.00894595
R18934 VPWR.n4955 VPWR.n4951 0.00894595
R18935 VPWR.n5805 VPWR.n5804 0.00894595
R18936 VPWR.n4965 VPWR.n4964 0.00894595
R18937 VPWR.n6569 VPWR.n6568 0.00894595
R18938 VPWR.n2277 VPWR.n2269 0.00894595
R18939 VPWR.n2362 VPWR.n2361 0.00894595
R18940 VPWR.n2744 VPWR.n2743 0.00894595
R18941 VPWR.n2996 VPWR.n2995 0.00894595
R18942 VPWR.n3491 VPWR.n3488 0.00894595
R18943 VPWR.n3519 VPWR.n3515 0.00894595
R18944 VPWR.n3501 VPWR.n3500 0.00894595
R18945 VPWR.n2481 VPWR.n2478 0.00894595
R18946 VPWR.n3027 VPWR.n3026 0.00894595
R18947 VPWR.n3014 VPWR.n3013 0.00894595
R18948 VPWR.n2813 VPWR.n2812 0.00894595
R18949 VPWR.n2469 VPWR.n2464 0.00894595
R18950 VPWR.n3041 VPWR.n3040 0.00894595
R18951 VPWR.n3062 VPWR.n3061 0.00894595
R18952 VPWR.n3071 VPWR.n3070 0.00894595
R18953 VPWR.n5790 VPWR.n5786 0.00894595
R18954 VPWR.n5775 VPWR.n5774 0.00894595
R18955 VPWR.n5759 VPWR.n5758 0.00894595
R18956 VPWR.n5820 VPWR.n5819 0.00894595
R18957 VPWR.n3162 VPWR.n3161 0.00894595
R18958 VPWR.n2402 VPWR.n2398 0.00894595
R18959 VPWR.n3207 VPWR.n3204 0.00894595
R18960 VPWR.n6084 VPWR.n6083 0.00894595
R18961 VPWR.n6076 VPWR.n6075 0.00894595
R18962 VPWR.n7806 VPWR.n7803 0.00894595
R18963 VPWR.n6448 VPWR.n6446 0.00894595
R18964 VPWR.n6457 VPWR.n6456 0.00894595
R18965 VPWR.n5712 VPWR.n5710 0.00894595
R18966 VPWR.n6353 VPWR.n6352 0.00894595
R18967 VPWR.n3369 VPWR.n3364 0.00894595
R18968 VPWR.n2375 VPWR.n2374 0.00894595
R18969 VPWR.n6025 VPWR.n6024 0.00894595
R18970 VPWR.n5992 VPWR.n5991 0.00894595
R18971 VPWR.n2488 VPWR.n2487 0.00837842
R18972 VPWR.n2368 VPWR.n2367 0.00837842
R18973 VPWR.n2370 VPWR.n2369 0.00837842
R18974 VPWR.n6693 VPWR.n6692 0.0083125
R18975 VPWR.n6610 VPWR 0.0083125
R18976 VPWR.n7603 VPWR.n7602 0.0083125
R18977 VPWR.n5487 VPWR.n5486 0.0083125
R18978 VPWR.n7022 VPWR.n7018 0.0083125
R18979 VPWR.n7213 VPWR 0.0083125
R18980 VPWR.n701 VPWR.n694 0.0083125
R18981 VPWR VPWR.n716 0.0083125
R18982 VPWR.n1116 VPWR.n1115 0.0083125
R18983 VPWR.n4608 VPWR.n4606 0.0083125
R18984 VPWR.n1403 VPWR.n1402 0.0083125
R18985 VPWR.n2024 VPWR.n1460 0.0083125
R18986 VPWR.n4126 VPWR.n4124 0.0083125
R18987 VPWR.n4121 VPWR 0.0083125
R18988 VPWR.n2100 VPWR.n2099 0.0083125
R18989 VPWR.n3580 VPWR.n3578 0.0083125
R18990 VPWR.n2834 VPWR.n2832 0.0083125
R18991 VPWR.n3457 VPWR.n3455 0.0083125
R18992 VPWR.n6544 VPWR.n6541 0.0083125
R18993 VPWR.n7730 VPWR.n7728 0.0083125
R18994 VPWR.n3098 VPWR.n3097 0.0083125
R18995 VPWR.n3213 VPWR.n3211 0.0083125
R18996 VPWR.n6200 VPWR.n6199 0.0083125
R18997 VPWR.n6869 VPWR.n6867 0.00757276
R18998 VPWR.n7215 VPWR.n7214 0.00757276
R18999 VPWR.n886 VPWR.n585 0.00757276
R19000 VPWR.n3805 VPWR.n3804 0.00757276
R19001 VPWR.n5836 VPWR.n5835 0.00757276
R19002 VPWR.n6908 VPWR.n6905 0.00739914
R19003 VPWR.n7769 VPWR.n7768 0.00725676
R19004 VPWR.n7749 VPWR.n7748 0.00725676
R19005 VPWR.n7626 VPWR.n152 0.00725676
R19006 VPWR.n139 VPWR.n138 0.00725676
R19007 VPWR.n6680 VPWR.n6679 0.00725676
R19008 VPWR.n6885 VPWR.n6884 0.00725676
R19009 VPWR.n4931 VPWR.n4930 0.00725676
R19010 VPWR.n4889 VPWR.n4888 0.00725676
R19011 VPWR.n7178 VPWR.n7177 0.00725676
R19012 VPWR.n7165 VPWR.n7154 0.00725676
R19013 VPWR.n7041 VPWR.n7040 0.00725676
R19014 VPWR.n855 VPWR.n854 0.00725676
R19015 VPWR.n841 VPWR.n836 0.00725676
R19016 VPWR.n710 VPWR.n709 0.00725676
R19017 VPWR.n4591 VPWR.n4590 0.00725676
R19018 VPWR.n4577 VPWR.n4576 0.00725676
R19019 VPWR.n1108 VPWR.n1107 0.00725676
R19020 VPWR.n3788 VPWR.n3787 0.00725676
R19021 VPWR.n4305 VPWR.n4304 0.00725676
R19022 VPWR.n4401 VPWR.n4400 0.00725676
R19023 VPWR.n4154 VPWR.n4153 0.00725676
R19024 VPWR.n4140 VPWR.n4139 0.00725676
R19025 VPWR.n4251 VPWR.n4250 0.00725676
R19026 VPWR.n2169 VPWR.n2168 0.00725676
R19027 VPWR.n2179 VPWR.n2178 0.00725676
R19028 VPWR.n2058 VPWR.n2057 0.00725676
R19029 VPWR.n5807 VPWR.n5806 0.00725676
R19030 VPWR.n2194 VPWR.n2193 0.00725676
R19031 VPWR.n2202 VPWR.n2201 0.00725676
R19032 VPWR.n3029 VPWR.n3028 0.00725676
R19033 VPWR.n3053 VPWR.n3052 0.00725676
R19034 VPWR.n5777 VPWR.n5776 0.00725676
R19035 VPWR.n2410 VPWR.n2409 0.00725676
R19036 VPWR.n3195 VPWR.n3194 0.00725676
R19037 VPWR.n6071 VPWR.n6070 0.00725676
R19038 VPWR.n6065 VPWR.n6064 0.00725676
R19039 VPWR VPWR.n5674 0.00701042
R19040 VPWR.n6692 VPWR.n6685 0.00701042
R19041 VPWR VPWR.n7617 0.00701042
R19042 VPWR.n5486 VPWR.n5485 0.00701042
R19043 VPWR VPWR.n5328 0.00701042
R19044 VPWR.n7023 VPWR.n7022 0.00701042
R19045 VPWR VPWR.n7312 0.00701042
R19046 VPWR VPWR.n471 0.00701042
R19047 VPWR.n702 VPWR.n701 0.00701042
R19048 VPWR.n4781 VPWR 0.00701042
R19049 VPWR.n1115 VPWR.n1113 0.00701042
R19050 VPWR.n4458 VPWR 0.00701042
R19051 VPWR.n1297 VPWR 0.00701042
R19052 VPWR.n1402 VPWR.n1401 0.00701042
R19053 VPWR.n4248 VPWR.n1460 0.00701042
R19054 VPWR VPWR.n1818 0.00701042
R19055 VPWR.n1592 VPWR 0.00701042
R19056 VPWR.n2099 VPWR.n2097 0.00701042
R19057 VPWR.n2782 VPWR 0.00701042
R19058 VPWR.n2835 VPWR.n2834 0.00701042
R19059 VPWR.n2330 VPWR 0.00701042
R19060 VPWR VPWR.n6418 0.00701042
R19061 VPWR.n6545 VPWR.n6544 0.00701042
R19062 VPWR.n3097 VPWR.n3095 0.00701042
R19063 VPWR.n3191 VPWR 0.00701042
R19064 VPWR.n6199 VPWR.n6197 0.00701042
R19065 VPWR VPWR.n6086 0.00701042
R19066 VPWR.n2371 VPWR.n2370 0.00696227
R19067 VPWR.n6702 VPWR.n6701 0.00693178
R19068 VPWR.n5495 VPWR.n5494 0.00693178
R19069 VPWR.n1422 VPWR.n1421 0.00693178
R19070 VPWR.n3002 VPWR.n2488 0.00657697
R19071 VPWR.n2367 VPWR.n2206 0.00657697
R19072 VPWR.n2366 VPWR.n2365 0.00648266
R19073 VPWR.n2998 VPWR.n2685 0.00648266
R19074 VPWR.n3494 VPWR.n3493 0.00648266
R19075 VPWR.n3504 VPWR.n3503 0.00648266
R19076 VPWR.n2486 VPWR.n2485 0.00648266
R19077 VPWR.n126 VPWR.n117 0.00619697
R19078 VPWR.n7654 VPWR.n7641 0.00619697
R19079 VPWR.n254 VPWR.n253 0.00619697
R19080 VPWR.n7511 VPWR.n7499 0.00619697
R19081 VPWR.n7631 VPWR.n146 0.00619697
R19082 VPWR.n142 VPWR.n141 0.00619697
R19083 VPWR.n5684 VPWR.n5683 0.00619697
R19084 VPWR.n5679 VPWR.n5678 0.00619697
R19085 VPWR.n6674 VPWR.n6673 0.00619697
R19086 VPWR.n6669 VPWR.n6668 0.00619697
R19087 VPWR.n7494 VPWR.n270 0.00619697
R19088 VPWR.n266 VPWR.n265 0.00619697
R19089 VPWR.n6891 VPWR.n6890 0.00619697
R19090 VPWR.n6896 VPWR.n6895 0.00619697
R19091 VPWR.n5653 VPWR.n5652 0.00619697
R19092 VPWR.n5648 VPWR.n5647 0.00619697
R19093 VPWR.n4907 VPWR.n4906 0.00619697
R19094 VPWR.n4902 VPWR.n4901 0.00619697
R19095 VPWR.n7394 VPWR.n7383 0.00619697
R19096 VPWR.n7379 VPWR.n7378 0.00619697
R19097 VPWR.n7173 VPWR.n7172 0.00619697
R19098 VPWR.n7168 VPWR.n7167 0.00619697
R19099 VPWR.n5421 VPWR.n5420 0.00619697
R19100 VPWR.n5416 VPWR.n5415 0.00619697
R19101 VPWR.n7059 VPWR.n7058 0.00619697
R19102 VPWR.n7054 VPWR.n7053 0.00619697
R19103 VPWR.n4853 VPWR.n315 0.00619697
R19104 VPWR.n311 VPWR.n310 0.00619697
R19105 VPWR.n849 VPWR.n848 0.00619697
R19106 VPWR.n844 VPWR.n843 0.00619697
R19107 VPWR.n547 VPWR.n546 0.00619697
R19108 VPWR.n542 VPWR.n541 0.00619697
R19109 VPWR.n731 VPWR.n730 0.00619697
R19110 VPWR.n726 VPWR.n725 0.00619697
R19111 VPWR.n4753 VPWR.n4742 0.00619697
R19112 VPWR.n4738 VPWR.n4737 0.00619697
R19113 VPWR.n4585 VPWR.n4584 0.00619697
R19114 VPWR.n4580 VPWR.n4579 0.00619697
R19115 VPWR.n1006 VPWR.n1005 0.00619697
R19116 VPWR.n1001 VPWR.n1000 0.00619697
R19117 VPWR.n4447 VPWR.n4446 0.00619697
R19118 VPWR.n4452 VPWR.n4451 0.00619697
R19119 VPWR.n3761 VPWR.n3750 0.00619697
R19120 VPWR.n3746 VPWR.n3745 0.00619697
R19121 VPWR.n4313 VPWR.n4312 0.00619697
R19122 VPWR.n4308 VPWR.n4307 0.00619697
R19123 VPWR.n1286 VPWR.n1285 0.00619697
R19124 VPWR.n1291 VPWR.n1290 0.00619697
R19125 VPWR.n4419 VPWR.n4418 0.00619697
R19126 VPWR.n4414 VPWR.n4413 0.00619697
R19127 VPWR.n3985 VPWR.n3974 0.00619697
R19128 VPWR.n3970 VPWR.n3969 0.00619697
R19129 VPWR.n4148 VPWR.n4147 0.00619697
R19130 VPWR.n4143 VPWR.n4142 0.00619697
R19131 VPWR.n1917 VPWR.n1916 0.00619697
R19132 VPWR.n1912 VPWR.n1911 0.00619697
R19133 VPWR.n4269 VPWR.n4268 0.00619697
R19134 VPWR.n4264 VPWR.n4263 0.00619697
R19135 VPWR.n1828 VPWR.n1827 0.00619697
R19136 VPWR.n1823 VPWR.n1822 0.00619697
R19137 VPWR.n2187 VPWR.n2186 0.00619697
R19138 VPWR.n2182 VPWR.n2181 0.00619697
R19139 VPWR.n3731 VPWR.n3721 0.00619697
R19140 VPWR.n1564 VPWR.n1552 0.00619697
R19141 VPWR.n2063 VPWR.n2052 0.00619697
R19142 VPWR.n2048 VPWR.n2047 0.00619697
R19143 VPWR.n5812 VPWR.n5801 0.00619697
R19144 VPWR.n3410 VPWR.n3409 0.00619697
R19145 VPWR.n2287 VPWR.n2285 0.00619697
R19146 VPWR.n2737 VPWR.n2726 0.00619697
R19147 VPWR.n2774 VPWR.n2771 0.00619697
R19148 VPWR.n3520 VPWR.n3510 0.00619697
R19149 VPWR.n2204 VPWR.n2190 0.00619697
R19150 VPWR.n3034 VPWR.n3022 0.00619697
R19151 VPWR.n3016 VPWR.n3005 0.00619697
R19152 VPWR.n3047 VPWR.n3046 0.00619697
R19153 VPWR.n3065 VPWR.n3051 0.00619697
R19154 VPWR.n5782 VPWR.n5771 0.00619697
R19155 VPWR.n2404 VPWR.n2403 0.00619697
R19156 VPWR.n3199 VPWR.n2408 0.00619697
R19157 VPWR.n9 VPWR.n8 0.00619697
R19158 VPWR.n14 VPWR.n13 0.00619697
R19159 VPWR.n7757 VPWR.n7756 0.00619697
R19160 VPWR.n7763 VPWR.n7761 0.00619697
R19161 VPWR.n6376 VPWR.n6375 0.00619697
R19162 VPWR.n5708 VPWR.n5696 0.00619697
R19163 VPWR.n2676 VPWR.n2664 0.00619697
R19164 VPWR.n2660 VPWR.n2659 0.00619697
R19165 VPWR.n3380 VPWR.n3379 0.00619697
R19166 VPWR.n3398 VPWR.n3384 0.00619697
R19167 VPWR.n6019 VPWR.n6010 0.00619697
R19168 VPWR.n6006 VPWR.n6005 0.00619697
R19169 VPWR.n2684 VPWR.n2683 0.00590801
R19170 VPWR.n5675 VPWR 0.00570833
R19171 VPWR.n6682 VPWR.n6681 0.00570833
R19172 VPWR.n6763 VPWR 0.00570833
R19173 VPWR.n7625 VPWR.n7624 0.00570833
R19174 VPWR.n7621 VPWR.n7620 0.00570833
R19175 VPWR.n5482 VPWR.n5481 0.00570833
R19176 VPWR.n6903 VPWR.n6902 0.00570833
R19177 VPWR.n6791 VPWR.n6789 0.00570833
R19178 VPWR.n6793 VPWR 0.00570833
R19179 VPWR.n7039 VPWR.n7026 0.00570833
R19180 VPWR.n7148 VPWR.n7140 0.00570833
R19181 VPWR.n7164 VPWR.n7163 0.00570833
R19182 VPWR VPWR.n7160 0.00570833
R19183 VPWR.n562 VPWR 0.00570833
R19184 VPWR.n974 VPWR 0.00570833
R19185 VPWR.n711 VPWR.n705 0.00570833
R19186 VPWR.n856 VPWR.n823 0.00570833
R19187 VPWR.n840 VPWR.n839 0.00570833
R19188 VPWR VPWR.n4780 0.00570833
R19189 VPWR.n1110 VPWR.n1109 0.00570833
R19190 VPWR.n4593 VPWR.n4592 0.00570833
R19191 VPWR.n4598 VPWR.n4596 0.00570833
R19192 VPWR VPWR.n1296 0.00570833
R19193 VPWR.n1398 VPWR.n1397 0.00570833
R19194 VPWR.n3790 VPWR.n3789 0.00570833
R19195 VPWR.n3795 VPWR.n3793 0.00570833
R19196 VPWR.n4245 VPWR.n4244 0.00570833
R19197 VPWR.n4155 VPWR.n1488 0.00570833
R19198 VPWR.n1513 VPWR.n1511 0.00570833
R19199 VPWR.n1819 VPWR 0.00570833
R19200 VPWR.n2094 VPWR.n2093 0.00570833
R19201 VPWR.n3565 VPWR.n3564 0.00570833
R19202 VPWR.n3570 VPWR.n3568 0.00570833
R19203 VPWR VPWR.n2781 0.00570833
R19204 VPWR.n2839 VPWR.n2838 0.00570833
R19205 VPWR.n3470 VPWR.n3469 0.00570833
R19206 VPWR.n3466 VPWR.n3465 0.00570833
R19207 VPWR VPWR.n2270 0.00570833
R19208 VPWR.n2342 VPWR 0.00570833
R19209 VPWR.n6427 VPWR 0.00570833
R19210 VPWR.n6549 VPWR.n6548 0.00570833
R19211 VPWR.n7770 VPWR.n7745 0.00570833
R19212 VPWR.n7742 VPWR.n7741 0.00570833
R19213 VPWR.n3092 VPWR.n3091 0.00570833
R19214 VPWR.n3182 VPWR.n3181 0.00570833
R19215 VPWR.n3188 VPWR.n3185 0.00570833
R19216 VPWR.n6194 VPWR.n6193 0.00570833
R19217 VPWR.n6096 VPWR.n6095 0.00570833
R19218 VPWR.n6092 VPWR.n6091 0.00570833
R19219 VPWR.n3001 VPWR.n3000 0.005649
R19220 VPWR.n2673 VPWR.n2672 0.00556757
R19221 VPWR.n7644 VPWR.n7643 0.00556757
R19222 VPWR.n7753 VPWR.n7752 0.00556757
R19223 VPWR.n7735 VPWR.n7734 0.00556757
R19224 VPWR.n7733 VPWR.n28 0.00556757
R19225 VPWR.n7501 VPWR.n7500 0.00556757
R19226 VPWR.n7628 VPWR.n7627 0.00556757
R19227 VPWR.n7615 VPWR.n154 0.00556757
R19228 VPWR.n7613 VPWR.n7612 0.00556757
R19229 VPWR.n7606 VPWR.n156 0.00556757
R19230 VPWR.n5084 VPWR.n5083 0.00556757
R19231 VPWR.n6594 VPWR.n6593 0.00556757
R19232 VPWR.n6598 VPWR.n6597 0.00556757
R19233 VPWR.n6577 VPWR.n6576 0.00556757
R19234 VPWR.n7403 VPWR.n7402 0.00556757
R19235 VPWR.n6887 VPWR.n6886 0.00556757
R19236 VPWR.n6783 VPWR.n6782 0.00556757
R19237 VPWR.n6874 VPWR.n6785 0.00556757
R19238 VPWR.n6873 VPWR.n6787 0.00556757
R19239 VPWR.n5638 VPWR.n5637 0.00556757
R19240 VPWR.n7001 VPWR.n7000 0.00556757
R19241 VPWR.n7005 VPWR.n7004 0.00556757
R19242 VPWR.n4895 VPWR.n4894 0.00556757
R19243 VPWR.n7179 VPWR.n7176 0.00556757
R19244 VPWR.n7158 VPWR.n7156 0.00556757
R19245 VPWR.n7206 VPWR.n294 0.00556757
R19246 VPWR.n7209 VPWR.n7208 0.00556757
R19247 VPWR.n5406 VPWR.n5405 0.00556757
R19248 VPWR.n5327 VPWR.n5326 0.00556757
R19249 VPWR.n5297 VPWR.n5289 0.00556757
R19250 VPWR.n5296 VPWR.n5292 0.00556757
R19251 VPWR.n7047 VPWR.n7046 0.00556757
R19252 VPWR.n4762 VPWR.n4761 0.00556757
R19253 VPWR.n853 VPWR.n852 0.00556757
R19254 VPWR.n591 VPWR.n590 0.00556757
R19255 VPWR.n879 VPWR.n593 0.00556757
R19256 VPWR.n882 VPWR.n881 0.00556757
R19257 VPWR.n551 VPWR.n550 0.00556757
R19258 VPWR.n975 VPWR.n469 0.00556757
R19259 VPWR.n618 VPWR.n617 0.00556757
R19260 VPWR.n622 VPWR.n621 0.00556757
R19261 VPWR.n635 VPWR.n634 0.00556757
R19262 VPWR.n4685 VPWR.n4684 0.00556757
R19263 VPWR.n4589 VPWR.n4588 0.00556757
R19264 VPWR.n4561 VPWR.n4560 0.00556757
R19265 VPWR.n4567 VPWR.n4563 0.00556757
R19266 VPWR.n4566 VPWR.n4565 0.00556757
R19267 VPWR.n991 VPWR.n990 0.00556757
R19268 VPWR.n1207 VPWR.n1206 0.00556757
R19269 VPWR.n4427 VPWR.n4426 0.00556757
R19270 VPWR.n4431 VPWR.n4430 0.00556757
R19271 VPWR.n408 VPWR.n407 0.00556757
R19272 VPWR.n3786 VPWR.n3782 0.00556757
R19273 VPWR.n4289 VPWR.n4288 0.00556757
R19274 VPWR.n4295 VPWR.n4291 0.00556757
R19275 VPWR.n4294 VPWR.n4293 0.00556757
R19276 VPWR.n457 VPWR.n456 0.00556757
R19277 VPWR.n1416 VPWR.n1408 0.00556757
R19278 VPWR.n1415 VPWR.n1411 0.00556757
R19279 VPWR.n4407 VPWR.n4406 0.00556757
R19280 VPWR.n4057 VPWR.n4056 0.00556757
R19281 VPWR.n4152 VPWR.n4151 0.00556757
R19282 VPWR.n1518 VPWR.n1516 0.00556757
R19283 VPWR.n4130 VPWR.n1506 0.00556757
R19284 VPWR.n4129 VPWR.n1508 0.00556757
R19285 VPWR.n1921 VPWR.n1920 0.00556757
R19286 VPWR.n2029 VPWR.n1640 0.00556757
R19287 VPWR.n2033 VPWR.n2032 0.00556757
R19288 VPWR.n4257 VPWR.n4256 0.00556757
R19289 VPWR.n1666 VPWR.n1665 0.00556757
R19290 VPWR.n2171 VPWR.n2170 0.00556757
R19291 VPWR.n3530 VPWR.n3529 0.00556757
R19292 VPWR.n3536 VPWR.n3532 0.00556757
R19293 VPWR.n3535 VPWR.n3534 0.00556757
R19294 VPWR.n1556 VPWR.n1555 0.00556757
R19295 VPWR.n2106 VPWR.n2105 0.00556757
R19296 VPWR.n1591 VPWR.n1590 0.00556757
R19297 VPWR.n2041 VPWR.n2040 0.00556757
R19298 VPWR.n4951 VPWR.n4950 0.00556757
R19299 VPWR.n4955 VPWR.n4954 0.00556757
R19300 VPWR.n4961 VPWR.n4960 0.00556757
R19301 VPWR.n2351 VPWR.n2343 0.00556757
R19302 VPWR.n2734 VPWR.n2733 0.00556757
R19303 VPWR.n2995 VPWR.n2689 0.00556757
R19304 VPWR.n3517 VPWR.n3516 0.00556757
R19305 VPWR.n2199 VPWR.n2198 0.00556757
R19306 VPWR.n3501 VPWR.n3497 0.00556757
R19307 VPWR.n3500 VPWR.n3499 0.00556757
R19308 VPWR.n2478 VPWR.n2477 0.00556757
R19309 VPWR.n2481 VPWR.n2480 0.00556757
R19310 VPWR.n3024 VPWR.n3023 0.00556757
R19311 VPWR.n3007 VPWR.n3006 0.00556757
R19312 VPWR.n2464 VPWR.n2463 0.00556757
R19313 VPWR.n2469 VPWR.n2468 0.00556757
R19314 VPWR.n2466 VPWR.n2465 0.00556757
R19315 VPWR.n3055 VPWR.n3054 0.00556757
R19316 VPWR.n5786 VPWR.n5785 0.00556757
R19317 VPWR.n5790 VPWR.n5789 0.00556757
R19318 VPWR.n5755 VPWR.n5754 0.00556757
R19319 VPWR.n2400 VPWR.n2399 0.00556757
R19320 VPWR.n3204 VPWR.n2389 0.00556757
R19321 VPWR.n3207 VPWR.n3206 0.00556757
R19322 VPWR.n6073 VPWR.n6072 0.00556757
R19323 VPWR.n6062 VPWR.n6061 0.00556757
R19324 VPWR.n7803 VPWR.n2 0.00556757
R19325 VPWR.n7806 VPWR.n7805 0.00556757
R19326 VPWR.n6368 VPWR.n6367 0.00556757
R19327 VPWR.n5705 VPWR.n5704 0.00556757
R19328 VPWR.n3388 VPWR.n3387 0.00556757
R19329 VPWR.n6000 VPWR.n5999 0.00556757
R19330 VPWR.n2491 VPWR.n2490 0.00554564
R19331 VPWR.n6701 VPWR.n6699 0.00548035
R19332 VPWR.n5494 VPWR.n5493 0.00548035
R19333 VPWR.n1421 VPWR.n1419 0.00548035
R19334 VPWR.n2393 VPWR.n2205 0.00500002
R19335 VPWR.n3522 VPWR.n3521 0.00500002
R19336 VPWR.n3405 VPWR.n2284 0.00500002
R19337 VPWR.n3036 VPWR.n3035 0.00495986
R19338 VPWR.n6870 VPWR.n6869 0.00484057
R19339 VPWR.n7215 VPWR.n7212 0.00484057
R19340 VPWR.n886 VPWR.n885 0.00484057
R19341 VPWR.n3804 VPWR.n3802 0.00484057
R19342 VPWR.n5835 VPWR.n5833 0.00484057
R19343 VPWR.n2280 VPWR.n2279 0.00477273
R19344 VPWR.n2741 VPWR.n2740 0.00477273
R19345 VPWR.n5783 VPWR.n5764 0.00460158
R19346 VPWR.n5814 VPWR.n5813 0.00460158
R19347 VPWR.n6575 VPWR.n6574 0.00460158
R19348 VPWR.n6588 VPWR.n4908 0.00460158
R19349 VPWR.n7060 VPWR.n7009 0.00460158
R19350 VPWR.n732 VPWR.n626 0.00460158
R19351 VPWR.n4445 VPWR.n417 0.00460158
R19352 VPWR.n4421 VPWR.n4420 0.00460158
R19353 VPWR.n4271 VPWR.n4270 0.00460158
R19354 VPWR.n2064 VPWR.n2037 0.00460158
R19355 VPWR.n3066 VPWR.n3038 0.00460158
R19356 VPWR.n19 VPWR.n18 0.00460158
R19357 VPWR.n2188 VPWR.n2160 0.00460158
R19358 VPWR.n3200 VPWR.n2395 0.00460158
R19359 VPWR.n5709 VPWR.n5689 0.00460158
R19360 VPWR.n6377 VPWR.n6357 0.00460158
R19361 VPWR.n5686 VPWR.n5685 0.00460158
R19362 VPWR.n5655 VPWR.n5654 0.00460158
R19363 VPWR.n5423 VPWR.n5422 0.00460158
R19364 VPWR.n540 VPWR.n539 0.00460158
R19365 VPWR.n1007 VPWR.n980 0.00460158
R19366 VPWR.n1284 VPWR.n1212 0.00460158
R19367 VPWR.n1904 VPWR.n1654 0.00460158
R19368 VPWR.n1830 VPWR.n1829 0.00460158
R19369 VPWR.n5915 VPWR.n5910 0.00460158
R19370 VPWR.n5911 VPWR.n127 0.00460158
R19371 VPWR.n255 VPWR.n128 0.00460158
R19372 VPWR.n3400 VPWR.n3399 0.00460158
R19373 VPWR.n7512 VPWR.n7497 0.00460158
R19374 VPWR.n7655 VPWR.n7638 0.00460158
R19375 VPWR.n5132 VPWR.n5131 0.00440625
R19376 VPWR.n6698 VPWR.n6697 0.00440625
R19377 VPWR.n6695 VPWR.n6694 0.00440625
R19378 VPWR.n6607 VPWR.n4942 0.00440625
R19379 VPWR.n6756 VPWR.n6754 0.00440625
R19380 VPWR.n6752 VPWR.n153 0.00440625
R19381 VPWR.n7617 VPWR.n7616 0.00440625
R19382 VPWR.n7605 VPWR.n7604 0.00440625
R19383 VPWR.n224 VPWR.n223 0.00440625
R19384 VPWR VPWR.n234 0.00440625
R19385 VPWR.n5609 VPWR.n5608 0.00440625
R19386 VPWR.n5492 VPWR.n5491 0.00440625
R19387 VPWR.n5489 VPWR.n5488 0.00440625
R19388 VPWR.n5480 VPWR.n5479 0.00440625
R19389 VPWR.n6905 VPWR.n6904 0.00440625
R19390 VPWR.n6794 VPWR.n6793 0.00440625
R19391 VPWR.n6872 VPWR.n6871 0.00440625
R19392 VPWR.n278 VPWR.n276 0.00440625
R19393 VPWR.n7487 VPWR.n7486 0.00440625
R19394 VPWR.n7477 VPWR 0.00440625
R19395 VPWR.n5391 VPWR.n5216 0.00440625
R19396 VPWR.n5328 VPWR.n5217 0.00440625
R19397 VPWR.n5299 VPWR.n5298 0.00440625
R19398 VPWR.n7017 VPWR.n7016 0.00440625
R19399 VPWR.n7038 VPWR.n7037 0.00440625
R19400 VPWR.n7183 VPWR.n7182 0.00440625
R19401 VPWR.n7181 VPWR 0.00440625
R19402 VPWR.n7160 VPWR.n7159 0.00440625
R19403 VPWR.n7211 VPWR.n7210 0.00440625
R19404 VPWR.n7315 VPWR.n7313 0.00440625
R19405 VPWR.n530 VPWR.n529 0.00440625
R19406 VPWR.n974 VPWR.n973 0.00440625
R19407 VPWR.n690 VPWR.n689 0.00440625
R19408 VPWR.n693 VPWR.n692 0.00440625
R19409 VPWR.n713 VPWR.n712 0.00440625
R19410 VPWR.n858 VPWR.n857 0.00440625
R19411 VPWR.n588 VPWR.n587 0.00440625
R19412 VPWR.n884 VPWR.n883 0.00440625
R19413 VPWR.n323 VPWR.n318 0.00440625
R19414 VPWR.n4846 VPWR.n4845 0.00440625
R19415 VPWR.n1066 VPWR.n1065 0.00440625
R19416 VPWR.n1088 VPWR.n1087 0.00440625
R19417 VPWR.n1121 VPWR.n1120 0.00440625
R19418 VPWR.n1118 VPWR.n1117 0.00440625
R19419 VPWR.n1103 VPWR.n1102 0.00440625
R19420 VPWR VPWR.n4457 0.00440625
R19421 VPWR.n4538 VPWR.n4536 0.00440625
R19422 VPWR.n4534 VPWR.n379 0.00440625
R19423 VPWR.n4601 VPWR.n4600 0.00440625
R19424 VPWR.n4604 VPWR.n4603 0.00440625
R19425 VPWR.n4690 VPWR.n4689 0.00440625
R19426 VPWR.n4712 VPWR.n4711 0.00440625
R19427 VPWR.n1266 VPWR.n1265 0.00440625
R19428 VPWR.n1418 VPWR.n1417 0.00440625
R19429 VPWR.n1405 VPWR.n1404 0.00440625
R19430 VPWR.n1396 VPWR.n1395 0.00440625
R19431 VPWR.n1441 VPWR.n1439 0.00440625
R19432 VPWR.n3785 VPWR.n3784 0.00440625
R19433 VPWR.n3798 VPWR.n3797 0.00440625
R19434 VPWR.n3801 VPWR.n3800 0.00440625
R19435 VPWR.n3933 VPWR.n3932 0.00440625
R19436 VPWR.n1883 VPWR.n1650 0.00440625
R19437 VPWR.n2026 VPWR.n2025 0.00440625
R19438 VPWR.n4243 VPWR.n4242 0.00440625
R19439 VPWR.n4162 VPWR.n4160 0.00440625
R19440 VPWR.n4158 VPWR.n4156 0.00440625
R19441 VPWR VPWR.n1515 0.00440625
R19442 VPWR.n4128 VPWR.n4127 0.00440625
R19443 VPWR.n4062 VPWR.n4061 0.00440625
R19444 VPWR.n4039 VPWR.n4038 0.00440625
R19445 VPWR.n1724 VPWR.n1723 0.00440625
R19446 VPWR.n2104 VPWR.n1592 0.00440625
R19447 VPWR.n2102 VPWR.n2101 0.00440625
R19448 VPWR.n2092 VPWR.n2091 0.00440625
R19449 VPWR.n3560 VPWR.n3558 0.00440625
R19450 VPWR.n3563 VPWR.n3562 0.00440625
R19451 VPWR.n3573 VPWR.n3572 0.00440625
R19452 VPWR.n3576 VPWR.n3575 0.00440625
R19453 VPWR.n3694 VPWR.n3693 0.00440625
R19454 VPWR.n2756 VPWR.n2755 0.00440625
R19455 VPWR.n2828 VPWR.n2827 0.00440625
R19456 VPWR.n2831 VPWR.n2830 0.00440625
R19457 VPWR.n2841 VPWR.n2840 0.00440625
R19458 VPWR.n3477 VPWR.n3475 0.00440625
R19459 VPWR.n3473 VPWR.n3471 0.00440625
R19460 VPWR.n3462 VPWR.n3461 0.00440625
R19461 VPWR.n3459 VPWR.n3458 0.00440625
R19462 VPWR.n2352 VPWR.n2342 0.00440625
R19463 VPWR.n6437 VPWR.n6436 0.00440625
R19464 VPWR.n6537 VPWR.n6536 0.00440625
R19465 VPWR.n6540 VPWR.n6539 0.00440625
R19466 VPWR.n6552 VPWR.n6550 0.00440625
R19467 VPWR.n7772 VPWR.n7771 0.00440625
R19468 VPWR.n7738 VPWR 0.00440625
R19469 VPWR.n7732 VPWR.n7731 0.00440625
R19470 VPWR.n92 VPWR.n91 0.00440625
R19471 VPWR.n2626 VPWR.n2625 0.00440625
R19472 VPWR.n3103 VPWR.n3102 0.00440625
R19473 VPWR.n3100 VPWR.n3099 0.00440625
R19474 VPWR.n3090 VPWR.n3089 0.00440625
R19475 VPWR.n3178 VPWR.n3177 0.00440625
R19476 VPWR.n3180 VPWR.n3179 0.00440625
R19477 VPWR.n3191 VPWR.n3190 0.00440625
R19478 VPWR.n3209 VPWR.n3208 0.00440625
R19479 VPWR.n3342 VPWR.n3341 0.00440625
R19480 VPWR.n6329 VPWR.n6328 0.00440625
R19481 VPWR.n6205 VPWR.n6204 0.00440625
R19482 VPWR.n6202 VPWR.n6201 0.00440625
R19483 VPWR.n6192 VPWR.n6191 0.00440625
R19484 VPWR.n6100 VPWR.n6099 0.00440625
R19485 VPWR.n6098 VPWR.n6097 0.00440625
R19486 VPWR.n6086 VPWR.n0 0.00440625
R19487 VPWR.n7807 VPWR.n1 0.00440625
R19488 VPWR.n5979 VPWR.n5978 0.00440625
R19489 VPWR VPWR.n5989 0.00440625
R19490 VPWR.n6766 VPWR.n4934 0.00406061
R19491 VPWR.n5659 VPWR.n5658 0.00406061
R19492 VPWR.n6599 VPWR.n6590 0.00406061
R19493 VPWR.n7400 VPWR.n283 0.00406061
R19494 VPWR.n6777 VPWR.n6772 0.00406061
R19495 VPWR.n5583 VPWR.n5582 0.00406061
R19496 VPWR.n7006 VPWR.n6997 0.00406061
R19497 VPWR.n7294 VPWR.n7290 0.00406061
R19498 VPWR.n7201 VPWR.n4861 0.00406061
R19499 VPWR.n5228 VPWR.n5227 0.00406061
R19500 VPWR.n5295 VPWR.n5293 0.00406061
R19501 VPWR.n4759 VPWR.n328 0.00406061
R19502 VPWR.n874 VPWR.n599 0.00406061
R19503 VPWR.n977 VPWR.n464 0.00406061
R19504 VPWR.n623 VPWR.n614 0.00406061
R19505 VPWR.n4682 VPWR.n4680 0.00406061
R19506 VPWR.n4555 VPWR.n389 0.00406061
R19507 VPWR.n1209 VPWR.n1012 0.00406061
R19508 VPWR.n4432 VPWR.n4423 0.00406061
R19509 VPWR.n3956 VPWR.n3774 0.00406061
R19510 VPWR.n4283 VPWR.n4278 0.00406061
R19511 VPWR.n1223 VPWR.n1217 0.00406061
R19512 VPWR.n1414 VPWR.n1412 0.00406061
R19513 VPWR.n4054 VPWR.n1543 0.00406061
R19514 VPWR.n1501 VPWR.n1496 0.00406061
R19515 VPWR.n1841 VPWR.n1835 0.00406061
R19516 VPWR.n2034 VPWR.n1637 0.00406061
R19517 VPWR.n1809 VPWR.n1808 0.00406061
R19518 VPWR.n3537 VPWR.n3528 0.00406061
R19519 VPWR.n2072 VPWR.n2071 0.00406061
R19520 VPWR.n6570 VPWR.n4970 0.00406061
R19521 VPWR.n2278 VPWR.n2274 0.00406061
R19522 VPWR.n2363 VPWR.n2288 0.00406061
R19523 VPWR.n2997 VPWR.n2686 0.00406061
R19524 VPWR.n3492 VPWR.n2207 0.00406061
R19525 VPWR.n3502 VPWR.n3495 0.00406061
R19526 VPWR.n2811 VPWR.n2810 0.00406061
R19527 VPWR.n2470 VPWR.n2458 0.00406061
R19528 VPWR.n5818 VPWR.n5817 0.00406061
R19529 VPWR.n3160 VPWR.n3156 0.00406061
R19530 VPWR.n7802 VPWR.n7801 0.00406061
R19531 VPWR.n24 VPWR.n23 0.00406061
R19532 VPWR.n6455 VPWR.n6454 0.00406061
R19533 VPWR.n6354 VPWR.n5726 0.00406061
R19534 VPWR.n2498 VPWR.n2492 0.00406061
R19535 VPWR.n3370 VPWR.n2379 0.00406061
R19536 VPWR.n5993 VPWR.n5916 0.00406061
R19537 VPWR.n6600 VPWR.n6589 0.00393497
R19538 VPWR.n7008 VPWR.n7007 0.00393497
R19539 VPWR.n4881 VPWR.n4880 0.00393497
R19540 VPWR.n624 VPWR.n613 0.00393497
R19541 VPWR.n4433 VPWR.n4422 0.00393497
R19542 VPWR.n419 VPWR.n418 0.00393497
R19543 VPWR.n2036 VPWR.n2035 0.00393497
R19544 VPWR.n5816 VPWR.n5815 0.00393497
R19545 VPWR.n2471 VPWR.n2457 0.00393497
R19546 VPWR.n6572 VPWR.n6571 0.00393497
R19547 VPWR.n2070 VPWR.n2069 0.00393497
R19548 VPWR.n130 VPWR.n25 0.00393497
R19549 VPWR.n7633 VPWR.n7632 0.00393497
R19550 VPWR.n6768 VPWR.n6767 0.00393497
R19551 VPWR.n6878 VPWR.n6769 0.00393497
R19552 VPWR.n6778 VPWR.n6771 0.00393497
R19553 VPWR.n6770 VPWR.n298 0.00393497
R19554 VPWR.n7202 VPWR.n4860 0.00393497
R19555 VPWR.n597 VPWR.n299 0.00393497
R19556 VPWR.n875 VPWR.n598 0.00393497
R19557 VPWR.n4571 VPWR.n387 0.00393497
R19558 VPWR.n4556 VPWR.n388 0.00393497
R19559 VPWR.n4299 VPWR.n1450 0.00393497
R19560 VPWR.n4284 VPWR.n4277 0.00393497
R19561 VPWR.n4134 VPWR.n1451 0.00393497
R19562 VPWR.n2159 VPWR.n1502 0.00393497
R19563 VPWR.n3538 VPWR.n3524 0.00393497
R19564 VPWR.n7800 VPWR.n7799 0.00393497
R19565 VPWR.n2392 VPWR.n2391 0.00393497
R19566 VPWR.n7798 VPWR.n7797 0.00393497
R19567 VPWR.n6453 VPWR.n5688 0.00393497
R19568 VPWR.n5657 VPWR.n5656 0.00393497
R19569 VPWR.n5425 VPWR.n5424 0.00393497
R19570 VPWR.n5226 VPWR.n5225 0.00393497
R19571 VPWR.n979 VPWR.n978 0.00393497
R19572 VPWR.n1211 VPWR.n1210 0.00393497
R19573 VPWR.n1224 VPWR.n1213 0.00393497
R19574 VPWR.n1842 VPWR.n1831 0.00393497
R19575 VPWR.n1807 VPWR.n1806 0.00393497
R19576 VPWR.n2678 VPWR.n2677 0.00393497
R19577 VPWR.n6356 VPWR.n6355 0.00393497
R19578 VPWR.n2681 VPWR.n2680 0.00393497
R19579 VPWR.n7496 VPWR.n7495 0.00393497
R19580 VPWR.n7398 VPWR.n7397 0.00393497
R19581 VPWR.n7396 VPWR.n7395 0.00393497
R19582 VPWR.n7292 VPWR.n7291 0.00393497
R19583 VPWR.n4855 VPWR.n4854 0.00393497
R19584 VPWR.n4757 VPWR.n4756 0.00393497
R19585 VPWR.n4755 VPWR.n4754 0.00393497
R19586 VPWR.n3735 VPWR.n329 0.00393497
R19587 VPWR.n3762 VPWR.n3736 0.00393497
R19588 VPWR.n3958 VPWR.n3957 0.00393497
R19589 VPWR.n3986 VPWR.n3960 0.00393497
R19590 VPWR.n4052 VPWR.n3734 0.00393497
R19591 VPWR.n1565 VPWR.n1550 0.00393497
R19592 VPWR.n3371 VPWR.n2378 0.00393497
R19593 VPWR.n3733 VPWR.n3732 0.00393497
R19594 VPWR.n2666 VPWR.n2665 0.00387838
R19595 VPWR.n2669 VPWR.n2668 0.00387838
R19596 VPWR.n120 VPWR.n119 0.00387838
R19597 VPWR.n7650 VPWR.n7649 0.00387838
R19598 VPWR.n7647 VPWR.n7646 0.00387838
R19599 VPWR.n244 VPWR.n243 0.00387838
R19600 VPWR.n7507 VPWR.n7506 0.00387838
R19601 VPWR.n7504 VPWR.n7503 0.00387838
R19602 VPWR.n5077 VPWR.n5076 0.00387838
R19603 VPWR.n5080 VPWR.n5079 0.00387838
R19604 VPWR.n5090 VPWR.n5089 0.00387838
R19605 VPWR.n6657 VPWR.n6656 0.00387838
R19606 VPWR.n273 VPWR.n272 0.00387838
R19607 VPWR.n263 VPWR.n262 0.00387838
R19608 VPWR.n7428 VPWR.n7427 0.00387838
R19609 VPWR.n5631 VPWR.n5630 0.00387838
R19610 VPWR.n5634 VPWR.n5633 0.00387838
R19611 VPWR.n5644 VPWR.n5643 0.00387838
R19612 VPWR.n7386 VPWR.n7385 0.00387838
R19613 VPWR.n7376 VPWR.n7375 0.00387838
R19614 VPWR.n7318 VPWR.n7317 0.00387838
R19615 VPWR.n5395 VPWR.n5394 0.00387838
R19616 VPWR.n5396 VPWR.n5214 0.00387838
R19617 VPWR.n5412 VPWR.n5411 0.00387838
R19618 VPWR.n7067 VPWR.n7066 0.00387838
R19619 VPWR.n4778 VPWR.n4777 0.00387838
R19620 VPWR.n308 VPWR.n307 0.00387838
R19621 VPWR.n4788 VPWR.n4787 0.00387838
R19622 VPWR.n532 VPWR.n531 0.00387838
R19623 VPWR.n535 VPWR.n534 0.00387838
R19624 VPWR.n565 VPWR.n564 0.00387838
R19625 VPWR.n739 VPWR.n738 0.00387838
R19626 VPWR.n4745 VPWR.n4744 0.00387838
R19627 VPWR.n4735 VPWR.n4734 0.00387838
R19628 VPWR.n334 VPWR.n333 0.00387838
R19629 VPWR.n984 VPWR.n983 0.00387838
R19630 VPWR.n987 VPWR.n986 0.00387838
R19631 VPWR.n997 VPWR.n996 0.00387838
R19632 VPWR.n3753 VPWR.n3752 0.00387838
R19633 VPWR.n3743 VPWR.n3742 0.00387838
R19634 VPWR.n3767 VPWR.n3766 0.00387838
R19635 VPWR.n450 VPWR.n449 0.00387838
R19636 VPWR.n453 VPWR.n452 0.00387838
R19637 VPWR.n1294 VPWR.n1293 0.00387838
R19638 VPWR.n3977 VPWR.n3976 0.00387838
R19639 VPWR.n3967 VPWR.n3966 0.00387838
R19640 VPWR.n3991 VPWR.n3990 0.00387838
R19641 VPWR.n1887 VPWR.n1886 0.00387838
R19642 VPWR.n1888 VPWR.n1651 0.00387838
R19643 VPWR.n1908 VPWR.n1907 0.00387838
R19644 VPWR.n1659 VPWR.n1658 0.00387838
R19645 VPWR.n1662 VPWR.n1661 0.00387838
R19646 VPWR.n1672 VPWR.n1671 0.00387838
R19647 VPWR.n3724 VPWR.n3723 0.00387838
R19648 VPWR.n1562 VPWR.n1561 0.00387838
R19649 VPWR.n1559 VPWR.n1558 0.00387838
R19650 VPWR.n3414 VPWR.n3413 0.00387838
R19651 VPWR.n2348 VPWR.n2347 0.00387838
R19652 VPWR.n2345 VPWR.n2344 0.00387838
R19653 VPWR.n2729 VPWR.n2728 0.00387838
R19654 VPWR.n2732 VPWR.n2731 0.00387838
R19655 VPWR.n2779 VPWR.n2778 0.00387838
R19656 VPWR.n6361 VPWR.n6360 0.00387838
R19657 VPWR.n6364 VPWR.n6363 0.00387838
R19658 VPWR.n5698 VPWR.n5697 0.00387838
R19659 VPWR.n5701 VPWR.n5700 0.00387838
R19660 VPWR.n3374 VPWR.n3373 0.00387838
R19661 VPWR.n3394 VPWR.n3393 0.00387838
R19662 VPWR.n3391 VPWR.n3390 0.00387838
R19663 VPWR.n6014 VPWR.n6013 0.00387838
R19664 VPWR.n6003 VPWR.n6002 0.00387838
R19665 VPWR.n5919 VPWR.n5918 0.00387838
R19666 VPWR.n2742 VPWR.n2724 0.0033671
R19667 VPWR.n2482 VPWR.n2475 0.0033671
R19668 VPWR.n3017 VPWR.n2474 0.0032017
R19669 VPWR.n2474 VPWR.n2473 0.0032017
R19670 VPWR.n5913 VPWR.n5912 0.0032017
R19671 VPWR.n3404 VPWR.n3403 0.0032017
R19672 VPWR.n3403 VPWR.n3402 0.0032017
R19673 VPWR.n5914 VPWR.n5913 0.0032017
R19674 VPWR.n5126 VPWR.n5125 0.00310417
R19675 VPWR.n5127 VPWR.n5126 0.00310417
R19676 VPWR.n5130 VPWR.n5129 0.00310417
R19677 VPWR.n5674 VPWR.n5673 0.00310417
R19678 VPWR.n6609 VPWR.n6608 0.00310417
R19679 VPWR.n6664 VPWR 0.00310417
R19680 VPWR.n6605 VPWR.n6580 0.00310417
R19681 VPWR.n6750 VPWR.n6749 0.00310417
R19682 VPWR VPWR.n6762 0.00310417
R19683 VPWR.n7602 VPWR.n7601 0.00310417
R19684 VPWR.n213 VPWR.n212 0.00310417
R19685 VPWR.n221 VPWR.n218 0.00310417
R19686 VPWR.n226 VPWR.n225 0.00310417
R19687 VPWR.n231 VPWR.n230 0.00310417
R19688 VPWR.n5617 VPWR.n5616 0.00310417
R19689 VPWR.n5616 VPWR.n5615 0.00310417
R19690 VPWR.n5611 VPWR.n5610 0.00310417
R19691 VPWR.n5598 VPWR.n5597 0.00310417
R19692 VPWR.n6918 VPWR.n6917 0.00310417
R19693 VPWR.n7418 VPWR.n7417 0.00310417
R19694 VPWR.n7426 VPWR.n7423 0.00310417
R19695 VPWR.n7485 VPWR.n7484 0.00310417
R19696 VPWR.n7482 VPWR.n7479 0.00310417
R19697 VPWR.n5390 VPWR.n5389 0.00310417
R19698 VPWR.n5398 VPWR.n5390 0.00310417
R19699 VPWR.n5393 VPWR.n5392 0.00310417
R19700 VPWR.n5339 VPWR.n5338 0.00310417
R19701 VPWR.n5324 VPWR 0.00310417
R19702 VPWR.n7024 VPWR 0.00310417
R19703 VPWR.n7028 VPWR.n7027 0.00310417
R19704 VPWR.n7195 VPWR.n7190 0.00310417
R19705 VPWR.n7303 VPWR.n7302 0.00310417
R19706 VPWR.n7311 VPWR.n7309 0.00310417
R19707 VPWR.n7374 VPWR.n7316 0.00310417
R19708 VPWR.n7372 VPWR.n7370 0.00310417
R19709 VPWR.n518 VPWR 0.00310417
R19710 VPWR.n522 VPWR.n521 0.00310417
R19711 VPWR.n525 VPWR.n522 0.00310417
R19712 VPWR.n528 VPWR.n527 0.00310417
R19713 VPWR.n566 VPWR.n471 0.00310417
R19714 VPWR VPWR.n971 0.00310417
R19715 VPWR.n715 VPWR.n714 0.00310417
R19716 VPWR.n721 VPWR 0.00310417
R19717 VPWR.n742 VPWR.n741 0.00310417
R19718 VPWR.n868 VPWR.n866 0.00310417
R19719 VPWR.n4780 VPWR.n4779 0.00310417
R19720 VPWR.n4844 VPWR.n4843 0.00310417
R19721 VPWR.n4841 VPWR.n4839 0.00310417
R19722 VPWR.n1059 VPWR.n1058 0.00310417
R19723 VPWR.n1061 VPWR.n1059 0.00310417
R19724 VPWR.n1064 VPWR.n1063 0.00310417
R19725 VPWR.n1077 VPWR.n1076 0.00310417
R19726 VPWR.n1204 VPWR 0.00310417
R19727 VPWR.n1100 VPWR.n402 0.00310417
R19728 VPWR.n4549 VPWR.n4546 0.00310417
R19729 VPWR VPWR.n4544 0.00310417
R19730 VPWR.n4609 VPWR.n4608 0.00310417
R19731 VPWR.n4701 VPWR.n4700 0.00310417
R19732 VPWR.n4709 VPWR.n4706 0.00310417
R19733 VPWR.n4714 VPWR.n4713 0.00310417
R19734 VPWR.n4718 VPWR.n4717 0.00310417
R19735 VPWR.n1274 VPWR.n1273 0.00310417
R19736 VPWR.n1273 VPWR.n1272 0.00310417
R19737 VPWR.n1268 VPWR.n1267 0.00310417
R19738 VPWR.n1298 VPWR.n1297 0.00310417
R19739 VPWR.n1393 VPWR.n1391 0.00310417
R19740 VPWR.n4324 VPWR.n4322 0.00310417
R19741 VPWR VPWR.n4320 0.00310417
R19742 VPWR.n3944 VPWR.n3943 0.00310417
R19743 VPWR.n3938 VPWR.n3937 0.00310417
R19744 VPWR.n3931 VPWR.n3930 0.00310417
R19745 VPWR.n3928 VPWR.n3927 0.00310417
R19746 VPWR.n1894 VPWR.n1893 0.00310417
R19747 VPWR.n1893 VPWR.n1892 0.00310417
R19748 VPWR.n1885 VPWR.n1884 0.00310417
R19749 VPWR.n1934 VPWR.n1933 0.00310417
R19750 VPWR VPWR.n2023 0.00310417
R19751 VPWR.n4171 VPWR.n4170 0.00310417
R19752 VPWR VPWR.n4168 0.00310417
R19753 VPWR.n4124 VPWR.n4122 0.00310417
R19754 VPWR.n4031 VPWR.n4030 0.00310417
R19755 VPWR.n4041 VPWR.n4040 0.00310417
R19756 VPWR.n4044 VPWR.n4043 0.00310417
R19757 VPWR.n1719 VPWR.n1718 0.00310417
R19758 VPWR.n1722 VPWR.n1721 0.00310417
R19759 VPWR.n1818 VPWR.n1817 0.00310417
R19760 VPWR.n2089 VPWR.n2087 0.00310417
R19761 VPWR.n3549 VPWR.n3548 0.00310417
R19762 VPWR.n3581 VPWR.n3580 0.00310417
R19763 VPWR.n3702 VPWR.n3701 0.00310417
R19764 VPWR.n3697 VPWR.n3696 0.00310417
R19765 VPWR.n3692 VPWR.n3691 0.00310417
R19766 VPWR.n3689 VPWR.n3686 0.00310417
R19767 VPWR.n2748 VPWR.n2747 0.00310417
R19768 VPWR.n2751 VPWR.n2748 0.00310417
R19769 VPWR.n2754 VPWR.n2753 0.00310417
R19770 VPWR.n2783 VPWR.n2782 0.00310417
R19771 VPWR.n2994 VPWR 0.00310417
R19772 VPWR VPWR.n2991 0.00310417
R19773 VPWR.n3486 VPWR.n3485 0.00310417
R19774 VPWR.n3455 VPWR.n3453 0.00310417
R19775 VPWR.n3415 VPWR.n2270 0.00310417
R19776 VPWR.n2337 VPWR.n2334 0.00310417
R19777 VPWR.n2354 VPWR.n2353 0.00310417
R19778 VPWR.n2357 VPWR.n2356 0.00310417
R19779 VPWR.n6443 VPWR.n6442 0.00310417
R19780 VPWR.n6442 VPWR.n6441 0.00310417
R19781 VPWR.n6439 VPWR.n6438 0.00310417
R19782 VPWR.n6418 VPWR.n6417 0.00310417
R19783 VPWR.n6556 VPWR.n6554 0.00310417
R19784 VPWR.n7782 VPWR.n7781 0.00310417
R19785 VPWR VPWR.n7779 0.00310417
R19786 VPWR.n7728 VPWR.n7726 0.00310417
R19787 VPWR.n100 VPWR.n99 0.00310417
R19788 VPWR.n95 VPWR.n94 0.00310417
R19789 VPWR.n90 VPWR.n89 0.00310417
R19790 VPWR.n87 VPWR.n84 0.00310417
R19791 VPWR.n2619 VPWR.n2618 0.00310417
R19792 VPWR.n2621 VPWR.n2619 0.00310417
R19793 VPWR.n2624 VPWR.n2623 0.00310417
R19794 VPWR.n2637 VPWR.n2636 0.00310417
R19795 VPWR.n3087 VPWR.n3085 0.00310417
R19796 VPWR.n3170 VPWR.n3169 0.00310417
R19797 VPWR.n3214 VPWR.n3213 0.00310417
R19798 VPWR.n3353 VPWR.n3352 0.00310417
R19799 VPWR.n3347 VPWR.n3346 0.00310417
R19800 VPWR.n3340 VPWR.n3339 0.00310417
R19801 VPWR.n3337 VPWR.n3334 0.00310417
R19802 VPWR.n6322 VPWR.n6321 0.00310417
R19803 VPWR.n6324 VPWR.n6322 0.00310417
R19804 VPWR.n6327 VPWR.n6326 0.00310417
R19805 VPWR.n6340 VPWR.n6339 0.00310417
R19806 VPWR.n6189 VPWR.n6187 0.00310417
R19807 VPWR.n6108 VPWR.n6107 0.00310417
R19808 VPWR.n5968 VPWR.n5967 0.00310417
R19809 VPWR.n5976 VPWR.n5973 0.00310417
R19810 VPWR.n5981 VPWR.n5980 0.00310417
R19811 VPWR.n5986 VPWR.n5985 0.00310417
R19812 VPWR.n5794 VPWR.n5783 0.0028004
R19813 VPWR.n3067 VPWR.n3066 0.0028004
R19814 VPWR.n5813 VPWR.n4959 0.0028004
R19815 VPWR.n4270 VPWR.n1453 0.0028004
R19816 VPWR.n4420 VPWR.n4393 0.0028004
R19817 VPWR.n4445 VPWR.n4444 0.0028004
R19818 VPWR.n733 VPWR.n732 0.0028004
R19819 VPWR.n7061 VPWR.n7060 0.0028004
R19820 VPWR.n6996 VPWR.n4908 0.0028004
R19821 VPWR.n6601 VPWR.n6575 0.0028004
R19822 VPWR.n2068 VPWR.n2064 0.0028004
R19823 VPWR.n20 VPWR.n19 0.0028004
R19824 VPWR.n3201 VPWR.n3200 0.0028004
R19825 VPWR.n3539 VPWR.n2188 0.0028004
R19826 VPWR.n6452 VPWR.n6377 0.0028004
R19827 VPWR.n5685 VPWR.n5073 0.0028004
R19828 VPWR.n5654 VPWR.n5627 0.0028004
R19829 VPWR.n5422 VPWR.n5211 0.0028004
R19830 VPWR.n540 VPWR.n460 0.0028004
R19831 VPWR.n1008 VPWR.n1007 0.0028004
R19832 VPWR.n1284 VPWR.n1283 0.0028004
R19833 VPWR.n1904 VPWR.n1903 0.0028004
R19834 VPWR.n1829 VPWR.n1655 0.0028004
R19835 VPWR.n5716 VPWR.n5709 0.0028004
R19836 VPWR.n7513 VPWR.n7512 0.0028004
R19837 VPWR.n7513 VPWR.n255 0.0028004
R19838 VPWR.n7656 VPWR.n127 0.0028004
R19839 VPWR.n7656 VPWR.n7655 0.0028004
R19840 VPWR.n3399 VPWR.n3372 0.0028004
R19841 VPWR.n5915 VPWR.n5914 0.0028004
R19842 VPWR.n6023 VPWR.n5909 0.00277474
R19843 VPWR.n7659 VPWR.n7657 0.00251462
R19844 VPWR.n7516 VPWR.n7514 0.00251462
R19845 VPWR.n5120 VPWR.n5118 0.00251462
R19846 VPWR.n5626 VPWR.n5625 0.00251462
R19847 VPWR.n5384 VPWR.n5382 0.00251462
R19848 VPWR.n514 VPWR.n512 0.00251462
R19849 VPWR.n1051 VPWR.n1049 0.00251462
R19850 VPWR.n1282 VPWR.n1281 0.00251462
R19851 VPWR.n1902 VPWR.n1901 0.00251462
R19852 VPWR.n1712 VPWR.n1710 0.00251462
R19853 VPWR.n3542 VPWR.n3540 0.00251462
R19854 VPWR.n3715 VPWR.n3714 0.00251462
R19855 VPWR.n2067 VPWR.n2066 0.00251462
R19856 VPWR.n1471 VPWR.n1470 0.00251462
R19857 VPWR.n4392 VPWR.n4391 0.00251462
R19858 VPWR.n4443 VPWR.n4442 0.00251462
R19859 VPWR.n735 VPWR.n734 0.00251462
R19860 VPWR.n7063 VPWR.n7062 0.00251462
R19861 VPWR.n6995 VPWR.n6994 0.00251462
R19862 VPWR.n6603 VPWR.n6602 0.00251462
R19863 VPWR.n6451 VPWR.n6450 0.00251462
R19864 VPWR.n239 VPWR.n238 0.00251462
R19865 VPWR.n1549 VPWR.n1548 0.00251462
R19866 VPWR.n113 VPWR.n112 0.00251462
R19867 VPWR.n2377 VPWR.n2376 0.00251462
R19868 VPWR.n5816 VPWR.n5794 0.00246749
R19869 VPWR.n6571 VPWR.n4959 0.00246749
R19870 VPWR.n2070 VPWR.n2068 0.00246749
R19871 VPWR.n3067 VPWR.n2471 0.00246749
R19872 VPWR.n2035 VPWR.n1453 0.00246749
R19873 VPWR.n4393 VPWR.n419 0.00246749
R19874 VPWR.n4444 VPWR.n4433 0.00246749
R19875 VPWR.n733 VPWR.n624 0.00246749
R19876 VPWR.n7061 VPWR.n4881 0.00246749
R19877 VPWR.n7007 VPWR.n6996 0.00246749
R19878 VPWR.n6601 VPWR.n6600 0.00246749
R19879 VPWR.n7800 VPWR.n20 0.00246749
R19880 VPWR.n7797 VPWR.n7796 0.00246749
R19881 VPWR.n3201 VPWR.n2392 0.00246749
R19882 VPWR.n3539 VPWR.n3538 0.00246749
R19883 VPWR.n4133 VPWR.n1502 0.00246749
R19884 VPWR.n4298 VPWR.n4284 0.00246749
R19885 VPWR.n4570 VPWR.n4556 0.00246749
R19886 VPWR.n876 VPWR.n875 0.00246749
R19887 VPWR.n7203 VPWR.n7202 0.00246749
R19888 VPWR.n6877 VPWR.n6778 0.00246749
R19889 VPWR.n6767 VPWR.n131 0.00246749
R19890 VPWR.n4134 VPWR.n4133 0.00246749
R19891 VPWR.n4299 VPWR.n4298 0.00246749
R19892 VPWR.n4571 VPWR.n4570 0.00246749
R19893 VPWR.n876 VPWR.n597 0.00246749
R19894 VPWR.n7203 VPWR.n298 0.00246749
R19895 VPWR.n6878 VPWR.n6877 0.00246749
R19896 VPWR.n7632 VPWR.n131 0.00246749
R19897 VPWR.n7796 VPWR.n25 0.00246749
R19898 VPWR.n6355 VPWR.n5716 0.00246749
R19899 VPWR.n2680 VPWR.n2679 0.00246749
R19900 VPWR.n6453 VPWR.n6452 0.00246749
R19901 VPWR.n5657 VPWR.n5073 0.00246749
R19902 VPWR.n5627 VPWR.n5425 0.00246749
R19903 VPWR.n5226 VPWR.n5211 0.00246749
R19904 VPWR.n978 VPWR.n460 0.00246749
R19905 VPWR.n1210 VPWR.n1008 0.00246749
R19906 VPWR.n1283 VPWR.n1224 0.00246749
R19907 VPWR.n1903 VPWR.n1842 0.00246749
R19908 VPWR.n1807 VPWR.n1655 0.00246749
R19909 VPWR.n2679 VPWR.n2678 0.00246749
R19910 VPWR.n3732 VPWR.n3716 0.00246749
R19911 VPWR.n3372 VPWR.n3371 0.00246749
R19912 VPWR.n7398 VPWR.n256 0.00246749
R19913 VPWR.n7292 VPWR.n284 0.00246749
R19914 VPWR.n4757 VPWR.n301 0.00246749
R19915 VPWR.n4728 VPWR.n329 0.00246749
R19916 VPWR.n3957 VPWR.n3773 0.00246749
R19917 VPWR.n4052 VPWR.n4051 0.00246749
R19918 VPWR.n4051 VPWR.n3986 0.00246749
R19919 VPWR.n3773 VPWR.n3762 0.00246749
R19920 VPWR.n4754 VPWR.n4728 0.00246749
R19921 VPWR.n4854 VPWR.n301 0.00246749
R19922 VPWR.n7395 VPWR.n284 0.00246749
R19923 VPWR.n7495 VPWR.n256 0.00246749
R19924 VPWR.n3716 VPWR.n1565 0.00246749
R19925 VPWR.n4786 VPWR.n4785 0.00228056
R19926 VPWR.n4036 VPWR.n4035 0.00228056
R19927 VPWR.n7765 VPWR.n7764 0.00218919
R19928 VPWR.n140 VPWR.n136 0.00218919
R19929 VPWR.n6676 VPWR.n6675 0.00218919
R19930 VPWR.n6658 VPWR.n6657 0.00218919
R19931 VPWR.n6898 VPWR.n6897 0.00218919
R19932 VPWR.n4893 VPWR.n4892 0.00218919
R19933 VPWR.n7166 VPWR.n7152 0.00218919
R19934 VPWR.n7045 VPWR.n7044 0.00218919
R19935 VPWR.n7066 VPWR.n7065 0.00218919
R19936 VPWR.n842 VPWR.n834 0.00218919
R19937 VPWR.n706 VPWR.n633 0.00218919
R19938 VPWR.n738 VPWR.n737 0.00218919
R19939 VPWR.n4578 VPWR.n4574 0.00218919
R19940 VPWR.n1104 VPWR.n416 0.00218919
R19941 VPWR.n4306 VPWR.n4302 0.00218919
R19942 VPWR.n4405 VPWR.n4404 0.00218919
R19943 VPWR.n4141 VPWR.n4137 0.00218919
R19944 VPWR.n4255 VPWR.n4254 0.00218919
R19945 VPWR.n2180 VPWR.n2176 0.00218919
R19946 VPWR.n2062 VPWR.n2061 0.00218919
R19947 VPWR.n5811 VPWR.n5810 0.00218919
R19948 VPWR.n2203 VPWR.n2197 0.00218919
R19949 VPWR.n3033 VPWR.n3032 0.00218919
R19950 VPWR.n3045 VPWR.n3044 0.00218919
R19951 VPWR.n5781 VPWR.n5780 0.00218919
R19952 VPWR.n3196 VPWR.n2413 0.00218919
R19953 VPWR.n6067 VPWR.n6066 0.00218919
R19954 VPWR.n4958 VPWR.n4957 0.00218193
R19955 VPWR.n3069 VPWR.n3068 0.00218193
R19956 VPWR.n5793 VPWR.n5792 0.00218193
R19957 VPWR.n3203 VPWR.n3202 0.00218193
R19958 VPWR.n4 VPWR.n3 0.00218193
R19959 VPWR.n4132 VPWR.n4131 0.00218193
R19960 VPWR.n4297 VPWR.n4296 0.00218193
R19961 VPWR.n4569 VPWR.n4568 0.00218193
R19962 VPWR.n878 VPWR.n877 0.00218193
R19963 VPWR.n7205 VPWR.n7204 0.00218193
R19964 VPWR.n6876 VPWR.n6875 0.00218193
R19965 VPWR.n7611 VPWR.n7610 0.00218193
R19966 VPWR.n7795 VPWR.n7794 0.00218193
R19967 VPWR.n5715 VPWR.n5714 0.00218193
R19968 VPWR.n2652 VPWR.n2651 0.00218193
R19969 VPWR.n4050 VPWR.n4049 0.00218193
R19970 VPWR.n3772 VPWR.n3771 0.00218193
R19971 VPWR.n4727 VPWR.n4726 0.00218193
R19972 VPWR.n4794 VPWR.n4793 0.00218193
R19973 VPWR.n7324 VPWR.n7323 0.00218193
R19974 VPWR.n7434 VPWR.n7433 0.00218193
R19975 VPWR.n2473 VPWR.n2472 0.00211562
R19976 VPWR.n3523 VPWR.n3522 0.00211562
R19977 VPWR.n2490 VPWR.n2489 0.00211562
R19978 VPWR.n2284 VPWR.n2283 0.00211562
R19979 VPWR.n2999 VPWR.n2491 0.00185526
R19980 VPWR.n5137 VPWR.n5136 0.00180208
R19981 VPWR VPWR.n5140 0.00180208
R19982 VPWR.n6661 VPWR 0.00180208
R19983 VPWR.n6659 VPWR.n6580 0.00180208
R19984 VPWR VPWR.n6606 0.00180208
R19985 VPWR.n6654 VPWR 0.00180208
R19986 VPWR.n232 VPWR.n231 0.00180208
R19987 VPWR.n235 VPWR 0.00180208
R19988 VPWR.n5606 VPWR.n5603 0.00180208
R19989 VPWR.n5601 VPWR 0.00180208
R19990 VPWR.n5469 VPWR.n4916 0.00180208
R19991 VPWR.n7405 VPWR 0.00180208
R19992 VPWR.n7479 VPWR.n7478 0.00180208
R19993 VPWR.n7475 VPWR 0.00180208
R19994 VPWR.n5402 VPWR.n5344 0.00180208
R19995 VPWR.n5302 VPWR.n5301 0.00180208
R19996 VPWR.n7029 VPWR.n7028 0.00180208
R19997 VPWR.n7370 VPWR.n7369 0.00180208
R19998 VPWR.n7365 VPWR 0.00180208
R19999 VPWR.n558 VPWR.n557 0.00180208
R20000 VPWR VPWR.n561 0.00180208
R20001 VPWR.n687 VPWR.n686 0.00180208
R20002 VPWR.n718 VPWR 0.00180208
R20003 VPWR.n742 VPWR.n605 0.00180208
R20004 VPWR.n857 VPWR 0.00180208
R20005 VPWR.n4764 VPWR 0.00180208
R20006 VPWR VPWR.n4774 0.00180208
R20007 VPWR.n4839 VPWR.n4838 0.00180208
R20008 VPWR.n4834 VPWR 0.00180208
R20009 VPWR.n1071 VPWR.n1070 0.00180208
R20010 VPWR.n1126 VPWR.n1125 0.00180208
R20011 VPWR.n404 VPWR 0.00180208
R20012 VPWR.n4461 VPWR.n400 0.00180208
R20013 VPWR VPWR.n4687 0.00180208
R20014 VPWR.n4720 VPWR.n4718 0.00180208
R20015 VPWR.n1263 VPWR.n1260 0.00180208
R20016 VPWR.n1258 VPWR 0.00180208
R20017 VPWR.n1382 VPWR.n428 0.00180208
R20018 VPWR.n3785 VPWR 0.00180208
R20019 VPWR.n3927 VPWR.n3926 0.00180208
R20020 VPWR.n1928 VPWR.n1926 0.00180208
R20021 VPWR VPWR.n1931 0.00180208
R20022 VPWR.n2020 VPWR.n2018 0.00180208
R20023 VPWR.n2028 VPWR 0.00180208
R20024 VPWR VPWR.n4247 0.00180208
R20025 VPWR.n4234 VPWR.n4233 0.00180208
R20026 VPWR VPWR.n4059 0.00180208
R20027 VPWR VPWR.n1730 0.00180208
R20028 VPWR.n2112 VPWR.n2111 0.00180208
R20029 VPWR.n2078 VPWR.n2077 0.00180208
R20030 VPWR.n3686 VPWR.n3685 0.00180208
R20031 VPWR.n2761 VPWR.n2760 0.00180208
R20032 VPWR VPWR.n2764 0.00180208
R20033 VPWR VPWR.n2993 0.00180208
R20034 VPWR.n2824 VPWR.n2822 0.00180208
R20035 VPWR.n2851 VPWR.n2849 0.00180208
R20036 VPWR.n3418 VPWR 0.00180208
R20037 VPWR.n2358 VPWR.n2357 0.00180208
R20038 VPWR.n6434 VPWR.n6431 0.00180208
R20039 VPWR.n6429 VPWR 0.00180208
R20040 VPWR.n6533 VPWR.n6531 0.00180208
R20041 VPWR.n6566 VPWR.n6564 0.00180208
R20042 VPWR.n84 VPWR.n83 0.00180208
R20043 VPWR.n2631 VPWR.n2630 0.00180208
R20044 VPWR.n3108 VPWR.n3107 0.00180208
R20045 VPWR.n3076 VPWR.n3075 0.00180208
R20046 VPWR.n3334 VPWR.n3333 0.00180208
R20047 VPWR.n6334 VPWR.n6333 0.00180208
R20048 VPWR.n6210 VPWR.n6209 0.00180208
R20049 VPWR.n6178 VPWR.n6177 0.00180208
R20050 VPWR.n5987 VPWR.n5986 0.00180208
R20051 VPWR.n5990 VPWR 0.00180208
R20052 VPWR.n1728 VPWR.n1726 0.00164032
R20053 VPWR.n2999 VPWR.n2684 0.0014919
R20054 VPWR.n3035 VPWR.n3017 0.00144128
R20055 VPWR.n3521 VPWR.n3505 0.00140106
R20056 VPWR.n3505 VPWR.n2205 0.00140106
R20057 VPWR.n3405 VPWR.n3404 0.00140106
R20058 trim[0] trim[0].n0 35.6343
R20059 trim[0].n0 trim[0] 19.2609
R20060 trim[0].n0 trim[0] 2.70819
R20061 ctlp[6].n1 ctlp[6] 89.5426
R20062 ctlp[6].n1 ctlp[6] 19.2609
R20063 ctlp[6] ctlp[6].n0 3.62598
R20064 ctlp[6] ctlp[6].n1 2.70819
R20065 ctlp[6].n0 ctlp[6] 0.154033
R20066 ctlp[6].n0 ctlp[6] 0.00363333
R20067 ctln[1].n0 ctln[1] 82.6354
R20068 ctln[1].n0 ctln[1] 7.38553
R20069 ctln[1] ctln[1].n0 2.82782
R20070 trim[1].n2 trim[1] 73.1612
R20071 trim[1].n2 trim[1].n1 9.3005
R20072 trim[1].n3 trim[1].n0 9.05196
R20073 trim[1].n1 trim[1].n0 9.01492
R20074 trim[1].n3 trim[1].n2 3.72602
R20075 trim[1] trim[1].n5 2.52311
R20076 trim[1].n5 trim[1].n4 2.24426
R20077 trim[1].n4 trim[1].n1 0.0365577
R20078 trim[1].n5 trim[1].n0 0.0141816
R20079 trim[1].n4 trim[1].n3 0.00292567
R20080 ctlp[7].n1 ctlp[7] 92.353
R20081 ctlp[7].n1 ctlp[7] 19.2609
R20082 ctlp[7] ctlp[7].n1 2.70819
R20083 ctlp[7] ctlp[7].n0 0.106146
R20084 ctlp[7].n0 ctlp[7] 0.0739375
R20085 ctlp[7].n0 ctlp[7] 0.0138097
R20086 ctln[4].n3 ctln[4] 81.7298
R20087 ctln[4].n3 ctln[4].n1 9.3005
R20088 ctln[4].n4 ctln[4].n3 9.3005
R20089 ctln[4].n4 ctln[4].n0 9.05098
R20090 ctln[4].n1 ctln[4].n0 9.01252
R20091 ctln[4].n5 ctln[4].n2 3.79439
R20092 ctln[4] ctln[4].n6 3.17386
R20093 ctln[4].n6 ctln[4].n5 2.24426
R20094 ctln[4].n2 ctln[4] 2.08974
R20095 ctln[4].n3 ctln[4].n2 2.03855
R20096 ctln[4].n7 ctln[4] 0.0747105
R20097 ctln[4].n5 ctln[4].n1 0.0389615
R20098 ctln[4].n6 ctln[4].n0 0.0141816
R20099 ctln[4] ctln[4].n7 0.0105337
R20100 ctln[4].n7 ctln[4] 0.00842135
R20101 ctln[4].n5 ctln[4].n4 0.00290385
R20102 ctln[2].n0 ctln[2] 82.6405
R20103 ctln[2].n0 ctln[2] 10.7299
R20104 ctln[2] ctln[2].n0 2.82364
R20105 trim[2].n2 trim[2] 27.08
R20106 trim[2].n3 trim[2].n1 9.3005
R20107 trim[2].n4 trim[2].n3 9.3005
R20108 trim[2].n4 trim[2].n0 9.04377
R20109 trim[2].n1 trim[2].n0 9.01973
R20110 trim[2].n5 trim[2].n2 4.25601
R20111 trim[2].n3 trim[2].n2 2.94352
R20112 trim[2] trim[2].n6 2.48707
R20113 trim[2].n6 trim[2].n5 2.24426
R20114 trim[2].n5 trim[2].n1 0.03175
R20115 trim[2].n6 trim[2].n0 0.0141816
R20116 trim[2].n5 trim[2].n4 0.0101154
R20117 result[0].n4 result[0].n3 593.188
R20118 result[0].n3 result[0] 79.5613
R20119 result[0] result[0].n2 10.4588
R20120 result[0].n5 result[0].n1 9.3005
R20121 result[0].n6 result[0].n5 9.3005
R20122 result[0].n6 result[0].n0 9.05098
R20123 result[0].n1 result[0].n0 9.01252
R20124 result[0].n3 result[0] 7.02795
R20125 result[0].n4 result[0] 3.93496
R20126 result[0].n7 result[0].n2 3.75172
R20127 result[0] result[0].n8 2.45104
R20128 result[0].n8 result[0].n7 2.24426
R20129 result[0].n5 result[0].n2 1.87152
R20130 result[0].n5 result[0].n4 0.0592523
R20131 result[0].n7 result[0].n1 0.0389615
R20132 result[0].n8 result[0].n0 0.0141816
R20133 result[0].n7 result[0].n6 0.00290385
R20134 ctln[5].n0 ctln[5] 82.6354
R20135 ctln[5].n0 ctln[5] 7.373
R20136 ctln[5] ctln[5].n0 2.82782
R20137 ctln[3].n0 ctln[3] 82.6354
R20138 ctln[3].n0 ctln[3] 7.38553
R20139 ctln[3] ctln[3].n0 2.82782
R20140 trim[3].n2 trim[3] 27.08
R20141 trim[3].n3 trim[3].n1 9.3005
R20142 trim[3].n4 trim[3].n3 9.3005
R20143 trim[3].n4 trim[3].n0 9.04377
R20144 trim[3].n1 trim[3].n0 9.01973
R20145 trim[3].n5 trim[3].n2 4.25601
R20146 trim[3].n3 trim[3].n2 2.94352
R20147 trim[3] trim[3].n6 2.48707
R20148 trim[3].n6 trim[3].n5 2.24426
R20149 trim[3].n5 trim[3].n1 0.03175
R20150 trim[3].n6 trim[3].n0 0.0141816
R20151 trim[3].n5 trim[3].n4 0.0101154
R20152 result[1].n4 result[1].n3 593.188
R20153 result[1].n3 result[1] 79.5613
R20154 result[1] result[1].n2 10.4588
R20155 result[1].n5 result[1].n1 9.3005
R20156 result[1].n6 result[1].n5 9.3005
R20157 result[1].n6 result[1].n0 9.05098
R20158 result[1].n1 result[1].n0 9.01252
R20159 result[1].n3 result[1] 7.02795
R20160 result[1].n4 result[1] 3.93496
R20161 result[1].n7 result[1].n2 3.75172
R20162 result[1] result[1].n8 3.05818
R20163 result[1].n8 result[1].n7 2.24426
R20164 result[1].n5 result[1].n2 1.87152
R20165 result[1].n5 result[1].n4 0.0592523
R20166 result[1].n7 result[1].n1 0.0389615
R20167 result[1].n8 result[1].n0 0.0141816
R20168 result[1].n7 result[1].n6 0.00290385
R20169 ctln[6].n6 ctln[6].n5 65.4043
R20170 ctln[6].n6 ctln[6] 9.00791
R20171 ctln[6].n5 ctln[6].n4 4.57357
R20172 ctln[6].n1 ctln[6] 4.21294
R20173 ctln[6].n3 ctln[6].n1 2.24426
R20174 ctln[6] ctln[6].n6 1.73877
R20175 ctln[6].n3 ctln[6].n2 0.0365577
R20176 ctln[6].n1 ctln[6].n0 0.0141816
R20177 ctln[6].n4 ctln[6].n3 0.00336382
R20178 trim[4].n2 trim[4] 27.08
R20179 trim[4].n3 trim[4].n1 9.3005
R20180 trim[4].n4 trim[4].n3 9.3005
R20181 trim[4].n4 trim[4].n0 9.04377
R20182 trim[4].n1 trim[4].n0 9.01973
R20183 trim[4].n5 trim[4].n2 4.25601
R20184 trim[4].n3 trim[4].n2 2.94352
R20185 trim[4] trim[4].n6 2.48707
R20186 trim[4].n6 trim[4].n5 2.24426
R20187 trim[4].n5 trim[4].n1 0.03175
R20188 trim[4].n6 trim[4].n0 0.0141816
R20189 trim[4].n5 trim[4].n4 0.0101154
R20190 result[2].n0 result[2] 8.05976
R20191 result[2] result[2].n0 6.41086
R20192 result[2].n0 result[2] 2.68692
R20193 ctln[7].n0 ctln[7] 78.348
R20194 ctln[7].n0 ctln[7] 9.00791
R20195 ctln[7] ctln[7].n0 1.73877
R20196 trimb[0].n2 trimb[0] 11.1817
R20197 trimb[0].n3 trimb[0].n1 9.3005
R20198 trimb[0].n4 trimb[0].n3 9.3005
R20199 trimb[0].n4 trimb[0].n0 9.04377
R20200 trimb[0].n1 trimb[0].n0 9.01973
R20201 trimb[0].n5 trimb[0].n2 4.19732
R20202 trimb[0].n3 trimb[0].n2 3.00661
R20203 trimb[0] trimb[0].n6 2.29709
R20204 trimb[0].n6 trimb[0].n5 2.24426
R20205 trimb[0].n5 trimb[0].n1 0.03175
R20206 trimb[0].n6 trimb[0].n0 0.0141816
R20207 trimb[0].n5 trimb[0].n4 0.0101154
R20208 result[3].n5 result[3] 81.7298
R20209 result[3].n5 result[3].n4 9.3005
R20210 result[3].n6 result[3].n5 9.3005
R20211 result[3].n7 result[3].n6 9.05098
R20212 result[3].n4 result[3].n0 9.04085
R20213 result[3].n3 result[3].n2 3.79439
R20214 result[3].n8 result[3].n7 3.41895
R20215 result[3].n3 result[3] 2.08974
R20216 result[3].n5 result[3].n3 2.03855
R20217 result[3].n2 result[3].n1 1.35818
R20218 result[3].n8 result[3].n0 0.868169
R20219 result[3] result[3].n8 0.129323
R20220 result[3].n4 result[3].n2 0.0389615
R20221 result[3].n7 result[3].n1 0.0376622
R20222 result[3].n1 result[3].n0 0.0103621
R20223 result[3].n6 result[3].n2 0.00290385
R20224 ctlp[0].n7 ctlp[0].n6 32.7416
R20225 ctlp[0].n7 ctlp[0] 19.2609
R20226 ctlp[0].n6 ctlp[0].n4 4.25601
R20227 ctlp[0].n0 ctlp[0] 3.38228
R20228 ctlp[0].n6 ctlp[0].n5 2.94352
R20229 ctlp[0] ctlp[0].n7 2.70819
R20230 ctlp[0].n2 ctlp[0].n1 2.25561
R20231 ctlp[0].n1 ctlp[0].n0 0.0509808
R20232 ctlp[0].n4 ctlp[0].n3 0.03175
R20233 ctlp[0].n4 ctlp[0].n2 0.00339788
R20234 trimb[1].n2 trimb[1] 27.08
R20235 trimb[1].n3 trimb[1].n1 9.3005
R20236 trimb[1].n4 trimb[1].n3 9.3005
R20237 trimb[1].n4 trimb[1].n0 9.04377
R20238 trimb[1].n1 trimb[1].n0 9.01973
R20239 trimb[1].n5 trimb[1].n2 4.25601
R20240 trimb[1].n3 trimb[1].n2 2.94352
R20241 trimb[1] trimb[1].n6 2.48707
R20242 trimb[1].n6 trimb[1].n5 2.24426
R20243 trimb[1].n5 trimb[1].n1 0.03175
R20244 trimb[1].n6 trimb[1].n0 0.0141816
R20245 trimb[1].n5 trimb[1].n4 0.0101154
R20246 result[4].n3 result[4] 81.7298
R20247 result[4].n3 result[4].n1 9.3005
R20248 result[4].n4 result[4].n3 9.3005
R20249 result[4].n4 result[4].n0 9.05098
R20250 result[4].n1 result[4].n0 9.01252
R20251 result[4].n5 result[4].n2 3.79439
R20252 result[4] result[4].n6 2.45104
R20253 result[4].n6 result[4].n5 2.24426
R20254 result[4].n2 result[4] 2.08974
R20255 result[4].n3 result[4].n2 2.03855
R20256 result[4].n5 result[4].n1 0.0389615
R20257 result[4].n6 result[4].n0 0.0141816
R20258 result[4].n5 result[4].n4 0.00290385
R20259 ctlp[1].n0 ctlp[1] 16.6059
R20260 ctlp[1].n1 ctlp[1] 10.1205
R20261 ctlp[1] ctlp[1].n0 4.38347
R20262 ctlp[1].n1 ctlp[1] 0.131056
R20263 ctlp[1].n0 ctlp[1] 0.0672785
R20264 ctlp[1] ctlp[1].n1 0.00798673
R20265 trimb[2].n2 trimb[2] 27.08
R20266 trimb[2].n3 trimb[2].n1 9.3005
R20267 trimb[2].n4 trimb[2].n3 9.3005
R20268 trimb[2].n4 trimb[2].n0 9.04377
R20269 trimb[2].n1 trimb[2].n0 9.01973
R20270 trimb[2].n5 trimb[2].n2 4.25601
R20271 trimb[2].n3 trimb[2].n2 2.94352
R20272 trimb[2] trimb[2].n6 2.48707
R20273 trimb[2].n6 trimb[2].n5 2.24426
R20274 trimb[2].n5 trimb[2].n1 0.03175
R20275 trimb[2].n6 trimb[2].n0 0.0141816
R20276 trimb[2].n5 trimb[2].n4 0.0101154
R20277 result[5].n3 result[5] 81.7298
R20278 result[5].n3 result[5].n1 9.3005
R20279 result[5].n4 result[5].n3 9.3005
R20280 result[5].n4 result[5].n0 9.05098
R20281 result[5].n1 result[5].n0 9.01252
R20282 result[5].n5 result[5].n2 3.79439
R20283 result[5] result[5].n6 3.05818
R20284 result[5].n6 result[5].n5 2.24426
R20285 result[5].n2 result[5] 2.08974
R20286 result[5].n3 result[5].n2 2.03855
R20287 result[5].n5 result[5].n1 0.0389615
R20288 result[5].n6 result[5].n0 0.0141816
R20289 result[5].n5 result[5].n4 0.00290385
R20290 ctlp[2].n1 ctlp[2] 16.6059
R20291 ctlp[2].n1 ctlp[2] 7.5522
R20292 ctlp[2] ctlp[2].n0 3.63219
R20293 ctlp[2].n0 ctlp[2] 0.0788333
R20294 ctlp[2] ctlp[2].n1 0.067306
R20295 ctlp[2].n0 ctlp[2] 0.0129779
R20296 clk.n0 clk.t7 184.768
R20297 clk.n1 clk.t3 184.768
R20298 clk.n2 clk.t0 184.768
R20299 clk.n3 clk.t1 184.768
R20300 clk.n0 clk.t4 146.208
R20301 clk.n1 clk.t2 146.208
R20302 clk.n2 clk.t5 146.208
R20303 clk.n3 clk.t6 146.208
R20304 clk clk.n3 97.6099
R20305 clk clk.n4 60.0555
R20306 clk.n1 clk.n0 40.6397
R20307 clk.n2 clk.n1 40.6397
R20308 clk.n3 clk.n2 40.6397
R20309 clk.n4 clk 10.3624
R20310 clk.n4 clk 3.45447
R20311 trimb[3] trimb[3].n0 35.6343
R20312 trimb[3].n0 trimb[3] 19.2609
R20313 trimb[3].n0 trimb[3] 2.70819
R20314 result[6] result[6].n0 10.0086
R20315 result[6].n0 result[6] 8.05976
R20316 result[6].n0 result[6] 2.68692
R20317 ctlp[3].n0 ctlp[3] 16.6059
R20318 ctlp[3].n0 ctlp[3] 7.85577
R20319 ctlp[3] ctlp[3].n0 0.067306
R20320 result[7].n3 result[7].n1 628.779
R20321 result[7].n3 result[7].n2 585
R20322 result[7] result[7].n4 574.529
R20323 result[7].n1 result[7] 85.0829
R20324 result[7].n4 result[7].n3 18.2412
R20325 result[7].n5 result[7] 12.2035
R20326 result[7].n4 result[7].n0 9.15497
R20327 result[7] result[7].n5 3.45106
R20328 result[7].n2 result[7] 1.50638
R20329 result[7] result[7].n1 1.50638
R20330 result[7].n2 result[7].n0 1.2554
R20331 result[7].n5 result[7].n0 1.10628
R20332 ctlp[4].n0 ctlp[4] 16.6059
R20333 ctlp[4].n1 ctlp[4] 10.132
R20334 ctlp[4] ctlp[4].n0 4.38347
R20335 ctlp[4].n1 ctlp[4] 0.0844286
R20336 ctlp[4].n0 ctlp[4] 0.0672785
R20337 ctlp[4] ctlp[4].n1 0.012146
R20338 ctlp[5].n0 ctlp[5] 16.6059
R20339 ctlp[5].n1 ctlp[5] 10.1093
R20340 ctlp[5] ctlp[5].n0 4.38347
R20341 ctlp[5].n1 ctlp[5] 0.0788333
R20342 ctlp[5].n0 ctlp[5] 0.0672785
R20343 ctlp[5] ctlp[5].n1 0.0129779
R20344 cal.n3 cal.t1 259.022
R20345 cal.n3 cal.t0 175.798
R20346 cal.n6 cal.n4 9.3005
R20347 cal.n7 cal.n6 9.3005
R20348 cal.n4 cal.n0 9.04669
R20349 cal.n8 cal.n7 9.04377
R20350 cal.n6 cal.n3 7.31035
R20351 cal.n5 cal.n2 3.98384
R20352 cal.n9 cal.n8 3.41895
R20353 cal.n5 cal 1.78438
R20354 cal.n6 cal.n5 1.74562
R20355 cal.n2 cal.n1 1.35824
R20356 cal.n9 cal.n0 0.867979
R20357 cal cal.n9 0.381556
R20358 cal.n8 cal.n1 0.0376622
R20359 cal.n4 cal.n2 0.03175
R20360 cal.n7 cal.n2 0.0101154
R20361 cal.n1 cal.n0 0.00974356
R20362 comp.n7 comp.t0 222.725
R20363 comp.n5 comp.t1 177.171
R20364 comp.n5 comp.n4 152
R20365 comp.n6 comp.n3 152
R20366 comp.n6 comp.n5 10.5442
R20367 comp.n9 comp.n8 9.3005
R20368 comp.n8 comp.n1 9.3005
R20369 comp.n9 comp.n0 9.05098
R20370 comp.n1 comp.n0 9.01252
R20371 comp.n8 comp.n7 8.76429
R20372 comp.n4 comp 5.51161
R20373 comp.n10 comp.n2 4.02719
R20374 comp comp.n11 3.39779
R20375 comp.n4 comp.n3 2.48939
R20376 comp.n7 comp.n6 2.25988
R20377 comp.n11 comp.n10 2.24426
R20378 comp.n2 comp 1.64775
R20379 comp.n8 comp.n2 1.61183
R20380 comp.n8 comp.n3 0.533833
R20381 comp.n10 comp.n1 0.0389615
R20382 comp.n11 comp.n0 0.0141816
R20383 comp.n10 comp.n9 0.00290385
R20384 en.n2 en.t1 259.027
R20385 en.n2 en.t0 175.782
R20386 en.n3 en.n1 9.3005
R20387 en.n6 en.n5 9.3005
R20388 en.n1 en.n0 9.04136
R20389 en.n6 en.n0 9.02214
R20390 en.n3 en.n2 7.31533
R20391 en.n7 en.n4 4.57427
R20392 en en.n8 3.02215
R20393 en.n5 en.n4 2.24915
R20394 en.n8 en.n7 2.24426
R20395 en.n4 en.n3 0.692392
R20396 en.n5 en 0.692392
R20397 en.n7 en.n6 0.03175
R20398 en.n8 en.n0 0.0141816
R20399 en.n7 en.n1 0.0101154
R20400 rstn.n3 rstn.t0 259.027
R20401 rstn.n3 rstn.t1 175.782
R20402 rstn.n5 rstn.n4 9.3005
R20403 rstn.n8 rstn.n7 9.3005
R20404 rstn.n4 rstn.n0 9.0697
R20405 rstn.n9 rstn.n8 9.02214
R20406 rstn.n5 rstn.n3 7.31533
R20407 rstn.n6 rstn.n2 4.57427
R20408 rstn.n10 rstn.n9 3.41895
R20409 rstn.n7 rstn.n6 2.24915
R20410 rstn.n2 rstn.n1 1.35818
R20411 rstn.n10 rstn.n0 0.868169
R20412 rstn.n6 rstn.n5 0.692392
R20413 rstn.n7 rstn 0.692392
R20414 rstn rstn.n10 0.0932894
R20415 rstn.n9 rstn.n1 0.0376622
R20416 rstn.n8 rstn.n2 0.03175
R20417 rstn.n1 rstn.n0 0.0103621
R20418 rstn.n4 rstn.n2 0.0101154
R20419 trimb[4].n2 trimb[4] 27.08
R20420 trimb[4].n3 trimb[4].n1 9.3005
R20421 trimb[4].n4 trimb[4].n3 9.3005
R20422 trimb[4].n4 trimb[4].n0 9.04377
R20423 trimb[4].n1 trimb[4].n0 9.01973
R20424 trimb[4].n5 trimb[4].n2 4.25601
R20425 trimb[4].n3 trimb[4].n2 2.94352
R20426 trimb[4] trimb[4].n6 2.48707
R20427 trimb[4].n6 trimb[4].n5 2.24426
R20428 trimb[4].n5 trimb[4].n1 0.03175
R20429 trimb[4].n6 trimb[4].n0 0.0141816
R20430 trimb[4].n5 trimb[4].n4 0.0101154
R20431 clkc.n4 clkc.n3 574.133
R20432 clkc.n3 clkc 80.894
R20433 clkc clkc.n2 11.0668
R20434 clkc.n5 clkc.n1 9.3005
R20435 clkc.n6 clkc.n5 9.3005
R20436 clkc.n6 clkc.n0 9.04617
R20437 clkc.n1 clkc.n0 9.01733
R20438 clkc.n7 clkc.n2 4.14532
R20439 clkc.n5 clkc.n2 2.97937
R20440 clkc.n3 clkc 2.84494
R20441 clkc clkc.n8 2.45104
R20442 clkc.n8 clkc.n7 2.24426
R20443 clkc.n4 clkc 1.83668
R20444 clkc.n5 clkc.n4 0.0512129
R20445 clkc.n7 clkc.n1 0.0341538
R20446 clkc.n8 clkc.n0 0.0141816
R20447 clkc.n7 clkc.n6 0.00771154
R20448 valid.n2 valid 25.6731
R20449 valid.n3 valid.n2 9.3005
R20450 valid.n3 valid.n0 9.01973
R20451 valid.n5 valid.n4 9.0005
R20452 valid.n2 valid.n1 4.5765
R20453 valid valid.n5 4.23171
R20454 valid.n1 valid.n0 2.25706
R20455 valid.n5 valid.n0 0.0509808
R20456 valid.n4 valid.n3 0.0341538
R20457 valid.n4 valid.n1 0.00200872
R20458 sample.n3 sample 27.08
R20459 sample.n5 sample.n4 9.3005
R20460 sample.n6 sample.n5 9.3005
R20461 sample.n4 sample.n0 9.0697
R20462 sample.n7 sample.n6 9.02214
R20463 sample.n3 sample.n2 4.25601
R20464 sample.n8 sample.n7 3.41895
R20465 sample.n5 sample.n3 2.94352
R20466 sample.n2 sample.n1 1.35818
R20467 sample.n8 sample.n0 0.868169
R20468 sample sample.n8 0.129323
R20469 sample.n7 sample.n1 0.0376622
R20470 sample.n6 sample.n2 0.03175
R20471 sample.n1 sample.n0 0.0103621
R20472 sample.n4 sample.n2 0.0101154
R20473 ctln[0].n0 ctln[0] 81.7298
R20474 ctln[0].n3 ctln[0] 4.18004
R20475 ctln[0].n6 ctln[0].n5 3.79439
R20476 ctln[0].n5 ctln[0].n3 2.24426
R20477 ctln[0] ctln[0].n6 2.08974
R20478 ctln[0].n6 ctln[0].n0 2.03855
R20479 ctln[0].n5 ctln[0].n1 0.0389615
R20480 ctln[0].n3 ctln[0].n2 0.0141816
R20481 ctln[0].n5 ctln[0].n4 0.00290385
X_294_ net2 cal_count\[2\] VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_0_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_277_ _117_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_1
X_200_ cal_itt\[1\] cal_itt\[0\] cal_itt\[2\] _062_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__a31o_1
X_329_ clknet_2_2__leaf_clk _026_ net46 VGND VGND VPWR VPWR trim_mask\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput31 net31 VGND VGND VPWR VPWR trim[0] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR ctlp[6] sky130_fd_sc_hd__clkbuf_4
Xoutput7 net7 VGND VGND VPWR VPWR ctln[1] sky130_fd_sc_hd__buf_2
X_293_ cal_count\[0\] _126_ _125_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_276_ _110_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ trim_mask\[3\] _104_ _064_ trim_mask\[4\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a22o_1
X_328_ clknet_2_2__leaf_clk _025_ net46 VGND VGND VPWR VPWR trim_mask\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput32 net32 VGND VGND VPWR VPWR trim[1] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 VGND VGND VPWR VPWR ctlp[7] sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR ctln[4] sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR ctln[2] sky130_fd_sc_hd__buf_2
X_292_ cal_count\[1\] _122_ _128_ _123_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_275_ trim_mask\[3\] net50 trim_val\[3\] VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_189_ _051_ _050_ _048_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand3b_2
X_258_ trim_mask\[2\] _104_ _064_ trim_mask\[3\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__a22o_1
X_327_ clknet_2_2__leaf_clk _024_ net46 VGND VGND VPWR VPWR trim_mask\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput33 net33 VGND VGND VPWR VPWR trim[2] sky130_fd_sc_hd__clkbuf_4
Xoutput22 net22 VGND VGND VPWR VPWR result[0] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR ctln[5] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR ctln[3] sky130_fd_sc_hd__buf_2
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ cal_count\[0\] _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_274_ _115_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ _061_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_257_ trim_mask\[1\] _104_ _064_ trim_mask\[2\] VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a22o_1
X_326_ clknet_2_1__leaf_clk _023_ net43 VGND VGND VPWR VPWR mask\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ clknet_2_1__leaf_clk _006_ net43 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput34 net34 VGND VGND VPWR VPWR trim[3] sky130_fd_sc_hd__clkbuf_4
Xoutput23 net23 VGND VGND VPWR VPWR result[1] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR ctln[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ _125_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and2b_1
X_273_ _110_ _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_20_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ clknet_2_3__leaf_clk en_co_clk VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__and2b_2
X_256_ trim_mask\[0\] _104_ _064_ trim_mask\[1\] VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a22o_1
X_325_ clknet_2_1__leaf_clk _022_ net43 VGND VGND VPWR VPWR mask\[6\] sky130_fd_sc_hd__dfrtp_1
X_239_ _050_ calibrate _048_ _051_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nor4b_2
X_308_ clknet_2_0__leaf_clk _005_ net43 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput35 net35 VGND VGND VPWR VPWR trim[4] sky130_fd_sc_hd__clkbuf_4
Xoutput24 net24 VGND VGND VPWR VPWR result[2] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR ctln[7] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ trim_mask\[2\] net48 trim_val\[2\] VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__a21o_1
X_341_ clknet_2_3__leaf_clk _038_ net46 VGND VGND VPWR VPWR cal_count\[3\] sky130_fd_sc_hd__dfrtp_1
X_186_ _059_ _060_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__nor2_1
X_255_ net30 _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand2_2
X_324_ clknet_2_1__leaf_clk _021_ net44 VGND VGND VPWR VPWR mask\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_169_ state\[1\] state\[2\] state\[0\] VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__and3b_2
X_238_ _097_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__clkbuf_1
X_307_ clknet_2_0__leaf_clk _004_ net45 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput36 net36 VGND VGND VPWR VPWR trimb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 VGND VGND VPWR VPWR result[3] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR ctlp[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_271_ _113_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__clkbuf_1
X_340_ clknet_2_3__leaf_clk _037_ net47 VGND VGND VPWR VPWR cal_count\[2\] sky130_fd_sc_hd__dfstp_1
X_185_ net54 state\[0\] VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__or2_1
X_254_ _092_ net42 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__nor2_1
X_323_ clknet_2_1__leaf_clk _020_ net47 VGND VGND VPWR VPWR mask\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_168_ _050_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__and2b_1
X_237_ _048_ _090_ _096_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__mux2_1
X_306_ clknet_2_0__leaf_clk _003_ net44 VGND VGND VPWR VPWR cal_itt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput37 net37 VGND VGND VPWR VPWR trimb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 VGND VGND VPWR VPWR result[4] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR ctlp[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _110_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__and2_1
X_322_ clknet_2_1__leaf_clk _019_ net44 VGND VGND VPWR VPWR mask\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ net55 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
X_253_ mask\[7\] _102_ _074_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_167_ state\[1\] VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__buf_6
X_236_ _092_ _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nor2_1
X_305_ clknet_2_1__leaf_clk _002_ net43 VGND VGND VPWR VPWR cal_itt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_219_ _074_ _083_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput38 net38 VGND VGND VPWR VPWR trimb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 VGND VGND VPWR VPWR result[5] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR ctlp[2] sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_183_ net35 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__inv_2
X_252_ net52 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__inv_2
X_321_ clknet_2_1__leaf_clk _018_ net43 VGND VGND VPWR VPWR mask\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_235_ net55 _094_ net54 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__o21a_1
X_304_ clknet_2_3__leaf_clk _001_ net47 VGND VGND VPWR VPWR cal_itt\[1\] sky130_fd_sc_hd__dfrtp_1
X_166_ state\[2\] VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ mask\[4\] net26 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__or2_1
X_218_ mask\[4\] _078_ net26 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput39 net39 VGND VGND VPWR VPWR trimb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 VGND VGND VPWR VPWR result[6] sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 VGND VGND VPWR VPWR ctlp[3] sky130_fd_sc_hd__buf_2
XFILLER_0_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ _058_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
X_251_ mask\[7\] net52 _101_ mask\[6\] VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a22o_1
X_320_ clknet_2_0__leaf_clk _017_ net44 VGND VGND VPWR VPWR mask\[1\] sky130_fd_sc_hd__dfrtp_1
X_165_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
X_234_ mask\[0\] _049_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__nor2_1
X_303_ clknet_2_3__leaf_clk _000_ net47 VGND VGND VPWR VPWR cal_itt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_148_ net17 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__inv_2
X_217_ _074_ _082_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput29 net29 VGND VGND VPWR VPWR result[7] sky130_fd_sc_hd__buf_2
Xoutput18 net18 VGND VGND VPWR VPWR ctlp[4] sky130_fd_sc_hd__buf_2
XFILLER_0_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ trim_val\[4\] trim_mask\[4\] VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or2_1
X_250_ mask\[6\] net53 _101_ mask\[5\] VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_164_ state\[0\] VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__buf_6
X_233_ calibrate _093_ _074_ net1 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a22o_1
X_302_ cal_count\[3\] _066_ _136_ _092_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_147_ _042_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
X_216_ mask\[3\] _078_ net25 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput19 net19 VGND VGND VPWR VPWR ctlp[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_180_ net34 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__inv_2
Xfanout43 net45 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_163_ net31 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__inv_2
X_232_ net54 _049_ _090_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__or4_4
X_301_ _134_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ mask\[3\] net25 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__or2_1
X_215_ _074_ _081_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout44 net45 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_162_ _047_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
X_231_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__buf_6
X_300_ cal_count\[3\] net2 VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 cal VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_145_ net16 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
X_214_ mask\[2\] _078_ net24 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout45 net4 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_161_ trim_val\[0\] trim_mask\[0\] VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or2_1
X_230_ _053_ _063_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 comp VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ _041_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_213_ _074_ _080_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout46 net4 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_160_ net21 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__inv_2
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_289_ net2 cal_count\[1\] VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 en VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_143_ mask\[2\] net24 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__or2_1
X_212_ mask\[1\] _078_ net23 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout47 net4 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_288_ net2 cal_count\[1\] VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__and2_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput4 rstn VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ net15 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__inv_2
X_211_ _074_ _079_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_287_ _124_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ _040_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
X_210_ mask\[0\] _078_ net22 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a21oi_1
X_339_ clknet_2_3__leaf_clk _036_ net47 VGND VGND VPWR VPWR cal_count\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_286_ _122_ _123_ cal_count\[0\] VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_140_ net23 mask\[1\] VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ trim_mask\[1\] net49 trim_val\[1\] VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__a21o_1
X_338_ clknet_2_3__leaf_clk _035_ net47 VGND VGND VPWR VPWR cal_count\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_285_ _053_ _063_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_199_ _065_ _069_ _070_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nor3_1
X_268_ _111_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
X_337_ clknet_2_0__leaf_clk _034_ net44 VGND VGND VPWR VPWR en_co_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_284_ _053_ _065_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_17_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_198_ cal_itt\[1\] cal_itt\[0\] _067_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__and3_1
X_267_ _109_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__and2_1
X_336_ clknet_2_2__leaf_clk _033_ net46 VGND VGND VPWR VPWR trim_val\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_319_ clknet_2_0__leaf_clk _016_ net43 VGND VGND VPWR VPWR mask\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_283_ _121_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_197_ cal_itt\[0\] _067_ cal_itt\[1\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__a21oi_1
X_266_ _048_ _106_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__or2_1
X_335_ clknet_2_2__leaf_clk _032_ net46 VGND VGND VPWR VPWR trim_val\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ mask\[5\] net53 _101_ mask\[4\] VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a22o_1
X_318_ clknet_2_0__leaf_clk _015_ net45 VGND VGND VPWR VPWR state\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ _065_ _120_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_334_ clknet_2_2__leaf_clk _031_ net46 VGND VGND VPWR VPWR trim_val\[2\] sky130_fd_sc_hd__dfrtp_1
X_196_ _068_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_265_ trim_mask\[0\] _108_ trim_val\[0\] VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_179_ _057_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
X_248_ mask\[4\] net53 _101_ mask\[3\] VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a22o_1
X_317_ clknet_2_0__leaf_clk _014_ net45 VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ _090_ _092_ _095_ en_co_clk VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ _062_ _067_ cal_itt\[0\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__mux2_1
X_264_ _106_ _107_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nor2_4
X_333_ clknet_2_2__leaf_clk _030_ net46 VGND VGND VPWR VPWR trim_val\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ mask\[3\] net52 _101_ mask\[2\] VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a22o_1
X_316_ clknet_2_0__leaf_clk _013_ net45 VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfrtp_1
X_178_ trim_val\[3\] trim_mask\[3\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _119_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ trim_mask\[0\] _064_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__a21oi_1
X_263_ net54 _059_ _048_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21a_1
X_332_ clknet_2_2__leaf_clk _029_ net46 VGND VGND VPWR VPWR trim_val\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_177_ net33 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__inv_2
X_246_ mask\[2\] net52 _101_ mask\[1\] VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a22o_1
X_315_ clknet_2_0__leaf_clk _012_ net45 VGND VGND VPWR VPWR calibrate sky130_fd_sc_hd__dfrtp_1
X_229_ _087_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_193_ _053_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__nor2_1
X_262_ _053_ _063_ _105_ net55 net42 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__a221o_1
X_331_ clknet_2_2__leaf_clk _028_ net45 VGND VGND VPWR VPWR trim_mask\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ _056_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
X_245_ mask\[1\] net52 _101_ mask\[0\] VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a22o_1
X_314_ clknet_2_1__leaf_clk _011_ net43 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_159_ _046_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
X_228_ _052_ _088_ _048_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__o21a_1
Xclone1 state\[2\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ net54 _050_ _048_ net3 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__and4bb_2
X_261_ _048_ cal_count\[3\] VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_1
X_330_ clknet_2_2__leaf_clk _027_ net46 VGND VGND VPWR VPWR trim_mask\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_175_ trim_val\[2\] trim_mask\[2\] VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__or2_1
X_244_ _065_ net51 VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nor2_2
X_313_ clknet_2_1__leaf_clk _010_ net43 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
X_158_ mask\[7\] net29 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__or2_1
X_227_ _051_ net55 trim_mask\[0\] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_260_ calibrate _049_ _052_ _104_ trim_mask\[4\] VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _062_ _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nor2_2
X_174_ net32 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__inv_2
X_243_ net55 _060_ _096_ _100_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a22o_1
X_312_ clknet_2_1__leaf_clk _009_ net44 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire42 _098_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
X_157_ net20 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__inv_2
X_226_ net3 _062_ _075_ _060_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_13_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_190_ cal_itt\[3\] cal_itt\[2\] cal_itt\[1\] cal_itt\[0\] VGND VGND VPWR VPWR _063_
+ sky130_fd_sc_hd__nand4b_2
XFILLER_0_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_173_ _055_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_242_ calibrate _048_ _052_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__o21a_1
X_311_ clknet_2_1__leaf_clk _008_ net44 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_156_ _045_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
X_225_ _074_ _086_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nor2_1
X_139_ net14 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__inv_2
X_208_ _065_ net2 _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ clknet_2_1__leaf_clk _007_ net43 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
X_172_ trim_val\[1\] trim_mask\[1\] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__or2_1
X_241_ _092_ _099_ _095_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ mask\[6\] net28 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__or2_1
X_224_ mask\[7\] _078_ net29 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_138_ _039_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_207_ _075_ _049_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_171_ _054_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
X_240_ _087_ _098_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer1 _108_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
X_223_ _074_ _085_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__nor2_1
X_154_ net19 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__inv_2
X_137_ net22 mask\[0\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__or2_1
X_206_ _050_ _051_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ _049_ _052_ _053_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21o_1
X_299_ _129_ _130_ _131_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 _108_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_153_ _044_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_222_ mask\[6\] _078_ net28 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone7 state\[1\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_205_ _065_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ cal_count\[2\] _122_ _133_ _123_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 _108_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_152_ mask\[5\] net27 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__or2_1
X_221_ _074_ _084_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__nor2_1
X_204_ _073_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_297_ _129_ _132_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__xnor2_1
Xrebuffer4 _076_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_151_ net18 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__inv_2
X_220_ mask\[5\] _078_ net27 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__a21oi_1
X_203_ cal_itt\[3\] _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ _130_ _131_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer5 net51 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_6
X_150_ _043_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ trim_val\[4\] _118_ _108_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ cal_itt\[2\] _070_ _072_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput40 net40 VGND VGND VPWR VPWR trimb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput5 net5 VGND VGND VPWR VPWR clkc sky130_fd_sc_hd__buf_1
X_295_ net2 cal_count\[2\] VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__nand2_1
Xrebuffer6 _076_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
X_278_ _062_ net40 net30 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__o21ai_1
X_201_ _067_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput41 net41 VGND VGND VPWR VPWR valid sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 VGND VGND VPWR VPWR sample sky130_fd_sc_hd__clkbuf_4
Xoutput6 net6 VGND VGND VPWR VPWR ctln[0] sky130_fd_sc_hd__buf_2
C17823 output6/a_27_47# VGND 0.454f
C17824 output30/a_27_47# VGND 0.775f
C17825 output41/a_27_47# VGND 0.71f
C17826 _201_/a_113_47# VGND 0.002f
C17827 _278_/a_27_47# VGND 0.215f
C17828 _278_/a_109_297# VGND 1.45e-19
C17829 rebuffer6/a_27_47# VGND 0.368f
C17830 _295_/a_113_47# VGND 0.0019f
C17831 output5/a_27_47# VGND 0.378f
C17832 output40/a_27_47# VGND 0.802f
C17833 _202_/a_297_47# VGND 0.209f
C17834 _202_/a_382_297# VGND 2.39e-19
C17835 _202_/a_79_21# VGND 0.289f
C17836 _279_/a_490_47# VGND 0.00768f
C17837 _279_/a_206_47# VGND 0.0126f
C17838 _279_/a_314_297# VGND 0.00636f
C17839 _279_/a_204_297# VGND 0.00643f
C17840 _279_/a_396_47# VGND 0.664f
C17841 _279_/a_27_47# VGND 0.253f
C17842 _150_/a_27_47# VGND 0.34f
C17843 rebuffer5/a_161_47# VGND 0.842f
C17844 _296_/a_113_47# VGND 0.00178f
C17845 _203_/a_145_75# VGND 0.00502f
C17846 _203_/a_59_75# VGND 0.296f
C17847 _220_/a_199_47# VGND 0.00418f
C17848 _220_/a_113_297# VGND 0.0381f
C17849 rebuffer4/a_27_47# VGND 0.353f
C17850 _297_/a_285_47# VGND 0.249f
C17851 _297_/a_129_47# VGND 0.00585f
C17852 _297_/a_377_297# VGND 0.00413f
C17853 _297_/a_47_47# VGND 0.417f
C17854 _204_/a_75_212# VGND 0.411f
C17855 _221_/a_109_297# VGND 4.76e-19
C17856 _152_/a_150_297# VGND 2.29e-19
C17857 _152_/a_68_297# VGND 0.297f
C17858 rebuffer3/a_75_212# VGND 0.365f
C17859 _298_/a_215_47# VGND 0.344f
C17860 _298_/a_493_297# VGND 3.11e-20
C17861 _298_/a_292_297# VGND 1.01e-19
C17862 _298_/a_78_199# VGND 0.226f
C17863 _205_/a_27_47# VGND 0.788f
C17864 clone7/a_27_47# VGND 0.464f
C17865 _222_/a_199_47# VGND 0.00399f
C17866 _222_/a_113_297# VGND 0.0432f
C17867 _153_/a_27_47# VGND 0.381f
C17868 rebuffer2/a_75_212# VGND 0.401f
C17869 _299_/a_382_47# VGND 0.00446f
C17870 _299_/a_298_297# VGND 0.0125f
C17871 _299_/a_215_297# VGND 0.431f
C17872 _299_/a_27_413# VGND 0.285f
C17873 _170_/a_384_47# VGND 0.0034f
C17874 _170_/a_299_297# VGND 0.0402f
C17875 _170_/a_81_21# VGND 0.319f
C17876 _206_/a_206_47# VGND 0.00474f
C17877 _206_/a_27_93# VGND 0.276f
C17878 _137_/a_150_297# VGND 3.36e-19
C17879 _137_/a_68_297# VGND 0.296f
C17880 _223_/a_109_297# VGND 9.28e-19
C17881 rebuffer1/a_75_212# VGND 0.351f
C17882 _240_/a_109_297# VGND 2.42e-19
C17883 _171_/a_27_47# VGND 0.487f
C17884 _207_/a_109_297# VGND 3.87e-19
C17885 _138_/a_27_47# VGND 0.354f
C17886 _224_/a_199_47# VGND 0.00384f
C17887 _224_/a_113_297# VGND 0.0407f
C17888 _155_/a_150_297# VGND 1.76e-19
C17889 _155_/a_68_297# VGND 0.269f
C17890 _241_/a_297_47# VGND 0.185f
C17891 _241_/a_388_297# VGND 0.00113f
C17892 _241_/a_105_352# VGND 0.238f
C17893 _172_/a_150_297# VGND 3.32e-19
C17894 _172_/a_68_297# VGND 0.281f
C17895 _310_/a_1462_47# VGND 0.00134f
C17896 _310_/a_1217_47# VGND 4.86e-19
C17897 _310_/a_805_47# VGND 0.00597f
C17898 _310_/a_639_47# VGND 0.00897f
C17899 _310_/a_1270_413# VGND 4.62e-20
C17900 _310_/a_651_413# VGND 0.00625f
C17901 _310_/a_448_47# VGND 0.0809f
C17902 _310_/a_1108_47# VGND 0.277f
C17903 _310_/a_1283_21# VGND 0.531f
C17904 _310_/a_543_47# VGND 0.301f
C17905 _310_/a_761_289# VGND 0.197f
C17906 _310_/a_193_47# VGND 0.343f
C17907 _310_/a_27_47# VGND 0.796f
C17908 clkbuf_2_3__f_clk/a_110_47# VGND 2.24f
C17909 _208_/a_439_47# VGND 0.00381f
C17910 _208_/a_218_47# VGND 0.00336f
C17911 _208_/a_535_374# VGND 0.00133f
C17912 _208_/a_218_374# VGND 5.68e-19
C17913 _208_/a_505_21# VGND 0.393f
C17914 _208_/a_76_199# VGND 0.311f
C17915 _225_/a_109_297# VGND 4.16e-19
C17916 _156_/a_27_47# VGND 0.379f
C17917 _311_/a_1462_47# VGND 0.00141f
C17918 _311_/a_1217_47# VGND 5.6e-19
C17919 _311_/a_805_47# VGND 0.0053f
C17920 _311_/a_639_47# VGND 0.00756f
C17921 _311_/a_1270_413# VGND 8.96e-20
C17922 _311_/a_651_413# VGND 0.00796f
C17923 _311_/a_448_47# VGND 0.0779f
C17924 _311_/a_1108_47# VGND 0.284f
C17925 _311_/a_1283_21# VGND 0.539f
C17926 _311_/a_543_47# VGND 0.299f
C17927 _311_/a_761_289# VGND 0.208f
C17928 _311_/a_193_47# VGND 0.374f
C17929 _311_/a_27_47# VGND 0.692f
C17930 _242_/a_297_47# VGND 0.159f
C17931 _242_/a_382_297# VGND 2.91e-19
C17932 _242_/a_79_21# VGND 0.302f
C17933 _173_/a_27_47# VGND 0.318f
C17934 _190_/a_655_47# VGND 0.206f
C17935 _190_/a_465_47# VGND 0.193f
C17936 _190_/a_215_47# VGND 0.177f
C17937 _190_/a_27_47# VGND 0.407f
C17938 _209_/a_27_47# VGND 0.612f
C17939 _226_/a_303_47# VGND 0.00334f
C17940 _226_/a_197_47# VGND 0.00333f
C17941 _226_/a_109_47# VGND 0.00162f
C17942 _226_/a_27_47# VGND 0.29f
C17943 wire42/a_75_212# VGND 0.351f
C17944 _312_/a_1462_47# VGND 0.00257f
C17945 _312_/a_1217_47# VGND 0.00115f
C17946 _312_/a_805_47# VGND 0.00634f
C17947 _312_/a_639_47# VGND 0.00977f
C17948 _312_/a_1270_413# VGND 1.66e-19
C17949 _312_/a_651_413# VGND 0.0118f
C17950 _312_/a_448_47# VGND 0.0868f
C17951 _312_/a_1108_47# VGND 0.306f
C17952 _312_/a_1283_21# VGND 0.564f
C17953 _312_/a_543_47# VGND 0.313f
C17954 _312_/a_761_289# VGND 0.221f
C17955 _312_/a_193_47# VGND 0.403f
C17956 _312_/a_27_47# VGND 0.815f
C17957 _243_/a_373_47# VGND 0.00263f
C17958 _243_/a_109_47# VGND 0.00627f
C17959 _243_/a_109_297# VGND 0.00357f
C17960 _243_/a_27_297# VGND 0.434f
C17961 _191_/a_27_297# VGND 0.0666f
C17962 _260_/a_584_47# VGND 0.00556f
C17963 _260_/a_346_47# VGND 0.00368f
C17964 _260_/a_256_47# VGND 0.00262f
C17965 _260_/a_250_297# VGND 0.0428f
C17966 _260_/a_93_21# VGND 0.388f
C17967 _227_/a_368_53# VGND 0.00252f
C17968 _227_/a_296_53# VGND 4.85e-19
C17969 _227_/a_209_311# VGND 0.258f
C17970 _227_/a_109_93# VGND 0.223f
C17971 _158_/a_150_297# VGND 5.09e-19
C17972 _158_/a_68_297# VGND 0.299f
C17973 _313_/a_1462_47# VGND 0.00137f
C17974 _313_/a_1217_47# VGND 5.28e-19
C17975 _313_/a_805_47# VGND 0.00526f
C17976 _313_/a_639_47# VGND 0.00748f
C17977 _313_/a_1270_413# VGND 1.18e-19
C17978 _313_/a_651_413# VGND 0.00836f
C17979 _313_/a_448_47# VGND 0.0799f
C17980 _313_/a_1108_47# VGND 0.287f
C17981 _313_/a_1283_21# VGND 0.54f
C17982 _313_/a_543_47# VGND 0.285f
C17983 _313_/a_761_289# VGND 0.195f
C17984 _313_/a_193_47# VGND 0.382f
C17985 _313_/a_27_47# VGND 0.641f
C17986 _244_/a_27_297# VGND 0.0668f
C17987 _175_/a_150_297# VGND 5.84e-19
C17988 _175_/a_68_297# VGND 0.292f
C17989 _330_/a_1462_47# VGND 0.00221f
C17990 _330_/a_1217_47# VGND 0.00104f
C17991 _330_/a_805_47# VGND 0.0053f
C17992 _330_/a_639_47# VGND 0.00754f
C17993 _330_/a_1270_413# VGND 2.57e-20
C17994 _330_/a_651_413# VGND 0.00807f
C17995 _330_/a_448_47# VGND 0.0763f
C17996 _330_/a_1108_47# VGND 0.284f
C17997 _330_/a_1283_21# VGND 0.54f
C17998 _330_/a_543_47# VGND 0.286f
C17999 _330_/a_761_289# VGND 0.206f
C18000 _330_/a_193_47# VGND 0.338f
C18001 _330_/a_27_47# VGND 0.637f
C18002 _261_/a_113_47# VGND 0.0019f
C18003 _192_/a_639_47# VGND 0.00355f
C18004 _192_/a_548_47# VGND 0.00342f
C18005 _192_/a_476_47# VGND 0.00184f
C18006 _192_/a_505_280# VGND 0.278f
C18007 _192_/a_27_47# VGND 0.291f
C18008 _192_/a_174_21# VGND 0.34f
C18009 clone1/a_27_47# VGND 0.408f
C18010 _228_/a_297_47# VGND 0.194f
C18011 _228_/a_382_297# VGND 2.68e-19
C18012 _228_/a_79_21# VGND 0.312f
C18013 _159_/a_27_47# VGND 0.342f
C18014 _314_/a_1462_47# VGND 0.00221f
C18015 _314_/a_1217_47# VGND 0.00107f
C18016 _314_/a_805_47# VGND 0.00605f
C18017 _314_/a_639_47# VGND 0.00911f
C18018 _314_/a_1270_413# VGND 1.18e-19
C18019 _314_/a_651_413# VGND 0.00755f
C18020 _314_/a_448_47# VGND 0.0837f
C18021 _314_/a_1108_47# VGND 0.309f
C18022 _314_/a_1283_21# VGND 0.591f
C18023 _314_/a_543_47# VGND 0.289f
C18024 _314_/a_761_289# VGND 0.2f
C18025 _314_/a_193_47# VGND 0.358f
C18026 _314_/a_27_47# VGND 0.75f
C18027 _245_/a_373_47# VGND 0.00382f
C18028 _245_/a_109_47# VGND 0.00649f
C18029 _245_/a_109_297# VGND 0.00637f
C18030 _245_/a_27_297# VGND 0.457f
C18031 _176_/a_27_47# VGND 0.372f
C18032 _331_/a_1462_47# VGND 0.00282f
C18033 _331_/a_1217_47# VGND 0.00122f
C18034 _331_/a_805_47# VGND 0.00648f
C18035 _331_/a_639_47# VGND 0.01f
C18036 _331_/a_1270_413# VGND 1.07e-19
C18037 _331_/a_651_413# VGND 0.00785f
C18038 _331_/a_448_47# VGND 0.0836f
C18039 _331_/a_1108_47# VGND 0.314f
C18040 _331_/a_1283_21# VGND 0.577f
C18041 _331_/a_543_47# VGND 0.297f
C18042 _331_/a_761_289# VGND 0.201f
C18043 _331_/a_193_47# VGND 0.37f
C18044 _331_/a_27_47# VGND 0.785f
C18045 _262_/a_465_47# VGND 0.00239f
C18046 _262_/a_205_47# VGND 0.00156f
C18047 _262_/a_193_297# VGND 0.00115f
C18048 _262_/a_109_297# VGND 8.69e-19
C18049 _262_/a_27_47# VGND 0.633f
C18050 _193_/a_109_297# VGND 5.61e-19
C18051 _229_/a_27_297# VGND 0.0661f
C18052 _315_/a_1462_47# VGND 0.00221f
C18053 _315_/a_1217_47# VGND 9.68e-19
C18054 _315_/a_805_47# VGND 0.00579f
C18055 _315_/a_639_47# VGND 0.00863f
C18056 _315_/a_1270_413# VGND 2.91e-20
C18057 _315_/a_651_413# VGND 0.00515f
C18058 _315_/a_448_47# VGND 0.0803f
C18059 _315_/a_1108_47# VGND 0.304f
C18060 _315_/a_1283_21# VGND 0.578f
C18061 _315_/a_543_47# VGND 0.281f
C18062 _315_/a_761_289# VGND 0.194f
C18063 _315_/a_193_47# VGND 0.355f
C18064 _315_/a_27_47# VGND 0.808f
C18065 _246_/a_373_47# VGND 0.00257f
C18066 _246_/a_109_47# VGND 0.00679f
C18067 _246_/a_109_297# VGND 0.0103f
C18068 _246_/a_27_297# VGND 0.451f
C18069 _332_/a_1462_47# VGND 0.00219f
C18070 _332_/a_1217_47# VGND 5.42e-19
C18071 _332_/a_805_47# VGND 0.00579f
C18072 _332_/a_639_47# VGND 0.00863f
C18073 _332_/a_1270_413# VGND 2.69e-19
C18074 _332_/a_651_413# VGND 0.00605f
C18075 _332_/a_448_47# VGND 0.0818f
C18076 _332_/a_1108_47# VGND 0.303f
C18077 _332_/a_1283_21# VGND 0.561f
C18078 _332_/a_543_47# VGND 0.302f
C18079 _332_/a_761_289# VGND 0.196f
C18080 _332_/a_193_47# VGND 0.375f
C18081 _332_/a_27_47# VGND 0.78f
C18082 _263_/a_297_47# VGND 0.191f
C18083 _263_/a_382_297# VGND 6.69e-20
C18084 _263_/a_79_21# VGND 0.269f
C18085 _194_/a_199_47# VGND 0.00434f
C18086 _194_/a_113_297# VGND 0.0429f
C18087 _280_/a_75_212# VGND 0.329f
C18088 _178_/a_150_297# VGND 1.44e-19
C18089 _178_/a_68_297# VGND 0.289f
C18090 _316_/a_1462_47# VGND 0.00146f
C18091 _316_/a_1217_47# VGND 5.91e-19
C18092 _316_/a_805_47# VGND 0.00649f
C18093 _316_/a_639_47# VGND 0.00909f
C18094 _316_/a_1270_413# VGND 1.17e-19
C18095 _316_/a_651_413# VGND 0.0147f
C18096 _316_/a_448_47# VGND 0.0785f
C18097 _316_/a_1108_47# VGND 0.287f
C18098 _316_/a_1283_21# VGND 0.553f
C18099 _316_/a_543_47# VGND 0.308f
C18100 _316_/a_761_289# VGND 0.215f
C18101 _316_/a_193_47# VGND 0.382f
C18102 _316_/a_27_47# VGND 0.672f
C18103 _247_/a_373_47# VGND 0.00218f
C18104 _247_/a_109_47# VGND 0.00675f
C18105 _247_/a_109_297# VGND 0.00485f
C18106 _247_/a_27_297# VGND 0.454f
C18107 _333_/a_1462_47# VGND 0.0025f
C18108 _333_/a_1217_47# VGND 0.0014f
C18109 _333_/a_805_47# VGND 0.00631f
C18110 _333_/a_639_47# VGND 0.0096f
C18111 _333_/a_1270_413# VGND 1.2e-19
C18112 _333_/a_651_413# VGND 0.00798f
C18113 _333_/a_448_47# VGND 0.0787f
C18114 _333_/a_1108_47# VGND 0.304f
C18115 _333_/a_1283_21# VGND 0.547f
C18116 _333_/a_543_47# VGND 0.296f
C18117 _333_/a_761_289# VGND 0.218f
C18118 _333_/a_193_47# VGND 0.367f
C18119 _333_/a_27_47# VGND 0.66f
C18120 _264_/a_27_297# VGND 0.0686f
C18121 _195_/a_439_47# VGND 0.00331f
C18122 _195_/a_218_47# VGND 0.00263f
C18123 _195_/a_535_374# VGND 2.7e-19
C18124 _195_/a_218_374# VGND 5.37e-20
C18125 _195_/a_505_21# VGND 0.375f
C18126 _195_/a_76_199# VGND 0.28f
C18127 _281_/a_253_47# VGND 0.211f
C18128 _281_/a_337_297# VGND 4e-19
C18129 _281_/a_253_297# VGND 2.75e-19
C18130 _281_/a_103_199# VGND 0.312f
C18131 clkbuf_2_2__f_clk/a_110_47# VGND 2.22f
C18132 _317_/a_1462_47# VGND 0.00276f
C18133 _317_/a_1217_47# VGND 0.00109f
C18134 _317_/a_805_47# VGND 0.00658f
C18135 _317_/a_639_47# VGND 0.0123f
C18136 _317_/a_1270_413# VGND 1.01e-19
C18137 _317_/a_651_413# VGND 0.0114f
C18138 _317_/a_448_47# VGND 0.0904f
C18139 _317_/a_1108_47# VGND 0.313f
C18140 _317_/a_1283_21# VGND 0.573f
C18141 _317_/a_543_47# VGND 0.323f
C18142 _317_/a_761_289# VGND 0.217f
C18143 _317_/a_193_47# VGND 0.395f
C18144 _317_/a_27_47# VGND 0.822f
C18145 _248_/a_373_47# VGND 0.00263f
C18146 _248_/a_109_47# VGND 0.00646f
C18147 _248_/a_109_297# VGND 0.00455f
C18148 _248_/a_27_297# VGND 0.437f
C18149 _179_/a_27_47# VGND 0.354f
C18150 _265_/a_384_47# VGND 0.00327f
C18151 _265_/a_299_297# VGND 0.044f
C18152 _265_/a_81_21# VGND 0.3f
C18153 _334_/a_1462_47# VGND 0.00405f
C18154 _334_/a_1217_47# VGND 0.00103f
C18155 _334_/a_805_47# VGND 0.00579f
C18156 _334_/a_639_47# VGND 0.00863f
C18157 _334_/a_1270_413# VGND 2.69e-19
C18158 _334_/a_651_413# VGND 0.00733f
C18159 _334_/a_448_47# VGND 0.08f
C18160 _334_/a_1108_47# VGND 0.319f
C18161 _334_/a_1283_21# VGND 0.576f
C18162 _334_/a_543_47# VGND 0.291f
C18163 _334_/a_761_289# VGND 0.212f
C18164 _334_/a_193_47# VGND 0.373f
C18165 _334_/a_27_47# VGND 0.738f
C18166 _282_/a_150_297# VGND 2.64e-19
C18167 _282_/a_68_297# VGND 0.269f
C18168 _318_/a_1462_47# VGND 0.00221f
C18169 _318_/a_1217_47# VGND 9.68e-19
C18170 _318_/a_805_47# VGND 0.00579f
C18171 _318_/a_639_47# VGND 0.00863f
C18172 _318_/a_651_413# VGND 0.00472f
C18173 _318_/a_448_47# VGND 0.0818f
C18174 _318_/a_1108_47# VGND 0.304f
C18175 _318_/a_1283_21# VGND 0.576f
C18176 _318_/a_543_47# VGND 0.298f
C18177 _318_/a_761_289# VGND 0.196f
C18178 _318_/a_193_47# VGND 0.374f
C18179 _318_/a_27_47# VGND 0.821f
C18180 _249_/a_373_47# VGND 0.00485f
C18181 _249_/a_109_47# VGND 0.0068f
C18182 _249_/a_109_297# VGND 0.0048f
C18183 _249_/a_27_297# VGND 0.485f
C18184 _335_/a_1462_47# VGND 0.00135f
C18185 _335_/a_1217_47# VGND 5.42e-19
C18186 _335_/a_805_47# VGND 0.0052f
C18187 _335_/a_639_47# VGND 0.00754f
C18188 _335_/a_1270_413# VGND 6.88e-20
C18189 _335_/a_651_413# VGND 0.0101f
C18190 _335_/a_448_47# VGND 0.0801f
C18191 _335_/a_1108_47# VGND 0.284f
C18192 _335_/a_1283_21# VGND 0.547f
C18193 _335_/a_543_47# VGND 0.289f
C18194 _335_/a_761_289# VGND 0.212f
C18195 _335_/a_193_47# VGND 0.364f
C18196 _335_/a_27_47# VGND 0.779f
C18197 _266_/a_150_297# VGND 9.13e-22
C18198 _266_/a_68_297# VGND 0.274f
C18199 _197_/a_199_47# VGND 0.00387f
C18200 _197_/a_113_297# VGND 0.0444f
C18201 _283_/a_75_212# VGND 0.333f
C18202 _319_/a_1462_47# VGND 0.00139f
C18203 _319_/a_1217_47# VGND 5.49e-19
C18204 _319_/a_805_47# VGND 0.00527f
C18205 _319_/a_639_47# VGND 0.0075f
C18206 _319_/a_1270_413# VGND 6.7e-20
C18207 _319_/a_651_413# VGND 0.00642f
C18208 _319_/a_448_47# VGND 0.0761f
C18209 _319_/a_1108_47# VGND 0.281f
C18210 _319_/a_1283_21# VGND 0.537f
C18211 _319_/a_543_47# VGND 0.278f
C18212 _319_/a_761_289# VGND 0.191f
C18213 _319_/a_193_47# VGND 0.336f
C18214 _319_/a_27_47# VGND 0.667f
C18215 _336_/a_1462_47# VGND 0.00127f
C18216 _336_/a_1217_47# VGND 4.65e-19
C18217 _336_/a_805_47# VGND 0.00513f
C18218 _336_/a_639_47# VGND 0.00719f
C18219 _336_/a_651_413# VGND 0.00587f
C18220 _336_/a_448_47# VGND 0.0747f
C18221 _336_/a_1108_47# VGND 0.277f
C18222 _336_/a_1283_21# VGND 0.526f
C18223 _336_/a_543_47# VGND 0.276f
C18224 _336_/a_761_289# VGND 0.19f
C18225 _336_/a_193_47# VGND 0.332f
C18226 _336_/a_27_47# VGND 0.649f
C18227 _267_/a_145_75# VGND 0.00339f
C18228 _267_/a_59_75# VGND 0.279f
C18229 _198_/a_181_47# VGND 0.00221f
C18230 _198_/a_109_47# VGND 8.26e-19
C18231 _198_/a_27_47# VGND 0.314f
C18232 _284_/a_150_297# VGND 2.82e-19
C18233 _284_/a_68_297# VGND 0.287f
C18234 _337_/a_1462_47# VGND 0.00248f
C18235 _337_/a_1217_47# VGND 0.00108f
C18236 _337_/a_805_47# VGND 0.00525f
C18237 _337_/a_639_47# VGND 0.0074f
C18238 _337_/a_1270_413# VGND 5.36e-20
C18239 _337_/a_651_413# VGND 0.00719f
C18240 _337_/a_448_47# VGND 0.0771f
C18241 _337_/a_1108_47# VGND 0.308f
C18242 _337_/a_1283_21# VGND 0.572f
C18243 _337_/a_543_47# VGND 0.282f
C18244 _337_/a_761_289# VGND 0.212f
C18245 _337_/a_193_47# VGND 0.367f
C18246 _337_/a_27_47# VGND 0.629f
C18247 _268_/a_75_212# VGND 0.366f
C18248 _199_/a_193_297# VGND 1.59e-20
C18249 _199_/a_109_297# VGND 2.46e-19
C18250 _285_/a_113_47# VGND 0.00209f
C18251 _338_/a_1296_47# VGND 0.00475f
C18252 _338_/a_1224_47# VGND 0.00121f
C18253 _338_/a_1056_47# VGND 0.00341f
C18254 _338_/a_796_47# VGND 0.00541f
C18255 _338_/a_586_47# VGND 8.36e-19
C18256 _338_/a_1140_413# VGND 3.5e-19
C18257 _338_/a_956_413# VGND 9.02e-19
C18258 _338_/a_562_413# VGND 5.72e-19
C18259 _338_/a_381_47# VGND 0.112f
C18260 _338_/a_1602_47# VGND 0.241f
C18261 _338_/a_1032_413# VGND 0.501f
C18262 _338_/a_1182_261# VGND 0.208f
C18263 _338_/a_476_47# VGND 0.5f
C18264 _338_/a_652_21# VGND 0.212f
C18265 _338_/a_193_47# VGND 0.447f
C18266 _338_/a_27_47# VGND 0.653f
C18267 _269_/a_384_47# VGND 0.00375f
C18268 _269_/a_299_297# VGND 0.0435f
C18269 _269_/a_81_21# VGND 0.308f
C18270 _140_/a_150_297# VGND 9.13e-22
C18271 _140_/a_68_297# VGND 0.267f
C18272 _286_/a_439_47# VGND 0.00328f
C18273 _286_/a_218_47# VGND 0.00302f
C18274 _286_/a_535_374# VGND 4.71e-19
C18275 _286_/a_218_374# VGND 6.4e-19
C18276 _286_/a_505_21# VGND 0.377f
C18277 _286_/a_76_199# VGND 0.306f
C18278 _339_/a_1296_47# VGND 0.00474f
C18279 _339_/a_1224_47# VGND 0.00119f
C18280 _339_/a_1056_47# VGND 0.00337f
C18281 _339_/a_796_47# VGND 0.00535f
C18282 _339_/a_586_47# VGND 8.52e-19
C18283 _339_/a_1140_413# VGND 6.77e-20
C18284 _339_/a_956_413# VGND 5.26e-19
C18285 _339_/a_562_413# VGND 1.7e-19
C18286 _339_/a_381_47# VGND 0.0985f
C18287 _339_/a_1602_47# VGND 0.21f
C18288 _339_/a_1032_413# VGND 0.458f
C18289 _339_/a_1182_261# VGND 0.187f
C18290 _339_/a_476_47# VGND 0.475f
C18291 _339_/a_652_21# VGND 0.211f
C18292 _339_/a_193_47# VGND 0.418f
C18293 _339_/a_27_47# VGND 0.611f
C18294 _210_/a_199_47# VGND 0.00411f
C18295 _210_/a_113_297# VGND 0.0442f
C18296 _141_/a_27_47# VGND 0.364f
C18297 _287_/a_75_212# VGND 0.331f
C18298 _211_/a_109_297# VGND 4.14e-19
C18299 clkbuf_2_1__f_clk/a_110_47# VGND 2.21f
C18300 _288_/a_145_75# VGND 0.00495f
C18301 _288_/a_59_75# VGND 0.33f
C18302 fanout47/a_27_47# VGND 0.53f
C18303 _212_/a_199_47# VGND 0.00379f
C18304 _212_/a_113_297# VGND 0.0375f
C18305 _143_/a_150_297# VGND 2.45e-19
C18306 _143_/a_68_297# VGND 0.286f
C18307 _289_/a_150_297# VGND 2.64e-19
C18308 _289_/a_68_297# VGND 0.288f
C18309 fanout46/a_27_47# VGND 0.705f
C18310 _144_/a_27_47# VGND 0.316f
C18311 _230_/a_145_75# VGND 0.00355f
C18312 _230_/a_59_75# VGND 0.281f
C18313 _161_/a_150_297# VGND 1.71e-19
C18314 _161_/a_68_297# VGND 0.266f
C18315 fanout45/a_27_47# VGND 0.458f
C18316 _214_/a_199_47# VGND 0.00523f
C18317 _214_/a_113_297# VGND 0.0494f
C18318 _300_/a_285_47# VGND 0.226f
C18319 _300_/a_129_47# VGND 0.0057f
C18320 _300_/a_377_297# VGND 4.18e-19
C18321 _300_/a_47_47# VGND 0.346f
C18322 _231_/a_161_47# VGND 0.855f
C18323 _162_/a_27_47# VGND 0.347f
C18324 fanout44/a_27_47# VGND 0.46f
C18325 _215_/a_109_297# VGND 0.00114f
C18326 _146_/a_150_297# VGND 1.78e-19
C18327 _146_/a_68_297# VGND 0.279f
C18328 _301_/a_285_47# VGND 0.225f
C18329 _301_/a_129_47# VGND 0.00565f
C18330 _301_/a_47_47# VGND 0.343f
C18331 _232_/a_304_297# VGND 4.88e-20
C18332 _232_/a_220_297# VGND 1.4e-19
C18333 _232_/a_114_297# VGND 2.21e-19
C18334 _232_/a_32_297# VGND 0.718f
C18335 fanout43/a_27_47# VGND 0.678f
C18336 output19/a_27_47# VGND 0.46f
C18337 _216_/a_199_47# VGND 0.00429f
C18338 _216_/a_113_297# VGND 0.0413f
C18339 _147_/a_27_47# VGND 0.386f
C18340 _302_/a_373_47# VGND 0.00231f
C18341 _302_/a_109_47# VGND 0.00653f
C18342 _302_/a_109_297# VGND 0.00732f
C18343 _302_/a_27_297# VGND 0.445f
C18344 _233_/a_373_47# VGND 0.00366f
C18345 _233_/a_109_47# VGND 0.00604f
C18346 _233_/a_109_297# VGND 0.00409f
C18347 _233_/a_27_297# VGND 0.46f
C18348 _164_/a_161_47# VGND 0.83f
C18349 _250_/a_373_47# VGND 0.00372f
C18350 _250_/a_109_47# VGND 0.00623f
C18351 _250_/a_109_297# VGND 0.00428f
C18352 _250_/a_27_297# VGND 0.443f
C18353 _181_/a_150_297# VGND 2.7e-19
C18354 _181_/a_68_297# VGND 0.283f
C18355 output18/a_27_47# VGND 0.464f
C18356 output29/a_27_47# VGND 0.457f
C18357 _217_/a_109_297# VGND 3.87e-19
C18358 _303_/a_1462_47# VGND 0.00242f
C18359 _303_/a_1217_47# VGND 0.00107f
C18360 _303_/a_805_47# VGND 0.00604f
C18361 _303_/a_639_47# VGND 0.00915f
C18362 _303_/a_1270_413# VGND 5.06e-20
C18363 _303_/a_651_413# VGND 0.00584f
C18364 _303_/a_448_47# VGND 0.0836f
C18365 _303_/a_1108_47# VGND 0.303f
C18366 _303_/a_1283_21# VGND 0.681f
C18367 _303_/a_543_47# VGND 0.285f
C18368 _303_/a_761_289# VGND 0.202f
C18369 _303_/a_193_47# VGND 0.363f
C18370 _303_/a_27_47# VGND 0.801f
C18371 _234_/a_109_297# VGND 9.65e-19
C18372 _320_/a_1462_47# VGND 0.00221f
C18373 _320_/a_1217_47# VGND 4.65e-19
C18374 _320_/a_805_47# VGND 0.00507f
C18375 _320_/a_639_47# VGND 0.00711f
C18376 _320_/a_1270_413# VGND 5.39e-20
C18377 _320_/a_651_413# VGND 0.00834f
C18378 _320_/a_448_47# VGND 0.0797f
C18379 _320_/a_1108_47# VGND 0.295f
C18380 _320_/a_1283_21# VGND 0.543f
C18381 _320_/a_543_47# VGND 0.296f
C18382 _320_/a_761_289# VGND 0.206f
C18383 _320_/a_193_47# VGND 0.356f
C18384 _320_/a_27_47# VGND 0.631f
C18385 _251_/a_373_47# VGND 0.00239f
C18386 _251_/a_109_47# VGND 0.00847f
C18387 _251_/a_109_297# VGND 0.00886f
C18388 _251_/a_27_297# VGND 0.453f
C18389 _182_/a_27_47# VGND 0.349f
C18390 clkbuf_2_0__f_clk/a_110_47# VGND 2.28f
C18391 output17/a_27_47# VGND 0.442f
C18392 output28/a_27_47# VGND 0.712f
C18393 output39/a_27_47# VGND 0.726f
C18394 _218_/a_199_47# VGND 0.00382f
C18395 _218_/a_113_297# VGND 0.0386f
C18396 _149_/a_150_297# VGND 1.18e-19
C18397 _149_/a_68_297# VGND 0.276f
C18398 _166_/a_161_47# VGND 0.903f
C18399 _304_/a_1462_47# VGND 0.00405f
C18400 _304_/a_1217_47# VGND 0.00116f
C18401 _304_/a_805_47# VGND 0.00622f
C18402 _304_/a_639_47# VGND 0.0094f
C18403 _304_/a_1270_413# VGND 1e-19
C18404 _304_/a_651_413# VGND 0.00897f
C18405 _304_/a_448_47# VGND 0.0817f
C18406 _304_/a_1108_47# VGND 0.32f
C18407 _304_/a_1283_21# VGND 0.588f
C18408 _304_/a_543_47# VGND 0.295f
C18409 _304_/a_761_289# VGND 0.213f
C18410 _304_/a_193_47# VGND 0.36f
C18411 _304_/a_27_47# VGND 0.749f
C18412 _235_/a_297_47# VGND 0.145f
C18413 _235_/a_79_21# VGND 0.269f
C18414 _321_/a_1462_47# VGND 0.00247f
C18415 _321_/a_1217_47# VGND 5.51e-19
C18416 _321_/a_805_47# VGND 0.00527f
C18417 _321_/a_639_47# VGND 0.00744f
C18418 _321_/a_1270_413# VGND 8.16e-20
C18419 _321_/a_651_413# VGND 0.00904f
C18420 _321_/a_448_47# VGND 0.0755f
C18421 _321_/a_1108_47# VGND 0.298f
C18422 _321_/a_1283_21# VGND 0.54f
C18423 _321_/a_543_47# VGND 0.297f
C18424 _321_/a_761_289# VGND 0.208f
C18425 _321_/a_193_47# VGND 0.355f
C18426 _321_/a_27_47# VGND 0.634f
C18427 output16/a_27_47# VGND 0.486f
C18428 output27/a_27_47# VGND 0.461f
C18429 output38/a_27_47# VGND 0.792f
C18430 _219_/a_109_297# VGND 1.66e-20
C18431 _305_/a_1462_47# VGND 0.00232f
C18432 _305_/a_1217_47# VGND 4.71e-19
C18433 _305_/a_805_47# VGND 0.00514f
C18434 _305_/a_639_47# VGND 0.00725f
C18435 _305_/a_1270_413# VGND 3.27e-20
C18436 _305_/a_651_413# VGND 0.00576f
C18437 _305_/a_448_47# VGND 0.0756f
C18438 _305_/a_1108_47# VGND 0.283f
C18439 _305_/a_1283_21# VGND 0.537f
C18440 _305_/a_543_47# VGND 0.281f
C18441 _305_/a_761_289# VGND 0.19f
C18442 _305_/a_193_47# VGND 0.339f
C18443 _305_/a_27_47# VGND 0.702f
C18444 _236_/a_109_297# VGND 5.53e-20
C18445 _167_/a_161_47# VGND 0.883f
C18446 _253_/a_384_47# VGND 0.0037f
C18447 _253_/a_299_297# VGND 0.0404f
C18448 _253_/a_81_21# VGND 0.316f
C18449 _322_/a_1462_47# VGND 0.00221f
C18450 _322_/a_1217_47# VGND 5.27e-19
C18451 _322_/a_805_47# VGND 0.00604f
C18452 _322_/a_639_47# VGND 0.00915f
C18453 _322_/a_1270_413# VGND 5.06e-20
C18454 _322_/a_651_413# VGND 0.00562f
C18455 _322_/a_448_47# VGND 0.0814f
C18456 _322_/a_1108_47# VGND 0.283f
C18457 _322_/a_1283_21# VGND 0.543f
C18458 _322_/a_543_47# VGND 0.301f
C18459 _322_/a_761_289# VGND 0.195f
C18460 _322_/a_193_47# VGND 0.35f
C18461 _322_/a_27_47# VGND 0.793f
C18462 _270_/a_145_75# VGND 0.0047f
C18463 _270_/a_59_75# VGND 0.327f
C18464 output15/a_27_47# VGND 0.458f
C18465 output26/a_27_47# VGND 0.461f
C18466 output37/a_27_47# VGND 0.737f
C18467 _306_/a_1462_47# VGND 0.00255f
C18468 _306_/a_1217_47# VGND 0.00115f
C18469 _306_/a_805_47# VGND 0.00723f
C18470 _306_/a_639_47# VGND 0.0132f
C18471 _306_/a_1270_413# VGND 9.17e-20
C18472 _306_/a_651_413# VGND 0.0132f
C18473 _306_/a_448_47# VGND 0.0838f
C18474 _306_/a_1108_47# VGND 0.294f
C18475 _306_/a_1283_21# VGND 0.542f
C18476 _306_/a_543_47# VGND 0.314f
C18477 _306_/a_761_289# VGND 0.212f
C18478 _306_/a_193_47# VGND 0.382f
C18479 _306_/a_27_47# VGND 0.787f
C18480 _237_/a_439_47# VGND 0.00301f
C18481 _237_/a_218_47# VGND 0.00264f
C18482 _237_/a_535_374# VGND 4.27e-19
C18483 _237_/a_218_374# VGND 4.4e-19
C18484 _237_/a_505_21# VGND 0.426f
C18485 _237_/a_76_199# VGND 0.292f
C18486 _168_/a_297_47# VGND 0.00547f
C18487 _168_/a_207_413# VGND 0.256f
C18488 _168_/a_27_413# VGND 0.292f
C18489 _323_/a_1462_47# VGND 0.00133f
C18490 _323_/a_1217_47# VGND 0.00103f
C18491 _323_/a_805_47# VGND 0.00595f
C18492 _323_/a_639_47# VGND 0.00896f
C18493 _323_/a_1270_413# VGND 2.27e-20
C18494 _323_/a_651_413# VGND 0.00734f
C18495 _323_/a_448_47# VGND 0.0814f
C18496 _323_/a_1108_47# VGND 0.304f
C18497 _323_/a_1283_21# VGND 0.537f
C18498 _323_/a_543_47# VGND 0.301f
C18499 _323_/a_761_289# VGND 0.211f
C18500 _323_/a_193_47# VGND 0.362f
C18501 _323_/a_27_47# VGND 0.757f
C18502 _254_/a_109_297# VGND 5.03e-19
C18503 _185_/a_150_297# VGND 1.36e-19
C18504 _185_/a_68_297# VGND 0.276f
C18505 _340_/a_1296_47# VGND 0.00523f
C18506 _340_/a_1224_47# VGND 0.00169f
C18507 _340_/a_1056_47# VGND 0.00386f
C18508 _340_/a_796_47# VGND 0.00583f
C18509 _340_/a_586_47# VGND 0.00172f
C18510 _340_/a_956_413# VGND 3.4e-19
C18511 _340_/a_381_47# VGND 0.101f
C18512 _340_/a_1602_47# VGND 0.229f
C18513 _340_/a_1032_413# VGND 0.463f
C18514 _340_/a_1182_261# VGND 0.191f
C18515 _340_/a_476_47# VGND 0.487f
C18516 _340_/a_652_21# VGND 0.212f
C18517 _340_/a_193_47# VGND 0.559f
C18518 _340_/a_27_47# VGND 0.634f
C18519 _271_/a_75_212# VGND 0.323f
C18520 output14/a_27_47# VGND 0.74f
C18521 output25/a_27_47# VGND 0.431f
C18522 output36/a_27_47# VGND 0.772f
C18523 _307_/a_1462_47# VGND 0.00248f
C18524 _307_/a_1217_47# VGND 0.00103f
C18525 _307_/a_805_47# VGND 0.00613f
C18526 _307_/a_639_47# VGND 0.00927f
C18527 _307_/a_1270_413# VGND 3.88e-20
C18528 _307_/a_651_413# VGND 0.00839f
C18529 _307_/a_448_47# VGND 0.0836f
C18530 _307_/a_1108_47# VGND 0.303f
C18531 _307_/a_1283_21# VGND 0.557f
C18532 _307_/a_543_47# VGND 0.296f
C18533 _307_/a_761_289# VGND 0.212f
C18534 _307_/a_193_47# VGND 0.363f
C18535 _307_/a_27_47# VGND 0.803f
C18536 _238_/a_75_212# VGND 0.345f
C18537 _169_/a_373_53# VGND 0.00247f
C18538 _169_/a_301_53# VGND 4.78e-19
C18539 _169_/a_109_53# VGND 0.218f
C18540 _169_/a_215_311# VGND 0.383f
C18541 _324_/a_1462_47# VGND 0.00233f
C18542 _324_/a_1217_47# VGND 0.00103f
C18543 _324_/a_805_47# VGND 0.00602f
C18544 _324_/a_639_47# VGND 0.00915f
C18545 _324_/a_1270_413# VGND 3.52e-20
C18546 _324_/a_651_413# VGND 0.0084f
C18547 _324_/a_448_47# VGND 0.084f
C18548 _324_/a_1108_47# VGND 0.292f
C18549 _324_/a_1283_21# VGND 0.554f
C18550 _324_/a_543_47# VGND 0.295f
C18551 _324_/a_761_289# VGND 0.21f
C18552 _324_/a_193_47# VGND 0.364f
C18553 _324_/a_27_47# VGND 0.766f
C18554 _255_/a_27_47# VGND 0.322f
C18555 _186_/a_109_297# VGND 9.13e-20
C18556 _341_/a_1462_47# VGND 0.00143f
C18557 _341_/a_1217_47# VGND 5.76e-19
C18558 _341_/a_805_47# VGND 0.00631f
C18559 _341_/a_639_47# VGND 0.00976f
C18560 _341_/a_1270_413# VGND 8.12e-20
C18561 _341_/a_651_413# VGND 0.00878f
C18562 _341_/a_448_47# VGND 0.0749f
C18563 _341_/a_1108_47# VGND 0.284f
C18564 _341_/a_1283_21# VGND 0.551f
C18565 _341_/a_543_47# VGND 0.309f
C18566 _341_/a_761_289# VGND 0.209f
C18567 _341_/a_193_47# VGND 0.374f
C18568 _341_/a_27_47# VGND 0.777f
C18569 _272_/a_384_47# VGND 0.00343f
C18570 _272_/a_299_297# VGND 0.0407f
C18571 _272_/a_81_21# VGND 0.319f
C18572 output13/a_27_47# VGND 0.797f
C18573 output24/a_27_47# VGND 0.755f
C18574 output35/a_27_47# VGND 0.764f
C18575 _308_/a_1462_47# VGND 0.00236f
C18576 _308_/a_1217_47# VGND 4.86e-19
C18577 _308_/a_805_47# VGND 0.00596f
C18578 _308_/a_639_47# VGND 0.00895f
C18579 _308_/a_1270_413# VGND 3.11e-20
C18580 _308_/a_651_413# VGND 0.00526f
C18581 _308_/a_448_47# VGND 0.0809f
C18582 _308_/a_1108_47# VGND 0.28f
C18583 _308_/a_1283_21# VGND 0.552f
C18584 _308_/a_543_47# VGND 0.283f
C18585 _308_/a_761_289# VGND 0.196f
C18586 _308_/a_193_47# VGND 0.34f
C18587 _308_/a_27_47# VGND 0.792f
C18588 _239_/a_474_297# VGND 0.0377f
C18589 _239_/a_277_297# VGND 0.0226f
C18590 _239_/a_27_297# VGND 0.0517f
C18591 _239_/a_694_21# VGND 0.44f
C18592 _325_/a_1462_47# VGND 0.00127f
C18593 _325_/a_1217_47# VGND 4.65e-19
C18594 _325_/a_805_47# VGND 0.00509f
C18595 _325_/a_639_47# VGND 0.00713f
C18596 _325_/a_651_413# VGND 0.00788f
C18597 _325_/a_448_47# VGND 0.075f
C18598 _325_/a_1108_47# VGND 0.28f
C18599 _325_/a_1283_21# VGND 0.555f
C18600 _325_/a_543_47# VGND 0.299f
C18601 _325_/a_761_289# VGND 0.205f
C18602 _325_/a_193_47# VGND 0.36f
C18603 _325_/a_27_47# VGND 0.702f
C18604 _256_/a_373_47# VGND 0.00282f
C18605 _256_/a_109_47# VGND 0.00645f
C18606 _256_/a_109_297# VGND 0.00531f
C18607 _256_/a_27_297# VGND 0.454f
C18608 _187_/a_297_47# VGND 0.00703f
C18609 _187_/a_212_413# VGND 0.422f
C18610 _187_/a_27_413# VGND 0.335f
C18611 _273_/a_145_75# VGND 0.00339f
C18612 _273_/a_59_75# VGND 0.284f
C18613 _290_/a_297_47# VGND 0.00528f
C18614 _290_/a_207_413# VGND 0.247f
C18615 _290_/a_27_413# VGND 0.282f
C18616 output12/a_27_47# VGND 0.824f
C18617 output23/a_27_47# VGND 0.453f
C18618 output34/a_27_47# VGND 0.75f
C18619 _309_/a_1462_47# VGND 0.00145f
C18620 _309_/a_1217_47# VGND 4.65e-19
C18621 _309_/a_805_47# VGND 0.00628f
C18622 _309_/a_639_47# VGND 0.00941f
C18623 _309_/a_651_413# VGND 0.008f
C18624 _309_/a_448_47# VGND 0.083f
C18625 _309_/a_1108_47# VGND 0.28f
C18626 _309_/a_1283_21# VGND 0.53f
C18627 _309_/a_543_47# VGND 0.306f
C18628 _309_/a_761_289# VGND 0.212f
C18629 _309_/a_193_47# VGND 0.355f
C18630 _309_/a_27_47# VGND 0.818f
C18631 _326_/a_1462_47# VGND 0.00221f
C18632 _326_/a_1217_47# VGND 9.68e-19
C18633 _326_/a_805_47# VGND 0.00579f
C18634 _326_/a_639_47# VGND 0.00863f
C18635 _326_/a_651_413# VGND 0.00471f
C18636 _326_/a_448_47# VGND 0.0818f
C18637 _326_/a_1108_47# VGND 0.3f
C18638 _326_/a_1283_21# VGND 0.557f
C18639 _326_/a_543_47# VGND 0.283f
C18640 _326_/a_761_289# VGND 0.194f
C18641 _326_/a_193_47# VGND 0.352f
C18642 _326_/a_27_47# VGND 0.752f
C18643 _257_/a_373_47# VGND 0.00244f
C18644 _257_/a_109_47# VGND 0.00755f
C18645 _257_/a_109_297# VGND 0.00581f
C18646 _257_/a_27_297# VGND 0.443f
C18647 _188_/a_27_47# VGND 0.382f
C18648 _274_/a_75_212# VGND 0.354f
C18649 _291_/a_285_47# VGND 0.00886f
C18650 _291_/a_285_297# VGND 0.0334f
C18651 _291_/a_117_297# VGND 0.00143f
C18652 _291_/a_35_297# VGND 0.467f
C18653 output9/a_27_47# VGND 0.439f
C18654 output11/a_27_47# VGND 0.465f
C18655 output22/a_27_47# VGND 0.464f
C18656 output33/a_27_47# VGND 0.729f
C18657 _327_/a_1462_47# VGND 0.00221f
C18658 _327_/a_1217_47# VGND 0.00102f
C18659 _327_/a_805_47# VGND 0.00596f
C18660 _327_/a_639_47# VGND 0.00901f
C18661 _327_/a_1270_413# VGND 4.68e-20
C18662 _327_/a_651_413# VGND 0.00866f
C18663 _327_/a_448_47# VGND 0.0816f
C18664 _327_/a_1108_47# VGND 0.304f
C18665 _327_/a_1283_21# VGND 0.687f
C18666 _327_/a_543_47# VGND 0.304f
C18667 _327_/a_761_289# VGND 0.212f
C18668 _327_/a_193_47# VGND 0.36f
C18669 _327_/a_27_47# VGND 0.813f
C18670 _258_/a_373_47# VGND 0.00224f
C18671 _258_/a_109_47# VGND 0.00652f
C18672 _258_/a_109_297# VGND 0.00582f
C18673 _258_/a_27_297# VGND 0.45f
C18674 _189_/a_408_47# VGND 0.283f
C18675 _189_/a_218_47# VGND 0.182f
C18676 _189_/a_27_47# VGND 0.422f
C18677 _275_/a_384_47# VGND 0.00344f
C18678 _275_/a_299_297# VGND 0.0408f
C18679 _275_/a_81_21# VGND 0.349f
C18680 _292_/a_215_47# VGND 0.327f
C18681 _292_/a_493_297# VGND 3.14e-20
C18682 _292_/a_292_297# VGND 1.8e-19
C18683 _292_/a_78_199# VGND 0.211f
C18684 output8/a_27_47# VGND 0.479f
C18685 output10/a_27_47# VGND 0.453f
C18686 output21/a_27_47# VGND 0.751f
C18687 output32/a_27_47# VGND 0.752f
C18688 _328_/a_1462_47# VGND 0.00135f
C18689 _328_/a_1217_47# VGND 4.73e-19
C18690 _328_/a_805_47# VGND 0.00613f
C18691 _328_/a_639_47# VGND 0.00936f
C18692 _328_/a_1270_413# VGND 5.15e-20
C18693 _328_/a_651_413# VGND 0.00863f
C18694 _328_/a_448_47# VGND 0.0839f
C18695 _328_/a_1108_47# VGND 0.283f
C18696 _328_/a_1283_21# VGND 0.536f
C18697 _328_/a_543_47# VGND 0.307f
C18698 _328_/a_761_289# VGND 0.213f
C18699 _328_/a_193_47# VGND 0.377f
C18700 _328_/a_27_47# VGND 0.733f
C18701 _259_/a_373_47# VGND 0.00363f
C18702 _259_/a_109_47# VGND 0.00717f
C18703 _259_/a_109_297# VGND 0.0119f
C18704 _259_/a_27_297# VGND 0.459f
C18705 _276_/a_145_75# VGND 0.00466f
C18706 _276_/a_59_75# VGND 0.314f
C18707 _293_/a_384_47# VGND 0.00472f
C18708 _293_/a_299_297# VGND 0.0577f
C18709 _293_/a_81_21# VGND 0.337f
C18710 output7/a_27_47# VGND 0.473f
C18711 output20/a_27_47# VGND 0.746f
C18712 output31/a_27_47# VGND 0.71f
C18713 _329_/a_1462_47# VGND 0.00257f
C18714 _329_/a_1217_47# VGND 0.00104f
C18715 _329_/a_805_47# VGND 0.00639f
C18716 _329_/a_639_47# VGND 0.00988f
C18717 _329_/a_1270_413# VGND 4.28e-20
C18718 _329_/a_651_413# VGND 0.00862f
C18719 _329_/a_448_47# VGND 0.0853f
C18720 _329_/a_1108_47# VGND 0.293f
C18721 _329_/a_1283_21# VGND 0.556f
C18722 _329_/a_543_47# VGND 0.296f
C18723 _329_/a_761_289# VGND 0.213f
C18724 _329_/a_193_47# VGND 0.38f
C18725 _329_/a_27_47# VGND 0.823f
C18726 _200_/a_303_47# VGND 0.00528f
C18727 _200_/a_209_47# VGND 0.00583f
C18728 _200_/a_209_297# VGND 0.00718f
C18729 _200_/a_80_21# VGND 0.405f
C18730 _277_/a_75_212# VGND 0.351f
C18731 _294_/a_150_297# VGND 2.53e-19
C18732 _294_/a_68_297# VGND 0.275f
.ends
