magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< metal3 >>
rect 9 72 211 80
rect 9 8 38 72
rect 102 8 118 72
rect 182 8 211 72
rect 9 0 211 8
<< via3 >>
rect 38 8 102 72
rect 118 8 182 72
<< metal4 >>
rect 9 72 211 88
rect 9 8 38 72
rect 102 8 118 72
rect 182 8 211 72
rect 9 -8 211 8
<< end >>
