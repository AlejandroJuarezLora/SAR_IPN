magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< metal1 >>
rect 20580 6473 20940 6519
rect 22734 6473 23094 6519
rect 21434 5633 21794 5679
rect 21880 4793 22240 4839
rect 20580 3953 20940 3999
rect 22734 3953 23094 3999
<< metal2 >>
rect 800 1156 900 9316
rect 1200 8206 1300 9316
rect 1200 8146 1456 8206
rect 1200 7366 1300 8146
rect 1200 7306 1456 7366
rect 1200 6526 1300 7306
rect 1200 6466 1456 6526
rect 1200 5686 1300 6466
rect 1200 5626 1456 5686
rect 1200 4846 1300 5626
rect 1200 4786 1456 4846
rect 1200 4006 1300 4786
rect 1200 3946 1456 4006
rect 1200 3166 1300 3946
rect 1200 3106 1456 3166
rect 1200 2326 1300 3106
rect 1200 2266 1456 2326
rect 1200 84 1300 2266
rect 2100 1156 2200 9316
rect 2500 8206 2600 9316
rect 2500 8146 2756 8206
rect 2500 7366 2600 8146
rect 2500 7306 2756 7366
rect 2500 6526 2600 7306
rect 2500 6466 2756 6526
rect 2500 5686 2600 6466
rect 2500 5626 2756 5686
rect 2500 4846 2600 5626
rect 2500 4786 2756 4846
rect 2500 4006 2600 4786
rect 2500 3946 2756 4006
rect 2500 3166 2600 3946
rect 2500 3106 2756 3166
rect 2500 2326 2600 3106
rect 2500 2266 2756 2326
rect 2500 244 2600 2266
rect 3400 1156 3500 9316
rect 3800 8206 3900 9316
rect 3800 8146 4056 8206
rect 3800 7366 3900 8146
rect 3800 7306 4056 7366
rect 3800 6526 3900 7306
rect 3800 6466 4056 6526
rect 3800 5686 3900 6466
rect 3800 5626 4056 5686
rect 3800 4846 3900 5626
rect 3800 4786 4056 4846
rect 3800 4006 3900 4786
rect 3800 3946 4056 4006
rect 3800 3166 3900 3946
rect 3800 3106 4056 3166
rect 3800 2326 3900 3106
rect 3800 2266 4056 2326
rect 3800 84 3900 2266
rect 4700 1156 4800 9316
rect 5100 8206 5200 9316
rect 5100 8146 5356 8206
rect 5100 7366 5200 8146
rect 5100 7306 5356 7366
rect 5100 6526 5200 7306
rect 5100 6466 5356 6526
rect 5100 5686 5200 6466
rect 5100 5626 5356 5686
rect 5100 4846 5200 5626
rect 5100 4786 5356 4846
rect 5100 4006 5200 4786
rect 5100 3946 5356 4006
rect 5100 3166 5200 3946
rect 5100 3106 5356 3166
rect 5100 2326 5200 3106
rect 5100 2266 5356 2326
rect 5100 84 5200 2266
rect 6000 1156 6100 9316
rect 6400 8206 6500 9316
rect 6400 8146 6656 8206
rect 6400 7366 6500 8146
rect 6400 7306 6656 7366
rect 6400 6526 6500 7306
rect 6400 6466 6656 6526
rect 6400 5686 6500 6466
rect 6400 5626 6656 5686
rect 6400 4846 6500 5626
rect 6400 4786 6656 4846
rect 6400 4006 6500 4786
rect 6400 3946 6656 4006
rect 6400 3166 6500 3946
rect 6400 3106 6656 3166
rect 6400 2326 6500 3106
rect 6400 2266 6656 2326
rect 6400 244 6500 2266
rect 7300 1156 7400 9316
rect 7700 8206 7800 9316
rect 7700 8146 7956 8206
rect 7700 7366 7800 8146
rect 7700 7306 7956 7366
rect 7700 6526 7800 7306
rect 7700 6466 7956 6526
rect 7700 5686 7800 6466
rect 7700 5626 7956 5686
rect 7700 4846 7800 5626
rect 7700 4786 7956 4846
rect 7700 4006 7800 4786
rect 7700 3946 7956 4006
rect 7700 3166 7800 3946
rect 7700 3106 7956 3166
rect 7700 2326 7800 3106
rect 7700 2266 7956 2326
rect 7700 84 7800 2266
rect 8600 1156 8700 9316
rect 9000 8206 9100 9316
rect 9000 8146 9256 8206
rect 9000 7366 9100 8146
rect 9000 7306 9256 7366
rect 9000 6526 9100 7306
rect 9000 6466 9256 6526
rect 9000 5686 9100 6466
rect 9000 5626 9256 5686
rect 9000 4846 9100 5626
rect 9000 4786 9256 4846
rect 9000 4006 9100 4786
rect 9000 3946 9256 4006
rect 9000 3166 9100 3946
rect 9000 3106 9256 3166
rect 9000 2326 9100 3106
rect 9000 2266 9256 2326
rect 9000 84 9100 2266
rect 9900 1156 10000 9316
rect 10300 8206 10400 9316
rect 10300 8146 10556 8206
rect 10300 7366 10400 8146
rect 10300 7306 10556 7366
rect 10300 6526 10400 7306
rect 10300 6466 10556 6526
rect 10300 5686 10400 6466
rect 10300 5626 10556 5686
rect 10300 4846 10400 5626
rect 10300 4786 10556 4846
rect 10300 4006 10400 4786
rect 10300 3946 10556 4006
rect 10300 3166 10400 3946
rect 10300 3106 10556 3166
rect 10300 2326 10400 3106
rect 10300 2266 10556 2326
rect 10300 324 10400 2266
rect 11200 1156 11300 9316
rect 11600 8206 11700 9316
rect 11600 8146 11856 8206
rect 11600 7366 11700 8146
rect 11600 7306 11856 7366
rect 11600 6526 11700 7306
rect 11600 6466 11856 6526
rect 11600 5686 11700 6466
rect 11600 5626 11856 5686
rect 11600 4846 11700 5626
rect 11600 4786 11856 4846
rect 11600 4006 11700 4786
rect 11600 3946 11856 4006
rect 11600 3166 11700 3946
rect 11600 3106 11856 3166
rect 11600 2326 11700 3106
rect 11600 2266 11856 2326
rect 11600 244 11700 2266
rect 12500 1156 12600 9316
rect 12900 8206 13000 9316
rect 12900 8146 13156 8206
rect 12900 7366 13000 8146
rect 12900 7306 13156 7366
rect 12900 6526 13000 7306
rect 12900 6466 13156 6526
rect 12900 5686 13000 6466
rect 12900 5626 13156 5686
rect 12900 4846 13000 5626
rect 12900 4786 13156 4846
rect 12900 4006 13000 4786
rect 12900 3946 13156 4006
rect 12900 3166 13000 3946
rect 12900 3106 13156 3166
rect 12900 2326 13000 3106
rect 12900 2266 13156 2326
rect 12900 84 13000 2266
rect 13800 1156 13900 9316
rect 14200 8206 14300 9316
rect 14200 8146 14456 8206
rect 14200 7366 14300 8146
rect 14200 7306 14456 7366
rect 14200 6526 14300 7306
rect 14200 6466 14456 6526
rect 14200 5686 14300 6466
rect 14200 5626 14456 5686
rect 14200 4846 14300 5626
rect 14200 4786 14456 4846
rect 14200 4006 14300 4786
rect 14200 3946 14456 4006
rect 14200 3166 14300 3946
rect 14200 3106 14456 3166
rect 14200 2326 14300 3106
rect 14200 2266 14456 2326
rect 14200 84 14300 2266
rect 15100 1156 15200 9316
rect 15500 8206 15600 9316
rect 15500 8146 15756 8206
rect 15500 7366 15600 8146
rect 15500 7306 15756 7366
rect 15500 6526 15600 7306
rect 15500 6466 15756 6526
rect 15500 5686 15600 6466
rect 15500 5626 15756 5686
rect 15500 4846 15600 5626
rect 15500 4786 15756 4846
rect 15500 4006 15600 4786
rect 15500 3946 15756 4006
rect 15500 3166 15600 3946
rect 15500 3106 15756 3166
rect 15500 2326 15600 3106
rect 15500 2266 15756 2326
rect 15500 404 15600 2266
rect 16400 1156 16500 9316
rect 16800 8206 16900 9316
rect 16800 8146 17056 8206
rect 16800 7366 16900 8146
rect 16800 7306 17056 7366
rect 16800 6526 16900 7306
rect 16800 6466 17056 6526
rect 16800 5686 16900 6466
rect 16800 5626 17056 5686
rect 16800 4846 16900 5626
rect 16800 4786 17056 4846
rect 16800 4006 16900 4786
rect 16800 3946 17056 4006
rect 16800 3166 16900 3946
rect 16800 3106 17056 3166
rect 16800 2326 16900 3106
rect 16800 2266 17056 2326
rect 16800 164 16900 2266
rect 17700 1156 17800 9316
rect 18100 8206 18200 9316
rect 18100 8146 18356 8206
rect 18100 7366 18200 8146
rect 18100 7306 18356 7366
rect 18100 6526 18200 7306
rect 18100 6466 18356 6526
rect 18100 5686 18200 6466
rect 18100 5626 18356 5686
rect 18100 4846 18200 5626
rect 18100 4786 18356 4846
rect 18100 4006 18200 4786
rect 18100 3946 18356 4006
rect 18100 3166 18200 3946
rect 18100 3106 18356 3166
rect 18100 2326 18200 3106
rect 18100 2266 18356 2326
rect 18100 84 18200 2266
rect 19000 1156 19100 9316
rect 19400 8206 19500 9316
rect 19400 8146 19656 8206
rect 19400 7366 19500 8146
rect 19400 7306 19656 7366
rect 19400 6526 19500 7306
rect 19400 6466 19656 6526
rect 19400 5686 19500 6466
rect 19400 5626 19656 5686
rect 19400 4846 19500 5626
rect 19400 4786 19656 4846
rect 19400 4006 19500 4786
rect 19400 3946 19656 4006
rect 19400 3166 19500 3946
rect 19400 3106 19656 3166
rect 19400 2326 19500 3106
rect 19400 2266 19656 2326
rect 19400 484 19500 2266
rect 20300 1156 20400 9316
rect 20700 8206 20800 9316
rect 20700 8146 20956 8206
rect 20700 7366 20800 8146
rect 20700 7306 20956 7366
rect 20700 3166 20800 7306
rect 21600 4846 21700 9316
rect 21444 4786 21700 4846
rect 20700 3106 20956 3166
rect 20700 2326 20800 3106
rect 20700 2266 20956 2326
rect 20700 644 20800 2266
rect 21600 1044 21700 4786
rect 22000 5685 22100 9316
rect 22900 8206 23000 9316
rect 22744 8146 23000 8206
rect 22900 7366 23000 8146
rect 22744 7306 23000 7366
rect 22000 5625 22256 5685
rect 22000 1044 22100 5625
rect 22900 3166 23000 7306
rect 22744 3106 23000 3166
rect 22900 2326 23000 3106
rect 22744 2266 23000 2326
rect 21300 -316 21400 1044
rect 21600 964 22100 1044
rect 21800 -156 21900 964
rect 22300 -476 22400 1044
rect 22900 644 23000 2266
rect 23300 1156 23400 9316
rect 24200 8206 24300 9316
rect 24044 8146 24300 8206
rect 24200 7366 24300 8146
rect 24044 7306 24300 7366
rect 24200 6526 24300 7306
rect 24044 6466 24300 6526
rect 24200 5686 24300 6466
rect 24044 5626 24300 5686
rect 24200 4846 24300 5626
rect 24044 4786 24300 4846
rect 24200 4006 24300 4786
rect 24044 3946 24300 4006
rect 24200 3166 24300 3946
rect 24044 3106 24300 3166
rect 24200 2326 24300 3106
rect 24044 2266 24300 2326
rect 24200 484 24300 2266
rect 24600 1156 24700 9316
rect 25500 8206 25600 9316
rect 25344 8146 25600 8206
rect 25500 7366 25600 8146
rect 25344 7306 25600 7366
rect 25500 6526 25600 7306
rect 25344 6466 25600 6526
rect 25500 5686 25600 6466
rect 25344 5626 25600 5686
rect 25500 4846 25600 5626
rect 25344 4786 25600 4846
rect 25500 4006 25600 4786
rect 25344 3946 25600 4006
rect 25500 3166 25600 3946
rect 25344 3106 25600 3166
rect 25500 2326 25600 3106
rect 25344 2266 25600 2326
rect 25500 54 25600 2266
rect 25900 1156 26000 9316
rect 26800 8206 26900 9316
rect 26644 8146 26900 8206
rect 26800 7366 26900 8146
rect 26644 7306 26900 7366
rect 26800 6526 26900 7306
rect 26644 6466 26900 6526
rect 26800 5686 26900 6466
rect 26644 5626 26900 5686
rect 26800 4846 26900 5626
rect 26644 4786 26900 4846
rect 26800 4006 26900 4786
rect 26644 3946 26900 4006
rect 26800 3166 26900 3946
rect 26644 3106 26900 3166
rect 26800 2326 26900 3106
rect 26644 2266 26900 2326
rect 26800 164 26900 2266
rect 27200 1156 27300 9316
rect 28100 8206 28200 9316
rect 27944 8146 28200 8206
rect 28100 7366 28200 8146
rect 27944 7306 28200 7366
rect 28100 6526 28200 7306
rect 27944 6466 28200 6526
rect 28100 5686 28200 6466
rect 27944 5626 28200 5686
rect 28100 4846 28200 5626
rect 27944 4786 28200 4846
rect 28100 4006 28200 4786
rect 27944 3946 28200 4006
rect 28100 3166 28200 3946
rect 27944 3106 28200 3166
rect 28100 2326 28200 3106
rect 27944 2266 28200 2326
rect 28100 324 28200 2266
rect 28500 1156 28600 9316
rect 29400 8206 29500 9316
rect 29244 8146 29500 8206
rect 29400 7366 29500 8146
rect 29244 7306 29500 7366
rect 29400 6526 29500 7306
rect 29244 6466 29500 6526
rect 29400 5686 29500 6466
rect 29244 5626 29500 5686
rect 29400 4846 29500 5626
rect 29244 4786 29500 4846
rect 29400 4006 29500 4786
rect 29244 3946 29500 4006
rect 29400 3166 29500 3946
rect 29244 3106 29500 3166
rect 29400 2326 29500 3106
rect 29244 2266 29500 2326
rect 25499 5 25600 54
rect 25500 4 25600 5
rect 29400 4 29500 2266
rect 29800 1156 29900 9316
rect 30700 8206 30800 9316
rect 30544 8146 30800 8206
rect 30700 7366 30800 8146
rect 30544 7306 30800 7366
rect 30700 6526 30800 7306
rect 30544 6466 30800 6526
rect 30700 5686 30800 6466
rect 30544 5626 30800 5686
rect 30700 4846 30800 5626
rect 30544 4786 30800 4846
rect 30700 4006 30800 4786
rect 30544 3946 30800 4006
rect 30700 3166 30800 3946
rect 30544 3106 30800 3166
rect 30700 2326 30800 3106
rect 30544 2266 30800 2326
rect 30700 4 30800 2266
rect 31100 1156 31200 9316
rect 32000 8206 32100 9316
rect 31844 8146 32100 8206
rect 32000 7366 32100 8146
rect 31844 7306 32100 7366
rect 32000 6526 32100 7306
rect 31844 6466 32100 6526
rect 32000 5686 32100 6466
rect 31844 5626 32100 5686
rect 32000 4846 32100 5626
rect 31844 4786 32100 4846
rect 32000 4006 32100 4786
rect 31844 3946 32100 4006
rect 32000 3166 32100 3946
rect 31844 3106 32100 3166
rect 32000 2326 32100 3106
rect 31844 2266 32100 2326
rect 32000 164 32100 2266
rect 32400 1156 32500 9316
rect 33300 8206 33400 9316
rect 33144 8146 33400 8206
rect 33300 7366 33400 8146
rect 33144 7306 33400 7366
rect 33300 6526 33400 7306
rect 33144 6466 33400 6526
rect 33300 5686 33400 6466
rect 33144 5626 33400 5686
rect 33300 4846 33400 5626
rect 33144 4786 33400 4846
rect 33300 4006 33400 4786
rect 33144 3946 33400 4006
rect 33300 3166 33400 3946
rect 33144 3106 33400 3166
rect 33300 2326 33400 3106
rect 33144 2266 33400 2326
rect 33300 324 33400 2266
rect 33700 1156 33800 9316
rect 34600 8206 34700 9316
rect 34444 8146 34700 8206
rect 34600 7366 34700 8146
rect 34444 7306 34700 7366
rect 34600 6526 34700 7306
rect 34444 6466 34700 6526
rect 34600 5686 34700 6466
rect 34444 5626 34700 5686
rect 34600 4846 34700 5626
rect 34444 4786 34700 4846
rect 34600 4006 34700 4786
rect 34444 3946 34700 4006
rect 34600 3166 34700 3946
rect 34444 3106 34700 3166
rect 34600 2326 34700 3106
rect 34444 2266 34700 2326
rect 34600 4 34700 2266
rect 35000 1156 35100 9316
rect 35900 8206 36000 9316
rect 35744 8146 36000 8206
rect 35900 7366 36000 8146
rect 35744 7306 36000 7366
rect 35900 6526 36000 7306
rect 35744 6466 36000 6526
rect 35900 5686 36000 6466
rect 35744 5626 36000 5686
rect 35900 4846 36000 5626
rect 35744 4786 36000 4846
rect 35900 4006 36000 4786
rect 35744 3946 36000 4006
rect 35900 3166 36000 3946
rect 35744 3106 36000 3166
rect 35900 2326 36000 3106
rect 35744 2266 36000 2326
rect 35900 4 36000 2266
rect 36300 1156 36400 9316
rect 37200 8206 37300 9316
rect 37044 8146 37300 8206
rect 37200 7366 37300 8146
rect 37044 7306 37300 7366
rect 37200 6526 37300 7306
rect 37044 6466 37300 6526
rect 37200 5686 37300 6466
rect 37044 5626 37300 5686
rect 37200 4846 37300 5626
rect 37044 4786 37300 4846
rect 37200 4006 37300 4786
rect 37044 3946 37300 4006
rect 37200 3166 37300 3946
rect 37044 3106 37300 3166
rect 37200 2326 37300 3106
rect 37044 2266 37300 2326
rect 37200 164 37300 2266
rect 37600 1156 37700 9316
rect 38500 8206 38600 9316
rect 38344 8146 38600 8206
rect 38500 7366 38600 8146
rect 38344 7306 38600 7366
rect 38500 6526 38600 7306
rect 38344 6466 38600 6526
rect 38500 5686 38600 6466
rect 38344 5626 38600 5686
rect 38500 4846 38600 5626
rect 38344 4786 38600 4846
rect 38500 4006 38600 4786
rect 38344 3946 38600 4006
rect 38500 3166 38600 3946
rect 38344 3106 38600 3166
rect 38500 2326 38600 3106
rect 38344 2266 38600 2326
rect 38500 4 38600 2266
rect 38900 1156 39000 9316
rect 39800 8206 39900 9316
rect 39644 8146 39900 8206
rect 39800 7366 39900 8146
rect 39644 7306 39900 7366
rect 39800 6526 39900 7306
rect 39644 6466 39900 6526
rect 39800 5686 39900 6466
rect 39644 5626 39900 5686
rect 39800 4846 39900 5626
rect 39644 4786 39900 4846
rect 39800 4006 39900 4786
rect 39644 3946 39900 4006
rect 39800 3166 39900 3946
rect 39644 3106 39900 3166
rect 39800 2326 39900 3106
rect 39644 2266 39900 2326
rect 39800 4 39900 2266
rect 40200 1156 40300 9316
rect 41100 8206 41200 9316
rect 40944 8146 41200 8206
rect 41100 7366 41200 8146
rect 40944 7306 41200 7366
rect 41100 6526 41200 7306
rect 40944 6466 41200 6526
rect 41100 5686 41200 6466
rect 40944 5626 41200 5686
rect 41100 4846 41200 5626
rect 40944 4786 41200 4846
rect 41100 4006 41200 4786
rect 40944 3946 41200 4006
rect 41100 3166 41200 3946
rect 40944 3106 41200 3166
rect 41100 2326 41200 3106
rect 40944 2266 41200 2326
rect 41100 164 41200 2266
rect 41500 1156 41600 9316
rect 42400 8206 42500 9316
rect 42244 8146 42500 8206
rect 42400 7366 42500 8146
rect 42244 7306 42500 7366
rect 42400 6526 42500 7306
rect 42244 6466 42500 6526
rect 42400 5686 42500 6466
rect 42244 5626 42500 5686
rect 42400 4846 42500 5626
rect 42244 4786 42500 4846
rect 42400 4006 42500 4786
rect 42244 3946 42500 4006
rect 42400 3166 42500 3946
rect 42244 3106 42500 3166
rect 42400 2326 42500 3106
rect 42244 2266 42500 2326
rect 42400 4 42500 2266
rect 42800 1156 42900 9316
<< metal3 >>
rect 900 1156 1000 9316
rect 1100 1156 1200 9316
rect 2200 1156 2300 9316
rect 2400 1156 2500 9316
rect 3500 1156 3600 9316
rect 3700 1156 3800 9316
rect 4800 1156 4900 9316
rect 5000 1156 5100 9316
rect 6100 1156 6200 9316
rect 6300 1156 6400 9316
rect 7400 1156 7500 9316
rect 7600 1156 7700 9316
rect 8700 1156 8800 9316
rect 8900 1156 9000 9316
rect 10000 1156 10100 9316
rect 10200 1156 10300 9316
rect 11300 1156 11400 9316
rect 11500 1156 11600 9316
rect 12600 1156 12700 9316
rect 12800 1156 12900 9316
rect 13900 1156 14000 9316
rect 14100 1156 14200 9316
rect 15200 1156 15300 9316
rect 15400 1156 15500 9316
rect 16500 1156 16600 9316
rect 16700 1156 16800 9316
rect 17800 1156 17900 9316
rect 18000 1156 18100 9316
rect 19100 1156 19200 9316
rect 19300 1156 19400 9316
rect 20400 1156 20500 9316
rect 20600 884 20700 9316
rect 21700 1044 21800 9316
rect 21460 964 21800 1044
rect 21900 1044 22000 9316
rect 21900 964 22240 1044
rect 23000 884 23100 9316
rect 23200 1156 23300 9316
rect 24300 1156 24400 9316
rect 24500 1156 24600 9316
rect 25600 1156 25700 9316
rect 25800 1156 25900 9316
rect 26900 1156 27000 9316
rect 27100 1156 27200 9316
rect 28200 1156 28300 9316
rect 28400 1156 28500 9316
rect 29500 1156 29600 9316
rect 29700 1156 29800 9316
rect 30800 1156 30900 9316
rect 31000 1156 31100 9316
rect 32100 1156 32200 9316
rect 32300 1156 32400 9316
rect 33400 1156 33500 9316
rect 33600 1156 33700 9316
rect 34700 1156 34800 9316
rect 34900 1156 35000 9316
rect 36000 1156 36100 9316
rect 36200 1156 36300 9316
rect 37300 1156 37400 9316
rect 37500 1156 37600 9316
rect 38600 1156 38700 9316
rect 38800 1156 38900 9316
rect 39900 1156 40000 9316
rect 40100 1156 40200 9316
rect 41200 1156 41300 9316
rect 41400 1156 41500 9316
rect 42500 1156 42600 9316
rect 42700 1156 42800 9316
rect 0 804 23100 884
rect 0 644 22840 724
rect 0 484 24140 564
rect 0 324 33400 404
rect 0 164 41191 244
rect 0 4 42490 84
rect 0 -156 21900 -76
rect 0 -316 21400 -236
rect 0 -476 22400 -396
<< metal4 >>
rect 352 9416 43700 9516
rect 352 1256 448 9416
rect 1652 1256 1748 9416
rect 2952 1256 3048 9416
rect 4252 1256 4348 9416
rect 5552 1256 5648 9416
rect 6852 1256 6948 9416
rect 8152 1256 8248 9416
rect 9452 1256 9548 9416
rect 10752 1256 10848 9416
rect 12052 1256 12148 9416
rect 13352 1256 13448 9416
rect 14652 1256 14748 9416
rect 15952 1256 16048 9416
rect 17252 1256 17348 9416
rect 18552 1256 18648 9416
rect 19852 1256 19948 9416
rect 21152 1256 21248 9416
rect 22452 1256 22548 9416
rect 23752 1256 23848 9416
rect 25052 1256 25148 9416
rect 26352 1256 26448 9416
rect 27652 1256 27748 9416
rect 28952 1256 29048 9416
rect 30252 1256 30348 9416
rect 31552 1256 31648 9416
rect 32852 1256 32948 9416
rect 34152 1256 34248 9416
rect 35452 1256 35548 9416
rect 36752 1256 36848 9416
rect 38052 1256 38148 9416
rect 39352 1256 39448 9416
rect 40652 1256 40748 9416
rect 41952 1256 42048 9416
rect 43252 1256 43348 9416
use C0_1  C0_1_0
timestamp 1696364841
transform 1 0 21250 0 1 5696
box -450 -340 350 260
use C1  C1_0
timestamp 1696364841
transform 1 0 21250 0 1 4856
box -450 -340 350 260
use C1  C1_1
timestamp 1696364841
transform 1 0 22550 0 1 5696
box -450 -340 350 260
use C2  C2_0
timestamp 1696364841
transform 1 0 21250 0 1 4016
box -450 -340 350 260
use C2  C2_1
timestamp 1696364841
transform 1 0 21250 0 1 6536
box -450 -340 350 260
use C2  C2_2
timestamp 1696364841
transform 1 0 22550 0 1 4016
box -450 -340 350 260
use C2  C2_3
timestamp 1696364841
transform 1 0 22550 0 1 6536
box -450 -340 350 260
use C3  C3_0
timestamp 1696364841
transform 1 0 21250 0 1 3176
box -450 -340 350 260
use C3  C3_1
timestamp 1696364841
transform 1 0 21250 0 1 2336
box -450 -340 350 260
use C3  C3_2
timestamp 1696364841
transform 1 0 21250 0 1 7376
box -450 -340 350 260
use C3  C3_3
timestamp 1696364841
transform 1 0 21250 0 1 8216
box -450 -340 350 260
use C3  C3_4
timestamp 1696364841
transform 1 0 22550 0 1 2336
box -450 -340 350 260
use C3  C3_5
timestamp 1696364841
transform 1 0 22550 0 1 3176
box -450 -340 350 260
use C3  C3_6
timestamp 1696364841
transform 1 0 22550 0 1 8216
box -450 -340 350 260
use C3  C3_7
timestamp 1696364841
transform 1 0 22550 0 1 7376
box -450 -340 350 260
use C4  C4_0
timestamp 1696364841
transform 1 0 19950 0 1 2336
box -450 -340 350 260
use C4  C4_1
timestamp 1696364841
transform 1 0 19950 0 1 3176
box -450 -340 350 260
use C4  C4_2
timestamp 1696364841
transform 1 0 19950 0 1 4016
box -450 -340 350 260
use C4  C4_3
timestamp 1696364841
transform 1 0 19950 0 1 5696
box -450 -340 350 260
use C4  C4_4
timestamp 1696364841
transform 1 0 19950 0 1 4856
box -450 -340 350 260
use C4  C4_5
timestamp 1696364841
transform 1 0 19950 0 1 6536
box -450 -340 350 260
use C4  C4_6
timestamp 1696364841
transform 1 0 19950 0 1 7376
box -450 -340 350 260
use C4  C4_7
timestamp 1696364841
transform 1 0 19950 0 1 8216
box -450 -340 350 260
use C4  C4_8
timestamp 1696364841
transform 1 0 23850 0 1 4016
box -450 -340 350 260
use C4  C4_9
timestamp 1696364841
transform 1 0 23850 0 1 2336
box -450 -340 350 260
use C4  C4_10
timestamp 1696364841
transform 1 0 23850 0 1 3176
box -450 -340 350 260
use C4  C4_11
timestamp 1696364841
transform 1 0 23850 0 1 4856
box -450 -340 350 260
use C4  C4_12
timestamp 1696364841
transform 1 0 23850 0 1 5696
box -450 -340 350 260
use C4  C4_13
timestamp 1696364841
transform 1 0 23850 0 1 6536
box -450 -340 350 260
use C4  C4_14
timestamp 1696364841
transform 1 0 23850 0 1 8216
box -450 -340 350 260
use C4  C4_15
timestamp 1696364841
transform 1 0 23850 0 1 7376
box -450 -340 350 260
use C5  C5_0
timestamp 1696364841
transform 1 0 16050 0 1 3176
box -450 -340 350 260
use C5  C5_1
timestamp 1696364841
transform 1 0 16050 0 1 2336
box -450 -340 350 260
use C5  C5_2
timestamp 1696364841
transform 1 0 16050 0 1 4016
box -450 -340 350 260
use C5  C5_3
timestamp 1696364841
transform 1 0 16050 0 1 8216
box -450 -340 350 260
use C5  C5_4
timestamp 1696364841
transform 1 0 16050 0 1 7376
box -450 -340 350 260
use C5  C5_5
timestamp 1696364841
transform 1 0 16050 0 1 4856
box -450 -340 350 260
use C5  C5_6
timestamp 1696364841
transform 1 0 16050 0 1 6536
box -450 -340 350 260
use C5  C5_7
timestamp 1696364841
transform 1 0 16050 0 1 5696
box -450 -340 350 260
use C5  C5_8
timestamp 1696364841
transform 1 0 10850 0 1 5696
box -450 -340 350 260
use C5  C5_9
timestamp 1696364841
transform 1 0 10850 0 1 6536
box -450 -340 350 260
use C5  C5_10
timestamp 1696364841
transform 1 0 10850 0 1 7376
box -450 -340 350 260
use C5  C5_11
timestamp 1696364841
transform 1 0 10850 0 1 8216
box -450 -340 350 260
use C5  C5_12
timestamp 1696364841
transform 1 0 10850 0 1 4016
box -450 -340 350 260
use C5  C5_13
timestamp 1696364841
transform 1 0 10850 0 1 3176
box -450 -340 350 260
use C5  C5_14
timestamp 1696364841
transform 1 0 10850 0 1 2336
box -450 -340 350 260
use C5  C5_15
timestamp 1696364841
transform 1 0 10850 0 1 4856
box -450 -340 350 260
use C5  C5_16
timestamp 1696364841
transform 1 0 27750 0 1 3176
box -450 -340 350 260
use C5  C5_17
timestamp 1696364841
transform 1 0 27750 0 1 2336
box -450 -340 350 260
use C5  C5_18
timestamp 1696364841
transform 1 0 27750 0 1 4016
box -450 -340 350 260
use C5  C5_19
timestamp 1696364841
transform 1 0 27750 0 1 7376
box -450 -340 350 260
use C5  C5_20
timestamp 1696364841
transform 1 0 27750 0 1 5696
box -450 -340 350 260
use C5  C5_21
timestamp 1696364841
transform 1 0 27750 0 1 6536
box -450 -340 350 260
use C5  C5_22
timestamp 1696364841
transform 1 0 27750 0 1 8216
box -450 -340 350 260
use C5  C5_23
timestamp 1696364841
transform 1 0 27750 0 1 4856
box -450 -340 350 260
use C5  C5_24
timestamp 1696364841
transform 1 0 32950 0 1 6536
box -450 -340 350 260
use C5  C5_25
timestamp 1696364841
transform 1 0 32950 0 1 5696
box -450 -340 350 260
use C5  C5_26
timestamp 1696364841
transform 1 0 32950 0 1 4016
box -450 -340 350 260
use C5  C5_27
timestamp 1696364841
transform 1 0 32950 0 1 3176
box -450 -340 350 260
use C5  C5_28
timestamp 1696364841
transform 1 0 32950 0 1 4856
box -450 -340 350 260
use C5  C5_29
timestamp 1696364841
transform 1 0 32950 0 1 2336
box -450 -340 350 260
use C5  C5_30
timestamp 1696364841
transform 1 0 32950 0 1 8216
box -450 -340 350 260
use C5  C5_31
timestamp 1696364841
transform 1 0 32950 0 1 7376
box -450 -340 350 260
use C6  C6_0
timestamp 1696364841
transform 1 0 12150 0 1 3176
box -450 -340 350 260
use C6  C6_1
timestamp 1696364841
transform 1 0 12150 0 1 4016
box -450 -340 350 260
use C6  C6_2
timestamp 1696364841
transform 1 0 12150 0 1 2336
box -450 -340 350 260
use C6  C6_3
timestamp 1696364841
transform 1 0 17350 0 1 2336
box -450 -340 350 260
use C6  C6_4
timestamp 1696364841
transform 1 0 17350 0 1 3176
box -450 -340 350 260
use C6  C6_5
timestamp 1696364841
transform 1 0 17350 0 1 4016
box -450 -340 350 260
use C6  C6_6
timestamp 1696364841
transform 1 0 3050 0 1 3176
box -450 -340 350 260
use C6  C6_7
timestamp 1696364841
transform 1 0 3050 0 1 4016
box -450 -340 350 260
use C6  C6_8
timestamp 1696364841
transform 1 0 3050 0 1 2336
box -450 -340 350 260
use C6  C6_9
timestamp 1696364841
transform 1 0 6950 0 1 4016
box -450 -340 350 260
use C6  C6_10
timestamp 1696364841
transform 1 0 6950 0 1 2336
box -450 -340 350 260
use C6  C6_11
timestamp 1696364841
transform 1 0 6950 0 1 3176
box -450 -340 350 260
use C6  C6_12
timestamp 1696364841
transform 1 0 6950 0 1 6536
box -450 -340 350 260
use C6  C6_13
timestamp 1696364841
transform 1 0 6950 0 1 4856
box -450 -340 350 260
use C6  C6_14
timestamp 1696364841
transform 1 0 6950 0 1 5696
box -450 -340 350 260
use C6  C6_15
timestamp 1696364841
transform 1 0 3050 0 1 4856
box -450 -340 350 260
use C6  C6_16
timestamp 1696364841
transform 1 0 3050 0 1 6536
box -450 -340 350 260
use C6  C6_17
timestamp 1696364841
transform 1 0 3050 0 1 5696
box -450 -340 350 260
use C6  C6_18
timestamp 1696364841
transform 1 0 3050 0 1 8216
box -450 -340 350 260
use C6  C6_19
timestamp 1696364841
transform 1 0 3050 0 1 7376
box -450 -340 350 260
use C6  C6_20
timestamp 1696364841
transform 1 0 6950 0 1 8216
box -450 -340 350 260
use C6  C6_21
timestamp 1696364841
transform 1 0 6950 0 1 7376
box -450 -340 350 260
use C6  C6_22
timestamp 1696364841
transform 1 0 17350 0 1 5696
box -450 -340 350 260
use C6  C6_23
timestamp 1696364841
transform 1 0 17350 0 1 4856
box -450 -340 350 260
use C6  C6_24
timestamp 1696364841
transform 1 0 17350 0 1 6536
box -450 -340 350 260
use C6  C6_25
timestamp 1696364841
transform 1 0 12150 0 1 4856
box -450 -340 350 260
use C6  C6_26
timestamp 1696364841
transform 1 0 12150 0 1 5696
box -450 -340 350 260
use C6  C6_27
timestamp 1696364841
transform 1 0 12150 0 1 6536
box -450 -340 350 260
use C6  C6_28
timestamp 1696364841
transform 1 0 12150 0 1 8216
box -450 -340 350 260
use C6  C6_29
timestamp 1696364841
transform 1 0 12150 0 1 7376
box -450 -340 350 260
use C6  C6_30
timestamp 1696364841
transform 1 0 17350 0 1 8216
box -450 -340 350 260
use C6  C6_31
timestamp 1696364841
transform 1 0 17350 0 1 7376
box -450 -340 350 260
use C6  C6_32
timestamp 1696364841
transform 1 0 36850 0 1 2336
box -450 -340 350 260
use C6  C6_33
timestamp 1696364841
transform 1 0 36850 0 1 4016
box -450 -340 350 260
use C6  C6_34
timestamp 1696364841
transform 1 0 36850 0 1 3176
box -450 -340 350 260
use C6  C6_35
timestamp 1696364841
transform 1 0 40750 0 1 4016
box -450 -340 350 260
use C6  C6_36
timestamp 1696364841
transform 1 0 40750 0 1 3176
box -450 -340 350 260
use C6  C6_37
timestamp 1696364841
transform 1 0 40750 0 1 2336
box -450 -340 350 260
use C6  C6_38
timestamp 1696364841
transform 1 0 26450 0 1 4016
box -450 -340 350 260
use C6  C6_39
timestamp 1696364841
transform 1 0 26450 0 1 2336
box -450 -340 350 260
use C6  C6_40
timestamp 1696364841
transform 1 0 26450 0 1 3176
box -450 -340 350 260
use C6  C6_41
timestamp 1696364841
transform 1 0 31650 0 1 4016
box -450 -340 350 260
use C6  C6_42
timestamp 1696364841
transform 1 0 31650 0 1 2336
box -450 -340 350 260
use C6  C6_43
timestamp 1696364841
transform 1 0 31650 0 1 3176
box -450 -340 350 260
use C6  C6_44
timestamp 1696364841
transform 1 0 31650 0 1 6536
box -450 -340 350 260
use C6  C6_45
timestamp 1696364841
transform 1 0 31650 0 1 4856
box -450 -340 350 260
use C6  C6_46
timestamp 1696364841
transform 1 0 31650 0 1 5696
box -450 -340 350 260
use C6  C6_47
timestamp 1696364841
transform 1 0 26450 0 1 6536
box -450 -340 350 260
use C6  C6_48
timestamp 1696364841
transform 1 0 26450 0 1 5696
box -450 -340 350 260
use C6  C6_49
timestamp 1696364841
transform 1 0 26450 0 1 4856
box -450 -340 350 260
use C6  C6_50
timestamp 1696364841
transform 1 0 26450 0 1 7376
box -450 -340 350 260
use C6  C6_51
timestamp 1696364841
transform 1 0 26450 0 1 8216
box -450 -340 350 260
use C6  C6_52
timestamp 1696364841
transform 1 0 31650 0 1 8216
box -450 -340 350 260
use C6  C6_53
timestamp 1696364841
transform 1 0 31650 0 1 7376
box -450 -340 350 260
use C6  C6_54
timestamp 1696364841
transform 1 0 40750 0 1 5696
box -450 -340 350 260
use C6  C6_55
timestamp 1696364841
transform 1 0 40750 0 1 4856
box -450 -340 350 260
use C6  C6_56
timestamp 1696364841
transform 1 0 40750 0 1 6536
box -450 -340 350 260
use C6  C6_57
timestamp 1696364841
transform 1 0 36850 0 1 6536
box -450 -340 350 260
use C6  C6_58
timestamp 1696364841
transform 1 0 36850 0 1 4856
box -450 -340 350 260
use C6  C6_59
timestamp 1696364841
transform 1 0 36850 0 1 5696
box -450 -340 350 260
use C6  C6_60
timestamp 1696364841
transform 1 0 36850 0 1 7376
box -450 -340 350 260
use C6  C6_61
timestamp 1696364841
transform 1 0 36850 0 1 8216
box -450 -340 350 260
use C6  C6_62
timestamp 1696364841
transform 1 0 40750 0 1 7376
box -450 -340 350 260
use C6  C6_63
timestamp 1696364841
transform 1 0 40750 0 1 8216
box -450 -340 350 260
use C7  C7_0
timestamp 1696364841
transform 1 0 14750 0 1 3176
box -450 -340 350 260
use C7  C7_1
timestamp 1696364841
transform 1 0 13450 0 1 3176
box -450 -340 350 260
use C7  C7_2
timestamp 1696364841
transform 1 0 14750 0 1 4016
box -450 -340 350 260
use C7  C7_3
timestamp 1696364841
transform 1 0 13450 0 1 4016
box -450 -340 350 260
use C7  C7_4
timestamp 1696364841
transform 1 0 14750 0 1 2336
box -450 -340 350 260
use C7  C7_5
timestamp 1696364841
transform 1 0 13450 0 1 2336
box -450 -340 350 260
use C7  C7_6
timestamp 1696364841
transform 1 0 18650 0 1 2336
box -450 -340 350 260
use C7  C7_7
timestamp 1696364841
transform 1 0 18650 0 1 3176
box -450 -340 350 260
use C7  C7_8
timestamp 1696364841
transform 1 0 18650 0 1 4016
box -450 -340 350 260
use C7  C7_9
timestamp 1696364841
transform 1 0 4350 0 1 4016
box -450 -340 350 260
use C7  C7_10
timestamp 1696364841
transform 1 0 4350 0 1 3176
box -450 -340 350 260
use C7  C7_11
timestamp 1696364841
transform 1 0 1750 0 1 3176
box -450 -340 350 260
use C7  C7_12
timestamp 1696364841
transform 1 0 1750 0 1 2336
box -450 -340 350 260
use C7  C7_13
timestamp 1696364841
transform 1 0 1750 0 1 4016
box -450 -340 350 260
use C7  C7_14
timestamp 1696364841
transform 1 0 4350 0 1 2336
box -450 -340 350 260
use C7  C7_15
timestamp 1696364841
transform 1 0 9550 0 1 4016
box -450 -340 350 260
use C7  C7_16
timestamp 1696364841
transform 1 0 8250 0 1 4016
box -450 -340 350 260
use C7  C7_17
timestamp 1696364841
transform 1 0 9550 0 1 2336
box -450 -340 350 260
use C7  C7_18
timestamp 1696364841
transform 1 0 8250 0 1 2336
box -450 -340 350 260
use C7  C7_19
timestamp 1696364841
transform 1 0 9550 0 1 3176
box -450 -340 350 260
use C7  C7_20
timestamp 1696364841
transform 1 0 8250 0 1 3176
box -450 -340 350 260
use C7  C7_21
timestamp 1696364841
transform 1 0 5650 0 1 3176
box -450 -340 350 260
use C7  C7_22
timestamp 1696364841
transform 1 0 5650 0 1 4016
box -450 -340 350 260
use C7  C7_23
timestamp 1696364841
transform 1 0 5650 0 1 2336
box -450 -340 350 260
use C7  C7_24
timestamp 1696364841
transform 1 0 9550 0 1 5696
box -450 -340 350 260
use C7  C7_25
timestamp 1696364841
transform 1 0 8250 0 1 5696
box -450 -340 350 260
use C7  C7_26
timestamp 1696364841
transform 1 0 9550 0 1 6536
box -450 -340 350 260
use C7  C7_27
timestamp 1696364841
transform 1 0 8250 0 1 6536
box -450 -340 350 260
use C7  C7_28
timestamp 1696364841
transform 1 0 9550 0 1 4856
box -450 -340 350 260
use C7  C7_29
timestamp 1696364841
transform 1 0 8250 0 1 4856
box -450 -340 350 260
use C7  C7_30
timestamp 1696364841
transform 1 0 4350 0 1 4856
box -450 -340 350 260
use C7  C7_31
timestamp 1696364841
transform 1 0 1750 0 1 4856
box -450 -340 350 260
use C7  C7_32
timestamp 1696364841
transform 1 0 1750 0 1 5696
box -450 -340 350 260
use C7  C7_33
timestamp 1696364841
transform 1 0 4350 0 1 6536
box -450 -340 350 260
use C7  C7_34
timestamp 1696364841
transform 1 0 1750 0 1 6536
box -450 -340 350 260
use C7  C7_35
timestamp 1696364841
transform 1 0 4350 0 1 5696
box -450 -340 350 260
use C7  C7_36
timestamp 1696364841
transform 1 0 1750 0 1 8216
box -450 -340 350 260
use C7  C7_37
timestamp 1696364841
transform 1 0 4350 0 1 8216
box -450 -340 350 260
use C7  C7_38
timestamp 1696364841
transform 1 0 1750 0 1 7376
box -450 -340 350 260
use C7  C7_39
timestamp 1696364841
transform 1 0 4350 0 1 7376
box -450 -340 350 260
use C7  C7_40
timestamp 1696364841
transform 1 0 9550 0 1 8216
box -450 -340 350 260
use C7  C7_41
timestamp 1696364841
transform 1 0 8250 0 1 8216
box -450 -340 350 260
use C7  C7_42
timestamp 1696364841
transform 1 0 9550 0 1 7376
box -450 -340 350 260
use C7  C7_43
timestamp 1696364841
transform 1 0 8250 0 1 7376
box -450 -340 350 260
use C7  C7_44
timestamp 1696364841
transform 1 0 5650 0 1 4856
box -450 -340 350 260
use C7  C7_45
timestamp 1696364841
transform 1 0 5650 0 1 8216
box -450 -340 350 260
use C7  C7_46
timestamp 1696364841
transform 1 0 5650 0 1 7376
box -450 -340 350 260
use C7  C7_47
timestamp 1696364841
transform 1 0 5650 0 1 6536
box -450 -340 350 260
use C7  C7_48
timestamp 1696364841
transform 1 0 5650 0 1 5696
box -450 -340 350 260
use C7  C7_49
timestamp 1696364841
transform 1 0 18650 0 1 4856
box -450 -340 350 260
use C7  C7_50
timestamp 1696364841
transform 1 0 18650 0 1 6536
box -450 -340 350 260
use C7  C7_51
timestamp 1696364841
transform 1 0 18650 0 1 5696
box -450 -340 350 260
use C7  C7_52
timestamp 1696364841
transform 1 0 14750 0 1 4856
box -450 -340 350 260
use C7  C7_53
timestamp 1696364841
transform 1 0 13450 0 1 4856
box -450 -340 350 260
use C7  C7_54
timestamp 1696364841
transform 1 0 14750 0 1 5696
box -450 -340 350 260
use C7  C7_55
timestamp 1696364841
transform 1 0 13450 0 1 5696
box -450 -340 350 260
use C7  C7_56
timestamp 1696364841
transform 1 0 14750 0 1 6536
box -450 -340 350 260
use C7  C7_57
timestamp 1696364841
transform 1 0 13450 0 1 6536
box -450 -340 350 260
use C7  C7_58
timestamp 1696364841
transform 1 0 14750 0 1 7376
box -450 -340 350 260
use C7  C7_59
timestamp 1696364841
transform 1 0 13450 0 1 7376
box -450 -340 350 260
use C7  C7_60
timestamp 1696364841
transform 1 0 13450 0 1 8216
box -450 -340 350 260
use C7  C7_61
timestamp 1696364841
transform 1 0 14750 0 1 8216
box -450 -340 350 260
use C7  C7_62
timestamp 1696364841
transform 1 0 18650 0 1 8216
box -450 -340 350 260
use C7  C7_63
timestamp 1696364841
transform 1 0 18650 0 1 7376
box -450 -340 350 260
use C7  C7_64
timestamp 1696364841
transform 1 0 35550 0 1 3176
box -450 -340 350 260
use C7  C7_65
timestamp 1696364841
transform 1 0 34250 0 1 2336
box -450 -340 350 260
use C7  C7_66
timestamp 1696364841
transform 1 0 35550 0 1 2336
box -450 -340 350 260
use C7  C7_67
timestamp 1696364841
transform 1 0 35550 0 1 4016
box -450 -340 350 260
use C7  C7_68
timestamp 1696364841
transform 1 0 34250 0 1 4016
box -450 -340 350 260
use C7  C7_69
timestamp 1696364841
transform 1 0 34250 0 1 3176
box -450 -340 350 260
use C7  C7_70
timestamp 1696364841
transform 1 0 42050 0 1 4016
box -450 -340 350 260
use C7  C7_71
timestamp 1696364841
transform 1 0 39450 0 1 4016
box -450 -340 350 260
use C7  C7_72
timestamp 1696364841
transform 1 0 42050 0 1 3176
box -450 -340 350 260
use C7  C7_73
timestamp 1696364841
transform 1 0 39450 0 1 2336
box -450 -340 350 260
use C7  C7_74
timestamp 1696364841
transform 1 0 42050 0 1 2336
box -450 -340 350 260
use C7  C7_75
timestamp 1696364841
transform 1 0 39450 0 1 3176
box -450 -340 350 260
use C7  C7_76
timestamp 1696364841
transform 1 0 38150 0 1 4016
box -450 -340 350 260
use C7  C7_77
timestamp 1696364841
transform 1 0 38150 0 1 3176
box -450 -340 350 260
use C7  C7_78
timestamp 1696364841
transform 1 0 38150 0 1 2336
box -450 -340 350 260
use C7  C7_79
timestamp 1696364841
transform 1 0 25150 0 1 4016
box -450 -340 350 260
use C7  C7_80
timestamp 1696364841
transform 1 0 25150 0 1 2336
box -450 -340 350 260
use C7  C7_81
timestamp 1696364841
transform 1 0 25150 0 1 3176
box -450 -340 350 260
use C7  C7_82
timestamp 1696364841
transform 1 0 29050 0 1 3176
box -450 -340 350 260
use C7  C7_83
timestamp 1696364841
transform 1 0 30350 0 1 4016
box -450 -340 350 260
use C7  C7_84
timestamp 1696364841
transform 1 0 29050 0 1 4016
box -450 -340 350 260
use C7  C7_85
timestamp 1696364841
transform 1 0 30350 0 1 3176
box -450 -340 350 260
use C7  C7_86
timestamp 1696364841
transform 1 0 30350 0 1 2336
box -450 -340 350 260
use C7  C7_87
timestamp 1696364841
transform 1 0 29050 0 1 2336
box -450 -340 350 260
use C7  C7_88
timestamp 1696364841
transform 1 0 30350 0 1 5696
box -450 -340 350 260
use C7  C7_89
timestamp 1696364841
transform 1 0 29050 0 1 5696
box -450 -340 350 260
use C7  C7_90
timestamp 1696364841
transform 1 0 30350 0 1 6536
box -450 -340 350 260
use C7  C7_91
timestamp 1696364841
transform 1 0 29050 0 1 6536
box -450 -340 350 260
use C7  C7_92
timestamp 1696364841
transform 1 0 30350 0 1 4856
box -450 -340 350 260
use C7  C7_93
timestamp 1696364841
transform 1 0 29050 0 1 4856
box -450 -340 350 260
use C7  C7_94
timestamp 1696364841
transform 1 0 25150 0 1 6536
box -450 -340 350 260
use C7  C7_95
timestamp 1696364841
transform 1 0 25150 0 1 5696
box -450 -340 350 260
use C7  C7_96
timestamp 1696364841
transform 1 0 25150 0 1 4856
box -450 -340 350 260
use C7  C7_97
timestamp 1696364841
transform 1 0 25150 0 1 8216
box -450 -340 350 260
use C7  C7_98
timestamp 1696364841
transform 1 0 25150 0 1 7376
box -450 -340 350 260
use C7  C7_99
timestamp 1696364841
transform 1 0 30350 0 1 8216
box -450 -340 350 260
use C7  C7_100
timestamp 1696364841
transform 1 0 29050 0 1 8216
box -450 -340 350 260
use C7  C7_101
timestamp 1696364841
transform 1 0 30350 0 1 7376
box -450 -340 350 260
use C7  C7_102
timestamp 1696364841
transform 1 0 29050 0 1 7376
box -450 -340 350 260
use C7  C7_103
timestamp 1696364841
transform 1 0 39450 0 1 6536
box -450 -340 350 260
use C7  C7_104
timestamp 1696364841
transform 1 0 42050 0 1 6536
box -450 -340 350 260
use C7  C7_105
timestamp 1696364841
transform 1 0 42050 0 1 5696
box -450 -340 350 260
use C7  C7_106
timestamp 1696364841
transform 1 0 42050 0 1 4856
box -450 -340 350 260
use C7  C7_107
timestamp 1696364841
transform 1 0 39450 0 1 4856
box -450 -340 350 260
use C7  C7_108
timestamp 1696364841
transform 1 0 39450 0 1 5696
box -450 -340 350 260
use C7  C7_109
timestamp 1696364841
transform 1 0 35550 0 1 6536
box -450 -340 350 260
use C7  C7_110
timestamp 1696364841
transform 1 0 34250 0 1 6536
box -450 -340 350 260
use C7  C7_111
timestamp 1696364841
transform 1 0 35550 0 1 4856
box -450 -340 350 260
use C7  C7_112
timestamp 1696364841
transform 1 0 34250 0 1 4856
box -450 -340 350 260
use C7  C7_113
timestamp 1696364841
transform 1 0 35550 0 1 5696
box -450 -340 350 260
use C7  C7_114
timestamp 1696364841
transform 1 0 34250 0 1 5696
box -450 -340 350 260
use C7  C7_115
timestamp 1696364841
transform 1 0 34250 0 1 8216
box -450 -340 350 260
use C7  C7_116
timestamp 1696364841
transform 1 0 35550 0 1 7376
box -450 -340 350 260
use C7  C7_117
timestamp 1696364841
transform 1 0 34250 0 1 7376
box -450 -340 350 260
use C7  C7_118
timestamp 1696364841
transform 1 0 35550 0 1 8216
box -450 -340 350 260
use C7  C7_119
timestamp 1696364841
transform 1 0 42050 0 1 7376
box -450 -340 350 260
use C7  C7_120
timestamp 1696364841
transform 1 0 39450 0 1 7376
box -450 -340 350 260
use C7  C7_121
timestamp 1696364841
transform 1 0 42050 0 1 8216
box -450 -340 350 260
use C7  C7_122
timestamp 1696364841
transform 1 0 39450 0 1 8216
box -450 -340 350 260
use C7  C7_123
timestamp 1696364841
transform 1 0 38150 0 1 8216
box -450 -340 350 260
use C7  C7_124
timestamp 1696364841
transform 1 0 38150 0 1 7376
box -450 -340 350 260
use C7  C7_125
timestamp 1696364841
transform 1 0 38150 0 1 5696
box -450 -340 350 260
use C7  C7_126
timestamp 1696364841
transform 1 0 38150 0 1 6536
box -450 -340 350 260
use C7  C7_127
timestamp 1696364841
transform 1 0 38150 0 1 4856
box -450 -340 350 260
use CDUM  CDUM_0
timestamp 1696364841
transform 1 0 22550 0 1 4856
box -450 -340 350 260
use DUMMY  DUMMY_0
timestamp 1696364841
transform 1 0 17350 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_1
timestamp 1696364841
transform 1 0 18650 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_2
timestamp 1696364841
transform 1 0 19950 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_3
timestamp 1696364841
transform 1 0 21250 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_4
timestamp 1696364841
transform 1 0 12150 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_5
timestamp 1696364841
transform 1 0 13450 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_6
timestamp 1696364841
transform 1 0 14750 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_7
timestamp 1696364841
transform 1 0 16050 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_8
timestamp 1696364841
transform 1 0 6950 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_9
timestamp 1696364841
transform 1 0 8250 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_10
timestamp 1696364841
transform 1 0 9550 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_11
timestamp 1696364841
transform 1 0 450 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_12
timestamp 1696364841
transform 1 0 1750 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_13
timestamp 1696364841
transform 1 0 3050 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_14
timestamp 1696364841
transform 1 0 4350 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_15
timestamp 1696364841
transform 1 0 450 0 1 3176
box -450 -340 350 260
use DUMMY  DUMMY_16
timestamp 1696364841
transform 1 0 450 0 1 4016
box -450 -340 350 260
use DUMMY  DUMMY_17
timestamp 1696364841
transform 1 0 450 0 1 2336
box -450 -340 350 260
use DUMMY  DUMMY_18
timestamp 1696364841
transform 1 0 5650 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_19
timestamp 1696364841
transform 1 0 450 0 1 5696
box -450 -340 350 260
use DUMMY  DUMMY_20
timestamp 1696364841
transform 1 0 450 0 1 4856
box -450 -340 350 260
use DUMMY  DUMMY_21
timestamp 1696364841
transform 1 0 450 0 1 6536
box -450 -340 350 260
use DUMMY  DUMMY_22
timestamp 1696364841
transform 1 0 450 0 1 8216
box -450 -340 350 260
use DUMMY  DUMMY_23
timestamp 1696364841
transform 1 0 450 0 1 7376
box -450 -340 350 260
use DUMMY  DUMMY_24
timestamp 1696364841
transform 1 0 1750 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_25
timestamp 1696364841
transform 1 0 450 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_26
timestamp 1696364841
transform 1 0 3050 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_27
timestamp 1696364841
transform 1 0 4350 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_28
timestamp 1696364841
transform 1 0 6950 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_29
timestamp 1696364841
transform 1 0 8250 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_30
timestamp 1696364841
transform 1 0 9550 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_31
timestamp 1696364841
transform 1 0 5650 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_32
timestamp 1696364841
transform 1 0 12150 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_33
timestamp 1696364841
transform 1 0 13450 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_34
timestamp 1696364841
transform 1 0 14750 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_35
timestamp 1696364841
transform 1 0 19950 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_36
timestamp 1696364841
transform 1 0 21250 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_37
timestamp 1696364841
transform 1 0 17350 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_38
timestamp 1696364841
transform 1 0 18650 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_39
timestamp 1696364841
transform 1 0 16050 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_40
timestamp 1696364841
transform 1 0 10850 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_41
timestamp 1696364841
transform 1 0 10850 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_42
timestamp 1696364841
transform 1 0 42050 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_43
timestamp 1696364841
transform 1 0 43350 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_44
timestamp 1696364841
transform 1 0 39450 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_45
timestamp 1696364841
transform 1 0 40750 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_46
timestamp 1696364841
transform 1 0 34250 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_47
timestamp 1696364841
transform 1 0 35550 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_48
timestamp 1696364841
transform 1 0 36850 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_49
timestamp 1696364841
transform 1 0 43350 0 1 4016
box -450 -340 350 260
use DUMMY  DUMMY_50
timestamp 1696364841
transform 1 0 43350 0 1 2336
box -450 -340 350 260
use DUMMY  DUMMY_51
timestamp 1696364841
transform 1 0 43350 0 1 3176
box -450 -340 350 260
use DUMMY  DUMMY_52
timestamp 1696364841
transform 1 0 38150 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_53
timestamp 1696364841
transform 1 0 29050 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_54
timestamp 1696364841
transform 1 0 31650 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_55
timestamp 1696364841
transform 1 0 30350 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_56
timestamp 1696364841
transform 1 0 26450 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_57
timestamp 1696364841
transform 1 0 22550 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_58
timestamp 1696364841
transform 1 0 23850 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_59
timestamp 1696364841
transform 1 0 25150 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_60
timestamp 1696364841
transform 1 0 27750 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_61
timestamp 1696364841
transform 1 0 23850 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_62
timestamp 1696364841
transform 1 0 25150 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_63
timestamp 1696364841
transform 1 0 26450 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_64
timestamp 1696364841
transform 1 0 22550 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_65
timestamp 1696364841
transform 1 0 30350 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_66
timestamp 1696364841
transform 1 0 31650 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_67
timestamp 1696364841
transform 1 0 29050 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_68
timestamp 1696364841
transform 1 0 27750 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_69
timestamp 1696364841
transform 1 0 43350 0 1 6536
box -450 -340 350 260
use DUMMY  DUMMY_70
timestamp 1696364841
transform 1 0 43350 0 1 5696
box -450 -340 350 260
use DUMMY  DUMMY_71
timestamp 1696364841
transform 1 0 43350 0 1 4856
box -450 -340 350 260
use DUMMY  DUMMY_72
timestamp 1696364841
transform 1 0 34250 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_73
timestamp 1696364841
transform 1 0 35550 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_74
timestamp 1696364841
transform 1 0 36850 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_75
timestamp 1696364841
transform 1 0 43350 0 1 8216
box -450 -340 350 260
use DUMMY  DUMMY_76
timestamp 1696364841
transform 1 0 43350 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_77
timestamp 1696364841
transform 1 0 43350 0 1 7376
box -450 -340 350 260
use DUMMY  DUMMY_78
timestamp 1696364841
transform 1 0 39450 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_79
timestamp 1696364841
transform 1 0 40750 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_80
timestamp 1696364841
transform 1 0 42050 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_81
timestamp 1696364841
transform 1 0 38150 0 1 9056
box -450 -340 350 260
use DUMMY  DUMMY_82
timestamp 1696364841
transform 1 0 32950 0 1 1496
box -450 -340 350 260
use DUMMY  DUMMY_83
timestamp 1696364841
transform 1 0 32950 0 1 9056
box -450 -340 350 260
use via23_4  via23_4_0
timestamp 1696364841
transform -1 0 21401 0 -1 -196
box 1 40 161 120
use via23_4  via23_4_1
timestamp 1696364841
transform 0 -1 20244 1 0 1375
box 1 40 161 120
use via23_4  via23_4_2
timestamp 1696364841
transform 0 -1 21544 1 0 1375
box 1 40 161 120
use via23_4  via23_4_3
timestamp 1696364841
transform 0 -1 17116 1 0 1375
box 1 40 161 120
use via23_4  via23_4_4
timestamp 1696364841
transform -1 0 16961 0 -1 284
box 1 40 161 120
use via23_4  via23_4_5
timestamp 1696364841
transform -1 0 18261 0 -1 124
box 1 40 161 120
use via23_4  via23_4_6
timestamp 1696364841
transform -1 0 19561 0 -1 604
box 1 40 161 120
use via23_4  via23_4_7
timestamp 1696364841
transform -1 0 20861 0 -1 764
box 1 40 161 120
use via23_4  via23_4_8
timestamp 1696364841
transform 1 0 21299 0 -1 1084
box 1 40 161 120
use via23_4  via23_4_9
timestamp 1696364841
transform 0 -1 18416 1 0 1375
box 1 40 161 120
use via23_4  via23_4_10
timestamp 1696364841
transform 0 -1 21016 1 0 1375
box 1 40 161 120
use via23_4  via23_4_11
timestamp 1696364841
transform 0 -1 18944 1 0 1375
box 1 40 161 120
use via23_4  via23_4_12
timestamp 1696364841
transform 0 -1 17644 1 0 1375
box 1 40 161 120
use via23_4  via23_4_13
timestamp 1696364841
transform 0 -1 19716 1 0 1375
box 1 40 161 120
use via23_4  via23_4_14
timestamp 1696364841
transform -1 0 11761 0 -1 284
box 1 40 161 120
use via23_4  via23_4_15
timestamp 1696364841
transform 0 -1 11144 1 0 1375
box 1 40 161 120
use via23_4  via23_4_16
timestamp 1696364841
transform 0 -1 11916 1 0 1375
box 1 40 161 120
use via23_4  via23_4_17
timestamp 1696364841
transform 0 -1 13216 1 0 1375
box 1 40 161 120
use via23_4  via23_4_18
timestamp 1696364841
transform 0 -1 15044 1 0 1375
box 1 40 161 120
use via23_4  via23_4_19
timestamp 1696364841
transform 0 -1 16344 1 0 1375
box 1 40 161 120
use via23_4  via23_4_20
timestamp 1696364841
transform 0 -1 12444 1 0 1375
box 1 40 161 120
use via23_4  via23_4_21
timestamp 1696364841
transform 0 -1 13744 1 0 1375
box 1 40 161 120
use via23_4  via23_4_22
timestamp 1696364841
transform 0 -1 14516 1 0 1375
box 1 40 161 120
use via23_4  via23_4_23
timestamp 1696364841
transform 0 -1 15816 1 0 1375
box 1 40 161 120
use via23_4  via23_4_24
timestamp 1696364841
transform -1 0 13061 0 -1 124
box 1 40 161 120
use via23_4  via23_4_25
timestamp 1696364841
transform -1 0 14361 0 -1 124
box 1 40 161 120
use via23_4  via23_4_26
timestamp 1696364841
transform -1 0 15661 0 -1 444
box 1 40 161 120
use via23_4  via23_4_27
timestamp 1696364841
transform 0 -1 11916 1 0 2215
box 1 40 161 120
use via23_4  via23_4_28
timestamp 1696364841
transform 0 -1 11144 1 0 3895
box 1 40 161 120
use via23_4  via23_4_29
timestamp 1696364841
transform 0 -1 15044 1 0 3055
box 1 40 161 120
use via23_4  via23_4_30
timestamp 1696364841
transform 0 -1 13744 1 0 3055
box 1 40 161 120
use via23_4  via23_4_31
timestamp 1696364841
transform 0 -1 15044 1 0 3895
box 1 40 161 120
use via23_4  via23_4_32
timestamp 1696364841
transform 0 -1 13744 1 0 3895
box 1 40 161 120
use via23_4  via23_4_33
timestamp 1696364841
transform 0 -1 12444 1 0 3895
box 1 40 161 120
use via23_4  via23_4_34
timestamp 1696364841
transform 0 -1 12444 1 0 3055
box 1 40 161 120
use via23_4  via23_4_35
timestamp 1696364841
transform 0 -1 16344 1 0 3895
box 1 40 161 120
use via23_4  via23_4_36
timestamp 1696364841
transform 0 -1 15816 1 0 3895
box 1 40 161 120
use via23_4  via23_4_37
timestamp 1696364841
transform 0 -1 14516 1 0 3895
box 1 40 161 120
use via23_4  via23_4_38
timestamp 1696364841
transform 0 -1 13216 1 0 3895
box 1 40 161 120
use via23_4  via23_4_39
timestamp 1696364841
transform 0 -1 11916 1 0 3895
box 1 40 161 120
use via23_4  via23_4_40
timestamp 1696364841
transform 0 -1 16344 1 0 3055
box 1 40 161 120
use via23_4  via23_4_41
timestamp 1696364841
transform 0 -1 15816 1 0 3055
box 1 40 161 120
use via23_4  via23_4_42
timestamp 1696364841
transform 0 -1 14516 1 0 3055
box 1 40 161 120
use via23_4  via23_4_43
timestamp 1696364841
transform 0 -1 13216 1 0 3055
box 1 40 161 120
use via23_4  via23_4_44
timestamp 1696364841
transform 0 -1 11916 1 0 3055
box 1 40 161 120
use via23_4  via23_4_45
timestamp 1696364841
transform 0 -1 11144 1 0 3055
box 1 40 161 120
use via23_4  via23_4_46
timestamp 1696364841
transform 0 -1 14516 1 0 2215
box 1 40 161 120
use via23_4  via23_4_47
timestamp 1696364841
transform 0 -1 13216 1 0 2215
box 1 40 161 120
use via23_4  via23_4_48
timestamp 1696364841
transform 0 -1 16344 1 0 2215
box 1 40 161 120
use via23_4  via23_4_49
timestamp 1696364841
transform 0 -1 15044 1 0 2215
box 1 40 161 120
use via23_4  via23_4_50
timestamp 1696364841
transform 0 -1 13744 1 0 2215
box 1 40 161 120
use via23_4  via23_4_51
timestamp 1696364841
transform 0 -1 15816 1 0 2215
box 1 40 161 120
use via23_4  via23_4_52
timestamp 1696364841
transform 0 -1 12444 1 0 2215
box 1 40 161 120
use via23_4  via23_4_53
timestamp 1696364841
transform 0 -1 11144 1 0 2215
box 1 40 161 120
use via23_4  via23_4_54
timestamp 1696364841
transform 0 -1 21016 1 0 2215
box 1 40 161 120
use via23_4  via23_4_55
timestamp 1696364841
transform 0 -1 21544 1 0 2215
box 1 40 161 120
use via23_4  via23_4_56
timestamp 1696364841
transform 0 -1 20244 1 0 3055
box 1 40 161 120
use via23_4  via23_4_57
timestamp 1696364841
transform 0 -1 21016 1 0 3055
box 1 40 161 120
use via23_4  via23_4_58
timestamp 1696364841
transform 0 -1 18944 1 0 3895
box 1 40 161 120
use via23_4  via23_4_59
timestamp 1696364841
transform 0 -1 17644 1 0 3895
box 1 40 161 120
use via23_4  via23_4_60
timestamp 1696364841
transform 0 -1 19716 1 0 3055
box 1 40 161 120
use via23_4  via23_4_61
timestamp 1696364841
transform 0 -1 20690 1 0 3895
box 1 40 161 120
use via23_4  via23_4_62
timestamp 1696364841
transform 0 -1 18416 1 0 3055
box 1 40 161 120
use via23_4  via23_4_63
timestamp 1696364841
transform 0 -1 17116 1 0 3055
box 1 40 161 120
use via23_4  via23_4_64
timestamp 1696364841
transform 0 -1 21016 1 0 3895
box 1 40 161 120
use via23_4  via23_4_65
timestamp 1696364841
transform 0 -1 18944 1 0 2215
box 1 40 161 120
use via23_4  via23_4_66
timestamp 1696364841
transform 0 -1 17644 1 0 2215
box 1 40 161 120
use via23_4  via23_4_67
timestamp 1696364841
transform 0 -1 18944 1 0 3055
box 1 40 161 120
use via23_4  via23_4_68
timestamp 1696364841
transform 0 -1 17644 1 0 3055
box 1 40 161 120
use via23_4  via23_4_69
timestamp 1696364841
transform 0 -1 21544 1 0 3895
box 1 40 161 120
use via23_4  via23_4_70
timestamp 1696364841
transform 0 -1 20244 1 0 3895
box 1 40 161 120
use via23_4  via23_4_71
timestamp 1696364841
transform 0 -1 21544 1 0 3055
box 1 40 161 120
use via23_4  via23_4_72
timestamp 1696364841
transform 0 -1 18416 1 0 2215
box 1 40 161 120
use via23_4  via23_4_73
timestamp 1696364841
transform 0 -1 19716 1 0 3895
box 1 40 161 120
use via23_4  via23_4_74
timestamp 1696364841
transform 0 -1 18416 1 0 3895
box 1 40 161 120
use via23_4  via23_4_75
timestamp 1696364841
transform 0 -1 17116 1 0 3895
box 1 40 161 120
use via23_4  via23_4_76
timestamp 1696364841
transform 0 -1 19716 1 0 2215
box 1 40 161 120
use via23_4  via23_4_77
timestamp 1696364841
transform 0 -1 17116 1 0 2215
box 1 40 161 120
use via23_4  via23_4_78
timestamp 1696364841
transform 0 -1 20244 1 0 2215
box 1 40 161 120
use via23_4  via23_4_79
timestamp 1696364841
transform 0 -1 5944 1 0 1375
box 1 40 161 120
use via23_4  via23_4_80
timestamp 1696364841
transform -1 0 9161 0 -1 124
box 1 40 161 120
use via23_4  via23_4_81
timestamp 1696364841
transform -1 0 7861 0 -1 124
box 1 40 161 120
use via23_4  via23_4_82
timestamp 1696364841
transform -1 0 10461 0 -1 444
box 1 40 161 120
use via23_4  via23_4_83
timestamp 1696364841
transform -1 0 6561 0 -1 284
box 1 40 161 120
use via23_4  via23_4_84
timestamp 1696364841
transform 0 -1 9844 1 0 1375
box 1 40 161 120
use via23_4  via23_4_85
timestamp 1696364841
transform 0 -1 6716 1 0 1375
box 1 40 161 120
use via23_4  via23_4_86
timestamp 1696364841
transform 0 -1 8016 1 0 1375
box 1 40 161 120
use via23_4  via23_4_87
timestamp 1696364841
transform 0 -1 7244 1 0 1375
box 1 40 161 120
use via23_4  via23_4_88
timestamp 1696364841
transform 0 -1 8544 1 0 1375
box 1 40 161 120
use via23_4  via23_4_89
timestamp 1696364841
transform 0 -1 10616 1 0 1375
box 1 40 161 120
use via23_4  via23_4_90
timestamp 1696364841
transform 0 -1 9316 1 0 1375
box 1 40 161 120
use via23_4  via23_4_91
timestamp 1696364841
transform 0 -1 3344 1 0 1375
box 1 40 161 120
use via23_4  via23_4_92
timestamp 1696364841
transform 0 -1 4644 1 0 1375
box 1 40 161 120
use via23_4  via23_4_93
timestamp 1696364841
transform 0 -1 744 1 0 1375
box 1 40 161 120
use via23_4  via23_4_94
timestamp 1696364841
transform 0 -1 4116 1 0 1375
box 1 40 161 120
use via23_4  via23_4_95
timestamp 1696364841
transform 0 -1 5416 1 0 1375
box 1 40 161 120
use via23_4  via23_4_96
timestamp 1696364841
transform 0 -1 216 1 0 1375
box 1 40 161 120
use via23_4  via23_4_97
timestamp 1696364841
transform -1 0 2661 0 -1 284
box 1 40 161 120
use via23_4  via23_4_98
timestamp 1696364841
transform -1 0 3961 0 -1 124
box 1 40 161 120
use via23_4  via23_4_99
timestamp 1696364841
transform -1 0 1361 0 -1 124
box 1 40 161 120
use via23_4  via23_4_100
timestamp 1696364841
transform -1 0 5261 0 -1 124
box 1 40 161 120
use via23_4  via23_4_101
timestamp 1696364841
transform 0 -1 2816 1 0 1375
box 1 40 161 120
use via23_4  via23_4_102
timestamp 1696364841
transform 0 -1 1516 1 0 1375
box 1 40 161 120
use via23_4  via23_4_103
timestamp 1696364841
transform 0 -1 2044 1 0 1375
box 1 40 161 120
use via23_4  via23_4_104
timestamp 1696364841
transform 0 -1 3344 1 0 3055
box 1 40 161 120
use via23_4  via23_4_105
timestamp 1696364841
transform 0 -1 216 1 0 3895
box 1 40 161 120
use via23_4  via23_4_106
timestamp 1696364841
transform 0 -1 216 1 0 3055
box 1 40 161 120
use via23_4  via23_4_107
timestamp 1696364841
transform 0 -1 2044 1 0 3055
box 1 40 161 120
use via23_4  via23_4_108
timestamp 1696364841
transform 0 -1 5416 1 0 3055
box 1 40 161 120
use via23_4  via23_4_109
timestamp 1696364841
transform 0 -1 4116 1 0 2215
box 1 40 161 120
use via23_4  via23_4_110
timestamp 1696364841
transform 0 -1 2816 1 0 2215
box 1 40 161 120
use via23_4  via23_4_111
timestamp 1696364841
transform 0 -1 744 1 0 3895
box 1 40 161 120
use via23_4  via23_4_112
timestamp 1696364841
transform 0 -1 4644 1 0 2215
box 1 40 161 120
use via23_4  via23_4_113
timestamp 1696364841
transform 0 -1 3344 1 0 2215
box 1 40 161 120
use via23_4  via23_4_114
timestamp 1696364841
transform 0 -1 5416 1 0 2215
box 1 40 161 120
use via23_4  via23_4_115
timestamp 1696364841
transform 0 -1 744 1 0 2215
box 1 40 161 120
use via23_4  via23_4_116
timestamp 1696364841
transform 0 -1 1516 1 0 2215
box 1 40 161 120
use via23_4  via23_4_117
timestamp 1696364841
transform 0 -1 744 1 0 3055
box 1 40 161 120
use via23_4  via23_4_118
timestamp 1696364841
transform 0 -1 4116 1 0 3055
box 1 40 161 120
use via23_4  via23_4_119
timestamp 1696364841
transform 0 -1 2816 1 0 3055
box 1 40 161 120
use via23_4  via23_4_120
timestamp 1696364841
transform 0 -1 1516 1 0 3055
box 1 40 161 120
use via23_4  via23_4_121
timestamp 1696364841
transform 0 -1 4644 1 0 3055
box 1 40 161 120
use via23_4  via23_4_122
timestamp 1696364841
transform 0 -1 4644 1 0 3895
box 1 40 161 120
use via23_4  via23_4_123
timestamp 1696364841
transform 0 -1 5416 1 0 3895
box 1 40 161 120
use via23_4  via23_4_124
timestamp 1696364841
transform 0 -1 4116 1 0 3895
box 1 40 161 120
use via23_4  via23_4_125
timestamp 1696364841
transform 0 -1 2816 1 0 3895
box 1 40 161 120
use via23_4  via23_4_126
timestamp 1696364841
transform 0 -1 3344 1 0 3895
box 1 40 161 120
use via23_4  via23_4_127
timestamp 1696364841
transform 0 -1 2044 1 0 3895
box 1 40 161 120
use via23_4  via23_4_128
timestamp 1696364841
transform 0 -1 216 1 0 2215
box 1 40 161 120
use via23_4  via23_4_129
timestamp 1696364841
transform 0 -1 2044 1 0 2215
box 1 40 161 120
use via23_4  via23_4_130
timestamp 1696364841
transform 0 -1 1516 1 0 3895
box 1 40 161 120
use via23_4  via23_4_131
timestamp 1696364841
transform 0 -1 6716 1 0 3055
box 1 40 161 120
use via23_4  via23_4_132
timestamp 1696364841
transform 0 -1 5944 1 0 2215
box 1 40 161 120
use via23_4  via23_4_133
timestamp 1696364841
transform 0 -1 10616 1 0 3895
box 1 40 161 120
use via23_4  via23_4_134
timestamp 1696364841
transform 0 -1 9316 1 0 3895
box 1 40 161 120
use via23_4  via23_4_135
timestamp 1696364841
transform 0 -1 6716 1 0 3895
box 1 40 161 120
use via23_4  via23_4_136
timestamp 1696364841
transform 0 -1 8016 1 0 3895
box 1 40 161 120
use via23_4  via23_4_137
timestamp 1696364841
transform 0 -1 7244 1 0 3895
box 1 40 161 120
use via23_4  via23_4_138
timestamp 1696364841
transform 0 -1 5944 1 0 3895
box 1 40 161 120
use via23_4  via23_4_139
timestamp 1696364841
transform 0 -1 9316 1 0 2215
box 1 40 161 120
use via23_4  via23_4_140
timestamp 1696364841
transform 0 -1 9844 1 0 3895
box 1 40 161 120
use via23_4  via23_4_141
timestamp 1696364841
transform 0 -1 9844 1 0 3055
box 1 40 161 120
use via23_4  via23_4_142
timestamp 1696364841
transform 0 -1 10616 1 0 2215
box 1 40 161 120
use via23_4  via23_4_143
timestamp 1696364841
transform 0 -1 9844 1 0 2215
box 1 40 161 120
use via23_4  via23_4_144
timestamp 1696364841
transform 0 -1 8544 1 0 2215
box 1 40 161 120
use via23_4  via23_4_145
timestamp 1696364841
transform 0 -1 10616 1 0 3055
box 1 40 161 120
use via23_4  via23_4_146
timestamp 1696364841
transform 0 -1 9316 1 0 3055
box 1 40 161 120
use via23_4  via23_4_147
timestamp 1696364841
transform 0 -1 8544 1 0 3895
box 1 40 161 120
use via23_4  via23_4_148
timestamp 1696364841
transform 0 -1 8016 1 0 3055
box 1 40 161 120
use via23_4  via23_4_149
timestamp 1696364841
transform 0 -1 7244 1 0 2215
box 1 40 161 120
use via23_4  via23_4_150
timestamp 1696364841
transform 0 -1 8016 1 0 2215
box 1 40 161 120
use via23_4  via23_4_151
timestamp 1696364841
transform 0 -1 6716 1 0 2215
box 1 40 161 120
use via23_4  via23_4_152
timestamp 1696364841
transform 0 -1 7244 1 0 3055
box 1 40 161 120
use via23_4  via23_4_153
timestamp 1696364841
transform 0 -1 5944 1 0 3055
box 1 40 161 120
use via23_4  via23_4_154
timestamp 1696364841
transform 0 -1 8544 1 0 3055
box 1 40 161 120
use via23_4  via23_4_155
timestamp 1696364841
transform 0 -1 6716 1 0 5575
box 1 40 161 120
use via23_4  via23_4_156
timestamp 1696364841
transform 0 -1 10616 1 0 6415
box 1 40 161 120
use via23_4  via23_4_157
timestamp 1696364841
transform 0 -1 6716 1 0 6415
box 1 40 161 120
use via23_4  via23_4_158
timestamp 1696364841
transform 0 -1 9844 1 0 5575
box 1 40 161 120
use via23_4  via23_4_159
timestamp 1696364841
transform 0 -1 8016 1 0 4735
box 1 40 161 120
use via23_4  via23_4_160
timestamp 1696364841
transform 0 -1 6716 1 0 4735
box 1 40 161 120
use via23_4  via23_4_161
timestamp 1696364841
transform 0 -1 9844 1 0 4735
box 1 40 161 120
use via23_4  via23_4_162
timestamp 1696364841
transform 0 -1 8544 1 0 4735
box 1 40 161 120
use via23_4  via23_4_163
timestamp 1696364841
transform 0 -1 7244 1 0 4735
box 1 40 161 120
use via23_4  via23_4_164
timestamp 1696364841
transform 0 -1 5944 1 0 4735
box 1 40 161 120
use via23_4  via23_4_165
timestamp 1696364841
transform 0 -1 7244 1 0 6415
box 1 40 161 120
use via23_4  via23_4_166
timestamp 1696364841
transform 0 -1 9316 1 0 5575
box 1 40 161 120
use via23_4  via23_4_167
timestamp 1696364841
transform 0 -1 8544 1 0 6415
box 1 40 161 120
use via23_4  via23_4_168
timestamp 1696364841
transform 0 -1 10616 1 0 4735
box 1 40 161 120
use via23_4  via23_4_169
timestamp 1696364841
transform 0 -1 9316 1 0 4735
box 1 40 161 120
use via23_4  via23_4_170
timestamp 1696364841
transform 0 -1 5944 1 0 6415
box 1 40 161 120
use via23_4  via23_4_171
timestamp 1696364841
transform 0 -1 8544 1 0 5575
box 1 40 161 120
use via23_4  via23_4_172
timestamp 1696364841
transform 0 -1 7244 1 0 5575
box 1 40 161 120
use via23_4  via23_4_173
timestamp 1696364841
transform 0 -1 10616 1 0 5575
box 1 40 161 120
use via23_4  via23_4_174
timestamp 1696364841
transform 0 -1 5944 1 0 5575
box 1 40 161 120
use via23_4  via23_4_175
timestamp 1696364841
transform 0 -1 9844 1 0 6415
box 1 40 161 120
use via23_4  via23_4_176
timestamp 1696364841
transform 0 -1 9316 1 0 6415
box 1 40 161 120
use via23_4  via23_4_177
timestamp 1696364841
transform 0 -1 8016 1 0 6415
box 1 40 161 120
use via23_4  via23_4_178
timestamp 1696364841
transform 0 -1 8016 1 0 5575
box 1 40 161 120
use via23_4  via23_4_179
timestamp 1696364841
transform 0 -1 216 1 0 6415
box 1 40 161 120
use via23_4  via23_4_180
timestamp 1696364841
transform 0 -1 216 1 0 5575
box 1 40 161 120
use via23_4  via23_4_181
timestamp 1696364841
transform 0 -1 3344 1 0 6415
box 1 40 161 120
use via23_4  via23_4_182
timestamp 1696364841
transform 0 -1 5416 1 0 5575
box 1 40 161 120
use via23_4  via23_4_183
timestamp 1696364841
transform 0 -1 4644 1 0 5575
box 1 40 161 120
use via23_4  via23_4_184
timestamp 1696364841
transform 0 -1 3344 1 0 5575
box 1 40 161 120
use via23_4  via23_4_185
timestamp 1696364841
transform 0 -1 2044 1 0 5575
box 1 40 161 120
use via23_4  via23_4_186
timestamp 1696364841
transform 0 -1 4116 1 0 5575
box 1 40 161 120
use via23_4  via23_4_187
timestamp 1696364841
transform 0 -1 2044 1 0 6415
box 1 40 161 120
use via23_4  via23_4_188
timestamp 1696364841
transform 0 -1 2816 1 0 5575
box 1 40 161 120
use via23_4  via23_4_189
timestamp 1696364841
transform 0 -1 5416 1 0 4735
box 1 40 161 120
use via23_4  via23_4_190
timestamp 1696364841
transform 0 -1 4116 1 0 4735
box 1 40 161 120
use via23_4  via23_4_191
timestamp 1696364841
transform 0 -1 3344 1 0 4735
box 1 40 161 120
use via23_4  via23_4_192
timestamp 1696364841
transform 0 -1 2044 1 0 4735
box 1 40 161 120
use via23_4  via23_4_193
timestamp 1696364841
transform 0 -1 2816 1 0 4735
box 1 40 161 120
use via23_4  via23_4_194
timestamp 1696364841
transform 0 -1 1516 1 0 5575
box 1 40 161 120
use via23_4  via23_4_195
timestamp 1696364841
transform 0 -1 4644 1 0 4735
box 1 40 161 120
use via23_4  via23_4_196
timestamp 1696364841
transform 0 -1 1516 1 0 4735
box 1 40 161 120
use via23_4  via23_4_197
timestamp 1696364841
transform 0 -1 744 1 0 4735
box 1 40 161 120
use via23_4  via23_4_198
timestamp 1696364841
transform 0 -1 744 1 0 6415
box 1 40 161 120
use via23_4  via23_4_199
timestamp 1696364841
transform 0 -1 216 1 0 4735
box 1 40 161 120
use via23_4  via23_4_200
timestamp 1696364841
transform 0 -1 744 1 0 5575
box 1 40 161 120
use via23_4  via23_4_201
timestamp 1696364841
transform 0 -1 4644 1 0 6415
box 1 40 161 120
use via23_4  via23_4_202
timestamp 1696364841
transform 0 -1 5416 1 0 6415
box 1 40 161 120
use via23_4  via23_4_203
timestamp 1696364841
transform 0 -1 4116 1 0 6415
box 1 40 161 120
use via23_4  via23_4_204
timestamp 1696364841
transform 0 -1 2816 1 0 6415
box 1 40 161 120
use via23_4  via23_4_205
timestamp 1696364841
transform 0 -1 1516 1 0 6415
box 1 40 161 120
use via23_4  via23_4_206
timestamp 1696364841
transform 0 -1 5416 1 0 7255
box 1 40 161 120
use via23_4  via23_4_207
timestamp 1696364841
transform 0 -1 4116 1 0 7255
box 1 40 161 120
use via23_4  via23_4_208
timestamp 1696364841
transform 0 -1 2816 1 0 7255
box 1 40 161 120
use via23_4  via23_4_209
timestamp 1696364841
transform 0 -1 2816 1 0 8095
box 1 40 161 120
use via23_4  via23_4_210
timestamp 1696364841
transform 0 -1 1516 1 0 8095
box 1 40 161 120
use via23_4  via23_4_211
timestamp 1696364841
transform 0 -1 4644 1 0 7255
box 1 40 161 120
use via23_4  via23_4_212
timestamp 1696364841
transform 0 -1 744 1 0 7255
box 1 40 161 120
use via23_4  via23_4_213
timestamp 1696364841
transform 0 -1 216 1 0 7255
box 1 40 161 120
use via23_4  via23_4_214
timestamp 1696364841
transform 0 -1 744 1 0 8095
box 1 40 161 120
use via23_4  via23_4_215
timestamp 1696364841
transform 0 -1 4644 1 0 8935
box 1 40 161 120
use via23_4  via23_4_216
timestamp 1696364841
transform 0 -1 1516 1 0 8935
box 1 40 161 120
use via23_4  via23_4_217
timestamp 1696364841
transform 0 -1 2816 1 0 8935
box 1 40 161 120
use via23_4  via23_4_218
timestamp 1696364841
transform 0 -1 4116 1 0 8935
box 1 40 161 120
use via23_4  via23_4_219
timestamp 1696364841
transform 0 -1 5416 1 0 8935
box 1 40 161 120
use via23_4  via23_4_220
timestamp 1696364841
transform 0 -1 216 1 0 8095
box 1 40 161 120
use via23_4  via23_4_221
timestamp 1696364841
transform 0 -1 1516 1 0 7255
box 1 40 161 120
use via23_4  via23_4_222
timestamp 1696364841
transform 0 -1 3344 1 0 7255
box 1 40 161 120
use via23_4  via23_4_223
timestamp 1696364841
transform 0 -1 2044 1 0 7255
box 1 40 161 120
use via23_4  via23_4_224
timestamp 1696364841
transform 0 -1 4644 1 0 8095
box 1 40 161 120
use via23_4  via23_4_225
timestamp 1696364841
transform 0 -1 3344 1 0 8095
box 1 40 161 120
use via23_4  via23_4_226
timestamp 1696364841
transform 0 -1 2044 1 0 8095
box 1 40 161 120
use via23_4  via23_4_227
timestamp 1696364841
transform 0 -1 744 1 0 8935
box 1 40 161 120
use via23_4  via23_4_228
timestamp 1696364841
transform 0 -1 216 1 0 8935
box 1 40 161 120
use via23_4  via23_4_229
timestamp 1696364841
transform 0 -1 2044 1 0 8935
box 1 40 161 120
use via23_4  via23_4_230
timestamp 1696364841
transform 0 -1 3344 1 0 8935
box 1 40 161 120
use via23_4  via23_4_231
timestamp 1696364841
transform 0 -1 5416 1 0 8095
box 1 40 161 120
use via23_4  via23_4_232
timestamp 1696364841
transform 0 -1 4116 1 0 8095
box 1 40 161 120
use via23_4  via23_4_233
timestamp 1696364841
transform 0 -1 9844 1 0 8935
box 1 40 161 120
use via23_4  via23_4_234
timestamp 1696364841
transform 0 -1 7244 1 0 8095
box 1 40 161 120
use via23_4  via23_4_235
timestamp 1696364841
transform 0 -1 10616 1 0 8095
box 1 40 161 120
use via23_4  via23_4_236
timestamp 1696364841
transform 0 -1 9316 1 0 8095
box 1 40 161 120
use via23_4  via23_4_237
timestamp 1696364841
transform 0 -1 8016 1 0 8095
box 1 40 161 120
use via23_4  via23_4_238
timestamp 1696364841
transform 0 -1 6716 1 0 8095
box 1 40 161 120
use via23_4  via23_4_239
timestamp 1696364841
transform 0 -1 5944 1 0 8095
box 1 40 161 120
use via23_4  via23_4_240
timestamp 1696364841
transform 0 -1 9844 1 0 8095
box 1 40 161 120
use via23_4  via23_4_241
timestamp 1696364841
transform 0 -1 8544 1 0 8095
box 1 40 161 120
use via23_4  via23_4_242
timestamp 1696364841
transform 0 -1 9844 1 0 7255
box 1 40 161 120
use via23_4  via23_4_243
timestamp 1696364841
transform 0 -1 8544 1 0 7255
box 1 40 161 120
use via23_4  via23_4_244
timestamp 1696364841
transform 0 -1 10616 1 0 8935
box 1 40 161 120
use via23_4  via23_4_245
timestamp 1696364841
transform 0 -1 5944 1 0 8935
box 1 40 161 120
use via23_4  via23_4_246
timestamp 1696364841
transform 0 -1 7244 1 0 8935
box 1 40 161 120
use via23_4  via23_4_247
timestamp 1696364841
transform 0 -1 8544 1 0 8935
box 1 40 161 120
use via23_4  via23_4_248
timestamp 1696364841
transform 0 -1 7244 1 0 7255
box 1 40 161 120
use via23_4  via23_4_249
timestamp 1696364841
transform 0 -1 6716 1 0 8935
box 1 40 161 120
use via23_4  via23_4_250
timestamp 1696364841
transform 0 -1 8016 1 0 8935
box 1 40 161 120
use via23_4  via23_4_251
timestamp 1696364841
transform 0 -1 9316 1 0 8935
box 1 40 161 120
use via23_4  via23_4_252
timestamp 1696364841
transform 0 -1 5944 1 0 7255
box 1 40 161 120
use via23_4  via23_4_253
timestamp 1696364841
transform 0 -1 10616 1 0 7255
box 1 40 161 120
use via23_4  via23_4_254
timestamp 1696364841
transform 0 -1 9316 1 0 7255
box 1 40 161 120
use via23_4  via23_4_255
timestamp 1696364841
transform 0 -1 8016 1 0 7255
box 1 40 161 120
use via23_4  via23_4_256
timestamp 1696364841
transform 0 -1 6716 1 0 7255
box 1 40 161 120
use via23_4  via23_4_257
timestamp 1696364841
transform 0 -1 21544 1 0 4735
box 1 40 161 120
use via23_4  via23_4_258
timestamp 1696364841
transform 0 -1 20244 1 0 4735
box 1 40 161 120
use via23_4  via23_4_259
timestamp 1696364841
transform 0 -1 18944 1 0 4735
box 1 40 161 120
use via23_4  via23_4_260
timestamp 1696364841
transform 0 -1 17644 1 0 4735
box 1 40 161 120
use via23_4  via23_4_261
timestamp 1696364841
transform 0 -1 21016 1 0 4735
box 1 40 161 120
use via23_4  via23_4_262
timestamp 1696364841
transform 0 -1 19716 1 0 4735
box 1 40 161 120
use via23_4  via23_4_263
timestamp 1696364841
transform 0 -1 18416 1 0 4735
box 1 40 161 120
use via23_4  via23_4_264
timestamp 1696364841
transform 0 -1 17116 1 0 4735
box 1 40 161 120
use via23_4  via23_4_265
timestamp 1696364841
transform 0 -1 20690 1 0 6415
box 1 40 161 120
use via23_4  via23_4_266
timestamp 1696364841
transform 0 -1 21544 1 0 5575
box 1 40 161 120
use via23_4  via23_4_267
timestamp 1696364841
transform 0 -1 20244 1 0 5575
box 1 40 161 120
use via23_4  via23_4_268
timestamp 1696364841
transform 0 -1 21544 1 0 6415
box 1 40 161 120
use via23_4  via23_4_269
timestamp 1696364841
transform 0 -1 21870 1 0 5575
box 1 40 161 120
use via23_4  via23_4_270
timestamp 1696364841
transform 0 -1 18944 1 0 5575
box 1 40 161 120
use via23_4  via23_4_271
timestamp 1696364841
transform 0 -1 21016 1 0 6415
box 1 40 161 120
use via23_4  via23_4_272
timestamp 1696364841
transform 0 -1 17644 1 0 5575
box 1 40 161 120
use via23_4  via23_4_273
timestamp 1696364841
transform 0 -1 20244 1 0 6415
box 1 40 161 120
use via23_4  via23_4_274
timestamp 1696364841
transform 0 -1 19716 1 0 6415
box 1 40 161 120
use via23_4  via23_4_275
timestamp 1696364841
transform 0 -1 18416 1 0 6415
box 1 40 161 120
use via23_4  via23_4_276
timestamp 1696364841
transform 0 -1 17116 1 0 6415
box 1 40 161 120
use via23_4  via23_4_277
timestamp 1696364841
transform 0 -1 21016 1 0 5575
box 1 40 161 120
use via23_4  via23_4_278
timestamp 1696364841
transform 0 -1 19716 1 0 5575
box 1 40 161 120
use via23_4  via23_4_279
timestamp 1696364841
transform 0 -1 18944 1 0 6415
box 1 40 161 120
use via23_4  via23_4_280
timestamp 1696364841
transform 0 -1 18416 1 0 5575
box 1 40 161 120
use via23_4  via23_4_281
timestamp 1696364841
transform 0 -1 17116 1 0 5575
box 1 40 161 120
use via23_4  via23_4_282
timestamp 1696364841
transform 0 -1 17644 1 0 6415
box 1 40 161 120
use via23_4  via23_4_283
timestamp 1696364841
transform 0 -1 12444 1 0 6415
box 1 40 161 120
use via23_4  via23_4_284
timestamp 1696364841
transform 0 -1 11144 1 0 6415
box 1 40 161 120
use via23_4  via23_4_285
timestamp 1696364841
transform 0 -1 13216 1 0 6415
box 1 40 161 120
use via23_4  via23_4_286
timestamp 1696364841
transform 0 -1 15044 1 0 4735
box 1 40 161 120
use via23_4  via23_4_287
timestamp 1696364841
transform 0 -1 15816 1 0 4735
box 1 40 161 120
use via23_4  via23_4_288
timestamp 1696364841
transform 0 -1 15816 1 0 6415
box 1 40 161 120
use via23_4  via23_4_289
timestamp 1696364841
transform 0 -1 14516 1 0 6415
box 1 40 161 120
use via23_4  via23_4_290
timestamp 1696364841
transform 0 -1 14516 1 0 4735
box 1 40 161 120
use via23_4  via23_4_291
timestamp 1696364841
transform 0 -1 13216 1 0 4735
box 1 40 161 120
use via23_4  via23_4_292
timestamp 1696364841
transform 0 -1 11916 1 0 6415
box 1 40 161 120
use via23_4  via23_4_293
timestamp 1696364841
transform 0 -1 16344 1 0 6415
box 1 40 161 120
use via23_4  via23_4_294
timestamp 1696364841
transform 0 -1 15044 1 0 6415
box 1 40 161 120
use via23_4  via23_4_295
timestamp 1696364841
transform 0 -1 11916 1 0 4735
box 1 40 161 120
use via23_4  via23_4_296
timestamp 1696364841
transform 0 -1 13744 1 0 4735
box 1 40 161 120
use via23_4  via23_4_297
timestamp 1696364841
transform 0 -1 12444 1 0 4735
box 1 40 161 120
use via23_4  via23_4_298
timestamp 1696364841
transform 0 -1 11144 1 0 4735
box 1 40 161 120
use via23_4  via23_4_299
timestamp 1696364841
transform 0 -1 16344 1 0 4735
box 1 40 161 120
use via23_4  via23_4_300
timestamp 1696364841
transform 0 -1 15816 1 0 5575
box 1 40 161 120
use via23_4  via23_4_301
timestamp 1696364841
transform 0 -1 14516 1 0 5575
box 1 40 161 120
use via23_4  via23_4_302
timestamp 1696364841
transform 0 -1 13216 1 0 5575
box 1 40 161 120
use via23_4  via23_4_303
timestamp 1696364841
transform 0 -1 16344 1 0 5575
box 1 40 161 120
use via23_4  via23_4_304
timestamp 1696364841
transform 0 -1 15044 1 0 5575
box 1 40 161 120
use via23_4  via23_4_305
timestamp 1696364841
transform 0 -1 13744 1 0 5575
box 1 40 161 120
use via23_4  via23_4_306
timestamp 1696364841
transform 0 -1 12444 1 0 5575
box 1 40 161 120
use via23_4  via23_4_307
timestamp 1696364841
transform 0 -1 11144 1 0 5575
box 1 40 161 120
use via23_4  via23_4_308
timestamp 1696364841
transform 0 -1 11916 1 0 5575
box 1 40 161 120
use via23_4  via23_4_309
timestamp 1696364841
transform 0 -1 13744 1 0 6415
box 1 40 161 120
use via23_4  via23_4_310
timestamp 1696364841
transform 0 -1 13216 1 0 7255
box 1 40 161 120
use via23_4  via23_4_311
timestamp 1696364841
transform 0 -1 11916 1 0 7255
box 1 40 161 120
use via23_4  via23_4_312
timestamp 1696364841
transform 0 -1 16344 1 0 8095
box 1 40 161 120
use via23_4  via23_4_313
timestamp 1696364841
transform 0 -1 13744 1 0 8095
box 1 40 161 120
use via23_4  via23_4_314
timestamp 1696364841
transform 0 -1 15816 1 0 8095
box 1 40 161 120
use via23_4  via23_4_315
timestamp 1696364841
transform 0 -1 14516 1 0 8095
box 1 40 161 120
use via23_4  via23_4_316
timestamp 1696364841
transform 0 -1 16344 1 0 7255
box 1 40 161 120
use via23_4  via23_4_317
timestamp 1696364841
transform 0 -1 13216 1 0 8095
box 1 40 161 120
use via23_4  via23_4_318
timestamp 1696364841
transform 0 -1 11916 1 0 8095
box 1 40 161 120
use via23_4  via23_4_319
timestamp 1696364841
transform 0 -1 15044 1 0 8095
box 1 40 161 120
use via23_4  via23_4_320
timestamp 1696364841
transform 0 -1 12444 1 0 8095
box 1 40 161 120
use via23_4  via23_4_321
timestamp 1696364841
transform 0 -1 15044 1 0 7255
box 1 40 161 120
use via23_4  via23_4_322
timestamp 1696364841
transform 0 -1 13744 1 0 7255
box 1 40 161 120
use via23_4  via23_4_323
timestamp 1696364841
transform 0 -1 12444 1 0 7255
box 1 40 161 120
use via23_4  via23_4_324
timestamp 1696364841
transform 0 -1 11144 1 0 8095
box 1 40 161 120
use via23_4  via23_4_325
timestamp 1696364841
transform 0 -1 11144 1 0 7255
box 1 40 161 120
use via23_4  via23_4_326
timestamp 1696364841
transform 0 -1 11144 1 0 8935
box 1 40 161 120
use via23_4  via23_4_327
timestamp 1696364841
transform 0 -1 12444 1 0 8935
box 1 40 161 120
use via23_4  via23_4_328
timestamp 1696364841
transform 0 -1 13744 1 0 8935
box 1 40 161 120
use via23_4  via23_4_329
timestamp 1696364841
transform 0 -1 15044 1 0 8935
box 1 40 161 120
use via23_4  via23_4_330
timestamp 1696364841
transform 0 -1 16344 1 0 8935
box 1 40 161 120
use via23_4  via23_4_331
timestamp 1696364841
transform 0 -1 11916 1 0 8935
box 1 40 161 120
use via23_4  via23_4_332
timestamp 1696364841
transform 0 -1 13216 1 0 8935
box 1 40 161 120
use via23_4  via23_4_333
timestamp 1696364841
transform 0 -1 14516 1 0 8935
box 1 40 161 120
use via23_4  via23_4_334
timestamp 1696364841
transform 0 -1 15816 1 0 8935
box 1 40 161 120
use via23_4  via23_4_335
timestamp 1696364841
transform 0 -1 15816 1 0 7255
box 1 40 161 120
use via23_4  via23_4_336
timestamp 1696364841
transform 0 -1 14516 1 0 7255
box 1 40 161 120
use via23_4  via23_4_337
timestamp 1696364841
transform 0 -1 20244 1 0 8095
box 1 40 161 120
use via23_4  via23_4_338
timestamp 1696364841
transform 0 -1 18944 1 0 8095
box 1 40 161 120
use via23_4  via23_4_339
timestamp 1696364841
transform 0 -1 21016 1 0 8095
box 1 40 161 120
use via23_4  via23_4_340
timestamp 1696364841
transform 0 -1 19716 1 0 8095
box 1 40 161 120
use via23_4  via23_4_341
timestamp 1696364841
transform 0 -1 17644 1 0 8095
box 1 40 161 120
use via23_4  via23_4_342
timestamp 1696364841
transform 0 -1 17644 1 0 8935
box 1 40 161 120
use via23_4  via23_4_343
timestamp 1696364841
transform 0 -1 18944 1 0 8935
box 1 40 161 120
use via23_4  via23_4_344
timestamp 1696364841
transform 0 -1 20244 1 0 8935
box 1 40 161 120
use via23_4  via23_4_345
timestamp 1696364841
transform 0 -1 17116 1 0 8935
box 1 40 161 120
use via23_4  via23_4_346
timestamp 1696364841
transform 0 -1 18416 1 0 8935
box 1 40 161 120
use via23_4  via23_4_347
timestamp 1696364841
transform 0 -1 19716 1 0 8935
box 1 40 161 120
use via23_4  via23_4_348
timestamp 1696364841
transform 0 -1 21016 1 0 7255
box 1 40 161 120
use via23_4  via23_4_349
timestamp 1696364841
transform 0 -1 19716 1 0 7255
box 1 40 161 120
use via23_4  via23_4_350
timestamp 1696364841
transform 0 -1 18416 1 0 7255
box 1 40 161 120
use via23_4  via23_4_351
timestamp 1696364841
transform 0 -1 17116 1 0 7255
box 1 40 161 120
use via23_4  via23_4_352
timestamp 1696364841
transform 0 -1 21544 1 0 7255
box 1 40 161 120
use via23_4  via23_4_353
timestamp 1696364841
transform 0 -1 21016 1 0 8935
box 1 40 161 120
use via23_4  via23_4_354
timestamp 1696364841
transform 0 -1 21544 1 0 8935
box 1 40 161 120
use via23_4  via23_4_355
timestamp 1696364841
transform 0 -1 20244 1 0 7255
box 1 40 161 120
use via23_4  via23_4_356
timestamp 1696364841
transform 0 -1 18944 1 0 7255
box 1 40 161 120
use via23_4  via23_4_357
timestamp 1696364841
transform 0 -1 17644 1 0 7255
box 1 40 161 120
use via23_4  via23_4_358
timestamp 1696364841
transform 0 -1 18416 1 0 8095
box 1 40 161 120
use via23_4  via23_4_359
timestamp 1696364841
transform 0 -1 17116 1 0 8095
box 1 40 161 120
use via23_4  via23_4_360
timestamp 1696364841
transform 0 -1 21544 1 0 8095
box 1 40 161 120
use via23_4  via23_4_361
timestamp 1696364841
transform 1 0 38439 0 -1 124
box 1 40 161 120
use via23_4  via23_4_362
timestamp 1696364841
transform 0 -1 39216 1 0 1375
box 1 40 161 120
use via23_4  via23_4_363
timestamp 1696364841
transform 0 -1 40516 1 0 1375
box 1 40 161 120
use via23_4  via23_4_364
timestamp 1696364841
transform 0 -1 41816 1 0 1375
box 1 40 161 120
use via23_4  via23_4_365
timestamp 1696364841
transform 0 -1 43116 1 0 1375
box 1 40 161 120
use via23_4  via23_4_366
timestamp 1696364841
transform 0 -1 42344 1 0 1375
box 1 40 161 120
use via23_4  via23_4_367
timestamp 1696364841
transform 0 -1 43644 1 0 1375
box 1 40 161 120
use via23_4  via23_4_368
timestamp 1696364841
transform 0 -1 39744 1 0 1375
box 1 40 161 120
use via23_4  via23_4_369
timestamp 1696364841
transform 0 -1 41044 1 0 1375
box 1 40 161 120
use via23_4  via23_4_370
timestamp 1696364841
transform 0 -1 38444 1 0 1375
box 1 40 161 120
use via23_4  via23_4_371
timestamp 1696364841
transform 1 0 41039 0 -1 284
box 1 40 161 120
use via23_4  via23_4_372
timestamp 1696364841
transform 1 0 42339 0 -1 124
box 1 40 161 120
use via23_4  via23_4_373
timestamp 1696364841
transform 1 0 39739 0 -1 124
box 1 40 161 120
use via23_4  via23_4_374
timestamp 1696364841
transform 1 0 33239 0 -1 444
box 1 40 161 120
use via23_4  via23_4_375
timestamp 1696364841
transform 0 -1 35844 1 0 1375
box 1 40 161 120
use via23_4  via23_4_376
timestamp 1696364841
transform 0 -1 37144 1 0 1375
box 1 40 161 120
use via23_4  via23_4_377
timestamp 1696364841
transform 0 -1 34544 1 0 1375
box 1 40 161 120
use via23_4  via23_4_378
timestamp 1696364841
transform 0 -1 34016 1 0 1375
box 1 40 161 120
use via23_4  via23_4_379
timestamp 1696364841
transform 0 -1 35316 1 0 1375
box 1 40 161 120
use via23_4  via23_4_380
timestamp 1696364841
transform 0 -1 36616 1 0 1375
box 1 40 161 120
use via23_4  via23_4_381
timestamp 1696364841
transform 0 -1 37916 1 0 1375
box 1 40 161 120
use via23_4  via23_4_382
timestamp 1696364841
transform 0 -1 33244 1 0 1375
box 1 40 161 120
use via23_4  via23_4_383
timestamp 1696364841
transform 1 0 37139 0 -1 284
box 1 40 161 120
use via23_4  via23_4_384
timestamp 1696364841
transform 1 0 35839 0 -1 124
box 1 40 161 120
use via23_4  via23_4_385
timestamp 1696364841
transform 1 0 34539 0 -1 124
box 1 40 161 120
use via23_4  via23_4_386
timestamp 1696364841
transform 0 -1 37144 1 0 3895
box 1 40 161 120
use via23_4  via23_4_387
timestamp 1696364841
transform 0 -1 37916 1 0 3055
box 1 40 161 120
use via23_4  via23_4_388
timestamp 1696364841
transform 0 -1 36616 1 0 3055
box 1 40 161 120
use via23_4  via23_4_389
timestamp 1696364841
transform 0 -1 35316 1 0 3055
box 1 40 161 120
use via23_4  via23_4_390
timestamp 1696364841
transform 0 -1 34016 1 0 3055
box 1 40 161 120
use via23_4  via23_4_391
timestamp 1696364841
transform 0 -1 37916 1 0 3895
box 1 40 161 120
use via23_4  via23_4_392
timestamp 1696364841
transform 0 -1 37144 1 0 3055
box 1 40 161 120
use via23_4  via23_4_393
timestamp 1696364841
transform 0 -1 35844 1 0 3055
box 1 40 161 120
use via23_4  via23_4_394
timestamp 1696364841
transform 0 -1 34016 1 0 2215
box 1 40 161 120
use via23_4  via23_4_395
timestamp 1696364841
transform 0 -1 36616 1 0 3895
box 1 40 161 120
use via23_4  via23_4_396
timestamp 1696364841
transform 0 -1 37916 1 0 2215
box 1 40 161 120
use via23_4  via23_4_397
timestamp 1696364841
transform 0 -1 36616 1 0 2215
box 1 40 161 120
use via23_4  via23_4_398
timestamp 1696364841
transform 0 -1 37144 1 0 2215
box 1 40 161 120
use via23_4  via23_4_399
timestamp 1696364841
transform 0 -1 35844 1 0 2215
box 1 40 161 120
use via23_4  via23_4_400
timestamp 1696364841
transform 0 -1 34544 1 0 2215
box 1 40 161 120
use via23_4  via23_4_401
timestamp 1696364841
transform 0 -1 33244 1 0 2215
box 1 40 161 120
use via23_4  via23_4_402
timestamp 1696364841
transform 0 -1 35316 1 0 2215
box 1 40 161 120
use via23_4  via23_4_403
timestamp 1696364841
transform 0 -1 35316 1 0 3895
box 1 40 161 120
use via23_4  via23_4_404
timestamp 1696364841
transform 0 -1 34016 1 0 3895
box 1 40 161 120
use via23_4  via23_4_405
timestamp 1696364841
transform 0 -1 35844 1 0 3895
box 1 40 161 120
use via23_4  via23_4_406
timestamp 1696364841
transform 0 -1 34544 1 0 3895
box 1 40 161 120
use via23_4  via23_4_407
timestamp 1696364841
transform 0 -1 34544 1 0 3055
box 1 40 161 120
use via23_4  via23_4_408
timestamp 1696364841
transform 0 -1 33244 1 0 3895
box 1 40 161 120
use via23_4  via23_4_409
timestamp 1696364841
transform 0 -1 33244 1 0 3055
box 1 40 161 120
use via23_4  via23_4_410
timestamp 1696364841
transform 0 -1 42344 1 0 3055
box 1 40 161 120
use via23_4  via23_4_411
timestamp 1696364841
transform 0 -1 40516 1 0 3055
box 1 40 161 120
use via23_4  via23_4_412
timestamp 1696364841
transform 0 -1 39216 1 0 3055
box 1 40 161 120
use via23_4  via23_4_413
timestamp 1696364841
transform 0 -1 43644 1 0 3055
box 1 40 161 120
use via23_4  via23_4_414
timestamp 1696364841
transform 0 -1 43116 1 0 3055
box 1 40 161 120
use via23_4  via23_4_415
timestamp 1696364841
transform 0 -1 41044 1 0 3055
box 1 40 161 120
use via23_4  via23_4_416
timestamp 1696364841
transform 0 -1 39744 1 0 3055
box 1 40 161 120
use via23_4  via23_4_417
timestamp 1696364841
transform 0 -1 38444 1 0 3055
box 1 40 161 120
use via23_4  via23_4_418
timestamp 1696364841
transform 0 -1 43116 1 0 3895
box 1 40 161 120
use via23_4  via23_4_419
timestamp 1696364841
transform 0 -1 43644 1 0 3895
box 1 40 161 120
use via23_4  via23_4_420
timestamp 1696364841
transform 0 -1 42344 1 0 3895
box 1 40 161 120
use via23_4  via23_4_421
timestamp 1696364841
transform 0 -1 41816 1 0 3055
box 1 40 161 120
use via23_4  via23_4_422
timestamp 1696364841
transform 0 -1 41816 1 0 2215
box 1 40 161 120
use via23_4  via23_4_423
timestamp 1696364841
transform 0 -1 42344 1 0 2215
box 1 40 161 120
use via23_4  via23_4_424
timestamp 1696364841
transform 0 -1 41044 1 0 2215
box 1 40 161 120
use via23_4  via23_4_425
timestamp 1696364841
transform 0 -1 41044 1 0 3895
box 1 40 161 120
use via23_4  via23_4_426
timestamp 1696364841
transform 0 -1 39744 1 0 3895
box 1 40 161 120
use via23_4  via23_4_427
timestamp 1696364841
transform 0 -1 43116 1 0 2215
box 1 40 161 120
use via23_4  via23_4_428
timestamp 1696364841
transform 0 -1 38444 1 0 3895
box 1 40 161 120
use via23_4  via23_4_429
timestamp 1696364841
transform 0 -1 43644 1 0 2215
box 1 40 161 120
use via23_4  via23_4_430
timestamp 1696364841
transform 0 -1 39744 1 0 2215
box 1 40 161 120
use via23_4  via23_4_431
timestamp 1696364841
transform 0 -1 38444 1 0 2215
box 1 40 161 120
use via23_4  via23_4_432
timestamp 1696364841
transform 0 -1 40516 1 0 2215
box 1 40 161 120
use via23_4  via23_4_433
timestamp 1696364841
transform 0 -1 39216 1 0 2215
box 1 40 161 120
use via23_4  via23_4_434
timestamp 1696364841
transform 0 -1 41816 1 0 3895
box 1 40 161 120
use via23_4  via23_4_435
timestamp 1696364841
transform 0 -1 40516 1 0 3895
box 1 40 161 120
use via23_4  via23_4_436
timestamp 1696364841
transform 0 -1 39216 1 0 3895
box 1 40 161 120
use via23_4  via23_4_437
timestamp 1696364841
transform 0 -1 27516 1 0 1375
box 1 40 161 120
use via23_4  via23_4_438
timestamp 1696364841
transform 0 -1 28816 1 0 1375
box 1 40 161 120
use via23_4  via23_4_439
timestamp 1696364841
transform 0 -1 32716 1 0 1375
box 1 40 161 120
use via23_4  via23_4_440
timestamp 1696364841
transform 1 0 29339 0 -1 124
box 1 40 161 120
use via23_4  via23_4_441
timestamp 1696364841
transform 1 0 28039 0 -1 444
box 1 40 161 120
use via23_4  via23_4_442
timestamp 1696364841
transform 1 0 31939 0 -1 284
box 1 40 161 120
use via23_4  via23_4_443
timestamp 1696364841
transform 1 0 30639 0 -1 124
box 1 40 161 120
use via23_4  via23_4_444
timestamp 1696364841
transform 0 -1 30644 1 0 1375
box 1 40 161 120
use via23_4  via23_4_445
timestamp 1696364841
transform 0 -1 31944 1 0 1375
box 1 40 161 120
use via23_4  via23_4_446
timestamp 1696364841
transform 0 -1 31416 1 0 1375
box 1 40 161 120
use via23_4  via23_4_447
timestamp 1696364841
transform 0 -1 30116 1 0 1375
box 1 40 161 120
use via23_4  via23_4_448
timestamp 1696364841
transform 0 -1 28044 1 0 1375
box 1 40 161 120
use via23_4  via23_4_449
timestamp 1696364841
transform 0 -1 29344 1 0 1375
box 1 40 161 120
use via23_4  via23_4_450
timestamp 1696364841
transform 1 0 25439 0 -1 124
box 1 40 161 120
use via23_4  via23_4_451
timestamp 1696364841
transform -1 0 22401 0 -1 1084
box 1 40 161 120
use via23_4  via23_4_452
timestamp 1696364841
transform -1 0 22401 0 -1 -356
box 1 40 161 120
use via23_4  via23_4_453
timestamp 1696364841
transform 0 -1 26744 1 0 1375
box 1 40 161 120
use via23_4  via23_4_454
timestamp 1696364841
transform 0 -1 22844 1 0 1375
box 1 40 161 120
use via23_4  via23_4_455
timestamp 1696364841
transform 0 -1 22316 1 0 1375
box 1 40 161 120
use via23_4  via23_4_456
timestamp 1696364841
transform 0 -1 23616 1 0 1375
box 1 40 161 120
use via23_4  via23_4_457
timestamp 1696364841
transform 0 -1 24916 1 0 1375
box 1 40 161 120
use via23_4  via23_4_458
timestamp 1696364841
transform 0 -1 26216 1 0 1375
box 1 40 161 120
use via23_4  via23_4_459
timestamp 1696364841
transform 0 -1 24144 1 0 1375
box 1 40 161 120
use via23_4  via23_4_460
timestamp 1696364841
transform 0 -1 25444 1 0 1375
box 1 40 161 120
use via23_4  via23_4_461
timestamp 1696364841
transform 1 0 22839 0 -1 764
box 1 40 161 120
use via23_4  via23_4_462
timestamp 1696364841
transform 1 0 24139 0 -1 604
box 1 40 161 120
use via23_4  via23_4_463
timestamp 1696364841
transform 1 0 26739 0 -1 284
box 1 40 161 120
use via23_4  via23_4_464
timestamp 1696364841
transform 0 -1 22844 1 0 2215
box 1 40 161 120
use via23_4  via23_4_465
timestamp 1696364841
transform 0 -1 26216 1 0 2215
box 1 40 161 120
use via23_4  via23_4_466
timestamp 1696364841
transform 0 -1 24916 1 0 2215
box 1 40 161 120
use via23_4  via23_4_467
timestamp 1696364841
transform 0 -1 23616 1 0 2215
box 1 40 161 120
use via23_4  via23_4_468
timestamp 1696364841
transform 0 -1 23170 1 0 3895
box 1 40 161 120
use via23_4  via23_4_469
timestamp 1696364841
transform 0 -1 26216 1 0 3055
box 1 40 161 120
use via23_4  via23_4_470
timestamp 1696364841
transform 0 -1 22316 1 0 3895
box 1 40 161 120
use via23_4  via23_4_471
timestamp 1696364841
transform 0 -1 22316 1 0 2215
box 1 40 161 120
use via23_4  via23_4_472
timestamp 1696364841
transform 0 -1 26744 1 0 3895
box 1 40 161 120
use via23_4  via23_4_473
timestamp 1696364841
transform 0 -1 23616 1 0 3895
box 1 40 161 120
use via23_4  via23_4_474
timestamp 1696364841
transform 0 -1 26216 1 0 3895
box 1 40 161 120
use via23_4  via23_4_475
timestamp 1696364841
transform 0 -1 23616 1 0 3055
box 1 40 161 120
use via23_4  via23_4_476
timestamp 1696364841
transform 0 -1 22844 1 0 3895
box 1 40 161 120
use via23_4  via23_4_477
timestamp 1696364841
transform 0 -1 22316 1 0 3055
box 1 40 161 120
use via23_4  via23_4_478
timestamp 1696364841
transform 0 -1 25444 1 0 3895
box 1 40 161 120
use via23_4  via23_4_479
timestamp 1696364841
transform 0 -1 26744 1 0 3055
box 1 40 161 120
use via23_4  via23_4_480
timestamp 1696364841
transform 0 -1 25444 1 0 3055
box 1 40 161 120
use via23_4  via23_4_481
timestamp 1696364841
transform 0 -1 24144 1 0 3055
box 1 40 161 120
use via23_4  via23_4_482
timestamp 1696364841
transform 0 -1 22844 1 0 3055
box 1 40 161 120
use via23_4  via23_4_483
timestamp 1696364841
transform 0 -1 24144 1 0 3895
box 1 40 161 120
use via23_4  via23_4_484
timestamp 1696364841
transform 0 -1 26744 1 0 2215
box 1 40 161 120
use via23_4  via23_4_485
timestamp 1696364841
transform 0 -1 24916 1 0 3055
box 1 40 161 120
use via23_4  via23_4_486
timestamp 1696364841
transform 0 -1 24916 1 0 3895
box 1 40 161 120
use via23_4  via23_4_487
timestamp 1696364841
transform 0 -1 25444 1 0 2215
box 1 40 161 120
use via23_4  via23_4_488
timestamp 1696364841
transform 0 -1 24144 1 0 2215
box 1 40 161 120
use via23_4  via23_4_489
timestamp 1696364841
transform 0 -1 28044 1 0 3895
box 1 40 161 120
use via23_4  via23_4_490
timestamp 1696364841
transform 0 -1 32716 1 0 3895
box 1 40 161 120
use via23_4  via23_4_491
timestamp 1696364841
transform 0 -1 27516 1 0 3895
box 1 40 161 120
use via23_4  via23_4_492
timestamp 1696364841
transform 0 -1 31944 1 0 3895
box 1 40 161 120
use via23_4  via23_4_493
timestamp 1696364841
transform 0 -1 30644 1 0 3895
box 1 40 161 120
use via23_4  via23_4_494
timestamp 1696364841
transform 0 -1 29344 1 0 3895
box 1 40 161 120
use via23_4  via23_4_495
timestamp 1696364841
transform 0 -1 31416 1 0 2215
box 1 40 161 120
use via23_4  via23_4_496
timestamp 1696364841
transform 0 -1 30116 1 0 2215
box 1 40 161 120
use via23_4  via23_4_497
timestamp 1696364841
transform 0 -1 28816 1 0 2215
box 1 40 161 120
use via23_4  via23_4_498
timestamp 1696364841
transform 0 -1 27516 1 0 2215
box 1 40 161 120
use via23_4  via23_4_499
timestamp 1696364841
transform 0 -1 27516 1 0 3055
box 1 40 161 120
use via23_4  via23_4_500
timestamp 1696364841
transform 0 -1 31944 1 0 3055
box 1 40 161 120
use via23_4  via23_4_501
timestamp 1696364841
transform 0 -1 32716 1 0 3055
box 1 40 161 120
use via23_4  via23_4_502
timestamp 1696364841
transform 0 -1 31416 1 0 3055
box 1 40 161 120
use via23_4  via23_4_503
timestamp 1696364841
transform 0 -1 30116 1 0 3055
box 1 40 161 120
use via23_4  via23_4_504
timestamp 1696364841
transform 0 -1 28816 1 0 3055
box 1 40 161 120
use via23_4  via23_4_505
timestamp 1696364841
transform 0 -1 31944 1 0 2215
box 1 40 161 120
use via23_4  via23_4_506
timestamp 1696364841
transform 0 -1 30644 1 0 2215
box 1 40 161 120
use via23_4  via23_4_507
timestamp 1696364841
transform 0 -1 29344 1 0 2215
box 1 40 161 120
use via23_4  via23_4_508
timestamp 1696364841
transform 0 -1 28044 1 0 2215
box 1 40 161 120
use via23_4  via23_4_509
timestamp 1696364841
transform 0 -1 32716 1 0 2215
box 1 40 161 120
use via23_4  via23_4_510
timestamp 1696364841
transform 0 -1 31416 1 0 3895
box 1 40 161 120
use via23_4  via23_4_511
timestamp 1696364841
transform 0 -1 30644 1 0 3055
box 1 40 161 120
use via23_4  via23_4_512
timestamp 1696364841
transform 0 -1 29344 1 0 3055
box 1 40 161 120
use via23_4  via23_4_513
timestamp 1696364841
transform 0 -1 28044 1 0 3055
box 1 40 161 120
use via23_4  via23_4_514
timestamp 1696364841
transform 0 -1 30116 1 0 3895
box 1 40 161 120
use via23_4  via23_4_515
timestamp 1696364841
transform 0 -1 28816 1 0 3895
box 1 40 161 120
use via23_4  via23_4_516
timestamp 1696364841
transform 0 -1 29344 1 0 6415
box 1 40 161 120
use via23_4  via23_4_517
timestamp 1696364841
transform 0 -1 31944 1 0 6415
box 1 40 161 120
use via23_4  via23_4_518
timestamp 1696364841
transform 0 -1 31944 1 0 5575
box 1 40 161 120
use via23_4  via23_4_519
timestamp 1696364841
transform 0 -1 30644 1 0 5575
box 1 40 161 120
use via23_4  via23_4_520
timestamp 1696364841
transform 0 -1 29344 1 0 5575
box 1 40 161 120
use via23_4  via23_4_521
timestamp 1696364841
transform 0 -1 28044 1 0 5575
box 1 40 161 120
use via23_4  via23_4_522
timestamp 1696364841
transform 0 -1 32716 1 0 5575
box 1 40 161 120
use via23_4  via23_4_523
timestamp 1696364841
transform 0 -1 31416 1 0 5575
box 1 40 161 120
use via23_4  via23_4_524
timestamp 1696364841
transform 0 -1 30116 1 0 5575
box 1 40 161 120
use via23_4  via23_4_525
timestamp 1696364841
transform 0 -1 28816 1 0 5575
box 1 40 161 120
use via23_4  via23_4_526
timestamp 1696364841
transform 0 -1 27516 1 0 5575
box 1 40 161 120
use via23_4  via23_4_527
timestamp 1696364841
transform 0 -1 31944 1 0 4735
box 1 40 161 120
use via23_4  via23_4_528
timestamp 1696364841
transform 0 -1 30644 1 0 4735
box 1 40 161 120
use via23_4  via23_4_529
timestamp 1696364841
transform 0 -1 29344 1 0 4735
box 1 40 161 120
use via23_4  via23_4_530
timestamp 1696364841
transform 0 -1 28044 1 0 4735
box 1 40 161 120
use via23_4  via23_4_531
timestamp 1696364841
transform 0 -1 32716 1 0 4735
box 1 40 161 120
use via23_4  via23_4_532
timestamp 1696364841
transform 0 -1 31416 1 0 4735
box 1 40 161 120
use via23_4  via23_4_533
timestamp 1696364841
transform 0 -1 30116 1 0 4735
box 1 40 161 120
use via23_4  via23_4_534
timestamp 1696364841
transform 0 -1 28816 1 0 4735
box 1 40 161 120
use via23_4  via23_4_535
timestamp 1696364841
transform 0 -1 27516 1 0 4735
box 1 40 161 120
use via23_4  via23_4_536
timestamp 1696364841
transform 0 -1 30644 1 0 6415
box 1 40 161 120
use via23_4  via23_4_537
timestamp 1696364841
transform 0 -1 32716 1 0 6415
box 1 40 161 120
use via23_4  via23_4_538
timestamp 1696364841
transform 0 -1 31416 1 0 6415
box 1 40 161 120
use via23_4  via23_4_539
timestamp 1696364841
transform 0 -1 30116 1 0 6415
box 1 40 161 120
use via23_4  via23_4_540
timestamp 1696364841
transform 0 -1 28816 1 0 6415
box 1 40 161 120
use via23_4  via23_4_541
timestamp 1696364841
transform 0 -1 27516 1 0 6415
box 1 40 161 120
use via23_4  via23_4_542
timestamp 1696364841
transform 0 -1 28044 1 0 6415
box 1 40 161 120
use via23_4  via23_4_543
timestamp 1696364841
transform 0 -1 23170 1 0 6415
box 1 40 161 120
use via23_4  via23_4_544
timestamp 1696364841
transform 0 -1 21990 1 0 4735
box 1 40 161 120
use via23_4  via23_4_545
timestamp 1696364841
transform 0 -1 24144 1 0 4735
box 1 40 161 120
use via23_4  via23_4_546
timestamp 1696364841
transform 0 -1 22844 1 0 4735
box 1 40 161 120
use via23_4  via23_4_547
timestamp 1696364841
transform 0 -1 24144 1 0 5575
box 1 40 161 120
use via23_4  via23_4_548
timestamp 1696364841
transform 0 -1 22844 1 0 5575
box 1 40 161 120
use via23_4  via23_4_549
timestamp 1696364841
transform 0 -1 26216 1 0 6415
box 1 40 161 120
use via23_4  via23_4_550
timestamp 1696364841
transform 0 -1 24916 1 0 6415
box 1 40 161 120
use via23_4  via23_4_551
timestamp 1696364841
transform 0 -1 23616 1 0 6415
box 1 40 161 120
use via23_4  via23_4_552
timestamp 1696364841
transform 0 -1 22316 1 0 6415
box 1 40 161 120
use via23_4  via23_4_553
timestamp 1696364841
transform 0 -1 26216 1 0 5575
box 1 40 161 120
use via23_4  via23_4_554
timestamp 1696364841
transform 0 -1 24916 1 0 5575
box 1 40 161 120
use via23_4  via23_4_555
timestamp 1696364841
transform 0 -1 26744 1 0 6415
box 1 40 161 120
use via23_4  via23_4_556
timestamp 1696364841
transform 0 -1 25444 1 0 6415
box 1 40 161 120
use via23_4  via23_4_557
timestamp 1696364841
transform 0 -1 24144 1 0 6415
box 1 40 161 120
use via23_4  via23_4_558
timestamp 1696364841
transform 0 -1 22844 1 0 6415
box 1 40 161 120
use via23_4  via23_4_559
timestamp 1696364841
transform 0 -1 23616 1 0 5575
box 1 40 161 120
use via23_4  via23_4_560
timestamp 1696364841
transform 0 -1 26744 1 0 5575
box 1 40 161 120
use via23_4  via23_4_561
timestamp 1696364841
transform 0 -1 25444 1 0 5575
box 1 40 161 120
use via23_4  via23_4_562
timestamp 1696364841
transform 0 -1 22316 1 0 5575
box 1 40 161 120
use via23_4  via23_4_563
timestamp 1696364841
transform 0 -1 26216 1 0 4735
box 1 40 161 120
use via23_4  via23_4_564
timestamp 1696364841
transform 0 -1 24916 1 0 4735
box 1 40 161 120
use via23_4  via23_4_565
timestamp 1696364841
transform 0 -1 23616 1 0 4735
box 1 40 161 120
use via23_4  via23_4_566
timestamp 1696364841
transform 0 -1 22316 1 0 4735
box 1 40 161 120
use via23_4  via23_4_567
timestamp 1696364841
transform 0 -1 26744 1 0 4735
box 1 40 161 120
use via23_4  via23_4_568
timestamp 1696364841
transform 0 -1 25444 1 0 4735
box 1 40 161 120
use via23_4  via23_4_569
timestamp 1696364841
transform 0 -1 26216 1 0 7255
box 1 40 161 120
use via23_4  via23_4_570
timestamp 1696364841
transform 0 -1 24916 1 0 7255
box 1 40 161 120
use via23_4  via23_4_571
timestamp 1696364841
transform 0 -1 23616 1 0 7255
box 1 40 161 120
use via23_4  via23_4_572
timestamp 1696364841
transform 0 -1 22844 1 0 8095
box 1 40 161 120
use via23_4  via23_4_573
timestamp 1696364841
transform 0 -1 23616 1 0 8095
box 1 40 161 120
use via23_4  via23_4_574
timestamp 1696364841
transform 0 -1 22316 1 0 8095
box 1 40 161 120
use via23_4  via23_4_575
timestamp 1696364841
transform 0 -1 26744 1 0 7255
box 1 40 161 120
use via23_4  via23_4_576
timestamp 1696364841
transform 0 -1 25444 1 0 7255
box 1 40 161 120
use via23_4  via23_4_577
timestamp 1696364841
transform 0 -1 24144 1 0 7255
box 1 40 161 120
use via23_4  via23_4_578
timestamp 1696364841
transform 0 -1 22844 1 0 7255
box 1 40 161 120
use via23_4  via23_4_579
timestamp 1696364841
transform 0 -1 22316 1 0 7255
box 1 40 161 120
use via23_4  via23_4_580
timestamp 1696364841
transform 0 -1 26744 1 0 8095
box 1 40 161 120
use via23_4  via23_4_581
timestamp 1696364841
transform 0 -1 25444 1 0 8095
box 1 40 161 120
use via23_4  via23_4_582
timestamp 1696364841
transform 0 -1 24144 1 0 8095
box 1 40 161 120
use via23_4  via23_4_583
timestamp 1696364841
transform 0 -1 22316 1 0 8935
box 1 40 161 120
use via23_4  via23_4_584
timestamp 1696364841
transform 0 -1 22844 1 0 8935
box 1 40 161 120
use via23_4  via23_4_585
timestamp 1696364841
transform 0 -1 24144 1 0 8935
box 1 40 161 120
use via23_4  via23_4_586
timestamp 1696364841
transform 0 -1 25444 1 0 8935
box 1 40 161 120
use via23_4  via23_4_587
timestamp 1696364841
transform 0 -1 26744 1 0 8935
box 1 40 161 120
use via23_4  via23_4_588
timestamp 1696364841
transform 0 -1 23616 1 0 8935
box 1 40 161 120
use via23_4  via23_4_589
timestamp 1696364841
transform 0 -1 24916 1 0 8935
box 1 40 161 120
use via23_4  via23_4_590
timestamp 1696364841
transform 0 -1 26216 1 0 8935
box 1 40 161 120
use via23_4  via23_4_591
timestamp 1696364841
transform 0 -1 26216 1 0 8095
box 1 40 161 120
use via23_4  via23_4_592
timestamp 1696364841
transform 0 -1 24916 1 0 8095
box 1 40 161 120
use via23_4  via23_4_593
timestamp 1696364841
transform 0 -1 27516 1 0 8935
box 1 40 161 120
use via23_4  via23_4_594
timestamp 1696364841
transform 0 -1 28816 1 0 8935
box 1 40 161 120
use via23_4  via23_4_595
timestamp 1696364841
transform 0 -1 30116 1 0 8935
box 1 40 161 120
use via23_4  via23_4_596
timestamp 1696364841
transform 0 -1 31416 1 0 8935
box 1 40 161 120
use via23_4  via23_4_597
timestamp 1696364841
transform 0 -1 32716 1 0 8935
box 1 40 161 120
use via23_4  via23_4_598
timestamp 1696364841
transform 0 -1 28044 1 0 8935
box 1 40 161 120
use via23_4  via23_4_599
timestamp 1696364841
transform 0 -1 29344 1 0 8935
box 1 40 161 120
use via23_4  via23_4_600
timestamp 1696364841
transform 0 -1 30644 1 0 8935
box 1 40 161 120
use via23_4  via23_4_601
timestamp 1696364841
transform 0 -1 31944 1 0 8935
box 1 40 161 120
use via23_4  via23_4_602
timestamp 1696364841
transform 0 -1 32716 1 0 7255
box 1 40 161 120
use via23_4  via23_4_603
timestamp 1696364841
transform 0 -1 31416 1 0 7255
box 1 40 161 120
use via23_4  via23_4_604
timestamp 1696364841
transform 0 -1 30116 1 0 7255
box 1 40 161 120
use via23_4  via23_4_605
timestamp 1696364841
transform 0 -1 28816 1 0 7255
box 1 40 161 120
use via23_4  via23_4_606
timestamp 1696364841
transform 0 -1 27516 1 0 7255
box 1 40 161 120
use via23_4  via23_4_607
timestamp 1696364841
transform 0 -1 31944 1 0 7255
box 1 40 161 120
use via23_4  via23_4_608
timestamp 1696364841
transform 0 -1 30644 1 0 7255
box 1 40 161 120
use via23_4  via23_4_609
timestamp 1696364841
transform 0 -1 29344 1 0 7255
box 1 40 161 120
use via23_4  via23_4_610
timestamp 1696364841
transform 0 -1 28044 1 0 7255
box 1 40 161 120
use via23_4  via23_4_611
timestamp 1696364841
transform 0 -1 32716 1 0 8095
box 1 40 161 120
use via23_4  via23_4_612
timestamp 1696364841
transform 0 -1 31416 1 0 8095
box 1 40 161 120
use via23_4  via23_4_613
timestamp 1696364841
transform 0 -1 30116 1 0 8095
box 1 40 161 120
use via23_4  via23_4_614
timestamp 1696364841
transform 0 -1 28816 1 0 8095
box 1 40 161 120
use via23_4  via23_4_615
timestamp 1696364841
transform 0 -1 27516 1 0 8095
box 1 40 161 120
use via23_4  via23_4_616
timestamp 1696364841
transform 0 -1 31944 1 0 8095
box 1 40 161 120
use via23_4  via23_4_617
timestamp 1696364841
transform 0 -1 30644 1 0 8095
box 1 40 161 120
use via23_4  via23_4_618
timestamp 1696364841
transform 0 -1 29344 1 0 8095
box 1 40 161 120
use via23_4  via23_4_619
timestamp 1696364841
transform 0 -1 28044 1 0 8095
box 1 40 161 120
use via23_4  via23_4_620
timestamp 1696364841
transform 0 -1 40516 1 0 5575
box 1 40 161 120
use via23_4  via23_4_621
timestamp 1696364841
transform 0 -1 39216 1 0 5575
box 1 40 161 120
use via23_4  via23_4_622
timestamp 1696364841
transform 0 -1 42344 1 0 6415
box 1 40 161 120
use via23_4  via23_4_623
timestamp 1696364841
transform 0 -1 41044 1 0 6415
box 1 40 161 120
use via23_4  via23_4_624
timestamp 1696364841
transform 0 -1 43644 1 0 6415
box 1 40 161 120
use via23_4  via23_4_625
timestamp 1696364841
transform 0 -1 42344 1 0 5575
box 1 40 161 120
use via23_4  via23_4_626
timestamp 1696364841
transform 0 -1 41044 1 0 5575
box 1 40 161 120
use via23_4  via23_4_627
timestamp 1696364841
transform 0 -1 39744 1 0 5575
box 1 40 161 120
use via23_4  via23_4_628
timestamp 1696364841
transform 0 -1 38444 1 0 5575
box 1 40 161 120
use via23_4  via23_4_629
timestamp 1696364841
transform 0 -1 41044 1 0 4735
box 1 40 161 120
use via23_4  via23_4_630
timestamp 1696364841
transform 0 -1 38444 1 0 4735
box 1 40 161 120
use via23_4  via23_4_631
timestamp 1696364841
transform 0 -1 39744 1 0 4735
box 1 40 161 120
use via23_4  via23_4_632
timestamp 1696364841
transform 0 -1 43644 1 0 5575
box 1 40 161 120
use via23_4  via23_4_633
timestamp 1696364841
transform 0 -1 39744 1 0 6415
box 1 40 161 120
use via23_4  via23_4_634
timestamp 1696364841
transform 0 -1 38444 1 0 6415
box 1 40 161 120
use via23_4  via23_4_635
timestamp 1696364841
transform 0 -1 43116 1 0 6415
box 1 40 161 120
use via23_4  via23_4_636
timestamp 1696364841
transform 0 -1 43116 1 0 4735
box 1 40 161 120
use via23_4  via23_4_637
timestamp 1696364841
transform 0 -1 42344 1 0 4735
box 1 40 161 120
use via23_4  via23_4_638
timestamp 1696364841
transform 0 -1 41816 1 0 4735
box 1 40 161 120
use via23_4  via23_4_639
timestamp 1696364841
transform 0 -1 40516 1 0 4735
box 1 40 161 120
use via23_4  via23_4_640
timestamp 1696364841
transform 0 -1 39216 1 0 4735
box 1 40 161 120
use via23_4  via23_4_641
timestamp 1696364841
transform 0 -1 43644 1 0 4735
box 1 40 161 120
use via23_4  via23_4_642
timestamp 1696364841
transform 0 -1 43116 1 0 5575
box 1 40 161 120
use via23_4  via23_4_643
timestamp 1696364841
transform 0 -1 41816 1 0 6415
box 1 40 161 120
use via23_4  via23_4_644
timestamp 1696364841
transform 0 -1 40516 1 0 6415
box 1 40 161 120
use via23_4  via23_4_645
timestamp 1696364841
transform 0 -1 39216 1 0 6415
box 1 40 161 120
use via23_4  via23_4_646
timestamp 1696364841
transform 0 -1 41816 1 0 5575
box 1 40 161 120
use via23_4  via23_4_647
timestamp 1696364841
transform 0 -1 35844 1 0 5575
box 1 40 161 120
use via23_4  via23_4_648
timestamp 1696364841
transform 0 -1 34544 1 0 5575
box 1 40 161 120
use via23_4  via23_4_649
timestamp 1696364841
transform 0 -1 33244 1 0 5575
box 1 40 161 120
use via23_4  via23_4_650
timestamp 1696364841
transform 0 -1 37916 1 0 5575
box 1 40 161 120
use via23_4  via23_4_651
timestamp 1696364841
transform 0 -1 36616 1 0 5575
box 1 40 161 120
use via23_4  via23_4_652
timestamp 1696364841
transform 0 -1 35316 1 0 5575
box 1 40 161 120
use via23_4  via23_4_653
timestamp 1696364841
transform 0 -1 34016 1 0 5575
box 1 40 161 120
use via23_4  via23_4_654
timestamp 1696364841
transform 0 -1 34544 1 0 4735
box 1 40 161 120
use via23_4  via23_4_655
timestamp 1696364841
transform 0 -1 33244 1 0 4735
box 1 40 161 120
use via23_4  via23_4_656
timestamp 1696364841
transform 0 -1 35316 1 0 6415
box 1 40 161 120
use via23_4  via23_4_657
timestamp 1696364841
transform 0 -1 36616 1 0 4735
box 1 40 161 120
use via23_4  via23_4_658
timestamp 1696364841
transform 0 -1 35316 1 0 4735
box 1 40 161 120
use via23_4  via23_4_659
timestamp 1696364841
transform 0 -1 34016 1 0 4735
box 1 40 161 120
use via23_4  via23_4_660
timestamp 1696364841
transform 0 -1 37144 1 0 4735
box 1 40 161 120
use via23_4  via23_4_661
timestamp 1696364841
transform 0 -1 34016 1 0 6415
box 1 40 161 120
use via23_4  via23_4_662
timestamp 1696364841
transform 0 -1 37916 1 0 6415
box 1 40 161 120
use via23_4  via23_4_663
timestamp 1696364841
transform 0 -1 37144 1 0 6415
box 1 40 161 120
use via23_4  via23_4_664
timestamp 1696364841
transform 0 -1 37916 1 0 4735
box 1 40 161 120
use via23_4  via23_4_665
timestamp 1696364841
transform 0 -1 35844 1 0 6415
box 1 40 161 120
use via23_4  via23_4_666
timestamp 1696364841
transform 0 -1 34544 1 0 6415
box 1 40 161 120
use via23_4  via23_4_667
timestamp 1696364841
transform 0 -1 33244 1 0 6415
box 1 40 161 120
use via23_4  via23_4_668
timestamp 1696364841
transform 0 -1 36616 1 0 6415
box 1 40 161 120
use via23_4  via23_4_669
timestamp 1696364841
transform 0 -1 35844 1 0 4735
box 1 40 161 120
use via23_4  via23_4_670
timestamp 1696364841
transform 0 -1 37144 1 0 5575
box 1 40 161 120
use via23_4  via23_4_671
timestamp 1696364841
transform 0 -1 34016 1 0 8935
box 1 40 161 120
use via23_4  via23_4_672
timestamp 1696364841
transform 0 -1 35316 1 0 8935
box 1 40 161 120
use via23_4  via23_4_673
timestamp 1696364841
transform 0 -1 36616 1 0 8935
box 1 40 161 120
use via23_4  via23_4_674
timestamp 1696364841
transform 0 -1 37916 1 0 8935
box 1 40 161 120
use via23_4  via23_4_675
timestamp 1696364841
transform 0 -1 33244 1 0 8935
box 1 40 161 120
use via23_4  via23_4_676
timestamp 1696364841
transform 0 -1 34544 1 0 8935
box 1 40 161 120
use via23_4  via23_4_677
timestamp 1696364841
transform 0 -1 35844 1 0 8935
box 1 40 161 120
use via23_4  via23_4_678
timestamp 1696364841
transform 0 -1 37144 1 0 8935
box 1 40 161 120
use via23_4  via23_4_679
timestamp 1696364841
transform 0 -1 36616 1 0 8095
box 1 40 161 120
use via23_4  via23_4_680
timestamp 1696364841
transform 0 -1 37144 1 0 8095
box 1 40 161 120
use via23_4  via23_4_681
timestamp 1696364841
transform 0 -1 35844 1 0 8095
box 1 40 161 120
use via23_4  via23_4_682
timestamp 1696364841
transform 0 -1 37144 1 0 7255
box 1 40 161 120
use via23_4  via23_4_683
timestamp 1696364841
transform 0 -1 35844 1 0 7255
box 1 40 161 120
use via23_4  via23_4_684
timestamp 1696364841
transform 0 -1 34544 1 0 7255
box 1 40 161 120
use via23_4  via23_4_685
timestamp 1696364841
transform 0 -1 33244 1 0 7255
box 1 40 161 120
use via23_4  via23_4_686
timestamp 1696364841
transform 0 -1 37916 1 0 7255
box 1 40 161 120
use via23_4  via23_4_687
timestamp 1696364841
transform 0 -1 36616 1 0 7255
box 1 40 161 120
use via23_4  via23_4_688
timestamp 1696364841
transform 0 -1 35316 1 0 7255
box 1 40 161 120
use via23_4  via23_4_689
timestamp 1696364841
transform 0 -1 34016 1 0 7255
box 1 40 161 120
use via23_4  via23_4_690
timestamp 1696364841
transform 0 -1 34544 1 0 8095
box 1 40 161 120
use via23_4  via23_4_691
timestamp 1696364841
transform 0 -1 33244 1 0 8095
box 1 40 161 120
use via23_4  via23_4_692
timestamp 1696364841
transform 0 -1 35316 1 0 8095
box 1 40 161 120
use via23_4  via23_4_693
timestamp 1696364841
transform 0 -1 37916 1 0 8095
box 1 40 161 120
use via23_4  via23_4_694
timestamp 1696364841
transform 0 -1 34016 1 0 8095
box 1 40 161 120
use via23_4  via23_4_695
timestamp 1696364841
transform 0 -1 43644 1 0 7255
box 1 40 161 120
use via23_4  via23_4_696
timestamp 1696364841
transform 0 -1 39744 1 0 8095
box 1 40 161 120
use via23_4  via23_4_697
timestamp 1696364841
transform 0 -1 38444 1 0 8095
box 1 40 161 120
use via23_4  via23_4_698
timestamp 1696364841
transform 0 -1 39216 1 0 8095
box 1 40 161 120
use via23_4  via23_4_699
timestamp 1696364841
transform 0 -1 41816 1 0 8095
box 1 40 161 120
use via23_4  via23_4_700
timestamp 1696364841
transform 0 -1 40516 1 0 8095
box 1 40 161 120
use via23_4  via23_4_701
timestamp 1696364841
transform 0 -1 43644 1 0 8935
box 1 40 161 120
use via23_4  via23_4_702
timestamp 1696364841
transform 0 -1 43116 1 0 8935
box 1 40 161 120
use via23_4  via23_4_703
timestamp 1696364841
transform 0 -1 43644 1 0 8095
box 1 40 161 120
use via23_4  via23_4_704
timestamp 1696364841
transform 0 -1 43116 1 0 8095
box 1 40 161 120
use via23_4  via23_4_705
timestamp 1696364841
transform 0 -1 43116 1 0 7255
box 1 40 161 120
use via23_4  via23_4_706
timestamp 1696364841
transform 0 -1 39216 1 0 8935
box 1 40 161 120
use via23_4  via23_4_707
timestamp 1696364841
transform 0 -1 40516 1 0 8935
box 1 40 161 120
use via23_4  via23_4_708
timestamp 1696364841
transform 0 -1 41816 1 0 8935
box 1 40 161 120
use via23_4  via23_4_709
timestamp 1696364841
transform 0 -1 38444 1 0 8935
box 1 40 161 120
use via23_4  via23_4_710
timestamp 1696364841
transform 0 -1 39744 1 0 8935
box 1 40 161 120
use via23_4  via23_4_711
timestamp 1696364841
transform 0 -1 41044 1 0 8935
box 1 40 161 120
use via23_4  via23_4_712
timestamp 1696364841
transform 0 -1 42344 1 0 8935
box 1 40 161 120
use via23_4  via23_4_713
timestamp 1696364841
transform 0 -1 42344 1 0 7255
box 1 40 161 120
use via23_4  via23_4_714
timestamp 1696364841
transform 0 -1 41044 1 0 7255
box 1 40 161 120
use via23_4  via23_4_715
timestamp 1696364841
transform 0 -1 39744 1 0 7255
box 1 40 161 120
use via23_4  via23_4_716
timestamp 1696364841
transform 0 -1 38444 1 0 7255
box 1 40 161 120
use via23_4  via23_4_717
timestamp 1696364841
transform 0 -1 41816 1 0 7255
box 1 40 161 120
use via23_4  via23_4_718
timestamp 1696364841
transform 0 -1 40516 1 0 7255
box 1 40 161 120
use via23_4  via23_4_719
timestamp 1696364841
transform 0 -1 39216 1 0 7255
box 1 40 161 120
use via23_4  via23_4_720
timestamp 1696364841
transform 0 -1 42344 1 0 8095
box 1 40 161 120
use via23_4  via23_4_721
timestamp 1696364841
transform 0 -1 41044 1 0 8095
box 1 40 161 120
use via23_4  via23_4_722
timestamp 1696364841
transform -1 0 21901 0 -1 -36
box 1 40 161 120
use via_M1_M2$1  via_M1_M2$1_0
timestamp 1696364841
transform 0 1 20896 -1 0 4046
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_1
timestamp 1696364841
transform 0 1 20570 -1 0 4046
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_2
timestamp 1696364841
transform 0 1 20896 -1 0 6566
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_3
timestamp 1696364841
transform 0 1 20570 -1 0 6566
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_4
timestamp 1696364841
transform 0 1 21750 -1 0 5726
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_5
timestamp 1696364841
transform 0 1 21424 -1 0 5726
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_6
timestamp 1696364841
transform 0 1 23050 -1 0 4046
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_7
timestamp 1696364841
transform 0 1 22724 -1 0 4046
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_8
timestamp 1696364841
transform 0 1 23050 -1 0 6566
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_9
timestamp 1696364841
transform 0 1 22724 -1 0 6566
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_10
timestamp 1696364841
transform 0 1 21870 -1 0 4886
box 0 0 140 80
use via_M1_M2$1  via_M1_M2$1_11
timestamp 1696364841
transform 0 1 22196 -1 0 4886
box 0 0 140 80
<< labels >>
flabel comment s 21650 5655 21650 5655 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel comment s 22096 4815 22096 4815 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel comment s 20796 6495 20796 6495 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel comment s 20796 3975 20796 3975 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel comment s 22950 6495 22950 6495 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel comment s 22950 3975 22950 3975 1 FreeSans 100 0 0 0 Replace with M3-M3 connection. DRC/PDK related
flabel metal2 s 28100 324 28200 374 2 FreeSans 44 0 0 0 n5
port 2 nsew
flabel metal2 s 25499 5 25599 54 2 FreeSans 44 0 0 0 n7
port 3 nsew
flabel metal2 s 16800 164 16900 214 2 FreeSans 44 0 0 0 n6
port 4 nsew
flabel metal3 s 0 804 40 884 1 FreeSans 96 0 0 0 n2
port 6 nsew
flabel metal3 s 0 644 40 724 1 FreeSans 96 0 0 0 n3
port 7 nsew
flabel metal3 s 0 484 40 564 1 FreeSans 96 0 0 0 n4
port 8 nsew
flabel metal3 s 0 324 40 404 1 FreeSans 96 0 0 0 n5
port 2 nsew
flabel metal3 s 0 164 40 244 1 FreeSans 96 0 0 0 n6
port 4 nsew
flabel metal3 s 0 4 40 84 1 FreeSans 96 0 0 0 n7
port 3 nsew
flabel metal3 s 0 -156 40 -76 1 FreeSans 96 0 0 0 n1
port 9 nsew
flabel metal3 s 0 -316 40 -236 1 FreeSans 96 0 0 0 n0
port 10 nsew
flabel metal3 s 0 -476 40 -396 1 FreeSans 96 0 0 0 ndum
port 11 nsew
flabel metal4 s 43650 9416 43700 9516 2 FreeSans 96 0 0 0 top
port 12 nsew
<< properties >>
string FIXED_BBOX 0 -476 43700 9516
string path 10.050 236.650 1091.250 236.650 
<< end >>
