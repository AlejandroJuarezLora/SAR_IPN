magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 590 542
<< pwell >>
rect 269 123 545 163
rect 4 -13 545 123
rect 29 -57 63 -13
rect 269 -19 545 -13
<< scnmos >>
rect 82 13 112 97
rect 166 13 196 97
rect 250 13 280 97
rect 348 7 378 137
rect 432 7 462 137
<< scpmoshvt >>
rect 82 257 112 341
rect 154 257 184 341
rect 250 257 280 341
rect 348 257 378 457
rect 432 257 462 457
<< ndiff >>
rect 295 97 348 137
rect 30 71 82 97
rect 30 37 38 71
rect 72 37 82 71
rect 30 13 82 37
rect 112 57 166 97
rect 112 23 122 57
rect 156 23 166 57
rect 112 13 166 23
rect 196 71 250 97
rect 196 37 206 71
rect 240 37 250 71
rect 196 13 250 37
rect 280 57 348 97
rect 280 23 300 57
rect 334 23 348 57
rect 280 13 348 23
rect 295 7 348 13
rect 378 95 432 137
rect 378 61 388 95
rect 422 61 432 95
rect 378 7 432 61
rect 462 125 519 137
rect 462 91 477 125
rect 511 91 519 125
rect 462 57 519 91
rect 462 23 477 57
rect 511 23 519 57
rect 462 7 519 23
<< pdiff >>
rect 295 445 348 457
rect 295 411 303 445
rect 337 411 348 445
rect 295 377 348 411
rect 295 343 303 377
rect 337 343 348 377
rect 295 341 348 343
rect 30 314 82 341
rect 30 280 38 314
rect 72 280 82 314
rect 30 257 82 280
rect 112 257 154 341
rect 184 257 250 341
rect 280 257 348 341
rect 378 414 432 457
rect 378 380 388 414
rect 422 380 432 414
rect 378 346 432 380
rect 378 312 388 346
rect 422 312 432 346
rect 378 257 432 312
rect 462 437 525 457
rect 462 403 477 437
rect 511 403 525 437
rect 462 369 525 403
rect 462 335 477 369
rect 511 335 525 369
rect 462 301 525 335
rect 462 267 477 301
rect 511 267 525 301
rect 462 257 525 267
<< ndiffc >>
rect 38 37 72 71
rect 122 23 156 57
rect 206 37 240 71
rect 300 23 334 57
rect 388 61 422 95
rect 477 91 511 125
rect 477 23 511 57
<< pdiffc >>
rect 303 411 337 445
rect 303 343 337 377
rect 38 280 72 314
rect 388 380 422 414
rect 388 312 422 346
rect 477 403 511 437
rect 477 335 511 369
rect 477 267 511 301
<< poly >>
rect 348 457 378 483
rect 432 457 462 483
rect 148 433 214 443
rect 148 399 164 433
rect 198 399 214 433
rect 148 389 214 399
rect 82 341 112 367
rect 154 341 184 389
rect 250 341 280 367
rect 82 225 112 257
rect 24 209 112 225
rect 24 175 34 209
rect 68 175 112 209
rect 24 159 112 175
rect 82 97 112 159
rect 154 142 184 257
rect 250 225 280 257
rect 348 225 378 257
rect 432 225 462 257
rect 235 209 289 225
rect 235 175 245 209
rect 279 175 289 209
rect 235 159 289 175
rect 331 209 462 225
rect 331 175 341 209
rect 375 175 462 209
rect 331 159 462 175
rect 154 112 196 142
rect 166 97 196 112
rect 250 97 280 159
rect 348 137 378 159
rect 432 137 462 159
rect 82 -13 112 13
rect 166 -13 196 13
rect 250 -13 280 13
rect 348 -19 378 7
rect 432 -19 462 7
<< polycont >>
rect 164 399 198 433
rect 34 175 68 209
rect 245 175 279 209
rect 341 175 375 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 290 445 346 487
rect 17 433 256 443
rect 17 399 164 433
rect 198 399 256 433
rect 17 385 256 399
rect 290 411 303 445
rect 337 411 346 445
rect 290 377 346 411
rect 21 317 254 351
rect 290 343 303 377
rect 337 343 346 377
rect 290 327 346 343
rect 388 414 443 453
rect 422 380 443 414
rect 388 346 443 380
rect 21 314 87 317
rect 21 280 38 314
rect 72 280 87 314
rect 220 293 254 317
rect 422 312 443 346
rect 21 259 87 280
rect 121 225 166 283
rect 220 259 354 293
rect 388 259 443 312
rect 320 225 354 259
rect 17 209 87 225
rect 17 175 34 209
rect 68 175 87 209
rect 17 159 87 175
rect 121 209 286 225
rect 121 175 245 209
rect 279 175 286 209
rect 121 159 286 175
rect 320 209 375 225
rect 320 175 341 209
rect 320 159 375 175
rect 320 125 354 159
rect 21 91 354 125
rect 409 112 443 259
rect 477 437 535 487
rect 511 403 535 437
rect 477 369 535 403
rect 511 335 535 369
rect 477 301 535 335
rect 511 267 535 301
rect 477 246 535 267
rect 388 95 443 112
rect 21 71 72 91
rect 21 37 38 71
rect 206 71 240 91
rect 21 21 72 37
rect 106 23 122 57
rect 156 23 172 57
rect 106 -23 172 23
rect 422 61 443 95
rect 206 21 240 37
rect 274 23 300 57
rect 334 23 350 57
rect 388 43 443 61
rect 477 125 535 143
rect 511 91 535 125
rect 477 57 535 91
rect 274 -23 350 23
rect 511 23 535 57
rect 477 -23 535 23
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
<< metal1 >>
rect 0 521 552 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 0 456 552 487
rect 0 -23 552 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
rect 0 -88 552 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or3_2
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 121 181 155 215 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 213 181 247 215 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 29 385 63 419 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 397 317 431 351 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 121 249 155 283 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 121 385 155 419 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 29 181 63 215 0 FreeSans 400 0 0 0 C
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 552 504
string path 0.000 -1.000 13.800 -1.000 
<< end >>
