magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1878 542
<< pwell >>
rect 1 -19 1822 117
rect 29 -57 63 -19
<< scnmos >>
rect 80 7 110 91
rect 166 7 196 91
rect 252 7 282 91
rect 338 7 368 91
rect 424 7 454 91
rect 510 7 540 91
rect 596 7 626 91
rect 682 7 712 91
rect 768 7 798 91
rect 854 7 884 91
rect 940 7 970 91
rect 1026 7 1056 91
rect 1111 7 1141 91
rect 1197 7 1227 91
rect 1283 7 1313 91
rect 1369 7 1399 91
rect 1455 7 1485 91
rect 1541 7 1571 91
rect 1627 7 1657 91
rect 1713 7 1743 91
<< scpmoshvt >>
rect 80 257 110 457
rect 166 257 196 457
rect 252 257 282 457
rect 338 257 368 457
rect 424 257 454 457
rect 510 257 540 457
rect 596 257 626 457
rect 682 257 712 457
rect 768 257 798 457
rect 854 257 884 457
rect 940 257 970 457
rect 1026 257 1056 457
rect 1111 257 1141 457
rect 1197 257 1227 457
rect 1283 257 1313 457
rect 1369 257 1399 457
rect 1455 257 1485 457
rect 1541 257 1571 457
rect 1627 257 1657 457
rect 1713 257 1743 457
<< ndiff >>
rect 27 53 80 91
rect 27 19 35 53
rect 69 19 80 53
rect 27 7 80 19
rect 110 66 166 91
rect 110 32 121 66
rect 155 32 166 66
rect 110 7 166 32
rect 196 66 252 91
rect 196 32 207 66
rect 241 32 252 66
rect 196 7 252 32
rect 282 66 338 91
rect 282 32 293 66
rect 327 32 338 66
rect 282 7 338 32
rect 368 66 424 91
rect 368 32 379 66
rect 413 32 424 66
rect 368 7 424 32
rect 454 66 510 91
rect 454 32 465 66
rect 499 32 510 66
rect 454 7 510 32
rect 540 57 596 91
rect 540 23 551 57
rect 585 23 596 57
rect 540 7 596 23
rect 626 66 682 91
rect 626 32 637 66
rect 671 32 682 66
rect 626 7 682 32
rect 712 57 768 91
rect 712 23 723 57
rect 757 23 768 57
rect 712 7 768 23
rect 798 66 854 91
rect 798 32 809 66
rect 843 32 854 66
rect 798 7 854 32
rect 884 57 940 91
rect 884 23 895 57
rect 929 23 940 57
rect 884 7 940 23
rect 970 66 1026 91
rect 970 32 981 66
rect 1015 32 1026 66
rect 970 7 1026 32
rect 1056 57 1111 91
rect 1056 23 1067 57
rect 1101 23 1111 57
rect 1056 7 1111 23
rect 1141 66 1197 91
rect 1141 32 1152 66
rect 1186 32 1197 66
rect 1141 7 1197 32
rect 1227 57 1283 91
rect 1227 23 1238 57
rect 1272 23 1283 57
rect 1227 7 1283 23
rect 1313 66 1369 91
rect 1313 32 1324 66
rect 1358 32 1369 66
rect 1313 7 1369 32
rect 1399 57 1455 91
rect 1399 23 1410 57
rect 1444 23 1455 57
rect 1399 7 1455 23
rect 1485 66 1541 91
rect 1485 32 1496 66
rect 1530 32 1541 66
rect 1485 7 1541 32
rect 1571 57 1627 91
rect 1571 23 1582 57
rect 1616 23 1627 57
rect 1571 7 1627 23
rect 1657 66 1713 91
rect 1657 32 1668 66
rect 1702 32 1713 66
rect 1657 7 1713 32
rect 1743 57 1796 91
rect 1743 23 1754 57
rect 1788 23 1796 57
rect 1743 7 1796 23
<< pdiff >>
rect 27 445 80 457
rect 27 411 35 445
rect 69 411 80 445
rect 27 377 80 411
rect 27 343 35 377
rect 69 343 80 377
rect 27 257 80 343
rect 110 437 166 457
rect 110 403 121 437
rect 155 403 166 437
rect 110 369 166 403
rect 110 335 121 369
rect 155 335 166 369
rect 110 257 166 335
rect 196 445 252 457
rect 196 411 207 445
rect 241 411 252 445
rect 196 377 252 411
rect 196 343 207 377
rect 241 343 252 377
rect 196 257 252 343
rect 282 429 338 457
rect 282 395 293 429
rect 327 395 338 429
rect 282 361 338 395
rect 282 327 293 361
rect 327 327 338 361
rect 282 257 338 327
rect 368 445 424 457
rect 368 411 379 445
rect 413 411 424 445
rect 368 377 424 411
rect 368 343 379 377
rect 413 343 424 377
rect 368 257 424 343
rect 454 401 510 457
rect 454 367 465 401
rect 499 367 510 401
rect 454 315 510 367
rect 454 281 465 315
rect 499 281 510 315
rect 454 257 510 281
rect 540 421 596 457
rect 540 387 551 421
rect 585 387 596 421
rect 540 257 596 387
rect 626 401 682 457
rect 626 367 637 401
rect 671 367 682 401
rect 626 315 682 367
rect 626 281 637 315
rect 671 281 682 315
rect 626 257 682 281
rect 712 421 768 457
rect 712 387 723 421
rect 757 387 768 421
rect 712 257 768 387
rect 798 401 854 457
rect 798 367 809 401
rect 843 367 854 401
rect 798 315 854 367
rect 798 281 809 315
rect 843 281 854 315
rect 798 257 854 281
rect 884 421 940 457
rect 884 387 895 421
rect 929 387 940 421
rect 884 257 940 387
rect 970 401 1026 457
rect 970 367 981 401
rect 1015 367 1026 401
rect 970 315 1026 367
rect 970 281 981 315
rect 1015 281 1026 315
rect 970 257 1026 281
rect 1056 421 1111 457
rect 1056 387 1067 421
rect 1101 387 1111 421
rect 1056 257 1111 387
rect 1141 401 1197 457
rect 1141 367 1152 401
rect 1186 367 1197 401
rect 1141 315 1197 367
rect 1141 281 1152 315
rect 1186 281 1197 315
rect 1141 257 1197 281
rect 1227 421 1283 457
rect 1227 387 1238 421
rect 1272 387 1283 421
rect 1227 257 1283 387
rect 1313 401 1369 457
rect 1313 367 1324 401
rect 1358 367 1369 401
rect 1313 315 1369 367
rect 1313 281 1324 315
rect 1358 281 1369 315
rect 1313 257 1369 281
rect 1399 421 1455 457
rect 1399 387 1410 421
rect 1444 387 1455 421
rect 1399 257 1455 387
rect 1485 401 1541 457
rect 1485 367 1496 401
rect 1530 367 1541 401
rect 1485 315 1541 367
rect 1485 281 1496 315
rect 1530 281 1541 315
rect 1485 257 1541 281
rect 1571 421 1627 457
rect 1571 387 1582 421
rect 1616 387 1627 421
rect 1571 257 1627 387
rect 1657 401 1713 457
rect 1657 367 1668 401
rect 1702 367 1713 401
rect 1657 315 1713 367
rect 1657 281 1668 315
rect 1702 281 1713 315
rect 1657 257 1713 281
rect 1743 421 1796 457
rect 1743 387 1754 421
rect 1788 387 1796 421
rect 1743 257 1796 387
<< ndiffc >>
rect 35 19 69 53
rect 121 32 155 66
rect 207 32 241 66
rect 293 32 327 66
rect 379 32 413 66
rect 465 32 499 66
rect 551 23 585 57
rect 637 32 671 66
rect 723 23 757 57
rect 809 32 843 66
rect 895 23 929 57
rect 981 32 1015 66
rect 1067 23 1101 57
rect 1152 32 1186 66
rect 1238 23 1272 57
rect 1324 32 1358 66
rect 1410 23 1444 57
rect 1496 32 1530 66
rect 1582 23 1616 57
rect 1668 32 1702 66
rect 1754 23 1788 57
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 121 403 155 437
rect 121 335 155 369
rect 207 411 241 445
rect 207 343 241 377
rect 293 395 327 429
rect 293 327 327 361
rect 379 411 413 445
rect 379 343 413 377
rect 465 367 499 401
rect 465 281 499 315
rect 551 387 585 421
rect 637 367 671 401
rect 637 281 671 315
rect 723 387 757 421
rect 809 367 843 401
rect 809 281 843 315
rect 895 387 929 421
rect 981 367 1015 401
rect 981 281 1015 315
rect 1067 387 1101 421
rect 1152 367 1186 401
rect 1152 281 1186 315
rect 1238 387 1272 421
rect 1324 367 1358 401
rect 1324 281 1358 315
rect 1410 387 1444 421
rect 1496 367 1530 401
rect 1496 281 1530 315
rect 1582 387 1616 421
rect 1668 367 1702 401
rect 1668 281 1702 315
rect 1754 387 1788 421
<< poly >>
rect 80 457 110 483
rect 166 457 196 483
rect 252 457 282 483
rect 338 457 368 483
rect 424 457 454 483
rect 510 457 540 483
rect 596 457 626 483
rect 682 457 712 483
rect 768 457 798 483
rect 854 457 884 483
rect 940 457 970 483
rect 1026 457 1056 483
rect 1111 457 1141 483
rect 1197 457 1227 483
rect 1283 457 1313 483
rect 1369 457 1399 483
rect 1455 457 1485 483
rect 1541 457 1571 483
rect 1627 457 1657 483
rect 1713 457 1743 483
rect 80 242 110 257
rect 166 242 196 257
rect 252 242 282 257
rect 338 242 368 257
rect 21 209 368 242
rect 21 175 37 209
rect 71 175 368 209
rect 21 140 368 175
rect 80 91 110 140
rect 166 91 196 140
rect 252 91 282 140
rect 338 91 368 140
rect 424 225 454 257
rect 510 225 540 257
rect 596 225 626 257
rect 682 225 712 257
rect 768 225 798 257
rect 854 225 884 257
rect 940 225 970 257
rect 1026 225 1056 257
rect 1111 225 1141 257
rect 1197 225 1227 257
rect 1283 225 1313 257
rect 1369 225 1399 257
rect 1455 225 1485 257
rect 1541 225 1571 257
rect 1627 225 1657 257
rect 1713 225 1743 257
rect 424 209 1743 225
rect 424 175 464 209
rect 498 175 532 209
rect 566 175 600 209
rect 634 175 668 209
rect 702 175 736 209
rect 770 175 804 209
rect 838 175 872 209
rect 906 175 940 209
rect 974 175 1008 209
rect 1042 175 1076 209
rect 1110 175 1144 209
rect 1178 175 1212 209
rect 1246 175 1280 209
rect 1314 175 1348 209
rect 1382 175 1416 209
rect 1450 175 1484 209
rect 1518 175 1743 209
rect 424 150 1743 175
rect 424 91 454 150
rect 510 91 540 150
rect 596 91 626 150
rect 682 91 712 150
rect 768 91 798 150
rect 854 91 884 150
rect 940 91 970 150
rect 1026 91 1056 150
rect 1111 91 1141 150
rect 1197 91 1227 150
rect 1283 91 1313 150
rect 1369 91 1399 150
rect 1455 91 1485 150
rect 1541 91 1571 150
rect 1627 91 1657 150
rect 1713 91 1743 150
rect 80 -19 110 7
rect 166 -19 196 7
rect 252 -19 282 7
rect 338 -19 368 7
rect 424 -19 454 7
rect 510 -19 540 7
rect 596 -19 626 7
rect 682 -19 712 7
rect 768 -19 798 7
rect 854 -19 884 7
rect 940 -19 970 7
rect 1026 -19 1056 7
rect 1111 -19 1141 7
rect 1197 -19 1227 7
rect 1283 -19 1313 7
rect 1369 -19 1399 7
rect 1455 -19 1485 7
rect 1541 -19 1571 7
rect 1627 -19 1657 7
rect 1713 -19 1743 7
<< polycont >>
rect 37 175 71 209
rect 464 175 498 209
rect 532 175 566 209
rect 600 175 634 209
rect 668 175 702 209
rect 736 175 770 209
rect 804 175 838 209
rect 872 175 906 209
rect 940 175 974 209
rect 1008 175 1042 209
rect 1076 175 1110 209
rect 1144 175 1178 209
rect 1212 175 1246 209
rect 1280 175 1314 209
rect 1348 175 1382 209
rect 1416 175 1450 209
rect 1484 175 1518 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1840 521
rect 19 445 78 487
rect 19 411 35 445
rect 69 411 78 445
rect 19 377 78 411
rect 19 343 35 377
rect 69 343 78 377
rect 19 325 78 343
rect 114 437 163 453
rect 114 403 121 437
rect 155 403 163 437
rect 114 369 163 403
rect 114 335 121 369
rect 155 335 163 369
rect 114 225 163 335
rect 198 445 250 487
rect 370 486 1625 487
rect 198 411 207 445
rect 241 411 250 445
rect 198 377 250 411
rect 198 343 207 377
rect 241 343 250 377
rect 198 325 250 343
rect 286 429 336 452
rect 286 395 293 429
rect 327 395 336 429
rect 286 361 336 395
rect 286 327 293 361
rect 327 327 336 361
rect 370 445 422 486
rect 370 411 379 445
rect 413 411 422 445
rect 370 377 422 411
rect 370 343 379 377
rect 413 343 422 377
rect 370 327 422 343
rect 456 401 508 452
rect 456 367 465 401
rect 499 367 508 401
rect 286 225 336 327
rect 456 315 508 367
rect 542 421 594 486
rect 542 387 551 421
rect 585 387 594 421
rect 542 341 594 387
rect 628 401 680 452
rect 628 367 637 401
rect 671 367 680 401
rect 456 281 465 315
rect 499 307 508 315
rect 628 315 680 367
rect 714 421 766 486
rect 714 387 723 421
rect 757 387 766 421
rect 714 341 766 387
rect 800 401 852 452
rect 800 367 809 401
rect 843 367 852 401
rect 628 307 637 315
rect 499 281 637 307
rect 671 307 680 315
rect 800 315 852 367
rect 886 421 938 486
rect 886 387 895 421
rect 929 387 938 421
rect 886 341 938 387
rect 972 401 1024 452
rect 972 367 981 401
rect 1015 367 1024 401
rect 800 307 809 315
rect 671 281 809 307
rect 843 307 852 315
rect 972 315 1024 367
rect 1058 421 1107 486
rect 1058 387 1067 421
rect 1101 387 1107 421
rect 1058 341 1107 387
rect 1141 401 1193 452
rect 1141 367 1152 401
rect 1186 367 1193 401
rect 972 307 981 315
rect 843 281 981 307
rect 1015 307 1024 315
rect 1141 315 1193 367
rect 1230 421 1279 486
rect 1230 387 1238 421
rect 1272 387 1279 421
rect 1230 341 1279 387
rect 1313 401 1365 452
rect 1313 367 1324 401
rect 1358 367 1365 401
rect 1141 307 1152 315
rect 1015 281 1152 307
rect 1186 307 1193 315
rect 1313 315 1365 367
rect 1402 421 1451 486
rect 1402 387 1410 421
rect 1444 387 1451 421
rect 1402 341 1451 387
rect 1485 401 1537 452
rect 1485 367 1496 401
rect 1530 367 1537 401
rect 1313 307 1324 315
rect 1186 281 1324 307
rect 1358 307 1365 315
rect 1485 315 1537 367
rect 1574 421 1625 486
rect 1574 387 1582 421
rect 1616 387 1625 421
rect 1574 341 1625 387
rect 1659 401 1717 452
rect 1659 367 1668 401
rect 1702 367 1717 401
rect 1485 307 1496 315
rect 1358 281 1496 307
rect 1530 304 1537 315
rect 1659 315 1717 367
rect 1751 421 1805 487
rect 1751 387 1754 421
rect 1788 387 1805 421
rect 1751 338 1805 387
rect 1659 304 1668 315
rect 1530 281 1668 304
rect 1702 304 1717 315
rect 1702 281 1805 304
rect 456 259 1805 281
rect 17 209 80 225
rect 17 175 37 209
rect 71 175 80 209
rect 17 113 80 175
rect 114 209 1538 225
rect 114 175 464 209
rect 498 175 532 209
rect 566 175 600 209
rect 634 175 668 209
rect 702 175 736 209
rect 770 175 804 209
rect 838 175 872 209
rect 906 175 940 209
rect 974 175 1008 209
rect 1042 175 1076 209
rect 1110 175 1144 209
rect 1178 175 1212 209
rect 1246 175 1280 209
rect 1314 175 1348 209
rect 1382 175 1416 209
rect 1450 175 1484 209
rect 1518 175 1538 209
rect 17 53 78 79
rect 17 19 35 53
rect 69 19 78 53
rect 17 -23 78 19
rect 114 66 164 175
rect 114 32 121 66
rect 155 32 164 66
rect 114 13 164 32
rect 198 66 250 82
rect 198 32 207 66
rect 241 32 250 66
rect 198 -23 250 32
rect 286 66 336 175
rect 1572 141 1805 259
rect 456 107 1805 141
rect 286 32 293 66
rect 327 32 336 66
rect 286 13 336 32
rect 370 66 422 89
rect 370 32 379 66
rect 413 32 422 66
rect 370 -23 422 32
rect 456 66 508 107
rect 456 32 465 66
rect 499 32 508 66
rect 456 16 508 32
rect 542 57 594 73
rect 542 23 551 57
rect 585 23 594 57
rect 542 -23 594 23
rect 628 66 680 107
rect 628 32 637 66
rect 671 32 680 66
rect 628 16 680 32
rect 714 57 766 73
rect 714 23 723 57
rect 757 23 766 57
rect 714 -23 766 23
rect 800 66 852 107
rect 800 32 809 66
rect 843 32 852 66
rect 800 16 852 32
rect 886 57 935 73
rect 886 23 895 57
rect 929 23 935 57
rect 886 -23 935 23
rect 969 66 1024 107
rect 969 32 981 66
rect 1015 32 1024 66
rect 969 16 1024 32
rect 1058 57 1107 73
rect 1058 23 1067 57
rect 1101 23 1107 57
rect 1058 -23 1107 23
rect 1141 66 1193 107
rect 1141 32 1152 66
rect 1186 32 1193 66
rect 1141 16 1193 32
rect 1229 57 1279 73
rect 1229 23 1238 57
rect 1272 23 1279 57
rect 1229 -23 1279 23
rect 1313 66 1365 107
rect 1313 32 1324 66
rect 1358 32 1365 66
rect 1313 16 1365 32
rect 1401 57 1451 73
rect 1401 23 1410 57
rect 1444 23 1451 57
rect 1401 -23 1451 23
rect 1485 66 1537 107
rect 1485 32 1496 66
rect 1530 32 1537 66
rect 1485 16 1537 32
rect 1573 57 1625 73
rect 1573 23 1582 57
rect 1616 23 1625 57
rect 1573 -23 1625 23
rect 1659 66 1711 107
rect 1659 32 1668 66
rect 1702 32 1711 66
rect 1659 16 1711 32
rect 1745 57 1805 73
rect 1745 23 1754 57
rect 1788 23 1805 57
rect 1745 -23 1805 23
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1840 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 1133 487 1167 521
rect 1225 487 1259 521
rect 1317 487 1351 521
rect 1409 487 1443 521
rect 1501 487 1535 521
rect 1593 487 1627 521
rect 1685 487 1719 521
rect 1777 487 1811 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
rect 1133 -57 1167 -23
rect 1225 -57 1259 -23
rect 1317 -57 1351 -23
rect 1409 -57 1443 -23
rect 1501 -57 1535 -23
rect 1593 -57 1627 -23
rect 1685 -57 1719 -23
rect 1777 -57 1811 -23
<< metal1 >>
rect 0 521 1840 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1840 521
rect 0 456 1840 487
rect 0 -23 1840 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1840 -23
rect 0 -88 1840 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 clkbuf_16
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel nwell s 46 504 46 504 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel pwell s 46 -40 46 -40 0 FreeSans 200 0 0 0 VNB
flabel locali s 1593 249 1627 283 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 1685 249 1719 283 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 1685 181 1719 215 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 1593 181 1627 215 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 1593 113 1627 147 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 1685 113 1719 147 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 29 113 63 147 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel locali s 29 181 63 215 0 FreeSans 200 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 1840 504
<< end >>
