magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< locali >>
rect 3893 10483 3927 10653
<< viali >>
rect 4905 12897 4939 12931
rect 12909 12897 12943 12931
rect 15025 12897 15059 12931
rect 949 12829 983 12863
rect 3249 12829 3283 12863
rect 3985 12829 4019 12863
rect 6929 12829 6963 12863
rect 9597 12829 9631 12863
rect 11253 12829 11287 12863
rect 14381 12829 14415 12863
rect 1133 12761 1167 12795
rect 1869 12761 1903 12795
rect 3433 12761 3467 12795
rect 4169 12761 4203 12795
rect 4813 12761 4847 12795
rect 5917 12761 5951 12795
rect 7113 12761 7147 12795
rect 8769 12761 8803 12795
rect 8953 12761 8987 12795
rect 9781 12761 9815 12795
rect 11437 12761 11471 12795
rect 12817 12761 12851 12795
rect 14197 12761 14231 12795
rect 14933 12761 14967 12795
rect 6101 12625 6135 12659
rect 1777 12557 1811 12591
rect 9137 12557 9171 12591
rect 9689 12353 9723 12387
rect 2329 12217 2363 12251
rect 6745 12217 6779 12251
rect 11437 12217 11471 12251
rect 581 12149 615 12183
rect 4353 12149 4387 12183
rect 4537 12149 4571 12183
rect 7205 12149 7239 12183
rect 8677 12149 8711 12183
rect 8769 12149 8803 12183
rect 8861 12149 8895 12183
rect 9137 12149 9171 12183
rect 857 12081 891 12115
rect 3525 12081 3559 12115
rect 3709 12081 3743 12115
rect 3893 12081 3927 12115
rect 6469 12081 6503 12115
rect 8979 12081 9013 12115
rect 11161 12081 11195 12115
rect 14933 12081 14967 12115
rect 15117 12081 15151 12115
rect 4445 12013 4479 12047
rect 4997 12013 5031 12047
rect 7297 12013 7331 12047
rect 8493 12013 8527 12047
rect 3525 11809 3559 11843
rect 4905 11809 4939 11843
rect 7941 11809 7975 11843
rect 10149 11809 10183 11843
rect 11161 11809 11195 11843
rect 14381 11809 14415 11843
rect 949 11741 983 11775
rect 2053 11741 2087 11775
rect 4537 11741 4571 11775
rect 8677 11741 8711 11775
rect 1777 11673 1811 11707
rect 4721 11673 4755 11707
rect 6193 11673 6227 11707
rect 11069 11673 11103 11707
rect 11253 11673 11287 11707
rect 14289 11673 14323 11707
rect 6469 11605 6503 11639
rect 8401 11605 8435 11639
rect 765 11537 799 11571
rect 2053 11265 2087 11299
rect 6929 11265 6963 11299
rect 8493 11265 8527 11299
rect 14289 11265 14323 11299
rect 3249 11197 3283 11231
rect 3985 11197 4019 11231
rect 4721 11129 4755 11163
rect 9873 11129 9907 11163
rect 949 11061 983 11095
rect 1869 11061 1903 11095
rect 2053 11061 2087 11095
rect 3249 11061 3283 11095
rect 3525 11061 3559 11095
rect 3985 11061 4019 11095
rect 4169 11061 4203 11095
rect 4261 11061 4295 11095
rect 6469 11061 6503 11095
rect 7114 11061 7148 11095
rect 7205 11061 7239 11095
rect 7573 11061 7607 11095
rect 8677 11061 8711 11095
rect 8861 11061 8895 11095
rect 8979 11061 9013 11095
rect 9137 11061 9171 11095
rect 14197 11061 14231 11095
rect 765 10993 799 11027
rect 3433 10993 3467 11027
rect 6193 10993 6227 11027
rect 7310 10993 7344 11027
rect 7435 10993 7469 11027
rect 8769 10993 8803 11027
rect 10149 10993 10183 11027
rect 14933 10993 14967 11027
rect 15117 10993 15151 11027
rect 11621 10925 11655 10959
rect 4169 10721 4203 10755
rect 5825 10721 5859 10755
rect 9413 10721 9447 10755
rect 11069 10721 11103 10755
rect 3341 10653 3375 10687
rect 3893 10653 3927 10687
rect 6101 10653 6135 10687
rect 11253 10653 11287 10687
rect 949 10585 983 10619
rect 3157 10585 3191 10619
rect 3433 10585 3467 10619
rect 1225 10517 1259 10551
rect 2697 10517 2731 10551
rect 3985 10585 4019 10619
rect 4721 10585 4755 10619
rect 6009 10585 6043 10619
rect 6239 10585 6273 10619
rect 6377 10585 6411 10619
rect 9321 10585 9355 10619
rect 9597 10585 9631 10619
rect 11437 10585 11471 10619
rect 12081 10585 12115 10619
rect 12541 10585 12575 10619
rect 15117 10585 15151 10619
rect 6837 10517 6871 10551
rect 7113 10517 7147 10551
rect 3893 10449 3927 10483
rect 9597 10449 9631 10483
rect 3157 10381 3191 10415
rect 4813 10381 4847 10415
rect 8585 10381 8619 10415
rect 11897 10381 11931 10415
rect 12725 10381 12759 10415
rect 14933 10381 14967 10415
rect 673 10177 707 10211
rect 1317 10177 1351 10211
rect 2237 10177 2271 10211
rect 8769 10177 8803 10211
rect 10241 10177 10275 10211
rect 14289 10177 14323 10211
rect 3525 10109 3559 10143
rect 9781 10109 9815 10143
rect 10977 10109 11011 10143
rect 489 9973 523 10007
rect 673 9973 707 10007
rect 1133 9973 1167 10007
rect 1317 9973 1351 10007
rect 6009 9973 6043 10007
rect 6469 9973 6503 10007
rect 8493 9973 8527 10007
rect 9505 9973 9539 10007
rect 10241 9973 10275 10007
rect 10425 9973 10459 10007
rect 11069 9973 11103 10007
rect 11529 9973 11563 10007
rect 12633 9973 12667 10007
rect 14381 9973 14415 10007
rect 2145 9905 2179 9939
rect 3341 9905 3375 9939
rect 5733 9905 5767 9939
rect 7297 9905 7331 9939
rect 8677 9905 8711 9939
rect 9784 9905 9818 9939
rect 14933 9905 14967 9939
rect 15117 9905 15151 9939
rect 4261 9837 4295 9871
rect 9597 9837 9631 9871
rect 11713 9837 11747 9871
rect 12725 9837 12759 9871
rect 5825 9633 5859 9667
rect 7205 9633 7239 9667
rect 12265 9633 12299 9667
rect 14749 9633 14783 9667
rect 949 9565 983 9599
rect 6331 9565 6365 9599
rect 1501 9497 1535 9531
rect 4261 9497 4295 9531
rect 4445 9497 4479 9531
rect 6010 9497 6044 9531
rect 6101 9497 6135 9531
rect 6206 9497 6240 9531
rect 7389 9497 7423 9531
rect 7481 9497 7515 9531
rect 7573 9497 7607 9531
rect 7711 9497 7745 9531
rect 8309 9497 8343 9531
rect 8493 9497 8527 9531
rect 9137 9497 9171 9531
rect 10149 9497 10183 9531
rect 11437 9497 11471 9531
rect 11529 9497 11563 9531
rect 11805 9497 11839 9531
rect 12265 9497 12299 9531
rect 12442 9497 12476 9531
rect 12909 9497 12943 9531
rect 13093 9497 13127 9531
rect 14013 9497 14047 9531
rect 14657 9497 14691 9531
rect 765 9429 799 9463
rect 1777 9429 1811 9463
rect 3249 9429 3283 9463
rect 6469 9429 6503 9463
rect 7849 9429 7883 9463
rect 4629 9361 4663 9395
rect 8309 9361 8343 9395
rect 9045 9293 9079 9327
rect 10057 9293 10091 9327
rect 11253 9293 11287 9327
rect 11713 9293 11747 9327
rect 13093 9293 13127 9327
rect 14105 9293 14139 9327
rect 1869 9089 1903 9123
rect 7481 9089 7515 9123
rect 3249 9021 3283 9055
rect 4721 8953 4755 8987
rect 6653 8953 6687 8987
rect 10425 8953 10459 8987
rect 10793 8953 10827 8987
rect 14197 8953 14231 8987
rect 949 8885 983 8919
rect 2145 8885 2179 8919
rect 3249 8885 3283 8919
rect 3433 8885 3467 8919
rect 3525 8885 3559 8919
rect 4077 8885 4111 8919
rect 4235 8885 4269 8919
rect 4445 8885 4479 8919
rect 4537 8885 4571 8919
rect 6929 8885 6963 8919
rect 7389 8885 7423 8919
rect 8769 8885 8803 8919
rect 9413 8885 9447 8919
rect 13921 8885 13955 8919
rect 14013 8885 14047 8919
rect 14289 8885 14323 8919
rect 765 8817 799 8851
rect 1869 8817 1903 8851
rect 4353 8817 4387 8851
rect 13737 8817 13771 8851
rect 14933 8817 14967 8851
rect 15117 8817 15151 8851
rect 2053 8749 2087 8783
rect 5181 8749 5215 8783
rect 8677 8749 8711 8783
rect 9321 8749 9355 8783
rect 12219 8749 12253 8783
rect 673 8545 707 8579
rect 9321 8545 9355 8579
rect 11161 8545 11195 8579
rect 2881 8477 2915 8511
rect 3065 8477 3099 8511
rect 4629 8477 4663 8511
rect 11989 8477 12023 8511
rect 12081 8477 12115 8511
rect 2421 8409 2455 8443
rect 4399 8409 4433 8443
rect 4537 8409 4571 8443
rect 4721 8409 4755 8443
rect 8125 8409 8159 8443
rect 8309 8409 8343 8443
rect 9505 8409 9539 8443
rect 9689 8409 9723 8443
rect 9965 8409 9999 8443
rect 11253 8409 11287 8443
rect 11897 8409 11931 8443
rect 12265 8409 12299 8443
rect 12725 8409 12759 8443
rect 2145 8341 2179 8375
rect 4261 8341 4295 8375
rect 4905 8341 4939 8375
rect 7389 8341 7423 8375
rect 7665 8341 7699 8375
rect 9781 8341 9815 8375
rect 13093 8341 13127 8375
rect 3249 8273 3283 8307
rect 9597 8273 9631 8307
rect 11713 8273 11747 8307
rect 5917 8205 5951 8239
rect 8217 8205 8251 8239
rect 14519 8205 14553 8239
rect 2053 8001 2087 8035
rect 4261 8001 4295 8035
rect 10241 8001 10275 8035
rect 11069 8001 11103 8035
rect 12817 8001 12851 8035
rect 1225 7933 1259 7967
rect 5365 7933 5399 7967
rect 14749 7933 14783 7967
rect 5917 7865 5951 7899
rect 7297 7865 7331 7899
rect 8769 7865 8803 7899
rect 11713 7865 11747 7899
rect 12173 7865 12207 7899
rect 14197 7865 14231 7899
rect 673 7797 707 7831
rect 1409 7797 1443 7831
rect 2329 7797 2363 7831
rect 3433 7797 3467 7831
rect 4077 7797 4111 7831
rect 5641 7797 5675 7831
rect 6745 7797 6779 7831
rect 7481 7797 7515 7831
rect 7573 7797 7607 7831
rect 8493 7797 8527 7831
rect 11253 7797 11287 7831
rect 11345 7797 11379 7831
rect 12541 7797 12575 7831
rect 12633 7797 12667 7831
rect 13904 7797 13938 7831
rect 14013 7797 14047 7831
rect 14289 7797 14323 7831
rect 14933 7797 14967 7831
rect 489 7729 523 7763
rect 1593 7729 1627 7763
rect 2053 7729 2087 7763
rect 6561 7729 6595 7763
rect 11621 7729 11655 7763
rect 12265 7729 12299 7763
rect 2237 7661 2271 7695
rect 3617 7661 3651 7695
rect 5825 7661 5859 7695
rect 7297 7661 7331 7695
rect 13737 7661 13771 7695
rect 3617 7457 3651 7491
rect 4077 7457 4111 7491
rect 9321 7457 9355 7491
rect 11069 7457 11103 7491
rect 1961 7389 1995 7423
rect 6837 7389 6871 7423
rect 7849 7389 7883 7423
rect 3157 7321 3191 7355
rect 3893 7321 3927 7355
rect 3985 7321 4019 7355
rect 5825 7321 5859 7355
rect 6009 7321 6043 7355
rect 6101 7321 6135 7355
rect 6360 7321 6394 7355
rect 7021 7321 7055 7355
rect 7573 7321 7607 7355
rect 9781 7321 9815 7355
rect 9965 7321 9999 7355
rect 11253 7321 11287 7355
rect 11529 7321 11563 7355
rect 11621 7321 11655 7355
rect 11805 7321 11839 7355
rect 12725 7321 12759 7355
rect 2237 7253 2271 7287
rect 4353 7253 4387 7287
rect 11437 7253 11471 7287
rect 13093 7253 13127 7287
rect 10057 7185 10091 7219
rect 489 7117 523 7151
rect 3065 7117 3099 7151
rect 4261 7117 4295 7151
rect 5825 7117 5859 7151
rect 6285 7117 6319 7151
rect 14519 7117 14553 7151
rect 3433 6913 3467 6947
rect 3617 6913 3651 6947
rect 7021 6913 7055 6947
rect 4445 6845 4479 6879
rect 14749 6845 14783 6879
rect 4537 6777 4571 6811
rect 9689 6777 9723 6811
rect 10149 6777 10183 6811
rect 11529 6777 11563 6811
rect 12081 6777 12115 6811
rect 14197 6777 14231 6811
rect 949 6709 983 6743
rect 1685 6709 1719 6743
rect 2145 6709 2179 6743
rect 2329 6709 2363 6743
rect 4629 6709 4663 6743
rect 4997 6709 5031 6743
rect 5089 6709 5123 6743
rect 5917 6709 5951 6743
rect 6377 6709 6411 6743
rect 6561 6709 6595 6743
rect 6656 6709 6690 6743
rect 6745 6709 6779 6743
rect 8861 6709 8895 6743
rect 9597 6709 9631 6743
rect 10057 6709 10091 6743
rect 10425 6709 10459 6743
rect 10609 6709 10643 6743
rect 11897 6709 11931 6743
rect 12817 6709 12851 6743
rect 13921 6709 13955 6743
rect 14013 6709 14047 6743
rect 14289 6709 14323 6743
rect 14933 6709 14967 6743
rect 765 6641 799 6675
rect 3249 6641 3283 6675
rect 3454 6641 3488 6675
rect 8493 6641 8527 6675
rect 8677 6641 8711 6675
rect 13737 6641 13771 6675
rect 1593 6573 1627 6607
rect 2329 6573 2363 6607
rect 11621 6573 11655 6607
rect 11713 6573 11747 6607
rect 12725 6573 12759 6607
rect 3341 6369 3375 6403
rect 3801 6369 3835 6403
rect 4905 6369 4939 6403
rect 7941 6369 7975 6403
rect 11529 6369 11563 6403
rect 13277 6369 13311 6403
rect 14381 6369 14415 6403
rect 949 6301 983 6335
rect 9781 6301 9815 6335
rect 12909 6301 12943 6335
rect 3709 6233 3743 6267
rect 4537 6233 4571 6267
rect 4721 6233 4755 6267
rect 6193 6233 6227 6267
rect 6653 6233 6687 6267
rect 8861 6233 8895 6267
rect 9045 6233 9079 6267
rect 11437 6233 11471 6267
rect 11621 6233 11655 6267
rect 12081 6233 12115 6267
rect 12725 6233 12759 6267
rect 13001 6233 13035 6267
rect 13093 6233 13127 6267
rect 14473 6233 14507 6267
rect 14933 6233 14967 6267
rect 15117 6233 15151 6267
rect 673 6165 707 6199
rect 2697 6165 2731 6199
rect 3985 6165 4019 6199
rect 12173 6165 12207 6199
rect 6101 6097 6135 6131
rect 9137 6097 9171 6131
rect 4537 6029 4571 6063
rect 9873 6029 9907 6063
rect 14933 6029 14967 6063
rect 857 5825 891 5859
rect 3525 5825 3559 5859
rect 5457 5825 5491 5859
rect 6653 5825 6687 5859
rect 8585 5825 8619 5859
rect 13829 5825 13863 5859
rect 1593 5757 1627 5791
rect 2329 5689 2363 5723
rect 6009 5689 6043 5723
rect 7113 5689 7147 5723
rect 12633 5689 12667 5723
rect 673 5621 707 5655
rect 857 5621 891 5655
rect 2145 5621 2179 5655
rect 4261 5621 4295 5655
rect 4353 5621 4387 5655
rect 4537 5621 4571 5655
rect 5825 5621 5859 5655
rect 5917 5621 5951 5655
rect 6837 5621 6871 5655
rect 6929 5621 6963 5655
rect 7205 5621 7239 5655
rect 8677 5621 8711 5655
rect 9229 5621 9263 5655
rect 11897 5621 11931 5655
rect 12541 5621 12575 5655
rect 13737 5621 13771 5655
rect 1409 5553 1443 5587
rect 3341 5553 3375 5587
rect 3525 5553 3559 5587
rect 4997 5553 5031 5587
rect 9505 5553 9539 5587
rect 14933 5553 14967 5587
rect 3709 5485 3743 5519
rect 10977 5485 11011 5519
rect 11989 5485 12023 5519
rect 15025 5485 15059 5519
rect 3065 5281 3099 5315
rect 5825 5281 5859 5315
rect 9413 5281 9447 5315
rect 9873 5281 9907 5315
rect 11069 5281 11103 5315
rect 11437 5281 11471 5315
rect 857 5213 891 5247
rect 2605 5213 2639 5247
rect 6193 5213 6227 5247
rect 12817 5213 12851 5247
rect 14933 5213 14967 5247
rect 15117 5213 15151 5247
rect 3249 5145 3283 5179
rect 3433 5145 3467 5179
rect 3985 5145 4019 5179
rect 4077 5145 4111 5179
rect 4261 5145 4295 5179
rect 6101 5145 6135 5179
rect 6285 5145 6319 5179
rect 7297 5145 7331 5179
rect 8309 5145 8343 5179
rect 8493 5145 8527 5179
rect 8769 5145 8803 5179
rect 9781 5145 9815 5179
rect 11529 5145 11563 5179
rect 14752 5145 14786 5179
rect 581 5077 615 5111
rect 3525 5077 3559 5111
rect 4721 5077 4755 5111
rect 6561 5077 6595 5111
rect 7113 5077 7147 5111
rect 7205 5077 7239 5111
rect 7389 5077 7423 5111
rect 7573 5077 7607 5111
rect 10057 5077 10091 5111
rect 11713 5077 11747 5111
rect 12541 5077 12575 5111
rect 14289 5077 14323 5111
rect 8953 5009 8987 5043
rect 6469 4941 6503 4975
rect 4997 4737 5031 4771
rect 11253 4737 11287 4771
rect 12817 4737 12851 4771
rect 14197 4737 14231 4771
rect 765 4669 799 4703
rect 11805 4669 11839 4703
rect 14749 4669 14783 4703
rect 1685 4601 1719 4635
rect 2145 4601 2179 4635
rect 3893 4601 3927 4635
rect 5641 4601 5675 4635
rect 6929 4601 6963 4635
rect 8769 4601 8803 4635
rect 949 4533 983 4567
rect 1777 4533 1811 4567
rect 3709 4533 3743 4567
rect 6837 4533 6871 4567
rect 7021 4533 7055 4567
rect 7113 4533 7147 4567
rect 11805 4533 11839 4567
rect 11989 4533 12023 4567
rect 12541 4533 12575 4567
rect 12633 4533 12667 4567
rect 14105 4533 14139 4567
rect 14749 4533 14783 4567
rect 14933 4533 14967 4567
rect 15025 4533 15059 4567
rect 2053 4465 2087 4499
rect 5457 4465 5491 4499
rect 9045 4465 9079 4499
rect 10977 4465 11011 4499
rect 11161 4465 11195 4499
rect 12817 4465 12851 4499
rect 13921 4465 13955 4499
rect 1501 4397 1535 4431
rect 3249 4397 3283 4431
rect 3617 4397 3651 4431
rect 5365 4397 5399 4431
rect 6653 4397 6687 4431
rect 10517 4397 10551 4431
rect 3157 4193 3191 4227
rect 4077 4193 4111 4227
rect 8217 4193 8251 4227
rect 9413 4193 9447 4227
rect 14289 4193 14323 4227
rect 7389 4125 7423 4159
rect 7573 4125 7607 4159
rect 8585 4125 8619 4159
rect 9781 4125 9815 4159
rect 14933 4125 14967 4159
rect 3341 4057 3375 4091
rect 4353 4057 4387 4091
rect 4445 4057 4479 4091
rect 4537 4057 4571 4091
rect 4721 4057 4755 4091
rect 6009 4057 6043 4091
rect 6193 4057 6227 4091
rect 9597 4057 9631 4091
rect 9689 4057 9723 4091
rect 9919 4057 9953 4091
rect 11069 4057 11103 4091
rect 11897 4057 11931 4091
rect 12081 4057 12115 4091
rect 12541 4057 12575 4091
rect 857 3989 891 4023
rect 1133 3989 1167 4023
rect 3617 3989 3651 4023
rect 8677 3989 8711 4023
rect 8861 3989 8895 4023
rect 10057 3989 10091 4023
rect 12817 3989 12851 4023
rect 15117 3989 15151 4023
rect 6377 3921 6411 3955
rect 7757 3921 7791 3955
rect 2605 3853 2639 3887
rect 3525 3853 3559 3887
rect 6193 3853 6227 3887
rect 11253 3853 11287 3887
rect 12081 3853 12115 3887
rect 857 3649 891 3683
rect 2237 3649 2271 3683
rect 3525 3649 3559 3683
rect 4261 3649 4295 3683
rect 5365 3649 5399 3683
rect 6837 3649 6871 3683
rect 14657 3649 14691 3683
rect 1685 3581 1719 3615
rect 11161 3581 11195 3615
rect 12817 3581 12851 3615
rect 13829 3581 13863 3615
rect 5273 3513 5307 3547
rect 5365 3513 5399 3547
rect 6009 3513 6043 3547
rect 11989 3513 12023 3547
rect 1501 3445 1535 3479
rect 2329 3445 2363 3479
rect 4169 3445 4203 3479
rect 5181 3445 5215 3479
rect 6193 3445 6227 3479
rect 7021 3445 7055 3479
rect 7205 3445 7239 3479
rect 9413 3445 9447 3479
rect 9597 3445 9631 3479
rect 9873 3445 9907 3479
rect 10425 3445 10459 3479
rect 11069 3445 11103 3479
rect 11897 3445 11931 3479
rect 12081 3445 12115 3479
rect 12541 3445 12575 3479
rect 14013 3445 14047 3479
rect 14841 3445 14875 3479
rect 14933 3445 14967 3479
rect 949 3377 983 3411
rect 3504 3377 3538 3411
rect 3709 3377 3743 3411
rect 5549 3377 5583 3411
rect 8677 3377 8711 3411
rect 9505 3377 9539 3411
rect 9735 3377 9769 3411
rect 12817 3377 12851 3411
rect 14197 3377 14231 3411
rect 14657 3377 14691 3411
rect 3341 3309 3375 3343
rect 8585 3309 8619 3343
rect 9229 3309 9263 3343
rect 10517 3309 10551 3343
rect 12633 3309 12667 3343
rect 3249 3105 3283 3139
rect 4261 3105 4295 3139
rect 5825 3105 5859 3139
rect 10149 3105 10183 3139
rect 14197 3105 14231 3139
rect 1225 3037 1259 3071
rect 4813 3037 4847 3071
rect 7021 3037 7055 3071
rect 7849 3037 7883 3071
rect 11345 3037 11379 3071
rect 12725 3037 12759 3071
rect 14933 3037 14967 3071
rect 3157 2969 3191 3003
rect 4077 2969 4111 3003
rect 4721 2969 4755 3003
rect 6009 2969 6043 3003
rect 6101 2969 6135 3003
rect 6193 2969 6227 3003
rect 6377 2969 6411 3003
rect 7665 2969 7699 3003
rect 8401 2969 8435 3003
rect 11253 2969 11287 3003
rect 11437 2969 11471 3003
rect 11575 2969 11609 3003
rect 949 2901 983 2935
rect 8677 2901 8711 2935
rect 11713 2901 11747 2935
rect 12449 2901 12483 2935
rect 15117 2833 15151 2867
rect 2697 2765 2731 2799
rect 6929 2765 6963 2799
rect 11069 2765 11103 2799
rect 1593 2561 1627 2595
rect 2329 2561 2363 2595
rect 9045 2561 9079 2595
rect 14013 2561 14047 2595
rect 15025 2561 15059 2595
rect 4261 2425 4295 2459
rect 10517 2425 10551 2459
rect 11897 2425 11931 2459
rect 1685 2357 1719 2391
rect 2145 2357 2179 2391
rect 2329 2357 2363 2391
rect 3985 2357 4019 2391
rect 4169 2357 4203 2391
rect 4721 2357 4755 2391
rect 7389 2357 7423 2391
rect 10793 2357 10827 2391
rect 11437 2357 11471 2391
rect 11621 2357 11655 2391
rect 12633 2357 12667 2391
rect 12817 2357 12851 2391
rect 13737 2357 13771 2391
rect 13921 2357 13955 2391
rect 14933 2357 14967 2391
rect 857 2289 891 2323
rect 4997 2289 5031 2323
rect 6745 2289 6779 2323
rect 7205 2289 7239 2323
rect 11529 2289 11563 2323
rect 11739 2289 11773 2323
rect 949 2221 983 2255
rect 3801 2221 3835 2255
rect 11253 2221 11287 2255
rect 12725 2221 12759 2255
rect 1133 2017 1167 2051
rect 6653 2017 6687 2051
rect 11713 2017 11747 2051
rect 4721 1949 4755 1983
rect 7573 1949 7607 1983
rect 8677 1949 8711 1983
rect 12633 1949 12667 1983
rect 14933 1949 14967 1983
rect 581 1881 615 1915
rect 1225 1881 1259 1915
rect 4629 1881 4663 1915
rect 4905 1881 4939 1915
rect 7389 1881 7423 1915
rect 7481 1881 7515 1915
rect 7757 1881 7791 1915
rect 11069 1881 11103 1915
rect 11897 1881 11931 1915
rect 1685 1813 1719 1847
rect 1961 1813 1995 1847
rect 4169 1813 4203 1847
rect 4261 1813 4295 1847
rect 6377 1813 6411 1847
rect 8401 1813 8435 1847
rect 10149 1813 10183 1847
rect 12357 1813 12391 1847
rect 489 1745 523 1779
rect 3433 1745 3467 1779
rect 5825 1745 5859 1779
rect 14105 1745 14139 1779
rect 15117 1745 15151 1779
rect 6193 1677 6227 1711
rect 6285 1677 6319 1711
rect 7205 1677 7239 1711
rect 11161 1677 11195 1711
rect 4721 1473 4755 1507
rect 10793 1473 10827 1507
rect 12081 1405 12115 1439
rect 5273 1337 5307 1371
rect 7021 1337 7055 1371
rect 9321 1337 9355 1371
rect 857 1269 891 1303
rect 2329 1269 2363 1303
rect 4261 1269 4295 1303
rect 4445 1269 4479 1303
rect 4537 1269 4571 1303
rect 4813 1269 4847 1303
rect 7297 1269 7331 1303
rect 9045 1269 9079 1303
rect 11437 1269 11471 1303
rect 11897 1269 11931 1303
rect 14289 1269 14323 1303
rect 14933 1269 14967 1303
rect 1501 1201 1535 1235
rect 3249 1201 3283 1235
rect 3433 1201 3467 1235
rect 765 1133 799 1167
rect 11253 1133 11287 1167
rect 14381 1133 14415 1167
rect 15117 1133 15151 1167
rect 5917 929 5951 963
rect 6837 929 6871 963
rect 9137 929 9171 963
rect 1133 861 1167 895
rect 3525 861 3559 895
rect 6069 861 6103 895
rect 6285 861 6319 895
rect 11437 861 11471 895
rect 12817 861 12851 895
rect 14197 861 14231 895
rect 14933 861 14967 895
rect 2145 793 2179 827
rect 6929 793 6963 827
rect 7481 793 7515 827
rect 9321 793 9355 827
rect 9413 793 9447 827
rect 9505 793 9539 827
rect 9689 793 9723 827
rect 10333 793 10367 827
rect 3249 725 3283 759
rect 949 657 983 691
rect 4997 657 5031 691
rect 7665 657 7699 691
rect 11253 657 11287 691
rect 14381 657 14415 691
rect 2237 589 2271 623
rect 6101 589 6135 623
rect 10149 589 10183 623
rect 12909 589 12943 623
rect 15025 589 15059 623
<< metal1 >>
rect 92 13042 15824 13064
rect 92 12990 5242 13042
rect 5294 12990 5306 13042
rect 5358 12990 5370 13042
rect 5422 12990 5434 13042
rect 5486 12990 10514 13042
rect 10566 12990 10578 13042
rect 10630 12990 10642 13042
rect 10694 12990 10706 13042
rect 10758 12990 15824 13042
rect 92 12968 15824 12990
rect 4890 12928 4896 12940
rect 4851 12900 4896 12928
rect 4890 12888 4896 12900
rect 4948 12888 4954 12940
rect 8938 12888 8944 12940
rect 8996 12928 9002 12940
rect 12894 12928 12900 12940
rect 8996 12900 9628 12928
rect 12855 12900 12900 12928
rect 8996 12888 9002 12900
rect 934 12860 940 12872
rect 895 12832 940 12860
rect 934 12820 940 12832
rect 992 12820 998 12872
rect 2866 12820 2872 12872
rect 2924 12860 2930 12872
rect 3237 12863 3295 12869
rect 3237 12860 3249 12863
rect 2924 12832 3249 12860
rect 2924 12820 2930 12832
rect 3237 12829 3249 12832
rect 3283 12829 3295 12863
rect 3970 12860 3976 12872
rect 3931 12832 3976 12860
rect 3237 12823 3295 12829
rect 3970 12820 3976 12832
rect 4028 12820 4034 12872
rect 6914 12820 6920 12872
rect 6972 12860 6978 12872
rect 9600 12869 9628 12900
rect 12894 12888 12900 12900
rect 12952 12888 12958 12940
rect 14918 12888 14924 12940
rect 14976 12928 14982 12940
rect 15013 12931 15071 12937
rect 15013 12928 15025 12931
rect 14976 12900 15025 12928
rect 14976 12888 14982 12900
rect 15013 12897 15025 12900
rect 15059 12897 15071 12931
rect 15013 12891 15071 12897
rect 9585 12863 9643 12869
rect 6972 12832 7017 12860
rect 6972 12820 6978 12832
rect 9585 12829 9597 12863
rect 9631 12829 9643 12863
rect 9585 12823 9643 12829
rect 10870 12820 10876 12872
rect 10928 12860 10934 12872
rect 11241 12863 11299 12869
rect 11241 12860 11253 12863
rect 10928 12832 11253 12860
rect 10928 12820 10934 12832
rect 11241 12829 11253 12832
rect 11287 12829 11299 12863
rect 14366 12860 14372 12872
rect 14327 12832 14372 12860
rect 11241 12823 11299 12829
rect 14366 12820 14372 12832
rect 14424 12820 14430 12872
rect 1118 12792 1124 12804
rect 1079 12764 1124 12792
rect 1118 12752 1124 12764
rect 1176 12752 1182 12804
rect 1854 12792 1860 12804
rect 1815 12764 1860 12792
rect 1854 12752 1860 12764
rect 1912 12752 1918 12804
rect 3418 12792 3424 12804
rect 3379 12764 3424 12792
rect 3418 12752 3424 12764
rect 3476 12752 3482 12804
rect 3510 12752 3516 12804
rect 3568 12792 3574 12804
rect 4157 12795 4215 12801
rect 4157 12792 4169 12795
rect 3568 12764 4169 12792
rect 3568 12752 3574 12764
rect 4157 12761 4169 12764
rect 4203 12761 4215 12795
rect 4157 12755 4215 12761
rect 4801 12795 4859 12801
rect 4801 12761 4813 12795
rect 4847 12792 4859 12795
rect 4890 12792 4896 12804
rect 4847 12764 4896 12792
rect 4847 12761 4859 12764
rect 4801 12755 4859 12761
rect 4890 12752 4896 12764
rect 4948 12752 4954 12804
rect 5905 12795 5963 12801
rect 5905 12761 5917 12795
rect 5951 12792 5963 12795
rect 7101 12795 7159 12801
rect 5951 12764 6914 12792
rect 5951 12761 5963 12764
rect 5905 12755 5963 12761
rect 6886 12724 6914 12764
rect 7101 12761 7113 12795
rect 7147 12792 7159 12795
rect 7190 12792 7196 12804
rect 7147 12764 7196 12792
rect 7147 12761 7159 12764
rect 7101 12755 7159 12761
rect 7190 12752 7196 12764
rect 7248 12752 7254 12804
rect 8754 12792 8760 12804
rect 8715 12764 8760 12792
rect 8754 12752 8760 12764
rect 8812 12752 8818 12804
rect 8938 12792 8944 12804
rect 8899 12764 8944 12792
rect 8938 12752 8944 12764
rect 8996 12752 9002 12804
rect 9122 12752 9128 12804
rect 9180 12792 9186 12804
rect 9769 12795 9827 12801
rect 9769 12792 9781 12795
rect 9180 12764 9781 12792
rect 9180 12752 9186 12764
rect 9769 12761 9781 12764
rect 9815 12761 9827 12795
rect 11422 12792 11428 12804
rect 11383 12764 11428 12792
rect 9769 12755 9827 12761
rect 11422 12752 11428 12764
rect 11480 12752 11486 12804
rect 12802 12792 12808 12804
rect 12763 12764 12808 12792
rect 12802 12752 12808 12764
rect 12860 12752 12866 12804
rect 14182 12792 14188 12804
rect 14143 12764 14188 12792
rect 14182 12752 14188 12764
rect 14240 12752 14246 12804
rect 14826 12752 14832 12804
rect 14884 12792 14890 12804
rect 14921 12795 14979 12801
rect 14921 12792 14933 12795
rect 14884 12764 14933 12792
rect 14884 12752 14890 12764
rect 14921 12761 14933 12764
rect 14967 12761 14979 12795
rect 14921 12755 14979 12761
rect 7742 12724 7748 12736
rect 6886 12696 7748 12724
rect 7742 12684 7748 12696
rect 7800 12684 7806 12736
rect 6089 12659 6147 12665
rect 6089 12625 6101 12659
rect 6135 12656 6147 12659
rect 12066 12656 12072 12668
rect 6135 12628 12072 12656
rect 6135 12625 6147 12628
rect 6089 12619 6147 12625
rect 12066 12616 12072 12628
rect 12124 12616 12130 12668
rect 1762 12588 1768 12600
rect 1723 12560 1768 12588
rect 1762 12548 1768 12560
rect 1820 12548 1826 12600
rect 9122 12588 9128 12600
rect 9083 12560 9128 12588
rect 9122 12548 9128 12560
rect 9180 12548 9186 12600
rect 92 12498 15824 12520
rect 92 12446 2606 12498
rect 2658 12446 2670 12498
rect 2722 12446 2734 12498
rect 2786 12446 2798 12498
rect 2850 12446 7878 12498
rect 7930 12446 7942 12498
rect 7994 12446 8006 12498
rect 8058 12446 8070 12498
rect 8122 12446 13150 12498
rect 13202 12446 13214 12498
rect 13266 12446 13278 12498
rect 13330 12446 13342 12498
rect 13394 12446 15824 12498
rect 92 12424 15824 12446
rect 934 12344 940 12396
rect 992 12384 998 12396
rect 8754 12384 8760 12396
rect 992 12356 8760 12384
rect 992 12344 998 12356
rect 8754 12344 8760 12356
rect 8812 12384 8818 12396
rect 9490 12384 9496 12396
rect 8812 12356 9496 12384
rect 8812 12344 8818 12356
rect 9490 12344 9496 12356
rect 9548 12384 9554 12396
rect 9677 12387 9735 12393
rect 9677 12384 9689 12387
rect 9548 12356 9689 12384
rect 9548 12344 9554 12356
rect 9677 12353 9689 12356
rect 9723 12353 9735 12387
rect 9677 12347 9735 12353
rect 2317 12251 2375 12257
rect 2317 12217 2329 12251
rect 2363 12217 2375 12251
rect 2317 12211 2375 12217
rect 566 12180 572 12192
rect 527 12152 572 12180
rect 566 12140 572 12152
rect 624 12140 630 12192
rect 2332 12180 2360 12211
rect 6454 12208 6460 12260
rect 6512 12248 6518 12260
rect 6733 12251 6791 12257
rect 6733 12248 6745 12251
rect 6512 12220 6745 12248
rect 6512 12208 6518 12220
rect 6733 12217 6745 12220
rect 6779 12217 6791 12251
rect 8938 12248 8944 12260
rect 6733 12211 6791 12217
rect 8772 12220 8944 12248
rect 4338 12180 4344 12192
rect 2332 12152 2774 12180
rect 4299 12152 4344 12180
rect 842 12112 848 12124
rect 803 12084 848 12112
rect 842 12072 848 12084
rect 900 12072 906 12124
rect 2498 12112 2504 12124
rect 2070 12084 2504 12112
rect 2498 12072 2504 12084
rect 2556 12072 2562 12124
rect 2746 12112 2774 12152
rect 4338 12140 4344 12152
rect 4396 12140 4402 12192
rect 4522 12180 4528 12192
rect 4483 12152 4528 12180
rect 4522 12140 4528 12152
rect 4580 12140 4586 12192
rect 7190 12180 7196 12192
rect 7151 12152 7196 12180
rect 7190 12140 7196 12152
rect 7248 12140 7254 12192
rect 8202 12140 8208 12192
rect 8260 12180 8266 12192
rect 8772 12189 8800 12220
rect 8938 12208 8944 12220
rect 8996 12248 9002 12260
rect 9398 12248 9404 12260
rect 8996 12220 9404 12248
rect 8996 12208 9002 12220
rect 9398 12208 9404 12220
rect 9456 12208 9462 12260
rect 9858 12208 9864 12260
rect 9916 12248 9922 12260
rect 11425 12251 11483 12257
rect 11425 12248 11437 12251
rect 9916 12220 11437 12248
rect 9916 12208 9922 12220
rect 11425 12217 11437 12220
rect 11471 12217 11483 12251
rect 11425 12211 11483 12217
rect 8665 12183 8723 12189
rect 8665 12180 8677 12183
rect 8260 12152 8677 12180
rect 8260 12140 8266 12152
rect 8665 12149 8677 12152
rect 8711 12149 8723 12183
rect 8665 12143 8723 12149
rect 8757 12183 8815 12189
rect 8757 12149 8769 12183
rect 8803 12149 8815 12183
rect 8757 12143 8815 12149
rect 8846 12140 8852 12192
rect 8904 12180 8910 12192
rect 9125 12183 9183 12189
rect 8904 12152 8949 12180
rect 8904 12140 8910 12152
rect 9125 12149 9137 12183
rect 9171 12180 9183 12183
rect 9582 12180 9588 12192
rect 9171 12152 9588 12180
rect 9171 12149 9183 12152
rect 9125 12143 9183 12149
rect 9582 12140 9588 12152
rect 9640 12140 9646 12192
rect 3234 12112 3240 12124
rect 2746 12084 3240 12112
rect 3234 12072 3240 12084
rect 3292 12112 3298 12124
rect 3510 12112 3516 12124
rect 3292 12084 3516 12112
rect 3292 12072 3298 12084
rect 3510 12072 3516 12084
rect 3568 12072 3574 12124
rect 3694 12112 3700 12124
rect 3655 12084 3700 12112
rect 3694 12072 3700 12084
rect 3752 12072 3758 12124
rect 3881 12115 3939 12121
rect 3881 12081 3893 12115
rect 3927 12112 3939 12115
rect 4798 12112 4804 12124
rect 3927 12084 4804 12112
rect 3927 12081 3939 12084
rect 3881 12075 3939 12081
rect 4798 12072 4804 12084
rect 4856 12072 4862 12124
rect 6457 12115 6515 12121
rect 5552 12056 5580 12098
rect 6457 12081 6469 12115
rect 6503 12112 6515 12115
rect 6914 12112 6920 12124
rect 6503 12084 6920 12112
rect 6503 12081 6515 12084
rect 6457 12075 6515 12081
rect 6914 12072 6920 12084
rect 6972 12072 6978 12124
rect 8938 12072 8944 12124
rect 8996 12121 9002 12124
rect 8996 12115 9025 12121
rect 9013 12081 9025 12115
rect 10870 12112 10876 12124
rect 10718 12084 10876 12112
rect 8996 12075 9025 12081
rect 8996 12072 9002 12075
rect 10870 12072 10876 12084
rect 10928 12072 10934 12124
rect 11146 12112 11152 12124
rect 11107 12084 11152 12112
rect 11146 12072 11152 12084
rect 11204 12072 11210 12124
rect 14274 12072 14280 12124
rect 14332 12112 14338 12124
rect 14921 12115 14979 12121
rect 14921 12112 14933 12115
rect 14332 12084 14933 12112
rect 14332 12072 14338 12084
rect 14921 12081 14933 12084
rect 14967 12081 14979 12115
rect 15102 12112 15108 12124
rect 15063 12084 15108 12112
rect 14921 12075 14979 12081
rect 15102 12072 15108 12084
rect 15160 12072 15166 12124
rect 4154 12004 4160 12056
rect 4212 12044 4218 12056
rect 4433 12047 4491 12053
rect 4433 12044 4445 12047
rect 4212 12016 4445 12044
rect 4212 12004 4218 12016
rect 4433 12013 4445 12016
rect 4479 12013 4491 12047
rect 4433 12007 4491 12013
rect 4706 12004 4712 12056
rect 4764 12044 4770 12056
rect 4985 12047 5043 12053
rect 4985 12044 4997 12047
rect 4764 12016 4997 12044
rect 4764 12004 4770 12016
rect 4985 12013 4997 12016
rect 5031 12013 5043 12047
rect 4985 12007 5043 12013
rect 5534 12004 5540 12056
rect 5592 12004 5598 12056
rect 7282 12044 7288 12056
rect 7243 12016 7288 12044
rect 7282 12004 7288 12016
rect 7340 12004 7346 12056
rect 8481 12047 8539 12053
rect 8481 12013 8493 12047
rect 8527 12044 8539 12047
rect 8662 12044 8668 12056
rect 8527 12016 8668 12044
rect 8527 12013 8539 12016
rect 8481 12007 8539 12013
rect 8662 12004 8668 12016
rect 8720 12004 8726 12056
rect 92 11954 15824 11976
rect 92 11902 5242 11954
rect 5294 11902 5306 11954
rect 5358 11902 5370 11954
rect 5422 11902 5434 11954
rect 5486 11902 10514 11954
rect 10566 11902 10578 11954
rect 10630 11902 10642 11954
rect 10694 11902 10706 11954
rect 10758 11902 15824 11954
rect 92 11880 15824 11902
rect 1854 11800 1860 11852
rect 1912 11840 1918 11852
rect 3513 11843 3571 11849
rect 3513 11840 3525 11843
rect 1912 11812 3525 11840
rect 1912 11800 1918 11812
rect 3513 11809 3525 11812
rect 3559 11840 3571 11843
rect 3970 11840 3976 11852
rect 3559 11812 3976 11840
rect 3559 11809 3571 11812
rect 3513 11803 3571 11809
rect 3970 11800 3976 11812
rect 4028 11840 4034 11852
rect 4893 11843 4951 11849
rect 4028 11812 4568 11840
rect 4028 11800 4034 11812
rect 934 11772 940 11784
rect 895 11744 940 11772
rect 934 11732 940 11744
rect 992 11732 998 11784
rect 1302 11732 1308 11784
rect 1360 11772 1366 11784
rect 2041 11775 2099 11781
rect 2041 11772 2053 11775
rect 1360 11744 2053 11772
rect 1360 11732 1366 11744
rect 2041 11741 2053 11744
rect 2087 11741 2099 11775
rect 2041 11735 2099 11741
rect 2498 11732 2504 11784
rect 2556 11732 2562 11784
rect 4540 11781 4568 11812
rect 4893 11809 4905 11843
rect 4939 11840 4951 11843
rect 7190 11840 7196 11852
rect 4939 11812 7196 11840
rect 4939 11809 4951 11812
rect 4893 11803 4951 11809
rect 7190 11800 7196 11812
rect 7248 11800 7254 11852
rect 7929 11843 7987 11849
rect 7929 11809 7941 11843
rect 7975 11840 7987 11843
rect 9398 11840 9404 11852
rect 7975 11812 9404 11840
rect 7975 11809 7987 11812
rect 7929 11803 7987 11809
rect 9398 11800 9404 11812
rect 9456 11800 9462 11852
rect 9582 11800 9588 11852
rect 9640 11840 9646 11852
rect 10137 11843 10195 11849
rect 10137 11840 10149 11843
rect 9640 11812 10149 11840
rect 9640 11800 9646 11812
rect 10137 11809 10149 11812
rect 10183 11809 10195 11843
rect 11146 11840 11152 11852
rect 11107 11812 11152 11840
rect 10137 11803 10195 11809
rect 11146 11800 11152 11812
rect 11204 11800 11210 11852
rect 14182 11800 14188 11852
rect 14240 11840 14246 11852
rect 14369 11843 14427 11849
rect 14369 11840 14381 11843
rect 14240 11812 14381 11840
rect 14240 11800 14246 11812
rect 14369 11809 14381 11812
rect 14415 11809 14427 11843
rect 14369 11803 14427 11809
rect 4525 11775 4583 11781
rect 4525 11741 4537 11775
rect 4571 11741 4583 11775
rect 6454 11772 6460 11784
rect 4525 11735 4583 11741
rect 6196 11744 6460 11772
rect 566 11664 572 11716
rect 624 11704 630 11716
rect 1765 11707 1823 11713
rect 1765 11704 1777 11707
rect 624 11676 1777 11704
rect 624 11664 630 11676
rect 1765 11673 1777 11676
rect 1811 11673 1823 11707
rect 4706 11704 4712 11716
rect 4667 11676 4712 11704
rect 1765 11667 1823 11673
rect 1780 11636 1808 11667
rect 4706 11664 4712 11676
rect 4764 11664 4770 11716
rect 6196 11713 6224 11744
rect 6454 11732 6460 11744
rect 6512 11732 6518 11784
rect 8386 11772 8392 11784
rect 7682 11744 8392 11772
rect 8386 11732 8392 11744
rect 8444 11732 8450 11784
rect 8662 11772 8668 11784
rect 8623 11744 8668 11772
rect 8662 11732 8668 11744
rect 8720 11732 8726 11784
rect 9950 11772 9956 11784
rect 9863 11744 9956 11772
rect 9950 11732 9956 11744
rect 10008 11772 10014 11784
rect 10870 11772 10876 11784
rect 10008 11744 10876 11772
rect 10008 11732 10014 11744
rect 10870 11732 10876 11744
rect 10928 11732 10934 11784
rect 6181 11707 6239 11713
rect 6181 11673 6193 11707
rect 6227 11673 6239 11707
rect 8294 11704 8300 11716
rect 6181 11667 6239 11673
rect 8220 11676 8300 11704
rect 6196 11636 6224 11667
rect 1780 11608 6224 11636
rect 6457 11639 6515 11645
rect 6457 11605 6469 11639
rect 6503 11636 6515 11639
rect 8220 11636 8248 11676
rect 8294 11664 8300 11676
rect 8352 11664 8358 11716
rect 11057 11707 11115 11713
rect 11057 11673 11069 11707
rect 11103 11704 11115 11707
rect 11146 11704 11152 11716
rect 11103 11676 11152 11704
rect 11103 11673 11115 11676
rect 11057 11667 11115 11673
rect 11146 11664 11152 11676
rect 11204 11664 11210 11716
rect 11241 11707 11299 11713
rect 11241 11673 11253 11707
rect 11287 11673 11299 11707
rect 11241 11667 11299 11673
rect 8386 11636 8392 11648
rect 6503 11608 8248 11636
rect 8347 11608 8392 11636
rect 6503 11605 6515 11608
rect 6457 11599 6515 11605
rect 8386 11596 8392 11608
rect 8444 11596 8450 11648
rect 9674 11636 9680 11648
rect 8496 11608 9680 11636
rect 750 11568 756 11580
rect 711 11540 756 11568
rect 750 11528 756 11540
rect 808 11528 814 11580
rect 8496 11568 8524 11608
rect 9674 11596 9680 11608
rect 9732 11596 9738 11648
rect 10042 11596 10048 11648
rect 10100 11636 10106 11648
rect 11256 11636 11284 11667
rect 13998 11664 14004 11716
rect 14056 11704 14062 11716
rect 14277 11707 14335 11713
rect 14277 11704 14289 11707
rect 14056 11676 14289 11704
rect 14056 11664 14062 11676
rect 14277 11673 14289 11676
rect 14323 11673 14335 11707
rect 14277 11667 14335 11673
rect 10100 11608 11284 11636
rect 10100 11596 10106 11608
rect 7484 11540 8524 11568
rect 3602 11460 3608 11512
rect 3660 11500 3666 11512
rect 7484 11500 7512 11540
rect 3660 11472 7512 11500
rect 3660 11460 3666 11472
rect 7558 11460 7564 11512
rect 7616 11500 7622 11512
rect 8846 11500 8852 11512
rect 7616 11472 8852 11500
rect 7616 11460 7622 11472
rect 8846 11460 8852 11472
rect 8904 11460 8910 11512
rect 92 11410 15824 11432
rect 92 11358 2606 11410
rect 2658 11358 2670 11410
rect 2722 11358 2734 11410
rect 2786 11358 2798 11410
rect 2850 11358 7878 11410
rect 7930 11358 7942 11410
rect 7994 11358 8006 11410
rect 8058 11358 8070 11410
rect 8122 11358 13150 11410
rect 13202 11358 13214 11410
rect 13266 11358 13278 11410
rect 13330 11358 13342 11410
rect 13394 11358 15824 11410
rect 92 11336 15824 11358
rect 842 11256 848 11308
rect 900 11296 906 11308
rect 2041 11299 2099 11305
rect 2041 11296 2053 11299
rect 900 11268 2053 11296
rect 900 11256 906 11268
rect 2041 11265 2053 11268
rect 2087 11265 2099 11299
rect 3602 11296 3608 11308
rect 2041 11259 2099 11265
rect 2148 11268 3608 11296
rect 2148 11160 2176 11268
rect 3602 11256 3608 11268
rect 3660 11256 3666 11308
rect 6914 11296 6920 11308
rect 6875 11268 6920 11296
rect 6914 11256 6920 11268
rect 6972 11256 6978 11308
rect 8294 11256 8300 11308
rect 8352 11296 8358 11308
rect 8481 11299 8539 11305
rect 8481 11296 8493 11299
rect 8352 11268 8493 11296
rect 8352 11256 8358 11268
rect 8481 11265 8493 11268
rect 8527 11265 8539 11299
rect 8481 11259 8539 11265
rect 8570 11256 8576 11308
rect 8628 11296 8634 11308
rect 9950 11296 9956 11308
rect 8628 11268 9956 11296
rect 8628 11256 8634 11268
rect 9950 11256 9956 11268
rect 10008 11256 10014 11308
rect 14274 11296 14280 11308
rect 14235 11268 14280 11296
rect 14274 11256 14280 11268
rect 14332 11256 14338 11308
rect 3237 11231 3295 11237
rect 3237 11228 3249 11231
rect 952 11132 2176 11160
rect 2746 11200 3249 11228
rect 952 11101 980 11132
rect 937 11095 995 11101
rect 937 11061 949 11095
rect 983 11061 995 11095
rect 1854 11092 1860 11104
rect 1815 11064 1860 11092
rect 937 11055 995 11061
rect 1854 11052 1860 11064
rect 1912 11052 1918 11104
rect 2041 11095 2099 11101
rect 2041 11061 2053 11095
rect 2087 11092 2099 11095
rect 2746 11092 2774 11200
rect 3237 11197 3249 11200
rect 3283 11197 3295 11231
rect 3237 11191 3295 11197
rect 3418 11188 3424 11240
rect 3476 11228 3482 11240
rect 3973 11231 4031 11237
rect 3973 11228 3985 11231
rect 3476 11200 3985 11228
rect 3476 11188 3482 11200
rect 3973 11197 3985 11200
rect 4019 11197 4031 11231
rect 3973 11191 4031 11197
rect 7024 11200 7420 11228
rect 3694 11120 3700 11172
rect 3752 11160 3758 11172
rect 4709 11163 4767 11169
rect 4709 11160 4721 11163
rect 3752 11132 4721 11160
rect 3752 11120 3758 11132
rect 4709 11129 4721 11132
rect 4755 11160 4767 11163
rect 6178 11160 6184 11172
rect 4755 11132 6184 11160
rect 4755 11129 4767 11132
rect 4709 11123 4767 11129
rect 6178 11120 6184 11132
rect 6236 11120 6242 11172
rect 3234 11092 3240 11104
rect 2087 11064 2774 11092
rect 3195 11064 3240 11092
rect 2087 11061 2099 11064
rect 2041 11055 2099 11061
rect 3234 11052 3240 11064
rect 3292 11052 3298 11104
rect 3510 11092 3516 11104
rect 3423 11064 3516 11092
rect 3510 11052 3516 11064
rect 3568 11092 3574 11104
rect 3970 11092 3976 11104
rect 3568 11064 3832 11092
rect 3931 11064 3976 11092
rect 3568 11052 3574 11064
rect 750 11024 756 11036
rect 711 10996 756 11024
rect 750 10984 756 10996
rect 808 10984 814 11036
rect 3421 11027 3479 11033
rect 3421 10993 3433 11027
rect 3467 11024 3479 11027
rect 3694 11024 3700 11036
rect 3467 10996 3700 11024
rect 3467 10993 3479 10996
rect 3421 10987 3479 10993
rect 3694 10984 3700 10996
rect 3752 10984 3758 11036
rect 3804 11024 3832 11064
rect 3970 11052 3976 11064
rect 4028 11052 4034 11104
rect 4062 11052 4068 11104
rect 4120 11092 4126 11104
rect 4157 11095 4215 11101
rect 4157 11092 4169 11095
rect 4120 11064 4169 11092
rect 4120 11052 4126 11064
rect 4157 11061 4169 11064
rect 4203 11061 4215 11095
rect 4157 11055 4215 11061
rect 4249 11095 4307 11101
rect 4249 11061 4261 11095
rect 4295 11092 4307 11095
rect 4430 11092 4436 11104
rect 4295 11064 4436 11092
rect 4295 11061 4307 11064
rect 4249 11055 4307 11061
rect 4264 11024 4292 11055
rect 4430 11052 4436 11064
rect 4488 11052 4494 11104
rect 6454 11052 6460 11104
rect 6512 11092 6518 11104
rect 6822 11092 6828 11104
rect 6512 11064 6828 11092
rect 6512 11052 6518 11064
rect 6822 11052 6828 11064
rect 6880 11052 6886 11104
rect 7024 11092 7052 11200
rect 7392 11172 7420 11200
rect 7466 11188 7472 11240
rect 7524 11228 7530 11240
rect 8938 11228 8944 11240
rect 7524 11200 8944 11228
rect 7524 11188 7530 11200
rect 8312 11172 8340 11200
rect 8938 11188 8944 11200
rect 8996 11188 9002 11240
rect 7374 11120 7380 11172
rect 7432 11160 7438 11172
rect 8202 11160 8208 11172
rect 7432 11132 8208 11160
rect 7432 11120 7438 11132
rect 8202 11120 8208 11132
rect 8260 11120 8266 11172
rect 8294 11120 8300 11172
rect 8352 11120 8358 11172
rect 8386 11120 8392 11172
rect 8444 11160 8450 11172
rect 9858 11160 9864 11172
rect 8444 11132 9864 11160
rect 8444 11120 8450 11132
rect 9858 11120 9864 11132
rect 9916 11120 9922 11172
rect 7102 11095 7160 11101
rect 7102 11092 7114 11095
rect 7024 11064 7114 11092
rect 7102 11061 7114 11064
rect 7148 11061 7160 11095
rect 7102 11055 7160 11061
rect 7190 11052 7196 11104
rect 7248 11092 7254 11104
rect 7561 11095 7619 11101
rect 7248 11064 7293 11092
rect 7248 11052 7254 11064
rect 7561 11061 7573 11095
rect 7607 11061 7619 11095
rect 8220 11092 8248 11120
rect 8665 11095 8723 11101
rect 8665 11092 8677 11095
rect 8220 11064 8677 11092
rect 7561 11055 7619 11061
rect 8665 11061 8677 11064
rect 8711 11061 8723 11095
rect 8846 11092 8852 11104
rect 8807 11064 8852 11092
rect 8665 11055 8723 11061
rect 3804 10996 4292 11024
rect 5534 10984 5540 11036
rect 5592 10984 5598 11036
rect 5902 10984 5908 11036
rect 5960 11024 5966 11036
rect 6181 11027 6239 11033
rect 6181 11024 6193 11027
rect 5960 10996 6193 11024
rect 5960 10984 5966 10996
rect 6181 10993 6193 10996
rect 6227 10993 6239 11027
rect 6181 10987 6239 10993
rect 6270 10984 6276 11036
rect 6328 11024 6334 11036
rect 7466 11033 7472 11036
rect 7298 11027 7356 11033
rect 7298 11024 7310 11027
rect 6328 10996 7310 11024
rect 6328 10984 6334 10996
rect 7298 10993 7310 10996
rect 7344 10993 7356 11027
rect 7298 10987 7356 10993
rect 7423 11027 7472 11033
rect 7423 10993 7435 11027
rect 7469 10993 7472 11027
rect 7423 10987 7472 10993
rect 7466 10984 7472 10987
rect 7524 10984 7530 11036
rect 7576 11024 7604 11055
rect 8846 11052 8852 11064
rect 8904 11052 8910 11104
rect 8938 11052 8944 11104
rect 8996 11101 9002 11104
rect 8996 11095 9025 11101
rect 9013 11061 9025 11095
rect 8996 11055 9025 11061
rect 9125 11095 9183 11101
rect 9125 11061 9137 11095
rect 9171 11092 9183 11095
rect 9398 11092 9404 11104
rect 9171 11064 9404 11092
rect 9171 11061 9183 11064
rect 9125 11055 9183 11061
rect 8996 11052 9002 11055
rect 9398 11052 9404 11064
rect 9456 11052 9462 11104
rect 13814 11052 13820 11104
rect 13872 11092 13878 11104
rect 14185 11095 14243 11101
rect 14185 11092 14197 11095
rect 13872 11064 14197 11092
rect 13872 11052 13878 11064
rect 14185 11061 14197 11064
rect 14231 11061 14243 11095
rect 14185 11055 14243 11061
rect 7650 11024 7656 11036
rect 7563 10996 7656 11024
rect 7650 10984 7656 10996
rect 7708 11024 7714 11036
rect 8757 11027 8815 11033
rect 8757 11024 8769 11027
rect 7708 10996 8769 11024
rect 7708 10984 7714 10996
rect 8757 10993 8769 10996
rect 8803 10993 8815 11027
rect 10134 11024 10140 11036
rect 10095 10996 10140 11024
rect 8757 10987 8815 10993
rect 10134 10984 10140 10996
rect 10192 10984 10198 11036
rect 10870 10984 10876 11036
rect 10928 10984 10934 11036
rect 14918 11024 14924 11036
rect 14879 10996 14924 11024
rect 14918 10984 14924 10996
rect 14976 10984 14982 11036
rect 15102 11024 15108 11036
rect 15063 10996 15108 11024
rect 15102 10984 15108 10996
rect 15160 10984 15166 11036
rect 10962 10916 10968 10968
rect 11020 10956 11026 10968
rect 11609 10959 11667 10965
rect 11609 10956 11621 10959
rect 11020 10928 11621 10956
rect 11020 10916 11026 10928
rect 11609 10925 11621 10928
rect 11655 10925 11667 10959
rect 11609 10919 11667 10925
rect 92 10866 15824 10888
rect 92 10814 5242 10866
rect 5294 10814 5306 10866
rect 5358 10814 5370 10866
rect 5422 10814 5434 10866
rect 5486 10814 10514 10866
rect 10566 10814 10578 10866
rect 10630 10814 10642 10866
rect 10694 10814 10706 10866
rect 10758 10814 15824 10866
rect 92 10792 15824 10814
rect 2498 10752 2504 10764
rect 1688 10724 2504 10752
rect 1486 10644 1492 10696
rect 1544 10684 1550 10696
rect 1688 10684 1716 10724
rect 2498 10712 2504 10724
rect 2556 10712 2562 10764
rect 4157 10755 4215 10761
rect 4157 10721 4169 10755
rect 4203 10752 4215 10755
rect 5813 10755 5871 10761
rect 4203 10724 5580 10752
rect 4203 10721 4215 10724
rect 4157 10715 4215 10721
rect 1544 10670 1716 10684
rect 3329 10687 3387 10693
rect 1544 10656 1702 10670
rect 1544 10644 1550 10656
rect 3329 10653 3341 10687
rect 3375 10684 3387 10687
rect 3881 10687 3939 10693
rect 3881 10684 3893 10687
rect 3375 10656 3893 10684
rect 3375 10653 3387 10656
rect 3329 10647 3387 10653
rect 3881 10653 3893 10656
rect 3927 10653 3939 10687
rect 4982 10684 4988 10696
rect 3881 10647 3939 10653
rect 3988 10656 4988 10684
rect 566 10576 572 10628
rect 624 10616 630 10628
rect 937 10619 995 10625
rect 937 10616 949 10619
rect 624 10588 949 10616
rect 624 10576 630 10588
rect 937 10585 949 10588
rect 983 10585 995 10619
rect 937 10579 995 10585
rect 3145 10619 3203 10625
rect 3145 10585 3157 10619
rect 3191 10585 3203 10619
rect 3145 10579 3203 10585
rect 3421 10619 3479 10625
rect 3421 10585 3433 10619
rect 3467 10616 3479 10619
rect 3510 10616 3516 10628
rect 3467 10588 3516 10616
rect 3467 10585 3479 10588
rect 3421 10579 3479 10585
rect 1210 10548 1216 10560
rect 1171 10520 1216 10548
rect 1210 10508 1216 10520
rect 1268 10508 1274 10560
rect 2685 10551 2743 10557
rect 2685 10548 2697 10551
rect 2424 10520 2697 10548
rect 934 10372 940 10424
rect 992 10412 998 10424
rect 2424 10412 2452 10520
rect 2685 10517 2697 10520
rect 2731 10548 2743 10551
rect 3160 10548 3188 10579
rect 3510 10576 3516 10588
rect 3568 10576 3574 10628
rect 3988 10625 4016 10656
rect 4982 10644 4988 10656
rect 5040 10644 5046 10696
rect 5552 10684 5580 10724
rect 5813 10721 5825 10755
rect 5859 10752 5871 10755
rect 5902 10752 5908 10764
rect 5859 10724 5908 10752
rect 5859 10721 5871 10724
rect 5813 10715 5871 10721
rect 5902 10712 5908 10724
rect 5960 10712 5966 10764
rect 7466 10712 7472 10764
rect 7524 10752 7530 10764
rect 9398 10752 9404 10764
rect 7524 10724 8340 10752
rect 9359 10724 9404 10752
rect 7524 10712 7530 10724
rect 6086 10684 6092 10696
rect 5552 10656 6092 10684
rect 6086 10644 6092 10656
rect 6144 10644 6150 10696
rect 7006 10684 7012 10696
rect 6656 10656 7012 10684
rect 3973 10619 4031 10625
rect 3973 10585 3985 10619
rect 4019 10585 4031 10619
rect 3973 10579 4031 10585
rect 4246 10576 4252 10628
rect 4304 10616 4310 10628
rect 4709 10619 4767 10625
rect 4709 10616 4721 10619
rect 4304 10588 4721 10616
rect 4304 10576 4310 10588
rect 4709 10585 4721 10588
rect 4755 10616 4767 10619
rect 4890 10616 4896 10628
rect 4755 10588 4896 10616
rect 4755 10585 4767 10588
rect 4709 10579 4767 10585
rect 4890 10576 4896 10588
rect 4948 10576 4954 10628
rect 5994 10616 6000 10628
rect 5955 10588 6000 10616
rect 5994 10576 6000 10588
rect 6052 10576 6058 10628
rect 6270 10625 6276 10628
rect 6227 10619 6276 10625
rect 6227 10585 6239 10619
rect 6273 10585 6276 10619
rect 6227 10579 6276 10585
rect 6270 10576 6276 10579
rect 6328 10576 6334 10628
rect 6365 10619 6423 10625
rect 6365 10585 6377 10619
rect 6411 10616 6423 10619
rect 6454 10616 6460 10628
rect 6411 10588 6460 10616
rect 6411 10585 6423 10588
rect 6365 10579 6423 10585
rect 6454 10576 6460 10588
rect 6512 10576 6518 10628
rect 6546 10548 6552 10560
rect 2731 10520 6552 10548
rect 2731 10517 2743 10520
rect 2685 10511 2743 10517
rect 6546 10508 6552 10520
rect 6604 10508 6610 10560
rect 3881 10483 3939 10489
rect 3881 10449 3893 10483
rect 3927 10480 3939 10483
rect 6656 10480 6684 10656
rect 7006 10644 7012 10656
rect 7064 10644 7070 10696
rect 8312 10684 8340 10724
rect 9398 10712 9404 10724
rect 9456 10712 9462 10764
rect 9582 10712 9588 10764
rect 9640 10712 9646 10764
rect 11054 10752 11060 10764
rect 10967 10724 11060 10752
rect 11054 10712 11060 10724
rect 11112 10752 11118 10764
rect 11422 10752 11428 10764
rect 11112 10724 11428 10752
rect 11112 10712 11118 10724
rect 11422 10712 11428 10724
rect 11480 10712 11486 10764
rect 8570 10684 8576 10696
rect 8312 10670 8576 10684
rect 8326 10656 8576 10670
rect 8570 10644 8576 10656
rect 8628 10644 8634 10696
rect 9600 10684 9628 10712
rect 11241 10687 11299 10693
rect 11241 10684 11253 10687
rect 9600 10656 11253 10684
rect 11241 10653 11253 10656
rect 11287 10653 11299 10687
rect 11241 10647 11299 10653
rect 9306 10616 9312 10628
rect 9267 10588 9312 10616
rect 9306 10576 9312 10588
rect 9364 10576 9370 10628
rect 9490 10576 9496 10628
rect 9548 10616 9554 10628
rect 9585 10619 9643 10625
rect 9585 10616 9597 10619
rect 9548 10588 9597 10616
rect 9548 10576 9554 10588
rect 9585 10585 9597 10588
rect 9631 10585 9643 10619
rect 9585 10579 9643 10585
rect 9674 10576 9680 10628
rect 9732 10616 9738 10628
rect 9950 10616 9956 10628
rect 9732 10588 9956 10616
rect 9732 10576 9738 10588
rect 9950 10576 9956 10588
rect 10008 10616 10014 10628
rect 10962 10616 10968 10628
rect 10008 10588 10968 10616
rect 10008 10576 10014 10588
rect 10962 10576 10968 10588
rect 11020 10616 11026 10628
rect 11425 10619 11483 10625
rect 11425 10616 11437 10619
rect 11020 10588 11437 10616
rect 11020 10576 11026 10588
rect 11425 10585 11437 10588
rect 11471 10585 11483 10619
rect 11425 10579 11483 10585
rect 11606 10576 11612 10628
rect 11664 10616 11670 10628
rect 12066 10616 12072 10628
rect 11664 10588 12072 10616
rect 11664 10576 11670 10588
rect 12066 10576 12072 10588
rect 12124 10576 12130 10628
rect 12529 10619 12587 10625
rect 12529 10616 12541 10619
rect 12406 10588 12541 10616
rect 6822 10548 6828 10560
rect 6735 10520 6828 10548
rect 6822 10508 6828 10520
rect 6880 10548 6886 10560
rect 7098 10548 7104 10560
rect 6880 10508 6914 10548
rect 7059 10520 7104 10548
rect 7098 10508 7104 10520
rect 7156 10508 7162 10560
rect 7742 10508 7748 10560
rect 7800 10548 7806 10560
rect 11514 10548 11520 10560
rect 7800 10520 11520 10548
rect 7800 10508 7806 10520
rect 11514 10508 11520 10520
rect 11572 10508 11578 10560
rect 11882 10508 11888 10560
rect 11940 10548 11946 10560
rect 12406 10548 12434 10588
rect 12529 10585 12541 10588
rect 12575 10585 12587 10619
rect 12529 10579 12587 10585
rect 15105 10619 15163 10625
rect 15105 10585 15117 10619
rect 15151 10616 15163 10619
rect 15562 10616 15568 10628
rect 15151 10588 15568 10616
rect 15151 10585 15163 10588
rect 15105 10579 15163 10585
rect 15562 10576 15568 10588
rect 15620 10576 15626 10628
rect 11940 10520 12434 10548
rect 11940 10508 11946 10520
rect 3927 10452 6684 10480
rect 3927 10449 3939 10452
rect 3881 10443 3939 10449
rect 3142 10412 3148 10424
rect 992 10384 2452 10412
rect 3103 10384 3148 10412
rect 992 10372 998 10384
rect 3142 10372 3148 10384
rect 3200 10372 3206 10424
rect 4706 10372 4712 10424
rect 4764 10412 4770 10424
rect 4801 10415 4859 10421
rect 4801 10412 4813 10415
rect 4764 10384 4813 10412
rect 4764 10372 4770 10384
rect 4801 10381 4813 10384
rect 4847 10381 4859 10415
rect 4801 10375 4859 10381
rect 4890 10372 4896 10424
rect 4948 10412 4954 10424
rect 6454 10412 6460 10424
rect 4948 10384 6460 10412
rect 4948 10372 4954 10384
rect 6454 10372 6460 10384
rect 6512 10372 6518 10424
rect 6886 10412 6914 10508
rect 9585 10483 9643 10489
rect 8128 10452 8708 10480
rect 8128 10412 8156 10452
rect 6886 10384 8156 10412
rect 8202 10372 8208 10424
rect 8260 10412 8266 10424
rect 8573 10415 8631 10421
rect 8573 10412 8585 10415
rect 8260 10384 8585 10412
rect 8260 10372 8266 10384
rect 8573 10381 8585 10384
rect 8619 10381 8631 10415
rect 8680 10412 8708 10452
rect 9585 10449 9597 10483
rect 9631 10480 9643 10483
rect 10042 10480 10048 10492
rect 9631 10452 10048 10480
rect 9631 10449 9643 10452
rect 9585 10443 9643 10449
rect 10042 10440 10048 10452
rect 10100 10440 10106 10492
rect 11885 10415 11943 10421
rect 11885 10412 11897 10415
rect 8680 10384 11897 10412
rect 8573 10375 8631 10381
rect 11885 10381 11897 10384
rect 11931 10381 11943 10415
rect 12710 10412 12716 10424
rect 12671 10384 12716 10412
rect 11885 10375 11943 10381
rect 12710 10372 12716 10384
rect 12768 10372 12774 10424
rect 14921 10415 14979 10421
rect 14921 10381 14933 10415
rect 14967 10412 14979 10415
rect 15010 10412 15016 10424
rect 14967 10384 15016 10412
rect 14967 10381 14979 10384
rect 14921 10375 14979 10381
rect 15010 10372 15016 10384
rect 15068 10372 15074 10424
rect 92 10322 15824 10344
rect 92 10270 2606 10322
rect 2658 10270 2670 10322
rect 2722 10270 2734 10322
rect 2786 10270 2798 10322
rect 2850 10270 7878 10322
rect 7930 10270 7942 10322
rect 7994 10270 8006 10322
rect 8058 10270 8070 10322
rect 8122 10270 13150 10322
rect 13202 10270 13214 10322
rect 13266 10270 13278 10322
rect 13330 10270 13342 10322
rect 13394 10270 15824 10322
rect 92 10248 15824 10270
rect 661 10211 719 10217
rect 661 10177 673 10211
rect 707 10208 719 10211
rect 1210 10208 1216 10220
rect 707 10180 1216 10208
rect 707 10177 719 10180
rect 661 10171 719 10177
rect 1210 10168 1216 10180
rect 1268 10168 1274 10220
rect 1302 10168 1308 10220
rect 1360 10208 1366 10220
rect 1360 10180 1405 10208
rect 1360 10168 1366 10180
rect 1854 10168 1860 10220
rect 1912 10208 1918 10220
rect 2225 10211 2283 10217
rect 2225 10208 2237 10211
rect 1912 10180 2237 10208
rect 1912 10168 1918 10180
rect 2225 10177 2237 10180
rect 2271 10208 2283 10211
rect 2271 10180 4660 10208
rect 2271 10177 2283 10180
rect 2225 10171 2283 10177
rect 2130 10100 2136 10152
rect 2188 10140 2194 10152
rect 3510 10140 3516 10152
rect 2188 10112 3372 10140
rect 3471 10112 3516 10140
rect 2188 10100 2194 10112
rect 3142 10072 3148 10084
rect 676 10044 3148 10072
rect 676 10013 704 10044
rect 3142 10032 3148 10044
rect 3200 10032 3206 10084
rect 3344 10072 3372 10112
rect 3510 10100 3516 10112
rect 3568 10100 3574 10152
rect 4522 10072 4528 10084
rect 3344 10044 4528 10072
rect 4522 10032 4528 10044
rect 4580 10032 4586 10084
rect 4632 10072 4660 10180
rect 4706 10168 4712 10220
rect 4764 10208 4770 10220
rect 8757 10211 8815 10217
rect 4764 10180 6960 10208
rect 4764 10168 4770 10180
rect 6932 10152 6960 10180
rect 8757 10177 8769 10211
rect 8803 10208 8815 10211
rect 8803 10180 10088 10208
rect 8803 10177 8815 10180
rect 8757 10171 8815 10177
rect 5994 10100 6000 10152
rect 6052 10140 6058 10152
rect 6822 10140 6828 10152
rect 6052 10112 6828 10140
rect 6052 10100 6058 10112
rect 6822 10100 6828 10112
rect 6880 10100 6886 10152
rect 6914 10100 6920 10152
rect 6972 10140 6978 10152
rect 7926 10140 7932 10152
rect 6972 10112 7932 10140
rect 6972 10100 6978 10112
rect 7926 10100 7932 10112
rect 7984 10140 7990 10152
rect 8294 10140 8300 10152
rect 7984 10112 8300 10140
rect 7984 10100 7990 10112
rect 8294 10100 8300 10112
rect 8352 10100 8358 10152
rect 9769 10143 9827 10149
rect 9769 10109 9781 10143
rect 9815 10109 9827 10143
rect 9769 10103 9827 10109
rect 4632 10044 9628 10072
rect 477 10007 535 10013
rect 477 9973 489 10007
rect 523 9973 535 10007
rect 477 9967 535 9973
rect 661 10007 719 10013
rect 661 9973 673 10007
rect 707 9973 719 10007
rect 661 9967 719 9973
rect 1121 10007 1179 10013
rect 1121 9973 1133 10007
rect 1167 9973 1179 10007
rect 1121 9967 1179 9973
rect 1305 10007 1363 10013
rect 1305 9973 1317 10007
rect 1351 10004 1363 10007
rect 3418 10004 3424 10016
rect 1351 9976 3424 10004
rect 1351 9973 1363 9976
rect 1305 9967 1363 9973
rect 492 9936 520 9967
rect 1136 9936 1164 9967
rect 3418 9964 3424 9976
rect 3476 9964 3482 10016
rect 5994 9964 6000 10016
rect 6052 10004 6058 10016
rect 6457 10007 6515 10013
rect 6052 9976 6097 10004
rect 6052 9964 6058 9976
rect 6457 9973 6469 10007
rect 6503 9973 6515 10007
rect 6457 9967 6515 9973
rect 1854 9936 1860 9948
rect 492 9908 1860 9936
rect 1854 9896 1860 9908
rect 1912 9896 1918 9948
rect 2130 9936 2136 9948
rect 2043 9908 2136 9936
rect 2130 9896 2136 9908
rect 2188 9896 2194 9948
rect 3329 9939 3387 9945
rect 3329 9905 3341 9939
rect 3375 9936 3387 9939
rect 3510 9936 3516 9948
rect 3375 9908 3516 9936
rect 3375 9905 3387 9908
rect 3329 9899 3387 9905
rect 3510 9896 3516 9908
rect 3568 9896 3574 9948
rect 5718 9936 5724 9948
rect 4172 9922 4554 9936
rect 4172 9908 4568 9922
rect 5679 9908 5724 9936
rect 1394 9828 1400 9880
rect 1452 9868 1458 9880
rect 2148 9868 2176 9896
rect 1452 9840 2176 9868
rect 1452 9828 1458 9840
rect 2590 9828 2596 9880
rect 2648 9868 2654 9880
rect 4172 9868 4200 9908
rect 2648 9840 4200 9868
rect 4249 9871 4307 9877
rect 2648 9828 2654 9840
rect 4249 9837 4261 9871
rect 4295 9868 4307 9871
rect 4430 9868 4436 9880
rect 4295 9840 4436 9868
rect 4295 9837 4307 9840
rect 4249 9831 4307 9837
rect 4430 9828 4436 9840
rect 4488 9828 4494 9880
rect 4540 9868 4568 9908
rect 5718 9896 5724 9908
rect 5776 9896 5782 9948
rect 6472 9936 6500 9967
rect 6546 9964 6552 10016
rect 6604 10004 6610 10016
rect 8481 10007 8539 10013
rect 8481 10004 8493 10007
rect 6604 9976 8493 10004
rect 6604 9964 6610 9976
rect 8481 9973 8493 9976
rect 8527 9973 8539 10007
rect 8481 9967 8539 9973
rect 9306 9964 9312 10016
rect 9364 10004 9370 10016
rect 9493 10007 9551 10013
rect 9493 10004 9505 10007
rect 9364 9976 9505 10004
rect 9364 9964 9370 9976
rect 9493 9973 9505 9976
rect 9539 9973 9551 10007
rect 9493 9967 9551 9973
rect 6104 9908 6500 9936
rect 7285 9939 7343 9945
rect 5534 9868 5540 9880
rect 4540 9840 5540 9868
rect 5534 9828 5540 9840
rect 5592 9868 5598 9880
rect 6104 9868 6132 9908
rect 7285 9905 7297 9939
rect 7331 9936 7343 9939
rect 7466 9936 7472 9948
rect 7331 9908 7472 9936
rect 7331 9905 7343 9908
rect 7285 9899 7343 9905
rect 7466 9896 7472 9908
rect 7524 9896 7530 9948
rect 8202 9896 8208 9948
rect 8260 9936 8266 9948
rect 8665 9939 8723 9945
rect 8665 9936 8677 9939
rect 8260 9908 8677 9936
rect 8260 9896 8266 9908
rect 8665 9905 8677 9908
rect 8711 9905 8723 9939
rect 9600 9936 9628 10044
rect 9784 10004 9812 10103
rect 10060 10072 10088 10180
rect 10134 10168 10140 10220
rect 10192 10208 10198 10220
rect 10229 10211 10287 10217
rect 10229 10208 10241 10211
rect 10192 10180 10241 10208
rect 10192 10168 10198 10180
rect 10229 10177 10241 10180
rect 10275 10177 10287 10211
rect 10229 10171 10287 10177
rect 14277 10211 14335 10217
rect 14277 10177 14289 10211
rect 14323 10208 14335 10211
rect 14918 10208 14924 10220
rect 14323 10180 14924 10208
rect 14323 10177 14335 10180
rect 14277 10171 14335 10177
rect 14918 10168 14924 10180
rect 14976 10168 14982 10220
rect 10965 10143 11023 10149
rect 10965 10109 10977 10143
rect 11011 10140 11023 10143
rect 12158 10140 12164 10152
rect 11011 10112 12164 10140
rect 11011 10109 11023 10112
rect 10965 10103 11023 10109
rect 12158 10100 12164 10112
rect 12216 10100 12222 10152
rect 12802 10072 12808 10084
rect 10060 10044 12808 10072
rect 10229 10007 10287 10013
rect 10229 10004 10241 10007
rect 9784 9976 10241 10004
rect 10229 9973 10241 9976
rect 10275 9973 10287 10007
rect 10229 9967 10287 9973
rect 10413 10007 10471 10013
rect 10413 9973 10425 10007
rect 10459 9973 10471 10007
rect 11054 10004 11060 10016
rect 11015 9976 11060 10004
rect 10413 9967 10471 9973
rect 9772 9939 9830 9945
rect 9600 9908 9720 9936
rect 8665 9899 8723 9905
rect 5592 9840 6132 9868
rect 5592 9828 5598 9840
rect 6178 9828 6184 9880
rect 6236 9868 6242 9880
rect 7558 9868 7564 9880
rect 6236 9840 7564 9868
rect 6236 9828 6242 9840
rect 7558 9828 7564 9840
rect 7616 9828 7622 9880
rect 7650 9828 7656 9880
rect 7708 9868 7714 9880
rect 9582 9868 9588 9880
rect 7708 9840 9588 9868
rect 7708 9828 7714 9840
rect 9582 9828 9588 9840
rect 9640 9828 9646 9880
rect 9692 9868 9720 9908
rect 9772 9905 9784 9939
rect 9818 9936 9830 9939
rect 9950 9936 9956 9948
rect 9818 9908 9956 9936
rect 9818 9905 9830 9908
rect 9772 9899 9830 9905
rect 9950 9896 9956 9908
rect 10008 9896 10014 9948
rect 10428 9936 10456 9967
rect 11054 9964 11060 9976
rect 11112 9964 11118 10016
rect 11514 10004 11520 10016
rect 11475 9976 11520 10004
rect 11514 9964 11520 9976
rect 11572 9964 11578 10016
rect 12636 10013 12664 10044
rect 12802 10032 12808 10044
rect 12860 10032 12866 10084
rect 12621 10007 12679 10013
rect 12621 9973 12633 10007
rect 12667 10004 12679 10007
rect 14369 10007 14427 10013
rect 12667 9976 12701 10004
rect 12667 9973 12679 9976
rect 12621 9967 12679 9973
rect 14369 9973 14381 10007
rect 14415 10004 14427 10007
rect 14734 10004 14740 10016
rect 14415 9976 14740 10004
rect 14415 9973 14427 9976
rect 14369 9967 14427 9973
rect 14734 9964 14740 9976
rect 14792 9964 14798 10016
rect 11146 9936 11152 9948
rect 10428 9908 11152 9936
rect 10428 9868 10456 9908
rect 11146 9896 11152 9908
rect 11204 9896 11210 9948
rect 14918 9936 14924 9948
rect 14879 9908 14924 9936
rect 14918 9896 14924 9908
rect 14976 9896 14982 9948
rect 15102 9936 15108 9948
rect 15063 9908 15108 9936
rect 15102 9896 15108 9908
rect 15160 9896 15166 9948
rect 9692 9840 10456 9868
rect 11701 9871 11759 9877
rect 11701 9837 11713 9871
rect 11747 9868 11759 9871
rect 11882 9868 11888 9880
rect 11747 9840 11888 9868
rect 11747 9837 11759 9840
rect 11701 9831 11759 9837
rect 11882 9828 11888 9840
rect 11940 9828 11946 9880
rect 12713 9871 12771 9877
rect 12713 9837 12725 9871
rect 12759 9868 12771 9871
rect 12802 9868 12808 9880
rect 12759 9840 12808 9868
rect 12759 9837 12771 9840
rect 12713 9831 12771 9837
rect 12802 9828 12808 9840
rect 12860 9828 12866 9880
rect 92 9778 15824 9800
rect 92 9726 5242 9778
rect 5294 9726 5306 9778
rect 5358 9726 5370 9778
rect 5422 9726 5434 9778
rect 5486 9726 10514 9778
rect 10566 9726 10578 9778
rect 10630 9726 10642 9778
rect 10694 9726 10706 9778
rect 10758 9726 15824 9778
rect 92 9704 15824 9726
rect 1486 9624 1492 9676
rect 1544 9664 1550 9676
rect 2590 9664 2596 9676
rect 1544 9636 2596 9664
rect 1544 9624 1550 9636
rect 934 9596 940 9608
rect 895 9568 940 9596
rect 934 9556 940 9568
rect 992 9556 998 9608
rect 2240 9582 2268 9636
rect 2590 9624 2596 9636
rect 2648 9624 2654 9676
rect 5718 9624 5724 9676
rect 5776 9664 5782 9676
rect 5813 9667 5871 9673
rect 5813 9664 5825 9667
rect 5776 9636 5825 9664
rect 5776 9624 5782 9636
rect 5813 9633 5825 9636
rect 5859 9633 5871 9667
rect 7006 9664 7012 9676
rect 5813 9627 5871 9633
rect 6104 9636 7012 9664
rect 4706 9556 4712 9608
rect 4764 9596 4770 9608
rect 4764 9568 6040 9596
rect 4764 9556 4770 9568
rect 566 9488 572 9540
rect 624 9528 630 9540
rect 1302 9528 1308 9540
rect 624 9500 1308 9528
rect 624 9488 630 9500
rect 1302 9488 1308 9500
rect 1360 9528 1366 9540
rect 1489 9531 1547 9537
rect 1489 9528 1501 9531
rect 1360 9500 1501 9528
rect 1360 9488 1366 9500
rect 1489 9497 1501 9500
rect 1535 9497 1547 9531
rect 4249 9531 4307 9537
rect 4249 9528 4261 9531
rect 1489 9491 1547 9497
rect 3252 9500 4261 9528
rect 3252 9472 3280 9500
rect 4249 9497 4261 9500
rect 4295 9497 4307 9531
rect 4430 9528 4436 9540
rect 4391 9500 4436 9528
rect 4249 9491 4307 9497
rect 4430 9488 4436 9500
rect 4488 9488 4494 9540
rect 6012 9537 6040 9568
rect 6104 9537 6132 9636
rect 7006 9624 7012 9636
rect 7064 9624 7070 9676
rect 7098 9624 7104 9676
rect 7156 9664 7162 9676
rect 7193 9667 7251 9673
rect 7193 9664 7205 9667
rect 7156 9636 7205 9664
rect 7156 9624 7162 9636
rect 7193 9633 7205 9636
rect 7239 9633 7251 9667
rect 12253 9667 12311 9673
rect 7193 9627 7251 9633
rect 7484 9636 7788 9664
rect 6319 9599 6377 9605
rect 6319 9565 6331 9599
rect 6365 9596 6377 9599
rect 6365 9568 6500 9596
rect 6365 9565 6377 9568
rect 6319 9559 6377 9565
rect 5998 9531 6056 9537
rect 5998 9497 6010 9531
rect 6044 9497 6056 9531
rect 5998 9491 6056 9497
rect 6089 9531 6147 9537
rect 6089 9497 6101 9531
rect 6135 9497 6147 9531
rect 6089 9491 6147 9497
rect 6194 9531 6252 9537
rect 6194 9497 6206 9531
rect 6240 9528 6252 9531
rect 6472 9528 6500 9568
rect 6546 9556 6552 9608
rect 6604 9596 6610 9608
rect 7484 9596 7512 9636
rect 6604 9568 7512 9596
rect 7760 9596 7788 9636
rect 12253 9633 12265 9667
rect 12299 9633 12311 9667
rect 12253 9627 12311 9633
rect 14737 9667 14795 9673
rect 14737 9633 14749 9667
rect 14783 9664 14795 9667
rect 14918 9664 14924 9676
rect 14783 9636 14924 9664
rect 14783 9633 14795 9636
rect 14737 9627 14795 9633
rect 12268 9596 12296 9627
rect 14918 9624 14924 9636
rect 14976 9624 14982 9676
rect 7760 9568 12296 9596
rect 6604 9556 6610 9568
rect 6914 9528 6920 9540
rect 6240 9500 6316 9528
rect 6472 9500 6920 9528
rect 6240 9497 6252 9500
rect 6194 9491 6252 9497
rect 750 9460 756 9472
rect 711 9432 756 9460
rect 750 9420 756 9432
rect 808 9420 814 9472
rect 1762 9460 1768 9472
rect 1723 9432 1768 9460
rect 1762 9420 1768 9432
rect 1820 9420 1826 9472
rect 3234 9420 3240 9472
rect 3292 9460 3298 9472
rect 3292 9432 3385 9460
rect 3292 9420 3298 9432
rect 5902 9420 5908 9472
rect 5960 9460 5966 9472
rect 6288 9460 6316 9500
rect 6914 9488 6920 9500
rect 6972 9488 6978 9540
rect 7374 9528 7380 9540
rect 7335 9500 7380 9528
rect 7374 9488 7380 9500
rect 7432 9488 7438 9540
rect 7469 9531 7527 9537
rect 7469 9497 7481 9531
rect 7515 9497 7527 9531
rect 7469 9491 7527 9497
rect 7561 9531 7619 9537
rect 7561 9497 7573 9531
rect 7607 9497 7619 9531
rect 7561 9491 7619 9497
rect 7699 9531 7757 9537
rect 7699 9497 7711 9531
rect 7745 9528 7757 9531
rect 7926 9528 7932 9540
rect 7745 9500 7932 9528
rect 7745 9497 7757 9500
rect 7699 9491 7757 9497
rect 5960 9432 6316 9460
rect 6457 9463 6515 9469
rect 5960 9420 5966 9432
rect 6457 9429 6469 9463
rect 6503 9460 6515 9463
rect 6638 9460 6644 9472
rect 6503 9432 6644 9460
rect 6503 9429 6515 9432
rect 6457 9423 6515 9429
rect 6638 9420 6644 9432
rect 6696 9420 6702 9472
rect 4617 9395 4675 9401
rect 4617 9361 4629 9395
rect 4663 9392 4675 9395
rect 7098 9392 7104 9404
rect 4663 9364 7104 9392
rect 4663 9361 4675 9364
rect 4617 9355 4675 9361
rect 7098 9352 7104 9364
rect 7156 9352 7162 9404
rect 4522 9284 4528 9336
rect 4580 9324 4586 9336
rect 6914 9324 6920 9336
rect 4580 9296 6920 9324
rect 4580 9284 4586 9296
rect 6914 9284 6920 9296
rect 6972 9284 6978 9336
rect 7484 9324 7512 9491
rect 7576 9404 7604 9491
rect 7926 9488 7932 9500
rect 7984 9488 7990 9540
rect 8297 9531 8355 9537
rect 8297 9497 8309 9531
rect 8343 9528 8355 9531
rect 8386 9528 8392 9540
rect 8343 9500 8392 9528
rect 8343 9497 8355 9500
rect 8297 9491 8355 9497
rect 8386 9488 8392 9500
rect 8444 9488 8450 9540
rect 8481 9531 8539 9537
rect 8481 9497 8493 9531
rect 8527 9528 8539 9531
rect 8662 9528 8668 9540
rect 8527 9500 8668 9528
rect 8527 9497 8539 9500
rect 8481 9491 8539 9497
rect 8662 9488 8668 9500
rect 8720 9488 8726 9540
rect 9122 9528 9128 9540
rect 9083 9500 9128 9528
rect 9122 9488 9128 9500
rect 9180 9488 9186 9540
rect 10134 9528 10140 9540
rect 10095 9500 10140 9528
rect 10134 9488 10140 9500
rect 10192 9488 10198 9540
rect 11425 9531 11483 9537
rect 11425 9497 11437 9531
rect 11471 9497 11483 9531
rect 11425 9491 11483 9497
rect 7837 9463 7895 9469
rect 7837 9429 7849 9463
rect 7883 9460 7895 9463
rect 8202 9460 8208 9472
rect 7883 9432 8208 9460
rect 7883 9429 7895 9432
rect 7837 9423 7895 9429
rect 8202 9420 8208 9432
rect 8260 9420 8266 9472
rect 8570 9460 8576 9472
rect 8312 9432 8576 9460
rect 7558 9352 7564 9404
rect 7616 9352 7622 9404
rect 8312 9401 8340 9432
rect 8570 9420 8576 9432
rect 8628 9420 8634 9472
rect 11440 9460 11468 9491
rect 11514 9488 11520 9540
rect 11572 9528 11578 9540
rect 11790 9528 11796 9540
rect 11572 9500 11617 9528
rect 11751 9500 11796 9528
rect 11572 9488 11578 9500
rect 11790 9488 11796 9500
rect 11848 9488 11854 9540
rect 12250 9488 12256 9540
rect 12308 9528 12314 9540
rect 12434 9537 12440 9540
rect 12308 9500 12353 9528
rect 12308 9488 12314 9500
rect 12430 9491 12440 9537
rect 12492 9528 12498 9540
rect 12492 9500 12530 9528
rect 12434 9488 12440 9491
rect 12492 9488 12498 9500
rect 12618 9488 12624 9540
rect 12676 9528 12682 9540
rect 12897 9531 12955 9537
rect 12897 9528 12909 9531
rect 12676 9500 12909 9528
rect 12676 9488 12682 9500
rect 12897 9497 12909 9500
rect 12943 9497 12955 9531
rect 12897 9491 12955 9497
rect 13081 9531 13139 9537
rect 13081 9497 13093 9531
rect 13127 9528 13139 9531
rect 13630 9528 13636 9540
rect 13127 9500 13636 9528
rect 13127 9497 13139 9500
rect 13081 9491 13139 9497
rect 13630 9488 13636 9500
rect 13688 9488 13694 9540
rect 13906 9488 13912 9540
rect 13964 9528 13970 9540
rect 14001 9531 14059 9537
rect 14001 9528 14013 9531
rect 13964 9500 14013 9528
rect 13964 9488 13970 9500
rect 14001 9497 14013 9500
rect 14047 9497 14059 9531
rect 14642 9528 14648 9540
rect 14603 9500 14648 9528
rect 14001 9491 14059 9497
rect 14642 9488 14648 9500
rect 14700 9488 14706 9540
rect 12066 9460 12072 9472
rect 11440 9432 12072 9460
rect 12066 9420 12072 9432
rect 12124 9420 12130 9472
rect 8297 9395 8355 9401
rect 8297 9361 8309 9395
rect 8343 9361 8355 9395
rect 8297 9355 8355 9361
rect 8386 9352 8392 9404
rect 8444 9392 8450 9404
rect 14458 9392 14464 9404
rect 8444 9364 14464 9392
rect 8444 9352 8450 9364
rect 14458 9352 14464 9364
rect 14516 9392 14522 9404
rect 14826 9392 14832 9404
rect 14516 9364 14832 9392
rect 14516 9352 14522 9364
rect 14826 9352 14832 9364
rect 14884 9352 14890 9404
rect 7650 9324 7656 9336
rect 7484 9296 7656 9324
rect 7650 9284 7656 9296
rect 7708 9284 7714 9336
rect 9030 9324 9036 9336
rect 8991 9296 9036 9324
rect 9030 9284 9036 9296
rect 9088 9284 9094 9336
rect 10042 9324 10048 9336
rect 10003 9296 10048 9324
rect 10042 9284 10048 9296
rect 10100 9284 10106 9336
rect 11241 9327 11299 9333
rect 11241 9293 11253 9327
rect 11287 9324 11299 9327
rect 11422 9324 11428 9336
rect 11287 9296 11428 9324
rect 11287 9293 11299 9296
rect 11241 9287 11299 9293
rect 11422 9284 11428 9296
rect 11480 9284 11486 9336
rect 11701 9327 11759 9333
rect 11701 9293 11713 9327
rect 11747 9324 11759 9327
rect 12250 9324 12256 9336
rect 11747 9296 12256 9324
rect 11747 9293 11759 9296
rect 11701 9287 11759 9293
rect 12250 9284 12256 9296
rect 12308 9284 12314 9336
rect 12526 9284 12532 9336
rect 12584 9324 12590 9336
rect 13081 9327 13139 9333
rect 13081 9324 13093 9327
rect 12584 9296 13093 9324
rect 12584 9284 12590 9296
rect 13081 9293 13093 9296
rect 13127 9293 13139 9327
rect 14090 9324 14096 9336
rect 14051 9296 14096 9324
rect 13081 9287 13139 9293
rect 14090 9284 14096 9296
rect 14148 9284 14154 9336
rect 92 9234 15824 9256
rect 92 9182 2606 9234
rect 2658 9182 2670 9234
rect 2722 9182 2734 9234
rect 2786 9182 2798 9234
rect 2850 9182 7878 9234
rect 7930 9182 7942 9234
rect 7994 9182 8006 9234
rect 8058 9182 8070 9234
rect 8122 9182 13150 9234
rect 13202 9182 13214 9234
rect 13266 9182 13278 9234
rect 13330 9182 13342 9234
rect 13394 9182 15824 9234
rect 92 9160 15824 9182
rect 1857 9123 1915 9129
rect 1857 9089 1869 9123
rect 1903 9120 1915 9123
rect 4338 9120 4344 9132
rect 1903 9092 4344 9120
rect 1903 9089 1915 9092
rect 1857 9083 1915 9089
rect 4338 9080 4344 9092
rect 4396 9080 4402 9132
rect 6454 9080 6460 9132
rect 6512 9120 6518 9132
rect 7469 9123 7527 9129
rect 7469 9120 7481 9123
rect 6512 9092 7481 9120
rect 6512 9080 6518 9092
rect 7469 9089 7481 9092
rect 7515 9089 7527 9123
rect 7469 9083 7527 9089
rect 2038 9012 2044 9064
rect 2096 9052 2102 9064
rect 3237 9055 3295 9061
rect 3237 9052 3249 9055
rect 2096 9024 3249 9052
rect 2096 9012 2102 9024
rect 3237 9021 3249 9024
rect 3283 9021 3295 9055
rect 3510 9052 3516 9064
rect 3237 9015 3295 9021
rect 3344 9024 3516 9052
rect 1302 8944 1308 8996
rect 1360 8984 1366 8996
rect 2498 8984 2504 8996
rect 1360 8956 2504 8984
rect 1360 8944 1366 8956
rect 2498 8944 2504 8956
rect 2556 8944 2562 8996
rect 3344 8984 3372 9024
rect 3510 9012 3516 9024
rect 3568 9012 3574 9064
rect 6914 9012 6920 9064
rect 6972 9052 6978 9064
rect 8662 9052 8668 9064
rect 6972 9024 8668 9052
rect 6972 9012 6978 9024
rect 8662 9012 8668 9024
rect 8720 9012 8726 9064
rect 4709 8987 4767 8993
rect 2976 8956 3372 8984
rect 3436 8956 4476 8984
rect 2976 8928 3004 8956
rect 937 8919 995 8925
rect 937 8885 949 8919
rect 983 8916 995 8919
rect 2133 8919 2191 8925
rect 983 8888 2084 8916
rect 983 8885 995 8888
rect 937 8879 995 8885
rect 750 8848 756 8860
rect 711 8820 756 8848
rect 750 8808 756 8820
rect 808 8808 814 8860
rect 1854 8848 1860 8860
rect 1815 8820 1860 8848
rect 1854 8808 1860 8820
rect 1912 8808 1918 8860
rect 2056 8848 2084 8888
rect 2133 8885 2145 8919
rect 2179 8916 2191 8919
rect 2958 8916 2964 8928
rect 2179 8888 2964 8916
rect 2179 8885 2191 8888
rect 2133 8879 2191 8885
rect 2958 8876 2964 8888
rect 3016 8876 3022 8928
rect 3234 8916 3240 8928
rect 3195 8888 3240 8916
rect 3234 8876 3240 8888
rect 3292 8876 3298 8928
rect 3436 8925 3464 8956
rect 4448 8928 4476 8956
rect 4709 8953 4721 8987
rect 4755 8984 4767 8987
rect 6641 8987 6699 8993
rect 6641 8984 6653 8987
rect 4755 8956 6653 8984
rect 4755 8953 4767 8956
rect 4709 8947 4767 8953
rect 6641 8953 6653 8956
rect 6687 8953 6699 8987
rect 6641 8947 6699 8953
rect 9858 8944 9864 8996
rect 9916 8984 9922 8996
rect 10413 8987 10471 8993
rect 10413 8984 10425 8987
rect 9916 8956 10425 8984
rect 9916 8944 9922 8956
rect 10413 8953 10425 8956
rect 10459 8953 10471 8987
rect 10413 8947 10471 8953
rect 10781 8987 10839 8993
rect 10781 8953 10793 8987
rect 10827 8984 10839 8987
rect 11054 8984 11060 8996
rect 10827 8956 11060 8984
rect 10827 8953 10839 8956
rect 10781 8947 10839 8953
rect 11054 8944 11060 8956
rect 11112 8944 11118 8996
rect 11532 8956 12112 8984
rect 3421 8919 3479 8925
rect 3421 8885 3433 8919
rect 3467 8885 3479 8919
rect 3421 8879 3479 8885
rect 3510 8876 3516 8928
rect 3568 8916 3574 8928
rect 4246 8925 4252 8928
rect 4065 8919 4123 8925
rect 3568 8888 3613 8916
rect 3568 8876 3574 8888
rect 4065 8885 4077 8919
rect 4111 8885 4123 8919
rect 4065 8879 4123 8885
rect 4223 8919 4252 8925
rect 4223 8885 4235 8919
rect 4223 8879 4252 8885
rect 3252 8848 3280 8876
rect 4080 8848 4108 8879
rect 4246 8876 4252 8879
rect 4304 8876 4310 8928
rect 4430 8916 4436 8928
rect 4391 8888 4436 8916
rect 4430 8876 4436 8888
rect 4488 8876 4494 8928
rect 4525 8919 4583 8925
rect 4525 8885 4537 8919
rect 4571 8916 4583 8919
rect 4614 8916 4620 8928
rect 4571 8888 4620 8916
rect 4571 8885 4583 8888
rect 4525 8879 4583 8885
rect 4614 8876 4620 8888
rect 4672 8876 4678 8928
rect 5534 8876 5540 8928
rect 5592 8876 5598 8928
rect 6914 8876 6920 8928
rect 6972 8916 6978 8928
rect 6972 8888 7017 8916
rect 6972 8876 6978 8888
rect 7190 8876 7196 8928
rect 7248 8916 7254 8928
rect 7377 8919 7435 8925
rect 7377 8916 7389 8919
rect 7248 8888 7389 8916
rect 7248 8876 7254 8888
rect 7377 8885 7389 8888
rect 7423 8885 7435 8919
rect 7377 8879 7435 8885
rect 8757 8919 8815 8925
rect 8757 8885 8769 8919
rect 8803 8916 8815 8919
rect 9306 8916 9312 8928
rect 8803 8888 9312 8916
rect 8803 8885 8815 8888
rect 8757 8879 8815 8885
rect 9306 8876 9312 8888
rect 9364 8876 9370 8928
rect 9398 8876 9404 8928
rect 9456 8916 9462 8928
rect 9456 8888 9501 8916
rect 9456 8876 9462 8888
rect 2056 8820 3280 8848
rect 3344 8820 4108 8848
rect 2041 8783 2099 8789
rect 2041 8749 2053 8783
rect 2087 8780 2099 8783
rect 3344 8780 3372 8820
rect 2087 8752 3372 8780
rect 4080 8780 4108 8820
rect 4341 8851 4399 8857
rect 4341 8817 4353 8851
rect 4387 8848 4399 8851
rect 4982 8848 4988 8860
rect 4387 8820 4988 8848
rect 4387 8817 4399 8820
rect 4341 8811 4399 8817
rect 4982 8808 4988 8820
rect 5040 8848 5046 8860
rect 5040 8820 5304 8848
rect 5040 8808 5046 8820
rect 4614 8780 4620 8792
rect 4080 8752 4620 8780
rect 2087 8749 2099 8752
rect 2041 8743 2099 8749
rect 4614 8740 4620 8752
rect 4672 8780 4678 8792
rect 5169 8783 5227 8789
rect 5169 8780 5181 8783
rect 4672 8752 5181 8780
rect 4672 8740 4678 8752
rect 5169 8749 5181 8752
rect 5215 8749 5227 8783
rect 5276 8780 5304 8820
rect 7208 8780 7236 8876
rect 5276 8752 7236 8780
rect 8665 8783 8723 8789
rect 5169 8743 5227 8749
rect 8665 8749 8677 8783
rect 8711 8780 8723 8783
rect 8754 8780 8760 8792
rect 8711 8752 8760 8780
rect 8711 8749 8723 8752
rect 8665 8743 8723 8749
rect 8754 8740 8760 8752
rect 8812 8740 8818 8792
rect 9309 8783 9367 8789
rect 9309 8749 9321 8783
rect 9355 8780 9367 8783
rect 9490 8780 9496 8792
rect 9355 8752 9496 8780
rect 9355 8749 9367 8752
rect 9309 8743 9367 8749
rect 9490 8740 9496 8752
rect 9548 8740 9554 8792
rect 9950 8740 9956 8792
rect 10008 8780 10014 8792
rect 10870 8780 10876 8792
rect 10008 8752 10876 8780
rect 10008 8740 10014 8752
rect 10870 8740 10876 8752
rect 10928 8780 10934 8792
rect 11164 8780 11192 8834
rect 11532 8780 11560 8956
rect 12084 8916 12112 8956
rect 12250 8944 12256 8996
rect 12308 8984 12314 8996
rect 14185 8987 14243 8993
rect 14185 8984 14197 8987
rect 12308 8956 14197 8984
rect 12308 8944 12314 8956
rect 14185 8953 14197 8956
rect 14231 8953 14243 8987
rect 14185 8947 14243 8953
rect 13446 8916 13452 8928
rect 12084 8888 13452 8916
rect 13446 8876 13452 8888
rect 13504 8876 13510 8928
rect 13909 8919 13967 8925
rect 13909 8885 13921 8919
rect 13955 8885 13967 8919
rect 13909 8879 13967 8885
rect 14001 8919 14059 8925
rect 14001 8885 14013 8919
rect 14047 8885 14059 8919
rect 14001 8879 14059 8885
rect 12066 8808 12072 8860
rect 12124 8848 12130 8860
rect 13725 8851 13783 8857
rect 13725 8848 13737 8851
rect 12124 8820 13737 8848
rect 12124 8808 12130 8820
rect 13725 8817 13737 8820
rect 13771 8817 13783 8851
rect 13725 8811 13783 8817
rect 10928 8752 11560 8780
rect 10928 8740 10934 8752
rect 11974 8740 11980 8792
rect 12032 8780 12038 8792
rect 12207 8783 12265 8789
rect 12207 8780 12219 8783
rect 12032 8752 12219 8780
rect 12032 8740 12038 8752
rect 12207 8749 12219 8752
rect 12253 8749 12265 8783
rect 13924 8780 13952 8879
rect 14016 8848 14044 8879
rect 14090 8876 14096 8928
rect 14148 8916 14154 8928
rect 14277 8919 14335 8925
rect 14277 8916 14289 8919
rect 14148 8888 14289 8916
rect 14148 8876 14154 8888
rect 14277 8885 14289 8888
rect 14323 8885 14335 8919
rect 14277 8879 14335 8885
rect 14182 8848 14188 8860
rect 14016 8820 14188 8848
rect 14182 8808 14188 8820
rect 14240 8808 14246 8860
rect 14918 8848 14924 8860
rect 14879 8820 14924 8848
rect 14918 8808 14924 8820
rect 14976 8808 14982 8860
rect 15102 8848 15108 8860
rect 15063 8820 15108 8848
rect 15102 8808 15108 8820
rect 15160 8808 15166 8860
rect 14274 8780 14280 8792
rect 13924 8752 14280 8780
rect 12207 8743 12265 8749
rect 14274 8740 14280 8752
rect 14332 8740 14338 8792
rect 92 8690 15824 8712
rect 92 8638 5242 8690
rect 5294 8638 5306 8690
rect 5358 8638 5370 8690
rect 5422 8638 5434 8690
rect 5486 8638 10514 8690
rect 10566 8638 10578 8690
rect 10630 8638 10642 8690
rect 10694 8638 10706 8690
rect 10758 8638 15824 8690
rect 92 8616 15824 8638
rect 658 8576 664 8588
rect 571 8548 664 8576
rect 658 8536 664 8548
rect 716 8576 722 8588
rect 716 8548 1900 8576
rect 716 8536 722 8548
rect 1872 8520 1900 8548
rect 5902 8536 5908 8588
rect 5960 8576 5966 8588
rect 9306 8576 9312 8588
rect 5960 8548 8340 8576
rect 9267 8548 9312 8576
rect 5960 8536 5966 8548
rect 1486 8468 1492 8520
rect 1544 8468 1550 8520
rect 1854 8468 1860 8520
rect 1912 8508 1918 8520
rect 2869 8511 2927 8517
rect 2869 8508 2881 8511
rect 1912 8480 2881 8508
rect 1912 8468 1918 8480
rect 2869 8477 2881 8480
rect 2915 8477 2927 8511
rect 2869 8471 2927 8477
rect 3053 8511 3111 8517
rect 3053 8477 3065 8511
rect 3099 8508 3111 8511
rect 4614 8508 4620 8520
rect 3099 8480 4620 8508
rect 3099 8477 3111 8480
rect 3053 8471 3111 8477
rect 4614 8468 4620 8480
rect 4672 8468 4678 8520
rect 5534 8468 5540 8520
rect 5592 8508 5598 8520
rect 5592 8480 6210 8508
rect 5592 8468 5598 8480
rect 7098 8468 7104 8520
rect 7156 8508 7162 8520
rect 7156 8480 8156 8508
rect 7156 8468 7162 8480
rect 2409 8443 2467 8449
rect 2409 8409 2421 8443
rect 2455 8440 2467 8443
rect 2498 8440 2504 8452
rect 2455 8412 2504 8440
rect 2455 8409 2467 8412
rect 2409 8403 2467 8409
rect 2498 8400 2504 8412
rect 2556 8400 2562 8452
rect 4338 8400 4344 8452
rect 4396 8449 4402 8452
rect 4396 8443 4445 8449
rect 4396 8409 4399 8443
rect 4433 8409 4445 8443
rect 4396 8403 4445 8409
rect 4525 8443 4583 8449
rect 4525 8409 4537 8443
rect 4571 8409 4583 8443
rect 4706 8440 4712 8452
rect 4667 8412 4712 8440
rect 4525 8403 4583 8409
rect 4396 8400 4402 8403
rect 2133 8375 2191 8381
rect 2133 8341 2145 8375
rect 2179 8372 2191 8375
rect 4154 8372 4160 8384
rect 2179 8344 4160 8372
rect 2179 8341 2191 8344
rect 2133 8335 2191 8341
rect 4154 8332 4160 8344
rect 4212 8332 4218 8384
rect 4249 8375 4307 8381
rect 4249 8341 4261 8375
rect 4295 8341 4307 8375
rect 4540 8372 4568 8403
rect 4706 8400 4712 8412
rect 4764 8400 4770 8452
rect 4982 8440 4988 8452
rect 4816 8412 4988 8440
rect 4816 8372 4844 8412
rect 4982 8400 4988 8412
rect 5040 8400 5046 8452
rect 8128 8449 8156 8480
rect 8312 8449 8340 8548
rect 9306 8536 9312 8548
rect 9364 8536 9370 8588
rect 11149 8579 11207 8585
rect 11149 8545 11161 8579
rect 11195 8576 11207 8579
rect 11790 8576 11796 8588
rect 11195 8548 11796 8576
rect 11195 8545 11207 8548
rect 11149 8539 11207 8545
rect 11790 8536 11796 8548
rect 11848 8576 11854 8588
rect 11848 8548 12112 8576
rect 11848 8536 11854 8548
rect 11974 8508 11980 8520
rect 11256 8480 11980 8508
rect 8113 8443 8171 8449
rect 8113 8409 8125 8443
rect 8159 8409 8171 8443
rect 8113 8403 8171 8409
rect 8297 8443 8355 8449
rect 8297 8409 8309 8443
rect 8343 8409 8355 8443
rect 8297 8403 8355 8409
rect 9493 8443 9551 8449
rect 9493 8409 9505 8443
rect 9539 8440 9551 8443
rect 9582 8440 9588 8452
rect 9539 8412 9588 8440
rect 9539 8409 9551 8412
rect 9493 8403 9551 8409
rect 9582 8400 9588 8412
rect 9640 8400 9646 8452
rect 9677 8443 9735 8449
rect 9677 8409 9689 8443
rect 9723 8440 9735 8443
rect 9953 8443 10011 8449
rect 9723 8412 9904 8440
rect 9723 8409 9735 8412
rect 9677 8403 9735 8409
rect 4540 8344 4844 8372
rect 4893 8375 4951 8381
rect 4249 8335 4307 8341
rect 4893 8341 4905 8375
rect 4939 8372 4951 8375
rect 7377 8375 7435 8381
rect 7377 8372 7389 8375
rect 4939 8344 7389 8372
rect 4939 8341 4951 8344
rect 4893 8335 4951 8341
rect 7377 8341 7389 8344
rect 7423 8341 7435 8375
rect 7650 8372 7656 8384
rect 7611 8344 7656 8372
rect 7377 8335 7435 8341
rect 3234 8304 3240 8316
rect 3195 8276 3240 8304
rect 3234 8264 3240 8276
rect 3292 8264 3298 8316
rect 3326 8264 3332 8316
rect 3384 8304 3390 8316
rect 4264 8304 4292 8335
rect 7650 8332 7656 8344
rect 7708 8332 7714 8384
rect 9766 8372 9772 8384
rect 9727 8344 9772 8372
rect 9766 8332 9772 8344
rect 9824 8332 9830 8384
rect 9876 8372 9904 8412
rect 9953 8409 9965 8443
rect 9999 8440 10011 8443
rect 10042 8440 10048 8452
rect 9999 8412 10048 8440
rect 9999 8409 10011 8412
rect 9953 8403 10011 8409
rect 10042 8400 10048 8412
rect 10100 8440 10106 8452
rect 10870 8440 10876 8452
rect 10100 8412 10876 8440
rect 10100 8400 10106 8412
rect 10870 8400 10876 8412
rect 10928 8400 10934 8452
rect 11256 8449 11284 8480
rect 11974 8468 11980 8480
rect 12032 8468 12038 8520
rect 12084 8517 12112 8548
rect 12069 8511 12127 8517
rect 12069 8477 12081 8511
rect 12115 8477 12127 8511
rect 12069 8471 12127 8477
rect 13446 8468 13452 8520
rect 13504 8468 13510 8520
rect 11241 8443 11299 8449
rect 11241 8409 11253 8443
rect 11287 8409 11299 8443
rect 11241 8403 11299 8409
rect 11330 8400 11336 8452
rect 11388 8440 11394 8452
rect 11885 8443 11943 8449
rect 11885 8440 11897 8443
rect 11388 8412 11897 8440
rect 11388 8400 11394 8412
rect 11885 8409 11897 8412
rect 11931 8409 11943 8443
rect 12250 8440 12256 8452
rect 12211 8412 12256 8440
rect 11885 8403 11943 8409
rect 12250 8400 12256 8412
rect 12308 8400 12314 8452
rect 12710 8440 12716 8452
rect 12671 8412 12716 8440
rect 12710 8400 12716 8412
rect 12768 8400 12774 8452
rect 11146 8372 11152 8384
rect 9876 8344 11152 8372
rect 11146 8332 11152 8344
rect 11204 8332 11210 8384
rect 11440 8344 12434 8372
rect 3384 8276 5948 8304
rect 3384 8264 3390 8276
rect 5920 8245 5948 8276
rect 8294 8264 8300 8316
rect 8352 8304 8358 8316
rect 9030 8304 9036 8316
rect 8352 8276 9036 8304
rect 8352 8264 8358 8276
rect 9030 8264 9036 8276
rect 9088 8264 9094 8316
rect 9585 8307 9643 8313
rect 9585 8273 9597 8307
rect 9631 8304 9643 8307
rect 9631 8276 9720 8304
rect 9631 8273 9643 8276
rect 9585 8267 9643 8273
rect 9692 8248 9720 8276
rect 9858 8264 9864 8316
rect 9916 8304 9922 8316
rect 11440 8304 11468 8344
rect 9916 8276 11468 8304
rect 9916 8264 9922 8276
rect 11514 8264 11520 8316
rect 11572 8304 11578 8316
rect 11701 8307 11759 8313
rect 11701 8304 11713 8307
rect 11572 8276 11713 8304
rect 11572 8264 11578 8276
rect 11701 8273 11713 8276
rect 11747 8273 11759 8307
rect 12406 8304 12434 8344
rect 12728 8304 12756 8400
rect 12894 8332 12900 8384
rect 12952 8372 12958 8384
rect 13081 8375 13139 8381
rect 13081 8372 13093 8375
rect 12952 8344 13093 8372
rect 12952 8332 12958 8344
rect 13081 8341 13093 8344
rect 13127 8341 13139 8375
rect 13081 8335 13139 8341
rect 12406 8276 12756 8304
rect 11701 8267 11759 8273
rect 5905 8239 5963 8245
rect 5905 8205 5917 8239
rect 5951 8236 5963 8239
rect 5994 8236 6000 8248
rect 5951 8208 6000 8236
rect 5951 8205 5963 8208
rect 5905 8199 5963 8205
rect 5994 8196 6000 8208
rect 6052 8196 6058 8248
rect 7190 8196 7196 8248
rect 7248 8236 7254 8248
rect 8205 8239 8263 8245
rect 8205 8236 8217 8239
rect 7248 8208 8217 8236
rect 7248 8196 7254 8208
rect 8205 8205 8217 8208
rect 8251 8205 8263 8239
rect 8205 8199 8263 8205
rect 9674 8196 9680 8248
rect 9732 8196 9738 8248
rect 13906 8196 13912 8248
rect 13964 8236 13970 8248
rect 14507 8239 14565 8245
rect 14507 8236 14519 8239
rect 13964 8208 14519 8236
rect 13964 8196 13970 8208
rect 14507 8205 14519 8208
rect 14553 8205 14565 8239
rect 14507 8199 14565 8205
rect 92 8146 15824 8168
rect 92 8094 2606 8146
rect 2658 8094 2670 8146
rect 2722 8094 2734 8146
rect 2786 8094 2798 8146
rect 2850 8094 7878 8146
rect 7930 8094 7942 8146
rect 7994 8094 8006 8146
rect 8058 8094 8070 8146
rect 8122 8094 13150 8146
rect 13202 8094 13214 8146
rect 13266 8094 13278 8146
rect 13330 8094 13342 8146
rect 13394 8094 15824 8146
rect 92 8072 15824 8094
rect 2041 8035 2099 8041
rect 2041 8001 2053 8035
rect 2087 8032 2099 8035
rect 2087 8004 2774 8032
rect 2087 8001 2099 8004
rect 2041 7995 2099 8001
rect 1118 7924 1124 7976
rect 1176 7964 1182 7976
rect 1213 7967 1271 7973
rect 1213 7964 1225 7967
rect 1176 7936 1225 7964
rect 1176 7924 1182 7936
rect 1213 7933 1225 7936
rect 1259 7933 1271 7967
rect 2746 7964 2774 8004
rect 4154 7992 4160 8044
rect 4212 8032 4218 8044
rect 4249 8035 4307 8041
rect 4249 8032 4261 8035
rect 4212 8004 4261 8032
rect 4212 7992 4218 8004
rect 4249 8001 4261 8004
rect 4295 8032 4307 8035
rect 5902 8032 5908 8044
rect 4295 8004 5908 8032
rect 4295 8001 4307 8004
rect 4249 7995 4307 8001
rect 5902 7992 5908 8004
rect 5960 7992 5966 8044
rect 7650 7992 7656 8044
rect 7708 8032 7714 8044
rect 9858 8032 9864 8044
rect 7708 8004 9864 8032
rect 7708 7992 7714 8004
rect 2746 7936 4384 7964
rect 1213 7927 1271 7933
rect 4356 7896 4384 7936
rect 4982 7924 4988 7976
rect 5040 7964 5046 7976
rect 5353 7967 5411 7973
rect 5353 7964 5365 7967
rect 5040 7936 5365 7964
rect 5040 7924 5046 7936
rect 5353 7933 5365 7936
rect 5399 7933 5411 7967
rect 8478 7964 8484 7976
rect 5353 7927 5411 7933
rect 5460 7936 8484 7964
rect 5460 7896 5488 7936
rect 8478 7924 8484 7936
rect 8536 7924 8542 7976
rect 5902 7896 5908 7908
rect 4356 7868 5488 7896
rect 5863 7868 5908 7896
rect 5902 7856 5908 7868
rect 5960 7856 5966 7908
rect 7190 7856 7196 7908
rect 7248 7896 7254 7908
rect 7285 7899 7343 7905
rect 7285 7896 7297 7899
rect 7248 7868 7297 7896
rect 7248 7856 7254 7868
rect 7285 7865 7297 7868
rect 7331 7865 7343 7899
rect 8588 7896 8616 8004
rect 9858 7992 9864 8004
rect 9916 7992 9922 8044
rect 10134 7992 10140 8044
rect 10192 8032 10198 8044
rect 10229 8035 10287 8041
rect 10229 8032 10241 8035
rect 10192 8004 10241 8032
rect 10192 7992 10198 8004
rect 10229 8001 10241 8004
rect 10275 8001 10287 8035
rect 11054 8032 11060 8044
rect 11015 8004 11060 8032
rect 10229 7995 10287 8001
rect 11054 7992 11060 8004
rect 11112 7992 11118 8044
rect 11330 7992 11336 8044
rect 11388 8032 11394 8044
rect 11698 8032 11704 8044
rect 11388 8004 11704 8032
rect 11388 7992 11394 8004
rect 11698 7992 11704 8004
rect 11756 7992 11762 8044
rect 12805 8035 12863 8041
rect 12805 8001 12817 8035
rect 12851 8032 12863 8035
rect 12894 8032 12900 8044
rect 12851 8004 12900 8032
rect 12851 8001 12863 8004
rect 12805 7995 12863 8001
rect 12894 7992 12900 8004
rect 12952 7992 12958 8044
rect 11238 7924 11244 7976
rect 11296 7964 11302 7976
rect 12250 7964 12256 7976
rect 11296 7936 12256 7964
rect 11296 7924 11302 7936
rect 12250 7924 12256 7936
rect 12308 7964 12314 7976
rect 14737 7967 14795 7973
rect 14737 7964 14749 7967
rect 12308 7936 14749 7964
rect 12308 7924 12314 7936
rect 14737 7933 14749 7936
rect 14783 7933 14795 7967
rect 14737 7927 14795 7933
rect 8754 7896 8760 7908
rect 7285 7859 7343 7865
rect 8496 7868 8616 7896
rect 8715 7868 8760 7896
rect 658 7828 664 7840
rect 619 7800 664 7828
rect 658 7788 664 7800
rect 716 7788 722 7840
rect 1397 7831 1455 7837
rect 1397 7797 1409 7831
rect 1443 7828 1455 7831
rect 2317 7831 2375 7837
rect 1443 7800 2268 7828
rect 1443 7797 1455 7800
rect 1397 7791 1455 7797
rect 474 7760 480 7772
rect 435 7732 480 7760
rect 474 7720 480 7732
rect 532 7720 538 7772
rect 1581 7763 1639 7769
rect 1581 7729 1593 7763
rect 1627 7760 1639 7763
rect 2041 7763 2099 7769
rect 2041 7760 2053 7763
rect 1627 7732 2053 7760
rect 1627 7729 1639 7732
rect 1581 7723 1639 7729
rect 2041 7729 2053 7732
rect 2087 7729 2099 7763
rect 2041 7723 2099 7729
rect 566 7652 572 7704
rect 624 7692 630 7704
rect 1596 7692 1624 7723
rect 2240 7701 2268 7800
rect 2317 7797 2329 7831
rect 2363 7797 2375 7831
rect 3418 7828 3424 7840
rect 3379 7800 3424 7828
rect 2317 7791 2375 7797
rect 2332 7760 2360 7791
rect 3418 7788 3424 7800
rect 3476 7788 3482 7840
rect 4062 7828 4068 7840
rect 4023 7800 4068 7828
rect 4062 7788 4068 7800
rect 4120 7788 4126 7840
rect 5629 7831 5687 7837
rect 5629 7797 5641 7831
rect 5675 7828 5687 7831
rect 6733 7831 6791 7837
rect 6733 7828 6745 7831
rect 5675 7800 6745 7828
rect 5675 7797 5687 7800
rect 5629 7791 5687 7797
rect 6733 7797 6745 7800
rect 6779 7797 6791 7831
rect 7466 7828 7472 7840
rect 7427 7800 7472 7828
rect 6733 7791 6791 7797
rect 2958 7760 2964 7772
rect 2332 7732 2964 7760
rect 2958 7720 2964 7732
rect 3016 7760 3022 7772
rect 3142 7760 3148 7772
rect 3016 7732 3148 7760
rect 3016 7720 3022 7732
rect 3142 7720 3148 7732
rect 3200 7720 3206 7772
rect 4706 7720 4712 7772
rect 4764 7760 4770 7772
rect 6549 7763 6607 7769
rect 6549 7760 6561 7763
rect 4764 7732 6561 7760
rect 4764 7720 4770 7732
rect 6549 7729 6561 7732
rect 6595 7760 6607 7763
rect 6638 7760 6644 7772
rect 6595 7732 6644 7760
rect 6595 7729 6607 7732
rect 6549 7723 6607 7729
rect 6638 7720 6644 7732
rect 6696 7720 6702 7772
rect 6748 7760 6776 7791
rect 7466 7788 7472 7800
rect 7524 7788 7530 7840
rect 8496 7837 8524 7868
rect 8754 7856 8760 7868
rect 8812 7856 8818 7908
rect 11701 7899 11759 7905
rect 11701 7865 11713 7899
rect 11747 7896 11759 7899
rect 11974 7896 11980 7908
rect 11747 7868 11980 7896
rect 11747 7865 11759 7868
rect 11701 7859 11759 7865
rect 11974 7856 11980 7868
rect 12032 7856 12038 7908
rect 12161 7899 12219 7905
rect 12161 7865 12173 7899
rect 12207 7896 12219 7899
rect 14185 7899 14243 7905
rect 12207 7868 13768 7896
rect 12207 7865 12219 7868
rect 12161 7859 12219 7865
rect 7561 7831 7619 7837
rect 7561 7797 7573 7831
rect 7607 7828 7619 7831
rect 8481 7831 8539 7837
rect 7607 7800 8064 7828
rect 7607 7797 7619 7800
rect 7561 7791 7619 7797
rect 7374 7760 7380 7772
rect 6748 7732 7380 7760
rect 7374 7720 7380 7732
rect 7432 7720 7438 7772
rect 624 7664 1624 7692
rect 2225 7695 2283 7701
rect 624 7652 630 7664
rect 2225 7661 2237 7695
rect 2271 7692 2283 7695
rect 3326 7692 3332 7704
rect 2271 7664 3332 7692
rect 2271 7661 2283 7664
rect 2225 7655 2283 7661
rect 3326 7652 3332 7664
rect 3384 7652 3390 7704
rect 3605 7695 3663 7701
rect 3605 7661 3617 7695
rect 3651 7692 3663 7695
rect 3786 7692 3792 7704
rect 3651 7664 3792 7692
rect 3651 7661 3663 7664
rect 3605 7655 3663 7661
rect 3786 7652 3792 7664
rect 3844 7652 3850 7704
rect 5718 7652 5724 7704
rect 5776 7692 5782 7704
rect 5813 7695 5871 7701
rect 5813 7692 5825 7695
rect 5776 7664 5825 7692
rect 5776 7652 5782 7664
rect 5813 7661 5825 7664
rect 5859 7692 5871 7695
rect 6822 7692 6828 7704
rect 5859 7664 6828 7692
rect 5859 7661 5871 7664
rect 5813 7655 5871 7661
rect 6822 7652 6828 7664
rect 6880 7652 6886 7704
rect 7285 7695 7343 7701
rect 7285 7661 7297 7695
rect 7331 7692 7343 7695
rect 7834 7692 7840 7704
rect 7331 7664 7840 7692
rect 7331 7661 7343 7664
rect 7285 7655 7343 7661
rect 7834 7652 7840 7664
rect 7892 7652 7898 7704
rect 8036 7692 8064 7800
rect 8481 7797 8493 7831
rect 8527 7797 8539 7831
rect 8481 7791 8539 7797
rect 11241 7831 11299 7837
rect 11241 7797 11253 7831
rect 11287 7797 11299 7831
rect 11241 7791 11299 7797
rect 10042 7760 10048 7772
rect 9982 7732 10048 7760
rect 10042 7720 10048 7732
rect 10100 7720 10106 7772
rect 11054 7720 11060 7772
rect 11112 7760 11118 7772
rect 11256 7760 11284 7791
rect 11330 7788 11336 7840
rect 11388 7828 11394 7840
rect 12526 7828 12532 7840
rect 11388 7800 11433 7828
rect 12487 7800 12532 7828
rect 11388 7788 11394 7800
rect 12526 7788 12532 7800
rect 12584 7788 12590 7840
rect 12621 7831 12679 7837
rect 12621 7797 12633 7831
rect 12667 7797 12679 7831
rect 13740 7828 13768 7868
rect 14185 7865 14197 7899
rect 14231 7896 14243 7899
rect 14366 7896 14372 7908
rect 14231 7868 14372 7896
rect 14231 7865 14243 7868
rect 14185 7859 14243 7865
rect 14366 7856 14372 7868
rect 14424 7896 14430 7908
rect 14424 7868 14964 7896
rect 14424 7856 14430 7868
rect 13906 7837 13912 7840
rect 13892 7831 13912 7837
rect 13892 7828 13904 7831
rect 13740 7800 13904 7828
rect 12621 7791 12679 7797
rect 13892 7797 13904 7800
rect 13892 7791 13912 7797
rect 11609 7763 11667 7769
rect 11609 7760 11621 7763
rect 11112 7732 11621 7760
rect 11112 7720 11118 7732
rect 11609 7729 11621 7732
rect 11655 7760 11667 7763
rect 12253 7763 12311 7769
rect 12253 7760 12265 7763
rect 11655 7732 12265 7760
rect 11655 7729 11667 7732
rect 11609 7723 11667 7729
rect 12253 7729 12265 7732
rect 12299 7760 12311 7763
rect 12636 7760 12664 7791
rect 13906 7788 13912 7791
rect 13964 7788 13970 7840
rect 14001 7831 14059 7837
rect 14001 7797 14013 7831
rect 14047 7797 14059 7831
rect 14001 7791 14059 7797
rect 12299 7732 12664 7760
rect 14016 7760 14044 7791
rect 14090 7788 14096 7840
rect 14148 7828 14154 7840
rect 14936 7837 14964 7868
rect 14277 7831 14335 7837
rect 14277 7828 14289 7831
rect 14148 7800 14289 7828
rect 14148 7788 14154 7800
rect 14277 7797 14289 7800
rect 14323 7797 14335 7831
rect 14277 7791 14335 7797
rect 14921 7831 14979 7837
rect 14921 7797 14933 7831
rect 14967 7797 14979 7831
rect 14921 7791 14979 7797
rect 14016 7732 14136 7760
rect 12299 7729 12311 7732
rect 12253 7723 12311 7729
rect 14108 7704 14136 7732
rect 9490 7692 9496 7704
rect 8036 7664 9496 7692
rect 9490 7652 9496 7664
rect 9548 7652 9554 7704
rect 13722 7692 13728 7704
rect 13683 7664 13728 7692
rect 13722 7652 13728 7664
rect 13780 7652 13786 7704
rect 14090 7652 14096 7704
rect 14148 7652 14154 7704
rect 92 7602 15824 7624
rect 92 7550 5242 7602
rect 5294 7550 5306 7602
rect 5358 7550 5370 7602
rect 5422 7550 5434 7602
rect 5486 7550 10514 7602
rect 10566 7550 10578 7602
rect 10630 7550 10642 7602
rect 10694 7550 10706 7602
rect 10758 7550 15824 7602
rect 92 7528 15824 7550
rect 3142 7448 3148 7500
rect 3200 7488 3206 7500
rect 3605 7491 3663 7497
rect 3605 7488 3617 7491
rect 3200 7460 3617 7488
rect 3200 7448 3206 7460
rect 3605 7457 3617 7460
rect 3651 7457 3663 7491
rect 3605 7451 3663 7457
rect 3970 7448 3976 7500
rect 4028 7488 4034 7500
rect 4065 7491 4123 7497
rect 4065 7488 4077 7491
rect 4028 7460 4077 7488
rect 4028 7448 4034 7460
rect 4065 7457 4077 7460
rect 4111 7457 4123 7491
rect 8570 7488 8576 7500
rect 4065 7451 4123 7457
rect 5552 7460 8576 7488
rect 1486 7380 1492 7432
rect 1544 7380 1550 7432
rect 1949 7423 2007 7429
rect 1949 7389 1961 7423
rect 1995 7420 2007 7423
rect 5552 7420 5580 7460
rect 8570 7448 8576 7460
rect 8628 7448 8634 7500
rect 9309 7491 9367 7497
rect 9309 7457 9321 7491
rect 9355 7488 9367 7491
rect 9398 7488 9404 7500
rect 9355 7460 9404 7488
rect 9355 7457 9367 7460
rect 9309 7451 9367 7457
rect 9398 7448 9404 7460
rect 9456 7448 9462 7500
rect 9950 7448 9956 7500
rect 10008 7448 10014 7500
rect 11057 7491 11115 7497
rect 11057 7457 11069 7491
rect 11103 7488 11115 7491
rect 11146 7488 11152 7500
rect 11103 7460 11152 7488
rect 11103 7457 11115 7460
rect 11057 7451 11115 7457
rect 11146 7448 11152 7460
rect 11204 7448 11210 7500
rect 1995 7392 5580 7420
rect 5920 7392 6132 7420
rect 1995 7389 2007 7392
rect 1949 7383 2007 7389
rect 2498 7312 2504 7364
rect 2556 7352 2562 7364
rect 3145 7355 3203 7361
rect 3145 7352 3157 7355
rect 2556 7324 3157 7352
rect 2556 7312 2562 7324
rect 3145 7321 3157 7324
rect 3191 7321 3203 7355
rect 3145 7315 3203 7321
rect 3510 7312 3516 7364
rect 3568 7352 3574 7364
rect 3881 7355 3939 7361
rect 3881 7352 3893 7355
rect 3568 7324 3893 7352
rect 3568 7312 3574 7324
rect 3881 7321 3893 7324
rect 3927 7321 3939 7355
rect 3881 7315 3939 7321
rect 3973 7355 4031 7361
rect 3973 7321 3985 7355
rect 4019 7321 4031 7355
rect 3973 7315 4031 7321
rect 2225 7287 2283 7293
rect 2225 7253 2237 7287
rect 2271 7253 2283 7287
rect 2225 7247 2283 7253
rect 477 7151 535 7157
rect 477 7117 489 7151
rect 523 7148 535 7151
rect 566 7148 572 7160
rect 523 7120 572 7148
rect 523 7117 535 7120
rect 477 7111 535 7117
rect 566 7108 572 7120
rect 624 7108 630 7160
rect 658 7108 664 7160
rect 716 7148 722 7160
rect 2240 7148 2268 7247
rect 3786 7176 3792 7228
rect 3844 7216 3850 7228
rect 3988 7216 4016 7315
rect 5534 7312 5540 7364
rect 5592 7352 5598 7364
rect 5813 7355 5871 7361
rect 5813 7352 5825 7355
rect 5592 7324 5825 7352
rect 5592 7312 5598 7324
rect 5813 7321 5825 7324
rect 5859 7321 5871 7355
rect 5813 7315 5871 7321
rect 4341 7287 4399 7293
rect 4341 7253 4353 7287
rect 4387 7284 4399 7287
rect 4982 7284 4988 7296
rect 4387 7256 4988 7284
rect 4387 7253 4399 7256
rect 4341 7247 4399 7253
rect 4982 7244 4988 7256
rect 5040 7244 5046 7296
rect 5074 7244 5080 7296
rect 5132 7284 5138 7296
rect 5920 7284 5948 7392
rect 6104 7361 6132 7392
rect 6454 7380 6460 7432
rect 6512 7420 6518 7432
rect 6825 7423 6883 7429
rect 6825 7420 6837 7423
rect 6512 7392 6837 7420
rect 6512 7380 6518 7392
rect 6825 7389 6837 7392
rect 6871 7389 6883 7423
rect 7834 7420 7840 7432
rect 7795 7392 7840 7420
rect 6825 7383 6883 7389
rect 7834 7380 7840 7392
rect 7892 7380 7898 7432
rect 9968 7420 9996 7448
rect 9062 7392 9996 7420
rect 10870 7380 10876 7432
rect 10928 7420 10934 7432
rect 10928 7392 11376 7420
rect 10928 7380 10934 7392
rect 5997 7355 6055 7361
rect 5997 7321 6009 7355
rect 6043 7321 6055 7355
rect 5997 7315 6055 7321
rect 6089 7355 6147 7361
rect 6089 7321 6101 7355
rect 6135 7321 6147 7355
rect 6089 7315 6147 7321
rect 6348 7355 6406 7361
rect 6348 7321 6360 7355
rect 6394 7352 6406 7355
rect 6730 7352 6736 7364
rect 6394 7324 6736 7352
rect 6394 7321 6406 7324
rect 6348 7315 6406 7321
rect 5132 7256 5948 7284
rect 6012 7284 6040 7315
rect 6730 7312 6736 7324
rect 6788 7312 6794 7364
rect 7006 7352 7012 7364
rect 6967 7324 7012 7352
rect 7006 7312 7012 7324
rect 7064 7312 7070 7364
rect 7558 7352 7564 7364
rect 7519 7324 7564 7352
rect 7558 7312 7564 7324
rect 7616 7312 7622 7364
rect 9490 7312 9496 7364
rect 9548 7352 9554 7364
rect 9769 7355 9827 7361
rect 9769 7352 9781 7355
rect 9548 7324 9781 7352
rect 9548 7312 9554 7324
rect 9769 7321 9781 7324
rect 9815 7321 9827 7355
rect 9769 7315 9827 7321
rect 9858 7312 9864 7364
rect 9916 7352 9922 7364
rect 9953 7355 10011 7361
rect 9953 7352 9965 7355
rect 9916 7324 9965 7352
rect 9916 7312 9922 7324
rect 9953 7321 9965 7324
rect 9999 7321 10011 7355
rect 11238 7352 11244 7364
rect 11199 7324 11244 7352
rect 9953 7315 10011 7321
rect 11238 7312 11244 7324
rect 11296 7312 11302 7364
rect 11348 7352 11376 7392
rect 11422 7380 11428 7432
rect 11480 7420 11486 7432
rect 11480 7392 11836 7420
rect 11480 7380 11486 7392
rect 11517 7355 11575 7361
rect 11517 7352 11529 7355
rect 11348 7324 11529 7352
rect 11517 7321 11529 7324
rect 11563 7321 11575 7355
rect 11517 7315 11575 7321
rect 11609 7355 11667 7361
rect 11609 7321 11621 7355
rect 11655 7352 11667 7355
rect 11698 7352 11704 7364
rect 11655 7324 11704 7352
rect 11655 7321 11667 7324
rect 11609 7315 11667 7321
rect 11698 7312 11704 7324
rect 11756 7312 11762 7364
rect 11808 7361 11836 7392
rect 13446 7380 13452 7432
rect 13504 7380 13510 7432
rect 11793 7355 11851 7361
rect 11793 7321 11805 7355
rect 11839 7321 11851 7355
rect 12710 7352 12716 7364
rect 12671 7324 12716 7352
rect 11793 7315 11851 7321
rect 12710 7312 12716 7324
rect 12768 7312 12774 7364
rect 6012 7256 6316 7284
rect 5132 7244 5138 7256
rect 6288 7216 6316 7256
rect 10134 7244 10140 7296
rect 10192 7284 10198 7296
rect 11425 7287 11483 7293
rect 11425 7284 11437 7287
rect 10192 7256 11437 7284
rect 10192 7244 10198 7256
rect 11425 7253 11437 7256
rect 11471 7253 11483 7287
rect 11425 7247 11483 7253
rect 12986 7244 12992 7296
rect 13044 7284 13050 7296
rect 13081 7287 13139 7293
rect 13081 7284 13093 7287
rect 13044 7256 13093 7284
rect 13044 7244 13050 7256
rect 13081 7253 13093 7256
rect 13127 7253 13139 7287
rect 14550 7284 14556 7296
rect 13081 7247 13139 7253
rect 13832 7256 14556 7284
rect 6822 7216 6828 7228
rect 3844 7188 6224 7216
rect 6288 7188 6828 7216
rect 3844 7176 3850 7188
rect 6196 7160 6224 7188
rect 6822 7176 6828 7188
rect 6880 7176 6886 7228
rect 10045 7219 10103 7225
rect 10045 7185 10057 7219
rect 10091 7216 10103 7219
rect 10091 7188 12434 7216
rect 10091 7185 10103 7188
rect 10045 7179 10103 7185
rect 3050 7148 3056 7160
rect 716 7120 2268 7148
rect 3011 7120 3056 7148
rect 716 7108 722 7120
rect 3050 7108 3056 7120
rect 3108 7108 3114 7160
rect 4249 7151 4307 7157
rect 4249 7117 4261 7151
rect 4295 7148 4307 7151
rect 5626 7148 5632 7160
rect 4295 7120 5632 7148
rect 4295 7117 4307 7120
rect 4249 7111 4307 7117
rect 5626 7108 5632 7120
rect 5684 7108 5690 7160
rect 5810 7148 5816 7160
rect 5771 7120 5816 7148
rect 5810 7108 5816 7120
rect 5868 7108 5874 7160
rect 6178 7108 6184 7160
rect 6236 7148 6242 7160
rect 6273 7151 6331 7157
rect 6273 7148 6285 7151
rect 6236 7120 6285 7148
rect 6236 7108 6242 7120
rect 6273 7117 6285 7120
rect 6319 7117 6331 7151
rect 12406 7148 12434 7188
rect 13832 7148 13860 7256
rect 14550 7244 14556 7256
rect 14608 7244 14614 7296
rect 12406 7120 13860 7148
rect 6273 7111 6331 7117
rect 13906 7108 13912 7160
rect 13964 7148 13970 7160
rect 14507 7151 14565 7157
rect 14507 7148 14519 7151
rect 13964 7120 14519 7148
rect 13964 7108 13970 7120
rect 14507 7117 14519 7120
rect 14553 7117 14565 7151
rect 14507 7111 14565 7117
rect 92 7058 15824 7080
rect 92 7006 2606 7058
rect 2658 7006 2670 7058
rect 2722 7006 2734 7058
rect 2786 7006 2798 7058
rect 2850 7006 7878 7058
rect 7930 7006 7942 7058
rect 7994 7006 8006 7058
rect 8058 7006 8070 7058
rect 8122 7006 13150 7058
rect 13202 7006 13214 7058
rect 13266 7006 13278 7058
rect 13330 7006 13342 7058
rect 13394 7006 15824 7058
rect 92 6984 15824 7006
rect 3142 6904 3148 6956
rect 3200 6944 3206 6956
rect 3418 6944 3424 6956
rect 3200 6916 3424 6944
rect 3200 6904 3206 6916
rect 3418 6904 3424 6916
rect 3476 6904 3482 6956
rect 3605 6947 3663 6953
rect 3605 6913 3617 6947
rect 3651 6944 3663 6947
rect 4062 6944 4068 6956
rect 3651 6916 4068 6944
rect 3651 6913 3663 6916
rect 3605 6907 3663 6913
rect 4062 6904 4068 6916
rect 4120 6904 4126 6956
rect 7009 6947 7067 6953
rect 6472 6916 6960 6944
rect 4154 6876 4160 6888
rect 2792 6848 4160 6876
rect 2792 6808 2820 6848
rect 4154 6836 4160 6848
rect 4212 6836 4218 6888
rect 4430 6876 4436 6888
rect 4391 6848 4436 6876
rect 4430 6836 4436 6848
rect 4488 6836 4494 6888
rect 5626 6836 5632 6888
rect 5684 6876 5690 6888
rect 6472 6876 6500 6916
rect 5684 6848 6500 6876
rect 5684 6836 5690 6848
rect 6638 6836 6644 6888
rect 6696 6876 6702 6888
rect 6932 6876 6960 6916
rect 7009 6913 7021 6947
rect 7055 6944 7067 6947
rect 7466 6944 7472 6956
rect 7055 6916 7472 6944
rect 7055 6913 7067 6916
rect 7009 6907 7067 6913
rect 7466 6904 7472 6916
rect 7524 6904 7530 6956
rect 11698 6876 11704 6888
rect 6696 6848 6776 6876
rect 6932 6848 11704 6876
rect 6696 6836 6702 6848
rect 4522 6808 4528 6820
rect 2148 6780 2820 6808
rect 2884 6780 3924 6808
rect 4483 6780 4528 6808
rect 566 6700 572 6752
rect 624 6740 630 6752
rect 2148 6749 2176 6780
rect 937 6743 995 6749
rect 937 6740 949 6743
rect 624 6712 949 6740
rect 624 6700 630 6712
rect 937 6709 949 6712
rect 983 6709 995 6743
rect 937 6703 995 6709
rect 1673 6743 1731 6749
rect 1673 6709 1685 6743
rect 1719 6709 1731 6743
rect 1673 6703 1731 6709
rect 2133 6743 2191 6749
rect 2133 6709 2145 6743
rect 2179 6709 2191 6743
rect 2314 6740 2320 6752
rect 2275 6712 2320 6740
rect 2133 6703 2191 6709
rect 750 6672 756 6684
rect 711 6644 756 6672
rect 750 6632 756 6644
rect 808 6632 814 6684
rect 1688 6672 1716 6703
rect 2314 6700 2320 6712
rect 2372 6700 2378 6752
rect 2884 6740 2912 6780
rect 2746 6712 2912 6740
rect 2746 6672 2774 6712
rect 2958 6700 2964 6752
rect 3016 6740 3022 6752
rect 3016 6712 3372 6740
rect 3016 6700 3022 6712
rect 1688 6644 2774 6672
rect 3050 6632 3056 6684
rect 3108 6672 3114 6684
rect 3237 6675 3295 6681
rect 3237 6672 3249 6675
rect 3108 6644 3249 6672
rect 3108 6632 3114 6644
rect 3237 6641 3249 6644
rect 3283 6641 3295 6675
rect 3344 6672 3372 6712
rect 3442 6675 3500 6681
rect 3442 6672 3454 6675
rect 3344 6644 3454 6672
rect 3237 6635 3295 6641
rect 3442 6641 3454 6644
rect 3488 6641 3500 6675
rect 3442 6635 3500 6641
rect 1394 6564 1400 6616
rect 1452 6604 1458 6616
rect 1578 6604 1584 6616
rect 1452 6576 1584 6604
rect 1452 6564 1458 6576
rect 1578 6564 1584 6576
rect 1636 6564 1642 6616
rect 1670 6564 1676 6616
rect 1728 6604 1734 6616
rect 1946 6604 1952 6616
rect 1728 6576 1952 6604
rect 1728 6564 1734 6576
rect 1946 6564 1952 6576
rect 2004 6564 2010 6616
rect 2317 6607 2375 6613
rect 2317 6573 2329 6607
rect 2363 6604 2375 6607
rect 3326 6604 3332 6616
rect 2363 6576 3332 6604
rect 2363 6573 2375 6576
rect 2317 6567 2375 6573
rect 3326 6564 3332 6576
rect 3384 6564 3390 6616
rect 3896 6604 3924 6780
rect 4522 6768 4528 6780
rect 4580 6768 4586 6820
rect 6270 6808 6276 6820
rect 4816 6780 6276 6808
rect 4617 6743 4675 6749
rect 4617 6709 4629 6743
rect 4663 6740 4675 6743
rect 4816 6740 4844 6780
rect 6270 6768 6276 6780
rect 6328 6808 6334 6820
rect 6328 6780 6687 6808
rect 6328 6768 6334 6780
rect 4982 6740 4988 6752
rect 4663 6712 4844 6740
rect 4943 6712 4988 6740
rect 4663 6709 4675 6712
rect 4617 6703 4675 6709
rect 4982 6700 4988 6712
rect 5040 6700 5046 6752
rect 5077 6743 5135 6749
rect 5077 6709 5089 6743
rect 5123 6709 5135 6743
rect 5077 6703 5135 6709
rect 5905 6743 5963 6749
rect 5905 6709 5917 6743
rect 5951 6709 5963 6743
rect 6362 6740 6368 6752
rect 6323 6712 6368 6740
rect 5905 6703 5963 6709
rect 3970 6632 3976 6684
rect 4028 6672 4034 6684
rect 5092 6672 5120 6703
rect 4028 6644 5120 6672
rect 5920 6672 5948 6703
rect 6362 6700 6368 6712
rect 6420 6700 6426 6752
rect 6454 6700 6460 6752
rect 6512 6740 6518 6752
rect 6659 6749 6687 6780
rect 6748 6749 6776 6848
rect 9674 6808 9680 6820
rect 9635 6780 9680 6808
rect 9674 6768 9680 6780
rect 9732 6768 9738 6820
rect 6549 6743 6607 6749
rect 6549 6740 6561 6743
rect 6512 6712 6561 6740
rect 6512 6700 6518 6712
rect 6549 6709 6561 6712
rect 6595 6709 6607 6743
rect 6549 6703 6607 6709
rect 6644 6743 6702 6749
rect 6644 6709 6656 6743
rect 6690 6709 6702 6743
rect 6644 6703 6702 6709
rect 6733 6743 6791 6749
rect 6733 6709 6745 6743
rect 6779 6709 6791 6743
rect 8849 6743 8907 6749
rect 8849 6740 8861 6743
rect 6733 6703 6791 6709
rect 8312 6712 8861 6740
rect 8312 6672 8340 6712
rect 8849 6709 8861 6712
rect 8895 6740 8907 6743
rect 9490 6740 9496 6752
rect 8895 6712 9496 6740
rect 8895 6709 8907 6712
rect 8849 6703 8907 6709
rect 9490 6700 9496 6712
rect 9548 6700 9554 6752
rect 9585 6743 9643 6749
rect 9585 6709 9597 6743
rect 9631 6709 9643 6743
rect 9968 6740 9996 6848
rect 11698 6836 11704 6848
rect 11756 6876 11762 6888
rect 14090 6876 14096 6888
rect 11756 6848 12434 6876
rect 11756 6836 11762 6848
rect 10134 6808 10140 6820
rect 10095 6780 10140 6808
rect 10134 6768 10140 6780
rect 10192 6768 10198 6820
rect 11238 6808 11244 6820
rect 10428 6780 11244 6808
rect 10428 6749 10456 6780
rect 11238 6768 11244 6780
rect 11296 6768 11302 6820
rect 11517 6811 11575 6817
rect 11517 6777 11529 6811
rect 11563 6808 11575 6811
rect 12066 6808 12072 6820
rect 11563 6780 12072 6808
rect 11563 6777 11575 6780
rect 11517 6771 11575 6777
rect 12066 6768 12072 6780
rect 12124 6768 12130 6820
rect 12406 6808 12434 6848
rect 13648 6848 14096 6876
rect 13648 6808 13676 6848
rect 14090 6836 14096 6848
rect 14148 6876 14154 6888
rect 14737 6879 14795 6885
rect 14737 6876 14749 6879
rect 14148 6848 14749 6876
rect 14148 6836 14154 6848
rect 14737 6845 14749 6848
rect 14783 6845 14795 6879
rect 14737 6839 14795 6845
rect 12406 6780 13676 6808
rect 13722 6768 13728 6820
rect 13780 6808 13786 6820
rect 14182 6808 14188 6820
rect 13780 6780 14044 6808
rect 14143 6780 14188 6808
rect 13780 6768 13786 6780
rect 10045 6743 10103 6749
rect 10045 6740 10057 6743
rect 9968 6712 10057 6740
rect 9585 6703 9643 6709
rect 10045 6709 10057 6712
rect 10091 6709 10103 6743
rect 10045 6703 10103 6709
rect 10413 6743 10471 6749
rect 10413 6709 10425 6743
rect 10459 6709 10471 6743
rect 10413 6703 10471 6709
rect 10597 6743 10655 6749
rect 10597 6709 10609 6743
rect 10643 6740 10655 6743
rect 10870 6740 10876 6752
rect 10643 6712 10876 6740
rect 10643 6709 10655 6712
rect 10597 6703 10655 6709
rect 8478 6672 8484 6684
rect 5920 6644 8340 6672
rect 8439 6644 8484 6672
rect 4028 6632 4034 6644
rect 8478 6632 8484 6644
rect 8536 6632 8542 6684
rect 8662 6672 8668 6684
rect 8623 6644 8668 6672
rect 8662 6632 8668 6644
rect 8720 6632 8726 6684
rect 9600 6672 9628 6703
rect 10870 6700 10876 6712
rect 10928 6700 10934 6752
rect 11885 6743 11943 6749
rect 11885 6740 11897 6743
rect 11624 6712 11897 6740
rect 11422 6672 11428 6684
rect 9600 6644 11428 6672
rect 11422 6632 11428 6644
rect 11480 6632 11486 6684
rect 7190 6604 7196 6616
rect 3896 6576 7196 6604
rect 7190 6564 7196 6576
rect 7248 6564 7254 6616
rect 11514 6564 11520 6616
rect 11572 6604 11578 6616
rect 11624 6613 11652 6712
rect 11885 6709 11897 6712
rect 11931 6709 11943 6743
rect 11885 6703 11943 6709
rect 12805 6743 12863 6749
rect 12805 6709 12817 6743
rect 12851 6740 12863 6743
rect 13906 6740 13912 6752
rect 12851 6712 13912 6740
rect 12851 6709 12863 6712
rect 12805 6703 12863 6709
rect 13906 6700 13912 6712
rect 13964 6700 13970 6752
rect 14016 6749 14044 6780
rect 14182 6768 14188 6780
rect 14240 6768 14246 6820
rect 14001 6743 14059 6749
rect 14001 6709 14013 6743
rect 14047 6709 14059 6743
rect 14274 6740 14280 6752
rect 14235 6712 14280 6740
rect 14001 6703 14059 6709
rect 14274 6700 14280 6712
rect 14332 6700 14338 6752
rect 14921 6743 14979 6749
rect 14921 6709 14933 6743
rect 14967 6740 14979 6743
rect 15010 6740 15016 6752
rect 14967 6712 15016 6740
rect 14967 6709 14979 6712
rect 14921 6703 14979 6709
rect 15010 6700 15016 6712
rect 15068 6700 15074 6752
rect 13630 6632 13636 6684
rect 13688 6672 13694 6684
rect 13725 6675 13783 6681
rect 13725 6672 13737 6675
rect 13688 6644 13737 6672
rect 13688 6632 13694 6644
rect 13725 6641 13737 6644
rect 13771 6641 13783 6675
rect 13725 6635 13783 6641
rect 11609 6607 11667 6613
rect 11609 6604 11621 6607
rect 11572 6576 11621 6604
rect 11572 6564 11578 6576
rect 11609 6573 11621 6576
rect 11655 6573 11667 6607
rect 11609 6567 11667 6573
rect 11698 6564 11704 6616
rect 11756 6604 11762 6616
rect 12713 6607 12771 6613
rect 11756 6576 11801 6604
rect 11756 6564 11762 6576
rect 12713 6573 12725 6607
rect 12759 6604 12771 6607
rect 12894 6604 12900 6616
rect 12759 6576 12900 6604
rect 12759 6573 12771 6576
rect 12713 6567 12771 6573
rect 12894 6564 12900 6576
rect 12952 6604 12958 6616
rect 14292 6604 14320 6700
rect 12952 6576 14320 6604
rect 12952 6564 12958 6576
rect 92 6514 15824 6536
rect 92 6462 5242 6514
rect 5294 6462 5306 6514
rect 5358 6462 5370 6514
rect 5422 6462 5434 6514
rect 5486 6462 10514 6514
rect 10566 6462 10578 6514
rect 10630 6462 10642 6514
rect 10694 6462 10706 6514
rect 10758 6462 15824 6514
rect 92 6440 15824 6462
rect 3329 6403 3387 6409
rect 3329 6400 3341 6403
rect 952 6372 3341 6400
rect 952 6341 980 6372
rect 3329 6369 3341 6372
rect 3375 6369 3387 6403
rect 3786 6400 3792 6412
rect 3747 6372 3792 6400
rect 3329 6363 3387 6369
rect 3786 6360 3792 6372
rect 3844 6360 3850 6412
rect 4893 6403 4951 6409
rect 4893 6369 4905 6403
rect 4939 6400 4951 6403
rect 7006 6400 7012 6412
rect 4939 6372 7012 6400
rect 4939 6369 4951 6372
rect 4893 6363 4951 6369
rect 7006 6360 7012 6372
rect 7064 6360 7070 6412
rect 7742 6360 7748 6412
rect 7800 6400 7806 6412
rect 7929 6403 7987 6409
rect 7929 6400 7941 6403
rect 7800 6372 7941 6400
rect 7800 6360 7806 6372
rect 7929 6369 7941 6372
rect 7975 6369 7987 6403
rect 7929 6363 7987 6369
rect 8662 6360 8668 6412
rect 8720 6400 8726 6412
rect 8846 6400 8852 6412
rect 8720 6372 8852 6400
rect 8720 6360 8726 6372
rect 8846 6360 8852 6372
rect 8904 6400 8910 6412
rect 8904 6372 9904 6400
rect 8904 6360 8910 6372
rect 937 6335 995 6341
rect 937 6301 949 6335
rect 983 6301 995 6335
rect 937 6295 995 6301
rect 1946 6292 1952 6344
rect 2004 6292 2010 6344
rect 6546 6332 6552 6344
rect 2240 6304 6552 6332
rect 566 6156 572 6208
rect 624 6196 630 6208
rect 661 6199 719 6205
rect 661 6196 673 6199
rect 624 6168 673 6196
rect 624 6156 630 6168
rect 661 6165 673 6168
rect 707 6165 719 6199
rect 661 6159 719 6165
rect 934 6156 940 6208
rect 992 6196 998 6208
rect 2240 6196 2268 6304
rect 6546 6292 6552 6304
rect 6604 6292 6610 6344
rect 6822 6292 6828 6344
rect 6880 6332 6886 6344
rect 6880 6304 9168 6332
rect 6880 6292 6886 6304
rect 3694 6264 3700 6276
rect 3655 6236 3700 6264
rect 3694 6224 3700 6236
rect 3752 6224 3758 6276
rect 4154 6224 4160 6276
rect 4212 6264 4218 6276
rect 4525 6267 4583 6273
rect 4525 6264 4537 6267
rect 4212 6236 4537 6264
rect 4212 6224 4218 6236
rect 4525 6233 4537 6236
rect 4571 6233 4583 6267
rect 4525 6227 4583 6233
rect 4709 6267 4767 6273
rect 4709 6233 4721 6267
rect 4755 6264 4767 6267
rect 4890 6264 4896 6276
rect 4755 6236 4896 6264
rect 4755 6233 4767 6236
rect 4709 6227 4767 6233
rect 4890 6224 4896 6236
rect 4948 6224 4954 6276
rect 5718 6224 5724 6276
rect 5776 6264 5782 6276
rect 6181 6267 6239 6273
rect 6181 6264 6193 6267
rect 5776 6236 6193 6264
rect 5776 6224 5782 6236
rect 6181 6233 6193 6236
rect 6227 6233 6239 6267
rect 6181 6227 6239 6233
rect 6454 6224 6460 6276
rect 6512 6264 6518 6276
rect 6641 6267 6699 6273
rect 6641 6264 6653 6267
rect 6512 6236 6653 6264
rect 6512 6224 6518 6236
rect 6641 6233 6653 6236
rect 6687 6233 6699 6267
rect 6641 6227 6699 6233
rect 8849 6267 8907 6273
rect 8849 6233 8861 6267
rect 8895 6233 8907 6267
rect 9030 6264 9036 6276
rect 8991 6236 9036 6264
rect 8849 6227 8907 6233
rect 992 6168 2268 6196
rect 2685 6199 2743 6205
rect 992 6156 998 6168
rect 2685 6165 2697 6199
rect 2731 6196 2743 6199
rect 3142 6196 3148 6208
rect 2731 6168 3148 6196
rect 2731 6165 2743 6168
rect 2685 6159 2743 6165
rect 3142 6156 3148 6168
rect 3200 6196 3206 6208
rect 3418 6196 3424 6208
rect 3200 6168 3424 6196
rect 3200 6156 3206 6168
rect 3418 6156 3424 6168
rect 3476 6156 3482 6208
rect 3973 6199 4031 6205
rect 3973 6165 3985 6199
rect 4019 6196 4031 6199
rect 4430 6196 4436 6208
rect 4019 6168 4436 6196
rect 4019 6165 4031 6168
rect 3973 6159 4031 6165
rect 4430 6156 4436 6168
rect 4488 6156 4494 6208
rect 8570 6156 8576 6208
rect 8628 6196 8634 6208
rect 8864 6196 8892 6227
rect 9030 6224 9036 6236
rect 9088 6224 9094 6276
rect 9140 6264 9168 6304
rect 9490 6292 9496 6344
rect 9548 6332 9554 6344
rect 9769 6335 9827 6341
rect 9769 6332 9781 6335
rect 9548 6304 9781 6332
rect 9548 6292 9554 6304
rect 9769 6301 9781 6304
rect 9815 6301 9827 6335
rect 9876 6332 9904 6372
rect 11330 6360 11336 6412
rect 11388 6400 11394 6412
rect 11517 6403 11575 6409
rect 11517 6400 11529 6403
rect 11388 6372 11529 6400
rect 11388 6360 11394 6372
rect 11517 6369 11529 6372
rect 11563 6369 11575 6403
rect 11517 6363 11575 6369
rect 12986 6360 12992 6412
rect 13044 6400 13050 6412
rect 13265 6403 13323 6409
rect 13265 6400 13277 6403
rect 13044 6372 13277 6400
rect 13044 6360 13050 6372
rect 13265 6369 13277 6372
rect 13311 6369 13323 6403
rect 14366 6400 14372 6412
rect 14327 6372 14372 6400
rect 13265 6363 13323 6369
rect 14366 6360 14372 6372
rect 14424 6360 14430 6412
rect 12894 6332 12900 6344
rect 9876 6304 12112 6332
rect 12855 6304 12900 6332
rect 9769 6295 9827 6301
rect 10134 6264 10140 6276
rect 9140 6236 10140 6264
rect 10134 6224 10140 6236
rect 10192 6224 10198 6276
rect 11422 6264 11428 6276
rect 11383 6236 11428 6264
rect 11422 6224 11428 6236
rect 11480 6224 11486 6276
rect 11609 6267 11667 6273
rect 11609 6233 11621 6267
rect 11655 6264 11667 6267
rect 11698 6264 11704 6276
rect 11655 6236 11704 6264
rect 11655 6233 11667 6236
rect 11609 6227 11667 6233
rect 11698 6224 11704 6236
rect 11756 6224 11762 6276
rect 12084 6273 12112 6304
rect 12894 6292 12900 6304
rect 12952 6292 12958 6344
rect 13906 6332 13912 6344
rect 13004 6304 13912 6332
rect 12069 6267 12127 6273
rect 12069 6233 12081 6267
rect 12115 6233 12127 6267
rect 12069 6227 12127 6233
rect 12250 6224 12256 6276
rect 12308 6264 12314 6276
rect 13004 6273 13032 6304
rect 13906 6292 13912 6304
rect 13964 6292 13970 6344
rect 15010 6332 15016 6344
rect 14476 6304 15016 6332
rect 14476 6273 14504 6304
rect 15010 6292 15016 6304
rect 15068 6292 15074 6344
rect 12713 6267 12771 6273
rect 12713 6264 12725 6267
rect 12308 6236 12725 6264
rect 12308 6224 12314 6236
rect 12713 6233 12725 6236
rect 12759 6233 12771 6267
rect 12713 6227 12771 6233
rect 12989 6267 13047 6273
rect 12989 6233 13001 6267
rect 13035 6233 13047 6267
rect 12989 6227 13047 6233
rect 13081 6267 13139 6273
rect 13081 6233 13093 6267
rect 13127 6233 13139 6267
rect 13081 6227 13139 6233
rect 14461 6267 14519 6273
rect 14461 6233 14473 6267
rect 14507 6233 14519 6267
rect 14921 6267 14979 6273
rect 14921 6264 14933 6267
rect 14461 6227 14519 6233
rect 14660 6236 14933 6264
rect 12161 6199 12219 6205
rect 12161 6196 12173 6199
rect 8628 6168 12173 6196
rect 8628 6156 8634 6168
rect 12161 6165 12173 6168
rect 12207 6165 12219 6199
rect 12618 6196 12624 6208
rect 12161 6159 12219 6165
rect 12406 6168 12624 6196
rect 2314 6088 2320 6140
rect 2372 6128 2378 6140
rect 5902 6128 5908 6140
rect 2372 6100 5908 6128
rect 2372 6088 2378 6100
rect 5902 6088 5908 6100
rect 5960 6128 5966 6140
rect 6089 6131 6147 6137
rect 6089 6128 6101 6131
rect 5960 6100 6101 6128
rect 5960 6088 5966 6100
rect 6089 6097 6101 6100
rect 6135 6097 6147 6131
rect 6089 6091 6147 6097
rect 9125 6131 9183 6137
rect 9125 6097 9137 6131
rect 9171 6128 9183 6131
rect 11606 6128 11612 6140
rect 9171 6100 11612 6128
rect 9171 6097 9183 6100
rect 9125 6091 9183 6097
rect 11606 6088 11612 6100
rect 11664 6088 11670 6140
rect 1578 6020 1584 6072
rect 1636 6060 1642 6072
rect 4338 6060 4344 6072
rect 1636 6032 4344 6060
rect 1636 6020 1642 6032
rect 4338 6020 4344 6032
rect 4396 6060 4402 6072
rect 4525 6063 4583 6069
rect 4525 6060 4537 6063
rect 4396 6032 4537 6060
rect 4396 6020 4402 6032
rect 4525 6029 4537 6032
rect 4571 6060 4583 6063
rect 4982 6060 4988 6072
rect 4571 6032 4988 6060
rect 4571 6029 4583 6032
rect 4525 6023 4583 6029
rect 4982 6020 4988 6032
rect 5040 6020 5046 6072
rect 5626 6020 5632 6072
rect 5684 6060 5690 6072
rect 9861 6063 9919 6069
rect 9861 6060 9873 6063
rect 5684 6032 9873 6060
rect 5684 6020 5690 6032
rect 9861 6029 9873 6032
rect 9907 6060 9919 6063
rect 11422 6060 11428 6072
rect 9907 6032 11428 6060
rect 9907 6029 9919 6032
rect 9861 6023 9919 6029
rect 11422 6020 11428 6032
rect 11480 6060 11486 6072
rect 12406 6060 12434 6168
rect 12618 6156 12624 6168
rect 12676 6196 12682 6208
rect 13096 6196 13124 6227
rect 12676 6168 13124 6196
rect 12676 6156 12682 6168
rect 13538 6088 13544 6140
rect 13596 6128 13602 6140
rect 14660 6128 14688 6236
rect 14921 6233 14933 6236
rect 14967 6233 14979 6267
rect 15102 6264 15108 6276
rect 15063 6236 15108 6264
rect 14921 6227 14979 6233
rect 15102 6224 15108 6236
rect 15160 6224 15166 6276
rect 13596 6100 14688 6128
rect 13596 6088 13602 6100
rect 11480 6032 12434 6060
rect 11480 6020 11486 6032
rect 13998 6020 14004 6072
rect 14056 6060 14062 6072
rect 14921 6063 14979 6069
rect 14921 6060 14933 6063
rect 14056 6032 14933 6060
rect 14056 6020 14062 6032
rect 14921 6029 14933 6032
rect 14967 6029 14979 6063
rect 14921 6023 14979 6029
rect 92 5970 15824 5992
rect 92 5918 2606 5970
rect 2658 5918 2670 5970
rect 2722 5918 2734 5970
rect 2786 5918 2798 5970
rect 2850 5918 7878 5970
rect 7930 5918 7942 5970
rect 7994 5918 8006 5970
rect 8058 5918 8070 5970
rect 8122 5918 13150 5970
rect 13202 5918 13214 5970
rect 13266 5918 13278 5970
rect 13330 5918 13342 5970
rect 13394 5918 15824 5970
rect 92 5896 15824 5918
rect 845 5859 903 5865
rect 845 5825 857 5859
rect 891 5856 903 5859
rect 1762 5856 1768 5868
rect 891 5828 1768 5856
rect 891 5825 903 5828
rect 845 5819 903 5825
rect 1762 5816 1768 5828
rect 1820 5816 1826 5868
rect 3418 5816 3424 5868
rect 3476 5856 3482 5868
rect 3513 5859 3571 5865
rect 3513 5856 3525 5859
rect 3476 5828 3525 5856
rect 3476 5816 3482 5828
rect 3513 5825 3525 5828
rect 3559 5825 3571 5859
rect 3513 5819 3571 5825
rect 1578 5788 1584 5800
rect 1539 5760 1584 5788
rect 1578 5748 1584 5760
rect 1636 5748 1642 5800
rect 3528 5788 3556 5819
rect 3694 5816 3700 5868
rect 3752 5856 3758 5868
rect 5445 5859 5503 5865
rect 5445 5856 5457 5859
rect 3752 5828 5457 5856
rect 3752 5816 3758 5828
rect 5445 5825 5457 5828
rect 5491 5825 5503 5859
rect 5445 5819 5503 5825
rect 6362 5816 6368 5868
rect 6420 5856 6426 5868
rect 6641 5859 6699 5865
rect 6641 5856 6653 5859
rect 6420 5828 6653 5856
rect 6420 5816 6426 5828
rect 6641 5825 6653 5828
rect 6687 5825 6699 5859
rect 6641 5819 6699 5825
rect 8478 5816 8484 5868
rect 8536 5856 8542 5868
rect 8573 5859 8631 5865
rect 8573 5856 8585 5859
rect 8536 5828 8585 5856
rect 8536 5816 8542 5828
rect 8573 5825 8585 5828
rect 8619 5825 8631 5859
rect 13817 5859 13875 5865
rect 8573 5819 8631 5825
rect 8680 5828 12756 5856
rect 3528 5760 4292 5788
rect 1394 5720 1400 5732
rect 676 5692 1400 5720
rect 676 5661 704 5692
rect 1394 5680 1400 5692
rect 1452 5680 1458 5732
rect 2317 5723 2375 5729
rect 2317 5689 2329 5723
rect 2363 5720 2375 5723
rect 3970 5720 3976 5732
rect 2363 5692 3976 5720
rect 2363 5689 2375 5692
rect 2317 5683 2375 5689
rect 3970 5680 3976 5692
rect 4028 5680 4034 5732
rect 4264 5664 4292 5760
rect 6914 5748 6920 5800
rect 6972 5748 6978 5800
rect 7006 5748 7012 5800
rect 7064 5788 7070 5800
rect 8680 5788 8708 5828
rect 7064 5760 8708 5788
rect 7064 5748 7070 5760
rect 11790 5748 11796 5800
rect 11848 5788 11854 5800
rect 12434 5788 12440 5800
rect 11848 5760 12440 5788
rect 11848 5748 11854 5760
rect 12434 5748 12440 5760
rect 12492 5748 12498 5800
rect 5994 5720 6000 5732
rect 5955 5692 6000 5720
rect 5994 5680 6000 5692
rect 6052 5680 6058 5732
rect 6932 5720 6960 5748
rect 7101 5723 7159 5729
rect 7101 5720 7113 5723
rect 6932 5692 7113 5720
rect 7101 5689 7113 5692
rect 7147 5720 7159 5723
rect 12621 5723 12679 5729
rect 12621 5720 12633 5723
rect 7147 5692 12633 5720
rect 7147 5689 7159 5692
rect 7101 5683 7159 5689
rect 12621 5689 12633 5692
rect 12667 5689 12679 5723
rect 12621 5683 12679 5689
rect 661 5655 719 5661
rect 661 5621 673 5655
rect 707 5621 719 5655
rect 661 5615 719 5621
rect 845 5655 903 5661
rect 845 5621 857 5655
rect 891 5652 903 5655
rect 2038 5652 2044 5664
rect 891 5624 2044 5652
rect 891 5621 903 5624
rect 845 5615 903 5621
rect 2038 5612 2044 5624
rect 2096 5612 2102 5664
rect 2133 5655 2191 5661
rect 2133 5621 2145 5655
rect 2179 5652 2191 5655
rect 2958 5652 2964 5664
rect 2179 5624 2964 5652
rect 2179 5621 2191 5624
rect 2133 5615 2191 5621
rect 2958 5612 2964 5624
rect 3016 5612 3022 5664
rect 4246 5652 4252 5664
rect 4207 5624 4252 5652
rect 4246 5612 4252 5624
rect 4304 5612 4310 5664
rect 4338 5612 4344 5664
rect 4396 5652 4402 5664
rect 4525 5655 4583 5661
rect 4396 5624 4441 5652
rect 4396 5612 4402 5624
rect 4525 5621 4537 5655
rect 4571 5652 4583 5655
rect 4890 5652 4896 5664
rect 4571 5624 4896 5652
rect 4571 5621 4583 5624
rect 4525 5615 4583 5621
rect 4890 5612 4896 5624
rect 4948 5612 4954 5664
rect 5810 5652 5816 5664
rect 5771 5624 5816 5652
rect 5810 5612 5816 5624
rect 5868 5612 5874 5664
rect 5902 5612 5908 5664
rect 5960 5652 5966 5664
rect 6822 5652 6828 5664
rect 5960 5624 6005 5652
rect 6783 5624 6828 5652
rect 5960 5612 5966 5624
rect 6822 5612 6828 5624
rect 6880 5612 6886 5664
rect 6914 5612 6920 5664
rect 6972 5652 6978 5664
rect 7193 5655 7251 5661
rect 6972 5624 7017 5652
rect 6972 5612 6978 5624
rect 7193 5621 7205 5655
rect 7239 5652 7251 5655
rect 8570 5652 8576 5664
rect 7239 5624 8576 5652
rect 7239 5621 7251 5624
rect 7193 5615 7251 5621
rect 8570 5612 8576 5624
rect 8628 5612 8634 5664
rect 8662 5612 8668 5664
rect 8720 5652 8726 5664
rect 9214 5652 9220 5664
rect 8720 5624 8765 5652
rect 9175 5624 9220 5652
rect 8720 5612 8726 5624
rect 9214 5612 9220 5624
rect 9272 5612 9278 5664
rect 11885 5655 11943 5661
rect 11885 5652 11897 5655
rect 10796 5624 11897 5652
rect 1397 5587 1455 5593
rect 1397 5553 1409 5587
rect 1443 5584 1455 5587
rect 3050 5584 3056 5596
rect 1443 5556 3056 5584
rect 1443 5553 1455 5556
rect 1397 5547 1455 5553
rect 3050 5544 3056 5556
rect 3108 5584 3114 5596
rect 3329 5587 3387 5593
rect 3329 5584 3341 5587
rect 3108 5556 3341 5584
rect 3108 5544 3114 5556
rect 3329 5553 3341 5556
rect 3375 5553 3387 5587
rect 3510 5584 3516 5596
rect 3471 5556 3516 5584
rect 3329 5547 3387 5553
rect 3510 5544 3516 5556
rect 3568 5544 3574 5596
rect 4985 5587 5043 5593
rect 4985 5553 4997 5587
rect 5031 5584 5043 5587
rect 6730 5584 6736 5596
rect 5031 5556 6736 5584
rect 5031 5553 5043 5556
rect 4985 5547 5043 5553
rect 6730 5544 6736 5556
rect 6788 5544 6794 5596
rect 9493 5587 9551 5593
rect 9493 5553 9505 5587
rect 9539 5553 9551 5587
rect 9493 5547 9551 5553
rect 3418 5476 3424 5528
rect 3476 5516 3482 5528
rect 3697 5519 3755 5525
rect 3697 5516 3709 5519
rect 3476 5488 3709 5516
rect 3476 5476 3482 5488
rect 3697 5485 3709 5488
rect 3743 5516 3755 5519
rect 9306 5516 9312 5528
rect 3743 5488 9312 5516
rect 3743 5485 3755 5488
rect 3697 5479 3755 5485
rect 9306 5476 9312 5488
rect 9364 5476 9370 5528
rect 9398 5476 9404 5528
rect 9456 5516 9462 5528
rect 9508 5516 9536 5547
rect 9766 5544 9772 5596
rect 9824 5544 9830 5596
rect 9950 5544 9956 5596
rect 10008 5544 10014 5596
rect 9456 5488 9536 5516
rect 9456 5476 9462 5488
rect 9582 5476 9588 5528
rect 9640 5516 9646 5528
rect 9784 5516 9812 5544
rect 10796 5516 10824 5624
rect 11885 5621 11897 5624
rect 11931 5652 11943 5655
rect 12250 5652 12256 5664
rect 11931 5624 12256 5652
rect 11931 5621 11943 5624
rect 11885 5615 11943 5621
rect 12250 5612 12256 5624
rect 12308 5612 12314 5664
rect 12529 5655 12587 5661
rect 12529 5621 12541 5655
rect 12575 5652 12587 5655
rect 12728 5652 12756 5828
rect 13817 5825 13829 5859
rect 13863 5856 13875 5859
rect 14182 5856 14188 5868
rect 13863 5828 14188 5856
rect 13863 5825 13875 5828
rect 13817 5819 13875 5825
rect 14182 5816 14188 5828
rect 14240 5816 14246 5868
rect 15102 5720 15108 5732
rect 13832 5692 15108 5720
rect 13722 5652 13728 5664
rect 12575 5624 12756 5652
rect 13683 5624 13728 5652
rect 12575 5621 12587 5624
rect 12529 5615 12587 5621
rect 13722 5612 13728 5624
rect 13780 5612 13786 5664
rect 11606 5544 11612 5596
rect 11664 5584 11670 5596
rect 13832 5584 13860 5692
rect 15102 5680 15108 5692
rect 15160 5680 15166 5732
rect 11664 5556 13860 5584
rect 11664 5544 11670 5556
rect 14182 5544 14188 5596
rect 14240 5584 14246 5596
rect 14921 5587 14979 5593
rect 14921 5584 14933 5587
rect 14240 5556 14933 5584
rect 14240 5544 14246 5556
rect 14921 5553 14933 5556
rect 14967 5584 14979 5587
rect 15102 5584 15108 5596
rect 14967 5556 15108 5584
rect 14967 5553 14979 5556
rect 14921 5547 14979 5553
rect 15102 5544 15108 5556
rect 15160 5544 15166 5596
rect 10962 5516 10968 5528
rect 9640 5488 10824 5516
rect 10923 5488 10968 5516
rect 9640 5476 9646 5488
rect 10962 5476 10968 5488
rect 11020 5476 11026 5528
rect 11054 5476 11060 5528
rect 11112 5516 11118 5528
rect 11977 5519 12035 5525
rect 11977 5516 11989 5519
rect 11112 5488 11989 5516
rect 11112 5476 11118 5488
rect 11977 5485 11989 5488
rect 12023 5485 12035 5519
rect 15010 5516 15016 5528
rect 14971 5488 15016 5516
rect 11977 5479 12035 5485
rect 15010 5476 15016 5488
rect 15068 5476 15074 5528
rect 92 5426 15824 5448
rect 92 5374 5242 5426
rect 5294 5374 5306 5426
rect 5358 5374 5370 5426
rect 5422 5374 5434 5426
rect 5486 5374 10514 5426
rect 10566 5374 10578 5426
rect 10630 5374 10642 5426
rect 10694 5374 10706 5426
rect 10758 5374 15824 5426
rect 92 5352 15824 5374
rect 3053 5315 3111 5321
rect 3053 5312 3065 5315
rect 860 5284 3065 5312
rect 860 5253 888 5284
rect 3053 5281 3065 5284
rect 3099 5281 3111 5315
rect 5626 5312 5632 5324
rect 3053 5275 3111 5281
rect 3252 5284 5632 5312
rect 845 5247 903 5253
rect 845 5213 857 5247
rect 891 5213 903 5247
rect 845 5207 903 5213
rect 2498 5204 2504 5256
rect 2556 5244 2562 5256
rect 2593 5247 2651 5253
rect 2593 5244 2605 5247
rect 2556 5216 2605 5244
rect 2556 5204 2562 5216
rect 2593 5213 2605 5216
rect 2639 5213 2651 5247
rect 2593 5207 2651 5213
rect 1946 5136 1952 5188
rect 2004 5136 2010 5188
rect 566 5108 572 5120
rect 527 5080 572 5108
rect 566 5068 572 5080
rect 624 5068 630 5120
rect 2608 5040 2636 5207
rect 3252 5185 3280 5284
rect 5626 5272 5632 5284
rect 5684 5272 5690 5324
rect 5813 5315 5871 5321
rect 5813 5281 5825 5315
rect 5859 5312 5871 5315
rect 5994 5312 6000 5324
rect 5859 5284 6000 5312
rect 5859 5281 5871 5284
rect 5813 5275 5871 5281
rect 5994 5272 6000 5284
rect 6052 5272 6058 5324
rect 6270 5312 6276 5324
rect 6104 5284 6276 5312
rect 4430 5244 4436 5256
rect 3436 5216 4436 5244
rect 3436 5185 3464 5216
rect 4430 5204 4436 5216
rect 4488 5204 4494 5256
rect 3237 5179 3295 5185
rect 3237 5145 3249 5179
rect 3283 5145 3295 5179
rect 3237 5139 3295 5145
rect 3421 5179 3479 5185
rect 3421 5145 3433 5179
rect 3467 5145 3479 5179
rect 3970 5176 3976 5188
rect 3931 5148 3976 5176
rect 3421 5139 3479 5145
rect 3970 5136 3976 5148
rect 4028 5136 4034 5188
rect 4065 5179 4123 5185
rect 4065 5145 4077 5179
rect 4111 5176 4123 5179
rect 4154 5176 4160 5188
rect 4111 5148 4160 5176
rect 4111 5145 4123 5148
rect 4065 5139 4123 5145
rect 4154 5136 4160 5148
rect 4212 5136 4218 5188
rect 4249 5179 4307 5185
rect 4249 5145 4261 5179
rect 4295 5176 4307 5179
rect 4295 5148 5580 5176
rect 4295 5145 4307 5148
rect 4249 5139 4307 5145
rect 3510 5108 3516 5120
rect 3471 5080 3516 5108
rect 3510 5068 3516 5080
rect 3568 5068 3574 5120
rect 4264 5108 4292 5139
rect 4172 5080 4292 5108
rect 4709 5111 4767 5117
rect 4172 5040 4200 5080
rect 4709 5077 4721 5111
rect 4755 5077 4767 5111
rect 5552 5108 5580 5148
rect 5902 5136 5908 5188
rect 5960 5176 5966 5188
rect 6104 5185 6132 5284
rect 6270 5272 6276 5284
rect 6328 5272 6334 5324
rect 9398 5312 9404 5324
rect 9359 5284 9404 5312
rect 9398 5272 9404 5284
rect 9456 5272 9462 5324
rect 9861 5315 9919 5321
rect 9861 5281 9873 5315
rect 9907 5312 9919 5315
rect 11057 5315 11115 5321
rect 11057 5312 11069 5315
rect 9907 5284 11069 5312
rect 9907 5281 9919 5284
rect 9861 5275 9919 5281
rect 11057 5281 11069 5284
rect 11103 5281 11115 5315
rect 11057 5275 11115 5281
rect 11238 5272 11244 5324
rect 11296 5312 11302 5324
rect 11425 5315 11483 5321
rect 11425 5312 11437 5315
rect 11296 5284 11437 5312
rect 11296 5272 11302 5284
rect 11425 5281 11437 5284
rect 11471 5312 11483 5315
rect 14182 5312 14188 5324
rect 11471 5284 14188 5312
rect 11471 5281 11483 5284
rect 11425 5275 11483 5281
rect 14182 5272 14188 5284
rect 14240 5272 14246 5324
rect 14734 5272 14740 5324
rect 14792 5312 14798 5324
rect 14792 5284 15148 5312
rect 14792 5272 14798 5284
rect 6181 5247 6239 5253
rect 6181 5213 6193 5247
rect 6227 5244 6239 5247
rect 6914 5244 6920 5256
rect 6227 5216 6920 5244
rect 6227 5213 6239 5216
rect 6181 5207 6239 5213
rect 6914 5204 6920 5216
rect 6972 5244 6978 5256
rect 6972 5216 8340 5244
rect 6972 5204 6978 5216
rect 6089 5179 6147 5185
rect 6089 5176 6101 5179
rect 5960 5148 6101 5176
rect 5960 5136 5966 5148
rect 6089 5145 6101 5148
rect 6135 5145 6147 5179
rect 6270 5176 6276 5188
rect 6231 5148 6276 5176
rect 6089 5139 6147 5145
rect 6270 5136 6276 5148
rect 6328 5136 6334 5188
rect 6730 5136 6736 5188
rect 6788 5176 6794 5188
rect 8312 5185 8340 5216
rect 8938 5204 8944 5256
rect 8996 5244 9002 5256
rect 8996 5216 11928 5244
rect 8996 5204 9002 5216
rect 7285 5179 7343 5185
rect 7285 5176 7297 5179
rect 6788 5148 7297 5176
rect 6788 5136 6794 5148
rect 7285 5145 7297 5148
rect 7331 5145 7343 5179
rect 7285 5139 7343 5145
rect 8297 5179 8355 5185
rect 8297 5145 8309 5179
rect 8343 5145 8355 5179
rect 8478 5176 8484 5188
rect 8439 5148 8484 5176
rect 8297 5139 8355 5145
rect 8478 5136 8484 5148
rect 8536 5136 8542 5188
rect 8757 5179 8815 5185
rect 8757 5145 8769 5179
rect 8803 5176 8815 5179
rect 9030 5176 9036 5188
rect 8803 5148 9036 5176
rect 8803 5145 8815 5148
rect 8757 5139 8815 5145
rect 6362 5108 6368 5120
rect 5552 5080 6368 5108
rect 4709 5071 4767 5077
rect 2608 5012 4200 5040
rect 4614 5000 4620 5052
rect 4672 5040 4678 5052
rect 4724 5040 4752 5071
rect 6362 5068 6368 5080
rect 6420 5108 6426 5120
rect 6549 5111 6607 5117
rect 6549 5108 6561 5111
rect 6420 5080 6561 5108
rect 6420 5068 6426 5080
rect 6549 5077 6561 5080
rect 6595 5108 6607 5111
rect 6638 5108 6644 5120
rect 6595 5080 6644 5108
rect 6595 5077 6607 5080
rect 6549 5071 6607 5077
rect 6638 5068 6644 5080
rect 6696 5068 6702 5120
rect 7098 5108 7104 5120
rect 7059 5080 7104 5108
rect 7098 5068 7104 5080
rect 7156 5068 7162 5120
rect 7193 5111 7251 5117
rect 7193 5077 7205 5111
rect 7239 5077 7251 5111
rect 7374 5108 7380 5120
rect 7335 5080 7380 5108
rect 7193 5071 7251 5077
rect 7208 5040 7236 5071
rect 7374 5068 7380 5080
rect 7432 5068 7438 5120
rect 7561 5111 7619 5117
rect 7561 5077 7573 5111
rect 7607 5108 7619 5111
rect 8772 5108 8800 5139
rect 9030 5136 9036 5148
rect 9088 5136 9094 5188
rect 9769 5179 9827 5185
rect 9769 5145 9781 5179
rect 9815 5176 9827 5179
rect 10962 5176 10968 5188
rect 9815 5148 10968 5176
rect 9815 5145 9827 5148
rect 9769 5139 9827 5145
rect 10962 5136 10968 5148
rect 11020 5136 11026 5188
rect 11517 5179 11575 5185
rect 11517 5145 11529 5179
rect 11563 5176 11575 5179
rect 11790 5176 11796 5188
rect 11563 5148 11796 5176
rect 11563 5145 11575 5148
rect 11517 5139 11575 5145
rect 11790 5136 11796 5148
rect 11848 5136 11854 5188
rect 7607 5080 8800 5108
rect 7607 5077 7619 5080
rect 7561 5071 7619 5077
rect 9122 5068 9128 5120
rect 9180 5108 9186 5120
rect 9858 5108 9864 5120
rect 9180 5080 9864 5108
rect 9180 5068 9186 5080
rect 9858 5068 9864 5080
rect 9916 5068 9922 5120
rect 10045 5111 10103 5117
rect 10045 5077 10057 5111
rect 10091 5077 10103 5111
rect 10045 5071 10103 5077
rect 11701 5111 11759 5117
rect 11701 5077 11713 5111
rect 11747 5108 11759 5111
rect 11900 5108 11928 5216
rect 12434 5204 12440 5256
rect 12492 5244 12498 5256
rect 12805 5247 12863 5253
rect 12805 5244 12817 5247
rect 12492 5216 12817 5244
rect 12492 5204 12498 5216
rect 12805 5213 12817 5216
rect 12851 5213 12863 5247
rect 12805 5207 12863 5213
rect 13446 5204 13452 5256
rect 13504 5204 13510 5256
rect 14826 5244 14832 5256
rect 14108 5216 14832 5244
rect 12342 5108 12348 5120
rect 11747 5080 12348 5108
rect 11747 5077 11759 5080
rect 11701 5071 11759 5077
rect 8846 5040 8852 5052
rect 4672 5012 8852 5040
rect 4672 5000 4678 5012
rect 8846 5000 8852 5012
rect 8904 5000 8910 5052
rect 8941 5043 8999 5049
rect 8941 5009 8953 5043
rect 8987 5040 8999 5043
rect 8987 5012 9352 5040
rect 8987 5009 8999 5012
rect 8941 5003 8999 5009
rect 6178 4932 6184 4984
rect 6236 4972 6242 4984
rect 6457 4975 6515 4981
rect 6457 4972 6469 4975
rect 6236 4944 6469 4972
rect 6236 4932 6242 4944
rect 6457 4941 6469 4944
rect 6503 4941 6515 4975
rect 6457 4935 6515 4941
rect 8754 4932 8760 4984
rect 8812 4972 8818 4984
rect 9214 4972 9220 4984
rect 8812 4944 9220 4972
rect 8812 4932 8818 4944
rect 9214 4932 9220 4944
rect 9272 4932 9278 4984
rect 9324 4972 9352 5012
rect 10060 4972 10088 5071
rect 12342 5068 12348 5080
rect 12400 5068 12406 5120
rect 12526 5108 12532 5120
rect 12487 5080 12532 5108
rect 12526 5068 12532 5080
rect 12584 5068 12590 5120
rect 14108 5108 14136 5216
rect 14826 5204 14832 5216
rect 14884 5244 14890 5256
rect 15120 5253 15148 5284
rect 14921 5247 14979 5253
rect 14921 5244 14933 5247
rect 14884 5216 14933 5244
rect 14884 5204 14890 5216
rect 14921 5213 14933 5216
rect 14967 5213 14979 5247
rect 14921 5207 14979 5213
rect 15105 5247 15163 5253
rect 15105 5213 15117 5247
rect 15151 5244 15163 5247
rect 15286 5244 15292 5256
rect 15151 5216 15292 5244
rect 15151 5213 15163 5216
rect 15105 5207 15163 5213
rect 15286 5204 15292 5216
rect 15344 5204 15350 5256
rect 14734 5176 14740 5188
rect 14292 5148 14740 5176
rect 14292 5117 14320 5148
rect 14734 5136 14740 5148
rect 14792 5136 14798 5188
rect 12636 5080 14136 5108
rect 14277 5111 14335 5117
rect 10134 5000 10140 5052
rect 10192 5040 10198 5052
rect 12636 5040 12664 5080
rect 14277 5077 14289 5111
rect 14323 5077 14335 5111
rect 14277 5071 14335 5077
rect 10192 5012 12664 5040
rect 10192 5000 10198 5012
rect 12342 4972 12348 4984
rect 9324 4944 12348 4972
rect 12342 4932 12348 4944
rect 12400 4932 12406 4984
rect 92 4882 15824 4904
rect 92 4830 2606 4882
rect 2658 4830 2670 4882
rect 2722 4830 2734 4882
rect 2786 4830 2798 4882
rect 2850 4830 7878 4882
rect 7930 4830 7942 4882
rect 7994 4830 8006 4882
rect 8058 4830 8070 4882
rect 8122 4830 13150 4882
rect 13202 4830 13214 4882
rect 13266 4830 13278 4882
rect 13330 4830 13342 4882
rect 13394 4830 15824 4882
rect 92 4808 15824 4830
rect 2148 4740 2774 4768
rect 750 4700 756 4712
rect 711 4672 756 4700
rect 750 4660 756 4672
rect 808 4660 814 4712
rect 1673 4635 1731 4641
rect 1673 4601 1685 4635
rect 1719 4632 1731 4635
rect 2038 4632 2044 4644
rect 1719 4604 2044 4632
rect 1719 4601 1731 4604
rect 1673 4595 1731 4601
rect 2038 4592 2044 4604
rect 2096 4592 2102 4644
rect 2148 4641 2176 4740
rect 2746 4700 2774 4740
rect 3510 4728 3516 4780
rect 3568 4768 3574 4780
rect 4985 4771 5043 4777
rect 4985 4768 4997 4771
rect 3568 4740 4997 4768
rect 3568 4728 3574 4740
rect 4985 4737 4997 4740
rect 5031 4737 5043 4771
rect 4985 4731 5043 4737
rect 5534 4728 5540 4780
rect 5592 4768 5598 4780
rect 6270 4768 6276 4780
rect 5592 4740 6276 4768
rect 5592 4728 5598 4740
rect 6270 4728 6276 4740
rect 6328 4728 6334 4780
rect 8478 4728 8484 4780
rect 8536 4768 8542 4780
rect 8536 4740 10272 4768
rect 8536 4728 8542 4740
rect 10244 4700 10272 4740
rect 10318 4728 10324 4780
rect 10376 4768 10382 4780
rect 11054 4768 11060 4780
rect 10376 4740 11060 4768
rect 10376 4728 10382 4740
rect 11054 4728 11060 4740
rect 11112 4728 11118 4780
rect 11238 4768 11244 4780
rect 11199 4740 11244 4768
rect 11238 4728 11244 4740
rect 11296 4728 11302 4780
rect 12805 4771 12863 4777
rect 12805 4737 12817 4771
rect 12851 4768 12863 4771
rect 13538 4768 13544 4780
rect 12851 4740 13544 4768
rect 12851 4737 12863 4740
rect 12805 4731 12863 4737
rect 13538 4728 13544 4740
rect 13596 4728 13602 4780
rect 14185 4771 14243 4777
rect 14185 4737 14197 4771
rect 14231 4768 14243 4771
rect 14642 4768 14648 4780
rect 14231 4740 14648 4768
rect 14231 4737 14243 4740
rect 14185 4731 14243 4737
rect 14642 4728 14648 4740
rect 14700 4728 14706 4780
rect 11793 4703 11851 4709
rect 11793 4700 11805 4703
rect 2746 4672 8892 4700
rect 10244 4672 11805 4700
rect 2133 4635 2191 4641
rect 2133 4601 2145 4635
rect 2179 4601 2191 4635
rect 2133 4595 2191 4601
rect 3881 4635 3939 4641
rect 3881 4601 3893 4635
rect 3927 4632 3939 4635
rect 4430 4632 4436 4644
rect 3927 4604 4436 4632
rect 3927 4601 3939 4604
rect 3881 4595 3939 4601
rect 4430 4592 4436 4604
rect 4488 4592 4494 4644
rect 5629 4635 5687 4641
rect 5629 4601 5641 4635
rect 5675 4632 5687 4635
rect 5994 4632 6000 4644
rect 5675 4604 6000 4632
rect 5675 4601 5687 4604
rect 5629 4595 5687 4601
rect 5994 4592 6000 4604
rect 6052 4592 6058 4644
rect 6917 4635 6975 4641
rect 6917 4601 6929 4635
rect 6963 4632 6975 4635
rect 8386 4632 8392 4644
rect 6963 4604 8392 4632
rect 6963 4601 6975 4604
rect 6917 4595 6975 4601
rect 8386 4592 8392 4604
rect 8444 4592 8450 4644
rect 8754 4632 8760 4644
rect 8715 4604 8760 4632
rect 8754 4592 8760 4604
rect 8812 4592 8818 4644
rect 8864 4632 8892 4672
rect 11793 4669 11805 4672
rect 11839 4669 11851 4703
rect 11793 4663 11851 4669
rect 13630 4660 13636 4712
rect 13688 4700 13694 4712
rect 14737 4703 14795 4709
rect 14737 4700 14749 4703
rect 13688 4672 14749 4700
rect 13688 4660 13694 4672
rect 14737 4669 14749 4672
rect 14783 4669 14795 4703
rect 14737 4663 14795 4669
rect 8864 4604 10272 4632
rect 934 4564 940 4576
rect 895 4536 940 4564
rect 934 4524 940 4536
rect 992 4524 998 4576
rect 1765 4567 1823 4573
rect 1765 4533 1777 4567
rect 1811 4564 1823 4567
rect 3142 4564 3148 4576
rect 1811 4536 3148 4564
rect 1811 4533 1823 4536
rect 1765 4527 1823 4533
rect 3142 4524 3148 4536
rect 3200 4524 3206 4576
rect 3697 4567 3755 4573
rect 3697 4533 3709 4567
rect 3743 4564 3755 4567
rect 3970 4564 3976 4576
rect 3743 4536 3976 4564
rect 3743 4533 3755 4536
rect 3697 4527 3755 4533
rect 3970 4524 3976 4536
rect 4028 4524 4034 4576
rect 6086 4524 6092 4576
rect 6144 4564 6150 4576
rect 6825 4567 6883 4573
rect 6825 4564 6837 4567
rect 6144 4536 6837 4564
rect 6144 4524 6150 4536
rect 6825 4533 6837 4536
rect 6871 4533 6883 4567
rect 6825 4527 6883 4533
rect 7009 4567 7067 4573
rect 7009 4533 7021 4567
rect 7055 4533 7067 4567
rect 7009 4527 7067 4533
rect 7101 4567 7159 4573
rect 7101 4533 7113 4567
rect 7147 4564 7159 4567
rect 10244 4564 10272 4604
rect 10870 4592 10876 4644
rect 10928 4632 10934 4644
rect 10928 4604 12020 4632
rect 10928 4592 10934 4604
rect 11790 4564 11796 4576
rect 7147 4536 8800 4564
rect 10244 4536 11284 4564
rect 11751 4536 11796 4564
rect 7147 4533 7159 4536
rect 7101 4527 7159 4533
rect 1394 4456 1400 4508
rect 1452 4496 1458 4508
rect 2041 4499 2099 4505
rect 2041 4496 2053 4499
rect 1452 4468 2053 4496
rect 1452 4456 1458 4468
rect 2041 4465 2053 4468
rect 2087 4465 2099 4499
rect 2041 4459 2099 4465
rect 4430 4456 4436 4508
rect 4488 4496 4494 4508
rect 5445 4499 5503 4505
rect 5445 4496 5457 4499
rect 4488 4468 5457 4496
rect 4488 4456 4494 4468
rect 5445 4465 5457 4468
rect 5491 4496 5503 4499
rect 5718 4496 5724 4508
rect 5491 4468 5724 4496
rect 5491 4465 5503 4468
rect 5445 4459 5503 4465
rect 5718 4456 5724 4468
rect 5776 4456 5782 4508
rect 7024 4496 7052 4527
rect 7190 4496 7196 4508
rect 7024 4468 7196 4496
rect 7190 4456 7196 4468
rect 7248 4456 7254 4508
rect 1210 4388 1216 4440
rect 1268 4428 1274 4440
rect 1489 4431 1547 4437
rect 1489 4428 1501 4431
rect 1268 4400 1501 4428
rect 1268 4388 1274 4400
rect 1489 4397 1501 4400
rect 1535 4397 1547 4431
rect 1489 4391 1547 4397
rect 1670 4388 1676 4440
rect 1728 4428 1734 4440
rect 3237 4431 3295 4437
rect 3237 4428 3249 4431
rect 1728 4400 3249 4428
rect 1728 4388 1734 4400
rect 3237 4397 3249 4400
rect 3283 4397 3295 4431
rect 3602 4428 3608 4440
rect 3563 4400 3608 4428
rect 3237 4391 3295 4397
rect 3602 4388 3608 4400
rect 3660 4388 3666 4440
rect 4706 4388 4712 4440
rect 4764 4428 4770 4440
rect 5353 4431 5411 4437
rect 5353 4428 5365 4431
rect 4764 4400 5365 4428
rect 4764 4388 4770 4400
rect 5353 4397 5365 4400
rect 5399 4397 5411 4431
rect 5353 4391 5411 4397
rect 6641 4431 6699 4437
rect 6641 4397 6653 4431
rect 6687 4428 6699 4431
rect 6730 4428 6736 4440
rect 6687 4400 6736 4428
rect 6687 4397 6699 4400
rect 6641 4391 6699 4397
rect 6730 4388 6736 4400
rect 6788 4388 6794 4440
rect 8772 4428 8800 4536
rect 9030 4496 9036 4508
rect 8991 4468 9036 4496
rect 9030 4456 9036 4468
rect 9088 4456 9094 4508
rect 9674 4456 9680 4508
rect 9732 4456 9738 4508
rect 10965 4499 11023 4505
rect 10965 4465 10977 4499
rect 11011 4465 11023 4499
rect 11146 4496 11152 4508
rect 11107 4468 11152 4496
rect 10965 4459 11023 4465
rect 10318 4428 10324 4440
rect 8772 4400 10324 4428
rect 10318 4388 10324 4400
rect 10376 4388 10382 4440
rect 10410 4388 10416 4440
rect 10468 4428 10474 4440
rect 10505 4431 10563 4437
rect 10505 4428 10517 4431
rect 10468 4400 10517 4428
rect 10468 4388 10474 4400
rect 10505 4397 10517 4400
rect 10551 4397 10563 4431
rect 10505 4391 10563 4397
rect 10870 4388 10876 4440
rect 10928 4428 10934 4440
rect 10980 4428 11008 4459
rect 11146 4456 11152 4468
rect 11204 4456 11210 4508
rect 11256 4496 11284 4536
rect 11790 4524 11796 4536
rect 11848 4524 11854 4576
rect 11992 4573 12020 4604
rect 11977 4567 12035 4573
rect 11977 4533 11989 4567
rect 12023 4533 12035 4567
rect 11977 4527 12035 4533
rect 12342 4524 12348 4576
rect 12400 4564 12406 4576
rect 12529 4567 12587 4573
rect 12529 4564 12541 4567
rect 12400 4536 12541 4564
rect 12400 4524 12406 4536
rect 12529 4533 12541 4536
rect 12575 4533 12587 4567
rect 12529 4527 12587 4533
rect 11698 4496 11704 4508
rect 11256 4468 11704 4496
rect 11698 4456 11704 4468
rect 11756 4456 11762 4508
rect 12544 4496 12572 4527
rect 12618 4524 12624 4576
rect 12676 4564 12682 4576
rect 14093 4567 14151 4573
rect 14093 4564 14105 4567
rect 12676 4536 14105 4564
rect 12676 4524 12682 4536
rect 14093 4533 14105 4536
rect 14139 4533 14151 4567
rect 14734 4564 14740 4576
rect 14695 4536 14740 4564
rect 14093 4527 14151 4533
rect 14734 4524 14740 4536
rect 14792 4524 14798 4576
rect 14826 4524 14832 4576
rect 14884 4564 14890 4576
rect 14921 4567 14979 4573
rect 14921 4564 14933 4567
rect 14884 4536 14933 4564
rect 14884 4524 14890 4536
rect 14921 4533 14933 4536
rect 14967 4533 14979 4567
rect 14921 4527 14979 4533
rect 15010 4524 15016 4576
rect 15068 4564 15074 4576
rect 15068 4536 15113 4564
rect 15068 4524 15074 4536
rect 12710 4496 12716 4508
rect 12544 4468 12716 4496
rect 12710 4456 12716 4468
rect 12768 4456 12774 4508
rect 12805 4499 12863 4505
rect 12805 4465 12817 4499
rect 12851 4496 12863 4499
rect 13909 4499 13967 4505
rect 13909 4496 13921 4499
rect 12851 4468 13921 4496
rect 12851 4465 12863 4468
rect 12805 4459 12863 4465
rect 13909 4465 13921 4468
rect 13955 4496 13967 4499
rect 14182 4496 14188 4508
rect 13955 4468 14188 4496
rect 13955 4465 13967 4468
rect 13909 4459 13967 4465
rect 14182 4456 14188 4468
rect 14240 4456 14246 4508
rect 10928 4400 11008 4428
rect 10928 4388 10934 4400
rect 14458 4388 14464 4440
rect 14516 4428 14522 4440
rect 14826 4428 14832 4440
rect 14516 4400 14832 4428
rect 14516 4388 14522 4400
rect 14826 4388 14832 4400
rect 14884 4388 14890 4440
rect 92 4338 15824 4360
rect 92 4286 5242 4338
rect 5294 4286 5306 4338
rect 5358 4286 5370 4338
rect 5422 4286 5434 4338
rect 5486 4286 10514 4338
rect 10566 4286 10578 4338
rect 10630 4286 10642 4338
rect 10694 4286 10706 4338
rect 10758 4286 15824 4338
rect 92 4264 15824 4286
rect 1946 4184 1952 4236
rect 2004 4184 2010 4236
rect 3142 4224 3148 4236
rect 3103 4196 3148 4224
rect 3142 4184 3148 4196
rect 3200 4184 3206 4236
rect 3602 4184 3608 4236
rect 3660 4224 3666 4236
rect 4065 4227 4123 4233
rect 4065 4224 4077 4227
rect 3660 4196 4077 4224
rect 3660 4184 3666 4196
rect 4065 4193 4077 4196
rect 4111 4193 4123 4227
rect 4065 4187 4123 4193
rect 4614 4184 4620 4236
rect 4672 4184 4678 4236
rect 4706 4184 4712 4236
rect 4764 4224 4770 4236
rect 7098 4224 7104 4236
rect 4764 4196 7104 4224
rect 4764 4184 4770 4196
rect 7098 4184 7104 4196
rect 7156 4224 7162 4236
rect 8205 4227 8263 4233
rect 8205 4224 8217 4227
rect 7156 4196 7420 4224
rect 7156 4184 7162 4196
rect 1964 4142 1992 4184
rect 4632 4156 4660 4184
rect 5902 4156 5908 4168
rect 4540 4128 4660 4156
rect 4724 4128 5908 4156
rect 3329 4091 3387 4097
rect 3329 4057 3341 4091
rect 3375 4088 3387 4091
rect 3418 4088 3424 4100
rect 3375 4060 3424 4088
rect 3375 4057 3387 4060
rect 3329 4051 3387 4057
rect 3418 4048 3424 4060
rect 3476 4048 3482 4100
rect 4540 4097 4568 4128
rect 4724 4097 4752 4128
rect 5902 4116 5908 4128
rect 5960 4116 5966 4168
rect 7392 4165 7420 4196
rect 7576 4196 8217 4224
rect 7576 4165 7604 4196
rect 8205 4193 8217 4196
rect 8251 4193 8263 4227
rect 8205 4187 8263 4193
rect 9030 4184 9036 4236
rect 9088 4224 9094 4236
rect 9401 4227 9459 4233
rect 9401 4224 9413 4227
rect 9088 4196 9413 4224
rect 9088 4184 9094 4196
rect 9401 4193 9413 4196
rect 9447 4193 9459 4227
rect 11790 4224 11796 4236
rect 9401 4187 9459 4193
rect 9600 4196 11796 4224
rect 7377 4159 7435 4165
rect 7377 4125 7389 4159
rect 7423 4125 7435 4159
rect 7377 4119 7435 4125
rect 7561 4159 7619 4165
rect 7561 4125 7573 4159
rect 7607 4125 7619 4159
rect 7561 4119 7619 4125
rect 8478 4116 8484 4168
rect 8536 4156 8542 4168
rect 8573 4159 8631 4165
rect 8573 4156 8585 4159
rect 8536 4128 8585 4156
rect 8536 4116 8542 4128
rect 8573 4125 8585 4128
rect 8619 4156 8631 4159
rect 8662 4156 8668 4168
rect 8619 4128 8668 4156
rect 8619 4125 8631 4128
rect 8573 4119 8631 4125
rect 8662 4116 8668 4128
rect 8720 4156 8726 4168
rect 9600 4156 9628 4196
rect 11790 4184 11796 4196
rect 11848 4184 11854 4236
rect 12618 4224 12624 4236
rect 12406 4196 12624 4224
rect 9766 4156 9772 4168
rect 8720 4128 9628 4156
rect 9727 4128 9772 4156
rect 8720 4116 8726 4128
rect 9766 4116 9772 4128
rect 9824 4156 9830 4168
rect 12406 4156 12434 4196
rect 12618 4184 12624 4196
rect 12676 4184 12682 4236
rect 14182 4184 14188 4236
rect 14240 4224 14246 4236
rect 14277 4227 14335 4233
rect 14277 4224 14289 4227
rect 14240 4196 14289 4224
rect 14240 4184 14246 4196
rect 14277 4193 14289 4196
rect 14323 4193 14335 4227
rect 14277 4187 14335 4193
rect 9824 4128 12434 4156
rect 9824 4116 9830 4128
rect 13446 4116 13452 4168
rect 13504 4116 13510 4168
rect 14642 4116 14648 4168
rect 14700 4156 14706 4168
rect 14921 4159 14979 4165
rect 14921 4156 14933 4159
rect 14700 4128 14933 4156
rect 14700 4116 14706 4128
rect 14921 4125 14933 4128
rect 14967 4125 14979 4159
rect 14921 4119 14979 4125
rect 4341 4091 4399 4097
rect 4341 4088 4353 4091
rect 3528 4060 4353 4088
rect 566 3980 572 4032
rect 624 4020 630 4032
rect 750 4020 756 4032
rect 624 3992 756 4020
rect 624 3980 630 3992
rect 750 3980 756 3992
rect 808 4020 814 4032
rect 845 4023 903 4029
rect 845 4020 857 4023
rect 808 3992 857 4020
rect 808 3980 814 3992
rect 845 3989 857 3992
rect 891 3989 903 4023
rect 1118 4020 1124 4032
rect 1079 3992 1124 4020
rect 845 3983 903 3989
rect 1118 3980 1124 3992
rect 1176 3980 1182 4032
rect 2130 3980 2136 4032
rect 2188 4020 2194 4032
rect 3528 4020 3556 4060
rect 4341 4057 4353 4060
rect 4387 4057 4399 4091
rect 4341 4051 4399 4057
rect 4433 4091 4491 4097
rect 4433 4057 4445 4091
rect 4479 4057 4491 4091
rect 4433 4051 4491 4057
rect 4525 4091 4583 4097
rect 4525 4057 4537 4091
rect 4571 4057 4583 4091
rect 4525 4051 4583 4057
rect 4709 4091 4767 4097
rect 4709 4057 4721 4091
rect 4755 4057 4767 4091
rect 4709 4051 4767 4057
rect 2188 3992 3556 4020
rect 3605 4023 3663 4029
rect 2188 3980 2194 3992
rect 3605 3989 3617 4023
rect 3651 4020 3663 4023
rect 3970 4020 3976 4032
rect 3651 3992 3976 4020
rect 3651 3989 3663 3992
rect 3605 3983 3663 3989
rect 3970 3980 3976 3992
rect 4028 3980 4034 4032
rect 4448 4020 4476 4051
rect 4890 4048 4896 4100
rect 4948 4088 4954 4100
rect 5997 4091 6055 4097
rect 5997 4088 6009 4091
rect 4948 4060 6009 4088
rect 4948 4048 4954 4060
rect 5997 4057 6009 4060
rect 6043 4088 6055 4091
rect 6086 4088 6092 4100
rect 6043 4060 6092 4088
rect 6043 4057 6055 4060
rect 5997 4051 6055 4057
rect 6086 4048 6092 4060
rect 6144 4048 6150 4100
rect 6181 4091 6239 4097
rect 6181 4057 6193 4091
rect 6227 4088 6239 4091
rect 6362 4088 6368 4100
rect 6227 4060 6368 4088
rect 6227 4057 6239 4060
rect 6181 4051 6239 4057
rect 6362 4048 6368 4060
rect 6420 4048 6426 4100
rect 9122 4088 9128 4100
rect 8680 4060 9128 4088
rect 6270 4020 6276 4032
rect 4448 3992 6276 4020
rect 6270 3980 6276 3992
rect 6328 4020 6334 4032
rect 8680 4029 8708 4060
rect 9122 4048 9128 4060
rect 9180 4048 9186 4100
rect 9306 4048 9312 4100
rect 9364 4088 9370 4100
rect 9585 4091 9643 4097
rect 9585 4088 9597 4091
rect 9364 4060 9597 4088
rect 9364 4048 9370 4060
rect 9585 4057 9597 4060
rect 9631 4057 9643 4091
rect 9585 4051 9643 4057
rect 9674 4048 9680 4100
rect 9732 4088 9738 4100
rect 9907 4091 9965 4097
rect 9732 4060 9777 4088
rect 9732 4048 9738 4060
rect 9907 4057 9919 4091
rect 9953 4088 9965 4091
rect 10134 4088 10140 4100
rect 9953 4060 10140 4088
rect 9953 4057 9965 4060
rect 9907 4051 9965 4057
rect 10134 4048 10140 4060
rect 10192 4048 10198 4100
rect 11057 4091 11115 4097
rect 11057 4057 11069 4091
rect 11103 4057 11115 4091
rect 11057 4051 11115 4057
rect 8665 4023 8723 4029
rect 8665 4020 8677 4023
rect 6328 3992 8677 4020
rect 6328 3980 6334 3992
rect 8665 3989 8677 3992
rect 8711 3989 8723 4023
rect 8665 3983 8723 3989
rect 8849 4023 8907 4029
rect 8849 3989 8861 4023
rect 8895 4020 8907 4023
rect 8938 4020 8944 4032
rect 8895 3992 8944 4020
rect 8895 3989 8907 3992
rect 8849 3983 8907 3989
rect 8938 3980 8944 3992
rect 8996 3980 9002 4032
rect 10045 4023 10103 4029
rect 10045 3989 10057 4023
rect 10091 4020 10103 4023
rect 10962 4020 10968 4032
rect 10091 3992 10968 4020
rect 10091 3989 10103 3992
rect 10045 3983 10103 3989
rect 10962 3980 10968 3992
rect 11020 3980 11026 4032
rect 11072 3964 11100 4051
rect 11606 4048 11612 4100
rect 11664 4088 11670 4100
rect 11885 4091 11943 4097
rect 11885 4088 11897 4091
rect 11664 4060 11897 4088
rect 11664 4048 11670 4060
rect 11885 4057 11897 4060
rect 11931 4057 11943 4091
rect 12066 4088 12072 4100
rect 12027 4060 12072 4088
rect 11885 4051 11943 4057
rect 12066 4048 12072 4060
rect 12124 4048 12130 4100
rect 12526 4088 12532 4100
rect 12487 4060 12532 4088
rect 12526 4048 12532 4060
rect 12584 4048 12590 4100
rect 12342 3980 12348 4032
rect 12400 4020 12406 4032
rect 12544 4020 12572 4048
rect 12400 3992 12572 4020
rect 12805 4023 12863 4029
rect 12400 3980 12406 3992
rect 12805 3989 12817 4023
rect 12851 4020 12863 4023
rect 13998 4020 14004 4032
rect 12851 3992 14004 4020
rect 12851 3989 12863 3992
rect 12805 3983 12863 3989
rect 13998 3980 14004 3992
rect 14056 3980 14062 4032
rect 15105 4023 15163 4029
rect 15105 3989 15117 4023
rect 15151 4020 15163 4023
rect 15470 4020 15476 4032
rect 15151 3992 15476 4020
rect 15151 3989 15163 3992
rect 15105 3983 15163 3989
rect 15470 3980 15476 3992
rect 15528 3980 15534 4032
rect 6365 3955 6423 3961
rect 6365 3921 6377 3955
rect 6411 3952 6423 3955
rect 7374 3952 7380 3964
rect 6411 3924 7380 3952
rect 6411 3921 6423 3924
rect 6365 3915 6423 3921
rect 7374 3912 7380 3924
rect 7432 3912 7438 3964
rect 7745 3955 7803 3961
rect 7745 3921 7757 3955
rect 7791 3952 7803 3955
rect 11054 3952 11060 3964
rect 7791 3924 11060 3952
rect 7791 3921 7803 3924
rect 7745 3915 7803 3921
rect 11054 3912 11060 3924
rect 11112 3912 11118 3964
rect 2593 3887 2651 3893
rect 2593 3853 2605 3887
rect 2639 3884 2651 3887
rect 3142 3884 3148 3896
rect 2639 3856 3148 3884
rect 2639 3853 2651 3856
rect 2593 3847 2651 3853
rect 3142 3844 3148 3856
rect 3200 3844 3206 3896
rect 3513 3887 3571 3893
rect 3513 3853 3525 3887
rect 3559 3884 3571 3887
rect 5902 3884 5908 3896
rect 3559 3856 5908 3884
rect 3559 3853 3571 3856
rect 3513 3847 3571 3853
rect 5902 3844 5908 3856
rect 5960 3844 5966 3896
rect 6178 3884 6184 3896
rect 6139 3856 6184 3884
rect 6178 3844 6184 3856
rect 6236 3844 6242 3896
rect 10962 3844 10968 3896
rect 11020 3884 11026 3896
rect 11241 3887 11299 3893
rect 11241 3884 11253 3887
rect 11020 3856 11253 3884
rect 11020 3844 11026 3856
rect 11241 3853 11253 3856
rect 11287 3853 11299 3887
rect 11241 3847 11299 3853
rect 12069 3887 12127 3893
rect 12069 3853 12081 3887
rect 12115 3884 12127 3887
rect 12250 3884 12256 3896
rect 12115 3856 12256 3884
rect 12115 3853 12127 3856
rect 12069 3847 12127 3853
rect 12250 3844 12256 3856
rect 12308 3844 12314 3896
rect 92 3794 15824 3816
rect 92 3742 2606 3794
rect 2658 3742 2670 3794
rect 2722 3742 2734 3794
rect 2786 3742 2798 3794
rect 2850 3742 7878 3794
rect 7930 3742 7942 3794
rect 7994 3742 8006 3794
rect 8058 3742 8070 3794
rect 8122 3742 13150 3794
rect 13202 3742 13214 3794
rect 13266 3742 13278 3794
rect 13330 3742 13342 3794
rect 13394 3742 15824 3794
rect 92 3720 15824 3742
rect 842 3680 848 3692
rect 803 3652 848 3680
rect 842 3640 848 3652
rect 900 3640 906 3692
rect 2038 3640 2044 3692
rect 2096 3680 2102 3692
rect 2225 3683 2283 3689
rect 2225 3680 2237 3683
rect 2096 3652 2237 3680
rect 2096 3640 2102 3652
rect 2225 3649 2237 3652
rect 2271 3649 2283 3683
rect 2225 3643 2283 3649
rect 3513 3683 3571 3689
rect 3513 3649 3525 3683
rect 3559 3680 3571 3683
rect 4154 3680 4160 3692
rect 3559 3652 4160 3680
rect 3559 3649 3571 3652
rect 3513 3643 3571 3649
rect 4154 3640 4160 3652
rect 4212 3680 4218 3692
rect 4249 3683 4307 3689
rect 4249 3680 4261 3683
rect 4212 3652 4261 3680
rect 4212 3640 4218 3652
rect 4249 3649 4261 3652
rect 4295 3649 4307 3683
rect 4249 3643 4307 3649
rect 5074 3640 5080 3692
rect 5132 3680 5138 3692
rect 5353 3683 5411 3689
rect 5353 3680 5365 3683
rect 5132 3652 5365 3680
rect 5132 3640 5138 3652
rect 5353 3649 5365 3652
rect 5399 3649 5411 3683
rect 5353 3643 5411 3649
rect 5902 3640 5908 3692
rect 5960 3680 5966 3692
rect 6825 3683 6883 3689
rect 6825 3680 6837 3683
rect 5960 3652 6837 3680
rect 5960 3640 5966 3652
rect 6825 3649 6837 3652
rect 6871 3649 6883 3683
rect 11330 3680 11336 3692
rect 6825 3643 6883 3649
rect 6932 3652 11336 3680
rect 1673 3615 1731 3621
rect 1673 3581 1685 3615
rect 1719 3612 1731 3615
rect 1719 3584 3485 3612
rect 1719 3581 1731 3584
rect 1673 3575 1731 3581
rect 3142 3544 3148 3556
rect 1504 3516 3148 3544
rect 1504 3485 1532 3516
rect 3142 3504 3148 3516
rect 3200 3504 3206 3556
rect 3457 3544 3485 3584
rect 4062 3572 4068 3624
rect 4120 3612 4126 3624
rect 6932 3612 6960 3652
rect 11330 3640 11336 3652
rect 11388 3640 11394 3692
rect 12066 3640 12072 3692
rect 12124 3680 12130 3692
rect 14645 3683 14703 3689
rect 14645 3680 14657 3683
rect 12124 3652 14657 3680
rect 12124 3640 12130 3652
rect 14645 3649 14657 3652
rect 14691 3649 14703 3683
rect 14645 3643 14703 3649
rect 4120 3584 6960 3612
rect 4120 3572 4126 3584
rect 7834 3572 7840 3624
rect 7892 3612 7898 3624
rect 8938 3612 8944 3624
rect 7892 3584 8944 3612
rect 7892 3572 7898 3584
rect 8938 3572 8944 3584
rect 8996 3572 9002 3624
rect 9306 3572 9312 3624
rect 9364 3612 9370 3624
rect 11149 3615 11207 3621
rect 11149 3612 11161 3615
rect 9364 3584 11161 3612
rect 9364 3572 9370 3584
rect 11149 3581 11161 3584
rect 11195 3612 11207 3615
rect 11238 3612 11244 3624
rect 11195 3584 11244 3612
rect 11195 3581 11207 3584
rect 11149 3575 11207 3581
rect 11238 3572 11244 3584
rect 11296 3572 11302 3624
rect 12434 3612 12440 3624
rect 11992 3584 12440 3612
rect 4890 3544 4896 3556
rect 3457 3516 4896 3544
rect 1489 3479 1547 3485
rect 1489 3445 1501 3479
rect 1535 3445 1547 3479
rect 1489 3439 1547 3445
rect 2222 3436 2228 3488
rect 2280 3476 2286 3488
rect 2317 3479 2375 3485
rect 2317 3476 2329 3479
rect 2280 3448 2329 3476
rect 2280 3436 2286 3448
rect 2317 3445 2329 3448
rect 2363 3445 2375 3479
rect 3457 3476 3485 3516
rect 4890 3504 4896 3516
rect 4948 3504 4954 3556
rect 4982 3504 4988 3556
rect 5040 3544 5046 3556
rect 5261 3547 5319 3553
rect 5261 3544 5273 3547
rect 5040 3516 5273 3544
rect 5040 3504 5046 3516
rect 5261 3513 5273 3516
rect 5307 3513 5319 3547
rect 5261 3507 5319 3513
rect 5353 3547 5411 3553
rect 5353 3513 5365 3547
rect 5399 3544 5411 3547
rect 5810 3544 5816 3556
rect 5399 3516 5816 3544
rect 5399 3513 5411 3516
rect 5353 3507 5411 3513
rect 5810 3504 5816 3516
rect 5868 3504 5874 3556
rect 5997 3547 6055 3553
rect 5997 3513 6009 3547
rect 6043 3544 6055 3547
rect 6270 3544 6276 3556
rect 6043 3516 6276 3544
rect 6043 3513 6055 3516
rect 5997 3507 6055 3513
rect 6270 3504 6276 3516
rect 6328 3504 6334 3556
rect 8386 3544 8392 3556
rect 7024 3516 8392 3544
rect 4157 3479 4215 3485
rect 3457 3448 3524 3476
rect 2317 3439 2375 3445
rect 3496 3417 3524 3448
rect 4157 3445 4169 3479
rect 4203 3476 4215 3479
rect 4246 3476 4252 3488
rect 4203 3448 4252 3476
rect 4203 3445 4215 3448
rect 4157 3439 4215 3445
rect 4246 3436 4252 3448
rect 4304 3436 4310 3488
rect 5169 3479 5227 3485
rect 5169 3445 5181 3479
rect 5215 3476 5227 3479
rect 5626 3476 5632 3488
rect 5215 3448 5632 3476
rect 5215 3445 5227 3448
rect 5169 3439 5227 3445
rect 5626 3436 5632 3448
rect 5684 3436 5690 3488
rect 5718 3436 5724 3488
rect 5776 3476 5782 3488
rect 6181 3479 6239 3485
rect 6181 3476 6193 3479
rect 5776 3448 6193 3476
rect 5776 3436 5782 3448
rect 6181 3445 6193 3448
rect 6227 3476 6239 3479
rect 6638 3476 6644 3488
rect 6227 3448 6644 3476
rect 6227 3445 6239 3448
rect 6181 3439 6239 3445
rect 6638 3436 6644 3448
rect 6696 3436 6702 3488
rect 7024 3485 7052 3516
rect 8386 3504 8392 3516
rect 8444 3504 8450 3556
rect 11992 3553 12020 3584
rect 12434 3572 12440 3584
rect 12492 3572 12498 3624
rect 12618 3572 12624 3624
rect 12676 3612 12682 3624
rect 12805 3615 12863 3621
rect 12805 3612 12817 3615
rect 12676 3584 12817 3612
rect 12676 3572 12682 3584
rect 12805 3581 12817 3584
rect 12851 3581 12863 3615
rect 13814 3612 13820 3624
rect 13775 3584 13820 3612
rect 12805 3575 12863 3581
rect 13814 3572 13820 3584
rect 13872 3572 13878 3624
rect 11977 3547 12035 3553
rect 8772 3516 10456 3544
rect 7009 3479 7067 3485
rect 7009 3445 7021 3479
rect 7055 3445 7067 3479
rect 7190 3476 7196 3488
rect 7103 3448 7196 3476
rect 7009 3439 7067 3445
rect 7190 3436 7196 3448
rect 7248 3476 7254 3488
rect 8772 3476 8800 3516
rect 10428 3488 10456 3516
rect 11977 3513 11989 3547
rect 12023 3513 12035 3547
rect 13630 3544 13636 3556
rect 11977 3507 12035 3513
rect 12406 3516 13636 3544
rect 7248 3448 8800 3476
rect 7248 3436 7254 3448
rect 9306 3436 9312 3488
rect 9364 3476 9370 3488
rect 9401 3479 9459 3485
rect 9401 3476 9413 3479
rect 9364 3448 9413 3476
rect 9364 3436 9370 3448
rect 9401 3445 9413 3448
rect 9447 3445 9459 3479
rect 9401 3439 9459 3445
rect 9585 3479 9643 3485
rect 9585 3445 9597 3479
rect 9631 3445 9643 3479
rect 9858 3476 9864 3488
rect 9819 3448 9864 3476
rect 9585 3439 9643 3445
rect 937 3411 995 3417
rect 937 3377 949 3411
rect 983 3408 995 3411
rect 3492 3411 3550 3417
rect 983 3380 2774 3408
rect 983 3377 995 3380
rect 937 3371 995 3377
rect 2746 3340 2774 3380
rect 3492 3377 3504 3411
rect 3538 3377 3550 3411
rect 3492 3371 3550 3377
rect 3697 3411 3755 3417
rect 3697 3377 3709 3411
rect 3743 3408 3755 3411
rect 4338 3408 4344 3420
rect 3743 3380 4344 3408
rect 3743 3377 3755 3380
rect 3697 3371 3755 3377
rect 4338 3368 4344 3380
rect 4396 3368 4402 3420
rect 5258 3368 5264 3420
rect 5316 3408 5322 3420
rect 5537 3411 5595 3417
rect 5537 3408 5549 3411
rect 5316 3380 5549 3408
rect 5316 3368 5322 3380
rect 5537 3377 5549 3380
rect 5583 3408 5595 3411
rect 5902 3408 5908 3420
rect 5583 3380 5908 3408
rect 5583 3377 5595 3380
rect 5537 3371 5595 3377
rect 5902 3368 5908 3380
rect 5960 3368 5966 3420
rect 8478 3408 8484 3420
rect 6012 3380 8484 3408
rect 3329 3343 3387 3349
rect 3329 3340 3341 3343
rect 2746 3312 3341 3340
rect 3329 3309 3341 3312
rect 3375 3309 3387 3343
rect 3329 3303 3387 3309
rect 4246 3300 4252 3352
rect 4304 3340 4310 3352
rect 6012 3340 6040 3380
rect 8478 3368 8484 3380
rect 8536 3368 8542 3420
rect 8662 3408 8668 3420
rect 8623 3380 8668 3408
rect 8662 3368 8668 3380
rect 8720 3368 8726 3420
rect 9122 3408 9128 3420
rect 8864 3380 9128 3408
rect 4304 3312 6040 3340
rect 4304 3300 4310 3312
rect 7742 3300 7748 3352
rect 7800 3340 7806 3352
rect 8573 3343 8631 3349
rect 8573 3340 8585 3343
rect 7800 3312 8585 3340
rect 7800 3300 7806 3312
rect 8573 3309 8585 3312
rect 8619 3340 8631 3343
rect 8864 3340 8892 3380
rect 9122 3368 9128 3380
rect 9180 3408 9186 3420
rect 9493 3411 9551 3417
rect 9493 3408 9505 3411
rect 9180 3380 9505 3408
rect 9180 3368 9186 3380
rect 9493 3377 9505 3380
rect 9539 3377 9551 3411
rect 9493 3371 9551 3377
rect 9600 3352 9628 3439
rect 9858 3436 9864 3448
rect 9916 3436 9922 3488
rect 10410 3476 10416 3488
rect 10371 3448 10416 3476
rect 10410 3436 10416 3448
rect 10468 3436 10474 3488
rect 11054 3476 11060 3488
rect 11015 3448 11060 3476
rect 11054 3436 11060 3448
rect 11112 3436 11118 3488
rect 11606 3436 11612 3488
rect 11664 3476 11670 3488
rect 11885 3479 11943 3485
rect 11885 3476 11897 3479
rect 11664 3448 11897 3476
rect 11664 3436 11670 3448
rect 11885 3445 11897 3448
rect 11931 3445 11943 3479
rect 11885 3439 11943 3445
rect 12069 3479 12127 3485
rect 12069 3445 12081 3479
rect 12115 3476 12127 3479
rect 12406 3476 12434 3516
rect 13630 3504 13636 3516
rect 13688 3504 13694 3556
rect 12526 3476 12532 3488
rect 12115 3448 12434 3476
rect 12487 3448 12532 3476
rect 12115 3445 12127 3448
rect 12069 3439 12127 3445
rect 12526 3436 12532 3448
rect 12584 3436 12590 3488
rect 14001 3479 14059 3485
rect 14001 3476 14013 3479
rect 12728 3448 14013 3476
rect 9723 3411 9781 3417
rect 9723 3377 9735 3411
rect 9769 3408 9781 3411
rect 9950 3408 9956 3420
rect 9769 3380 9956 3408
rect 9769 3377 9781 3380
rect 9723 3371 9781 3377
rect 9950 3368 9956 3380
rect 10008 3368 10014 3420
rect 11422 3368 11428 3420
rect 11480 3408 11486 3420
rect 11790 3408 11796 3420
rect 11480 3380 11796 3408
rect 11480 3368 11486 3380
rect 11790 3368 11796 3380
rect 11848 3408 11854 3420
rect 12728 3408 12756 3448
rect 14001 3445 14013 3448
rect 14047 3476 14059 3479
rect 14829 3479 14887 3485
rect 14829 3476 14841 3479
rect 14047 3448 14841 3476
rect 14047 3445 14059 3448
rect 14001 3439 14059 3445
rect 14829 3445 14841 3448
rect 14875 3445 14887 3479
rect 14829 3439 14887 3445
rect 14921 3479 14979 3485
rect 14921 3445 14933 3479
rect 14967 3476 14979 3479
rect 15010 3476 15016 3488
rect 14967 3448 15016 3476
rect 14967 3445 14979 3448
rect 14921 3439 14979 3445
rect 11848 3380 12756 3408
rect 12805 3411 12863 3417
rect 11848 3368 11854 3380
rect 12805 3377 12817 3411
rect 12851 3408 12863 3411
rect 13722 3408 13728 3420
rect 12851 3380 13728 3408
rect 12851 3377 12863 3380
rect 12805 3371 12863 3377
rect 13722 3368 13728 3380
rect 13780 3368 13786 3420
rect 14182 3408 14188 3420
rect 14095 3380 14188 3408
rect 14182 3368 14188 3380
rect 14240 3408 14246 3420
rect 14645 3411 14703 3417
rect 14645 3408 14657 3411
rect 14240 3380 14657 3408
rect 14240 3368 14246 3380
rect 14645 3377 14657 3380
rect 14691 3377 14703 3411
rect 14645 3371 14703 3377
rect 8619 3312 8892 3340
rect 8619 3309 8631 3312
rect 8573 3303 8631 3309
rect 8938 3300 8944 3352
rect 8996 3340 9002 3352
rect 9217 3343 9275 3349
rect 9217 3340 9229 3343
rect 8996 3312 9229 3340
rect 8996 3300 9002 3312
rect 9217 3309 9229 3312
rect 9263 3309 9275 3343
rect 9217 3303 9275 3309
rect 9582 3300 9588 3352
rect 9640 3300 9646 3352
rect 10134 3300 10140 3352
rect 10192 3340 10198 3352
rect 10505 3343 10563 3349
rect 10505 3340 10517 3343
rect 10192 3312 10517 3340
rect 10192 3300 10198 3312
rect 10505 3309 10517 3312
rect 10551 3309 10563 3343
rect 10505 3303 10563 3309
rect 12526 3300 12532 3352
rect 12584 3340 12590 3352
rect 12621 3343 12679 3349
rect 12621 3340 12633 3343
rect 12584 3312 12633 3340
rect 12584 3300 12590 3312
rect 12621 3309 12633 3312
rect 12667 3309 12679 3343
rect 12621 3303 12679 3309
rect 12710 3300 12716 3352
rect 12768 3340 12774 3352
rect 14936 3340 14964 3439
rect 15010 3436 15016 3448
rect 15068 3436 15074 3488
rect 12768 3312 14964 3340
rect 12768 3300 12774 3312
rect 92 3250 15824 3272
rect 92 3198 5242 3250
rect 5294 3198 5306 3250
rect 5358 3198 5370 3250
rect 5422 3198 5434 3250
rect 5486 3198 10514 3250
rect 10566 3198 10578 3250
rect 10630 3198 10642 3250
rect 10694 3198 10706 3250
rect 10758 3198 15824 3250
rect 92 3176 15824 3198
rect 2958 3096 2964 3148
rect 3016 3136 3022 3148
rect 3237 3139 3295 3145
rect 3237 3136 3249 3139
rect 3016 3108 3249 3136
rect 3016 3096 3022 3108
rect 3237 3105 3249 3108
rect 3283 3105 3295 3139
rect 4246 3136 4252 3148
rect 4207 3108 4252 3136
rect 3237 3099 3295 3105
rect 4246 3096 4252 3108
rect 4304 3096 4310 3148
rect 5810 3136 5816 3148
rect 5771 3108 5816 3136
rect 5810 3096 5816 3108
rect 5868 3096 5874 3148
rect 5902 3096 5908 3148
rect 5960 3136 5966 3148
rect 8846 3136 8852 3148
rect 5960 3108 6960 3136
rect 5960 3096 5966 3108
rect 1210 3068 1216 3080
rect 1171 3040 1216 3068
rect 1210 3028 1216 3040
rect 1268 3028 1274 3080
rect 1946 3028 1952 3080
rect 2004 3028 2010 3080
rect 4801 3071 4859 3077
rect 4801 3037 4813 3071
rect 4847 3068 4859 3071
rect 5626 3068 5632 3080
rect 4847 3040 5632 3068
rect 4847 3037 4859 3040
rect 4801 3031 4859 3037
rect 5626 3028 5632 3040
rect 5684 3068 5690 3080
rect 5684 3040 6224 3068
rect 5684 3028 5690 3040
rect 6196 3012 6224 3040
rect 3142 3000 3148 3012
rect 3103 2972 3148 3000
rect 3142 2960 3148 2972
rect 3200 2960 3206 3012
rect 4065 3003 4123 3009
rect 4065 2969 4077 3003
rect 4111 2969 4123 3003
rect 4065 2963 4123 2969
rect 750 2892 756 2944
rect 808 2932 814 2944
rect 937 2935 995 2941
rect 937 2932 949 2935
rect 808 2904 949 2932
rect 808 2892 814 2904
rect 937 2901 949 2904
rect 983 2932 995 2935
rect 1578 2932 1584 2944
rect 983 2904 1584 2932
rect 983 2901 995 2904
rect 937 2895 995 2901
rect 1578 2892 1584 2904
rect 1636 2892 1642 2944
rect 4080 2864 4108 2963
rect 4614 2960 4620 3012
rect 4672 3000 4678 3012
rect 4709 3003 4767 3009
rect 4709 3000 4721 3003
rect 4672 2972 4721 3000
rect 4672 2960 4678 2972
rect 4709 2969 4721 2972
rect 4755 2969 4767 3003
rect 5994 3000 6000 3012
rect 5955 2972 6000 3000
rect 4709 2963 4767 2969
rect 5994 2960 6000 2972
rect 6052 2960 6058 3012
rect 6089 3003 6147 3009
rect 6089 2969 6101 3003
rect 6135 2969 6147 3003
rect 6089 2963 6147 2969
rect 6104 2932 6132 2963
rect 6178 2960 6184 3012
rect 6236 3000 6242 3012
rect 6365 3003 6423 3009
rect 6236 2972 6281 3000
rect 6236 2960 6242 2972
rect 6365 2969 6377 3003
rect 6411 3000 6423 3003
rect 6822 3000 6828 3012
rect 6411 2972 6828 3000
rect 6411 2969 6423 2972
rect 6365 2963 6423 2969
rect 6822 2960 6828 2972
rect 6880 2960 6886 3012
rect 6932 3000 6960 3108
rect 7024 3108 8852 3136
rect 7024 3077 7052 3108
rect 8846 3096 8852 3108
rect 8904 3096 8910 3148
rect 9398 3096 9404 3148
rect 9456 3136 9462 3148
rect 9582 3136 9588 3148
rect 9456 3108 9588 3136
rect 9456 3096 9462 3108
rect 9582 3096 9588 3108
rect 9640 3136 9646 3148
rect 10137 3139 10195 3145
rect 10137 3136 10149 3139
rect 9640 3108 10149 3136
rect 9640 3096 9646 3108
rect 10137 3105 10149 3108
rect 10183 3136 10195 3139
rect 11146 3136 11152 3148
rect 10183 3108 11152 3136
rect 10183 3105 10195 3108
rect 10137 3099 10195 3105
rect 11146 3096 11152 3108
rect 11204 3096 11210 3148
rect 11606 3096 11612 3148
rect 11664 3136 11670 3148
rect 12894 3136 12900 3148
rect 11664 3108 12900 3136
rect 11664 3096 11670 3108
rect 12894 3096 12900 3108
rect 12952 3096 12958 3148
rect 14182 3136 14188 3148
rect 14143 3108 14188 3136
rect 14182 3096 14188 3108
rect 14240 3096 14246 3148
rect 7009 3071 7067 3077
rect 7009 3037 7021 3071
rect 7055 3037 7067 3071
rect 7834 3068 7840 3080
rect 7009 3031 7067 3037
rect 7589 3040 7840 3068
rect 7589 3000 7617 3040
rect 7834 3028 7840 3040
rect 7892 3028 7898 3080
rect 8570 3068 8576 3080
rect 8404 3040 8576 3068
rect 8404 3009 8432 3040
rect 8570 3028 8576 3040
rect 8628 3068 8634 3080
rect 8754 3068 8760 3080
rect 8628 3040 8760 3068
rect 8628 3028 8634 3040
rect 8754 3028 8760 3040
rect 8812 3028 8818 3080
rect 9214 3028 9220 3080
rect 9272 3028 9278 3080
rect 10870 3028 10876 3080
rect 10928 3068 10934 3080
rect 11333 3071 11391 3077
rect 11333 3068 11345 3071
rect 10928 3040 11345 3068
rect 10928 3028 10934 3040
rect 11333 3037 11345 3040
rect 11379 3037 11391 3071
rect 11333 3031 11391 3037
rect 12250 3028 12256 3080
rect 12308 3068 12314 3080
rect 12713 3071 12771 3077
rect 12713 3068 12725 3071
rect 12308 3040 12725 3068
rect 12308 3028 12314 3040
rect 12713 3037 12725 3040
rect 12759 3037 12771 3071
rect 12713 3031 12771 3037
rect 13446 3028 13452 3080
rect 13504 3028 13510 3080
rect 14921 3071 14979 3077
rect 14921 3037 14933 3071
rect 14967 3068 14979 3071
rect 15286 3068 15292 3080
rect 14967 3040 15292 3068
rect 14967 3037 14979 3040
rect 14921 3031 14979 3037
rect 15286 3028 15292 3040
rect 15344 3028 15350 3080
rect 6932 2972 7617 3000
rect 7653 3003 7711 3009
rect 7653 2969 7665 3003
rect 7699 2969 7711 3003
rect 7653 2963 7711 2969
rect 8389 3003 8447 3009
rect 8389 2969 8401 3003
rect 8435 2969 8447 3003
rect 11238 3000 11244 3012
rect 11199 2972 11244 3000
rect 8389 2963 8447 2969
rect 6270 2932 6276 2944
rect 6104 2904 6276 2932
rect 6270 2892 6276 2904
rect 6328 2892 6334 2944
rect 6914 2932 6920 2944
rect 6827 2904 6920 2932
rect 6914 2892 6920 2904
rect 6972 2932 6978 2944
rect 7668 2932 7696 2963
rect 11238 2960 11244 2972
rect 11296 2960 11302 3012
rect 11422 2960 11428 3012
rect 11480 3000 11486 3012
rect 11563 3003 11621 3009
rect 11480 2972 11525 3000
rect 11480 2960 11486 2972
rect 11563 2969 11575 3003
rect 11609 3000 11621 3003
rect 11609 2972 11836 3000
rect 11609 2969 11621 2972
rect 11563 2963 11621 2969
rect 8662 2932 8668 2944
rect 6972 2904 7696 2932
rect 8623 2904 8668 2932
rect 6972 2892 6978 2904
rect 8662 2892 8668 2904
rect 8720 2892 8726 2944
rect 9858 2892 9864 2944
rect 9916 2932 9922 2944
rect 10962 2932 10968 2944
rect 9916 2904 10968 2932
rect 9916 2892 9922 2904
rect 10962 2892 10968 2904
rect 11020 2932 11026 2944
rect 11698 2932 11704 2944
rect 11020 2904 11704 2932
rect 11020 2892 11026 2904
rect 11698 2892 11704 2904
rect 11756 2892 11762 2944
rect 6638 2864 6644 2876
rect 4080 2836 6644 2864
rect 6638 2824 6644 2836
rect 6696 2824 6702 2876
rect 2222 2756 2228 2808
rect 2280 2796 2286 2808
rect 2685 2799 2743 2805
rect 2685 2796 2697 2799
rect 2280 2768 2697 2796
rect 2280 2756 2286 2768
rect 2685 2765 2697 2768
rect 2731 2765 2743 2799
rect 2685 2759 2743 2765
rect 5902 2756 5908 2808
rect 5960 2796 5966 2808
rect 6932 2805 6960 2892
rect 9766 2824 9772 2876
rect 9824 2864 9830 2876
rect 11808 2864 11836 2972
rect 12434 2892 12440 2944
rect 12492 2932 12498 2944
rect 12492 2904 12537 2932
rect 12492 2892 12498 2904
rect 15102 2864 15108 2876
rect 9824 2836 11836 2864
rect 15063 2836 15108 2864
rect 9824 2824 9830 2836
rect 15102 2824 15108 2836
rect 15160 2824 15166 2876
rect 6917 2799 6975 2805
rect 6917 2796 6929 2799
rect 5960 2768 6929 2796
rect 5960 2756 5966 2768
rect 6917 2765 6929 2768
rect 6963 2765 6975 2799
rect 6917 2759 6975 2765
rect 9674 2756 9680 2808
rect 9732 2796 9738 2808
rect 10870 2796 10876 2808
rect 9732 2768 10876 2796
rect 9732 2756 9738 2768
rect 10870 2756 10876 2768
rect 10928 2756 10934 2808
rect 11054 2796 11060 2808
rect 11015 2768 11060 2796
rect 11054 2756 11060 2768
rect 11112 2756 11118 2808
rect 11146 2756 11152 2808
rect 11204 2796 11210 2808
rect 11330 2796 11336 2808
rect 11204 2768 11336 2796
rect 11204 2756 11210 2768
rect 11330 2756 11336 2768
rect 11388 2756 11394 2808
rect 92 2706 15824 2728
rect 92 2654 2606 2706
rect 2658 2654 2670 2706
rect 2722 2654 2734 2706
rect 2786 2654 2798 2706
rect 2850 2654 7878 2706
rect 7930 2654 7942 2706
rect 7994 2654 8006 2706
rect 8058 2654 8070 2706
rect 8122 2654 13150 2706
rect 13202 2654 13214 2706
rect 13266 2654 13278 2706
rect 13330 2654 13342 2706
rect 13394 2654 15824 2706
rect 92 2632 15824 2654
rect 1118 2552 1124 2604
rect 1176 2592 1182 2604
rect 1581 2595 1639 2601
rect 1581 2592 1593 2595
rect 1176 2564 1593 2592
rect 1176 2552 1182 2564
rect 1581 2561 1593 2564
rect 1627 2561 1639 2595
rect 1581 2555 1639 2561
rect 2317 2595 2375 2601
rect 2317 2561 2329 2595
rect 2363 2592 2375 2595
rect 4706 2592 4712 2604
rect 2363 2564 4712 2592
rect 2363 2561 2375 2564
rect 2317 2555 2375 2561
rect 4706 2552 4712 2564
rect 4764 2552 4770 2604
rect 5718 2592 5724 2604
rect 4816 2564 5724 2592
rect 4816 2524 4844 2564
rect 5718 2552 5724 2564
rect 5776 2552 5782 2604
rect 9033 2595 9091 2601
rect 9033 2561 9045 2595
rect 9079 2592 9091 2595
rect 9766 2592 9772 2604
rect 9079 2564 9772 2592
rect 9079 2561 9091 2564
rect 9033 2555 9091 2561
rect 9766 2552 9772 2564
rect 9824 2552 9830 2604
rect 9950 2552 9956 2604
rect 10008 2592 10014 2604
rect 12526 2592 12532 2604
rect 10008 2564 12532 2592
rect 10008 2552 10014 2564
rect 2332 2496 4844 2524
rect 1670 2388 1676 2400
rect 1631 2360 1676 2388
rect 1670 2348 1676 2360
rect 1728 2348 1734 2400
rect 2133 2391 2191 2397
rect 2133 2357 2145 2391
rect 2179 2388 2191 2391
rect 2222 2388 2228 2400
rect 2179 2360 2228 2388
rect 2179 2357 2191 2360
rect 2133 2351 2191 2357
rect 2222 2348 2228 2360
rect 2280 2348 2286 2400
rect 2332 2397 2360 2496
rect 4249 2459 4307 2465
rect 4249 2456 4261 2459
rect 2424 2428 4261 2456
rect 2317 2391 2375 2397
rect 2317 2357 2329 2391
rect 2363 2357 2375 2391
rect 2317 2351 2375 2357
rect 842 2320 848 2332
rect 803 2292 848 2320
rect 842 2280 848 2292
rect 900 2280 906 2332
rect 1210 2280 1216 2332
rect 1268 2320 1274 2332
rect 2424 2320 2452 2428
rect 4249 2425 4261 2428
rect 4295 2456 4307 2459
rect 5626 2456 5632 2468
rect 4295 2428 5632 2456
rect 4295 2425 4307 2428
rect 4249 2419 4307 2425
rect 5626 2416 5632 2428
rect 5684 2456 5690 2468
rect 6730 2456 6736 2468
rect 5684 2428 6736 2456
rect 5684 2416 5690 2428
rect 6730 2416 6736 2428
rect 6788 2416 6794 2468
rect 7190 2416 7196 2468
rect 7248 2456 7254 2468
rect 10505 2459 10563 2465
rect 7248 2428 7420 2456
rect 7248 2416 7254 2428
rect 3973 2391 4031 2397
rect 3973 2357 3985 2391
rect 4019 2357 4031 2391
rect 4154 2388 4160 2400
rect 4115 2360 4160 2388
rect 3973 2351 4031 2357
rect 3988 2320 4016 2351
rect 4154 2348 4160 2360
rect 4212 2348 4218 2400
rect 4706 2388 4712 2400
rect 4667 2360 4712 2388
rect 4706 2348 4712 2360
rect 4764 2348 4770 2400
rect 7282 2388 7288 2400
rect 6840 2360 7288 2388
rect 4522 2320 4528 2332
rect 1268 2292 2452 2320
rect 3620 2292 3924 2320
rect 3988 2292 4528 2320
rect 1268 2280 1274 2292
rect 937 2255 995 2261
rect 937 2221 949 2255
rect 983 2252 995 2255
rect 3620 2252 3648 2292
rect 3786 2252 3792 2264
rect 983 2224 3648 2252
rect 3747 2224 3792 2252
rect 983 2221 995 2224
rect 937 2215 995 2221
rect 3786 2212 3792 2224
rect 3844 2212 3850 2264
rect 3896 2252 3924 2292
rect 4522 2280 4528 2292
rect 4580 2280 4586 2332
rect 4985 2323 5043 2329
rect 4985 2289 4997 2323
rect 5031 2320 5043 2323
rect 5258 2320 5264 2332
rect 5031 2292 5264 2320
rect 5031 2289 5043 2292
rect 4985 2283 5043 2289
rect 5258 2280 5264 2292
rect 5316 2280 5322 2332
rect 5718 2280 5724 2332
rect 5776 2280 5782 2332
rect 6270 2280 6276 2332
rect 6328 2320 6334 2332
rect 6733 2323 6791 2329
rect 6733 2320 6745 2323
rect 6328 2292 6745 2320
rect 6328 2280 6334 2292
rect 6733 2289 6745 2292
rect 6779 2289 6791 2323
rect 6733 2283 6791 2289
rect 4430 2252 4436 2264
rect 3896 2224 4436 2252
rect 4430 2212 4436 2224
rect 4488 2212 4494 2264
rect 4890 2212 4896 2264
rect 4948 2252 4954 2264
rect 6840 2252 6868 2360
rect 7282 2348 7288 2360
rect 7340 2348 7346 2400
rect 7392 2397 7420 2428
rect 10505 2425 10517 2459
rect 10551 2456 10563 2459
rect 11054 2456 11060 2468
rect 10551 2428 11060 2456
rect 10551 2425 10563 2428
rect 10505 2419 10563 2425
rect 11054 2416 11060 2428
rect 11112 2416 11118 2468
rect 7377 2391 7435 2397
rect 7377 2357 7389 2391
rect 7423 2357 7435 2391
rect 7377 2351 7435 2357
rect 10781 2391 10839 2397
rect 10781 2357 10793 2391
rect 10827 2357 10839 2391
rect 10781 2351 10839 2357
rect 6914 2280 6920 2332
rect 6972 2320 6978 2332
rect 7193 2323 7251 2329
rect 7193 2320 7205 2323
rect 6972 2292 7205 2320
rect 6972 2280 6978 2292
rect 7193 2289 7205 2292
rect 7239 2289 7251 2323
rect 7193 2283 7251 2289
rect 9490 2280 9496 2332
rect 9548 2280 9554 2332
rect 4948 2224 6868 2252
rect 4948 2212 4954 2224
rect 8478 2212 8484 2264
rect 8536 2252 8542 2264
rect 10796 2252 10824 2351
rect 11238 2348 11244 2400
rect 11296 2388 11302 2400
rect 11425 2391 11483 2397
rect 11425 2388 11437 2391
rect 11296 2360 11437 2388
rect 11296 2348 11302 2360
rect 11425 2357 11437 2360
rect 11471 2357 11483 2391
rect 11532 2388 11560 2564
rect 12526 2552 12532 2564
rect 12584 2552 12590 2604
rect 13998 2592 14004 2604
rect 13959 2564 14004 2592
rect 13998 2552 14004 2564
rect 14056 2552 14062 2604
rect 14918 2552 14924 2604
rect 14976 2592 14982 2604
rect 15013 2595 15071 2601
rect 15013 2592 15025 2595
rect 14976 2564 15025 2592
rect 14976 2552 14982 2564
rect 15013 2561 15025 2564
rect 15059 2561 15071 2595
rect 15013 2555 15071 2561
rect 11698 2416 11704 2468
rect 11756 2456 11762 2468
rect 11885 2459 11943 2465
rect 11885 2456 11897 2459
rect 11756 2428 11897 2456
rect 11756 2416 11762 2428
rect 11885 2425 11897 2428
rect 11931 2425 11943 2459
rect 12544 2456 12572 2552
rect 12544 2428 13952 2456
rect 11885 2419 11943 2425
rect 11609 2391 11667 2397
rect 11609 2388 11621 2391
rect 11532 2360 11621 2388
rect 11425 2351 11483 2357
rect 11609 2357 11621 2360
rect 11655 2357 11667 2391
rect 12618 2388 12624 2400
rect 12579 2360 12624 2388
rect 11609 2351 11667 2357
rect 12618 2348 12624 2360
rect 12676 2348 12682 2400
rect 12805 2391 12863 2397
rect 12805 2357 12817 2391
rect 12851 2388 12863 2391
rect 12894 2388 12900 2400
rect 12851 2360 12900 2388
rect 12851 2357 12863 2360
rect 12805 2351 12863 2357
rect 12894 2348 12900 2360
rect 12952 2348 12958 2400
rect 13722 2388 13728 2400
rect 13683 2360 13728 2388
rect 13722 2348 13728 2360
rect 13780 2348 13786 2400
rect 13924 2397 13952 2428
rect 13909 2391 13967 2397
rect 13909 2357 13921 2391
rect 13955 2357 13967 2391
rect 13909 2351 13967 2357
rect 14921 2391 14979 2397
rect 14921 2357 14933 2391
rect 14967 2388 14979 2391
rect 15010 2388 15016 2400
rect 14967 2360 15016 2388
rect 14967 2357 14979 2360
rect 14921 2351 14979 2357
rect 15010 2348 15016 2360
rect 15068 2348 15074 2400
rect 10962 2280 10968 2332
rect 11020 2320 11026 2332
rect 11517 2323 11575 2329
rect 11517 2320 11529 2323
rect 11020 2292 11529 2320
rect 11020 2280 11026 2292
rect 11517 2289 11529 2292
rect 11563 2289 11575 2323
rect 11517 2283 11575 2289
rect 11698 2280 11704 2332
rect 11756 2329 11762 2332
rect 11756 2323 11785 2329
rect 11773 2289 11785 2323
rect 11756 2283 11785 2289
rect 11756 2280 11762 2283
rect 11238 2252 11244 2264
rect 8536 2224 10824 2252
rect 11199 2224 11244 2252
rect 8536 2212 8542 2224
rect 11238 2212 11244 2224
rect 11296 2212 11302 2264
rect 12618 2212 12624 2264
rect 12676 2252 12682 2264
rect 12713 2255 12771 2261
rect 12713 2252 12725 2255
rect 12676 2224 12725 2252
rect 12676 2212 12682 2224
rect 12713 2221 12725 2224
rect 12759 2221 12771 2255
rect 12713 2215 12771 2221
rect 92 2162 15824 2184
rect 92 2110 5242 2162
rect 5294 2110 5306 2162
rect 5358 2110 5370 2162
rect 5422 2110 5434 2162
rect 5486 2110 10514 2162
rect 10566 2110 10578 2162
rect 10630 2110 10642 2162
rect 10694 2110 10706 2162
rect 10758 2110 15824 2162
rect 92 2088 15824 2110
rect 1121 2051 1179 2057
rect 1121 2017 1133 2051
rect 1167 2048 1179 2051
rect 5074 2048 5080 2060
rect 1167 2020 5080 2048
rect 1167 2017 1179 2020
rect 1121 2011 1179 2017
rect 5074 2008 5080 2020
rect 5132 2008 5138 2060
rect 6638 2048 6644 2060
rect 6599 2020 6644 2048
rect 6638 2008 6644 2020
rect 6696 2008 6702 2060
rect 7282 2008 7288 2060
rect 7340 2048 7346 2060
rect 7340 2020 11100 2048
rect 7340 2008 7346 2020
rect 3510 1980 3516 1992
rect 3174 1952 3516 1980
rect 3510 1940 3516 1952
rect 3568 1940 3574 1992
rect 4154 1940 4160 1992
rect 4212 1980 4218 1992
rect 4706 1980 4712 1992
rect 4212 1952 4712 1980
rect 4212 1940 4218 1952
rect 4706 1940 4712 1952
rect 4764 1940 4770 1992
rect 6270 1980 6276 1992
rect 4816 1952 6276 1980
rect 569 1915 627 1921
rect 569 1881 581 1915
rect 615 1881 627 1915
rect 1210 1912 1216 1924
rect 1171 1884 1216 1912
rect 569 1875 627 1881
rect 584 1844 612 1875
rect 1210 1872 1216 1884
rect 1268 1872 1274 1924
rect 4614 1912 4620 1924
rect 4527 1884 4620 1912
rect 4614 1872 4620 1884
rect 4672 1912 4678 1924
rect 4816 1912 4844 1952
rect 6270 1940 6276 1952
rect 6328 1940 6334 1992
rect 6822 1940 6828 1992
rect 6880 1980 6886 1992
rect 7561 1983 7619 1989
rect 7561 1980 7573 1983
rect 6880 1952 7573 1980
rect 6880 1940 6886 1952
rect 7561 1949 7573 1952
rect 7607 1949 7619 1983
rect 7561 1943 7619 1949
rect 8665 1983 8723 1989
rect 8665 1949 8677 1983
rect 8711 1980 8723 1983
rect 8938 1980 8944 1992
rect 8711 1952 8944 1980
rect 8711 1949 8723 1952
rect 8665 1943 8723 1949
rect 8938 1940 8944 1952
rect 8996 1940 9002 1992
rect 9674 1940 9680 1992
rect 9732 1940 9738 1992
rect 4672 1884 4844 1912
rect 4893 1915 4951 1921
rect 4672 1872 4678 1884
rect 4893 1881 4905 1915
rect 4939 1912 4951 1915
rect 5902 1912 5908 1924
rect 4939 1884 5908 1912
rect 4939 1881 4951 1884
rect 4893 1875 4951 1881
rect 5902 1872 5908 1884
rect 5960 1872 5966 1924
rect 6730 1872 6736 1924
rect 6788 1912 6794 1924
rect 7377 1915 7435 1921
rect 7377 1912 7389 1915
rect 6788 1884 7389 1912
rect 6788 1872 6794 1884
rect 7377 1881 7389 1884
rect 7423 1881 7435 1915
rect 7377 1875 7435 1881
rect 7469 1915 7527 1921
rect 7469 1881 7481 1915
rect 7515 1881 7527 1915
rect 7742 1912 7748 1924
rect 7703 1884 7748 1912
rect 7469 1875 7527 1881
rect 1670 1844 1676 1856
rect 584 1816 1532 1844
rect 1631 1816 1676 1844
rect 477 1779 535 1785
rect 477 1745 489 1779
rect 523 1776 535 1779
rect 1302 1776 1308 1788
rect 523 1748 1308 1776
rect 523 1745 535 1748
rect 477 1739 535 1745
rect 1302 1736 1308 1748
rect 1360 1736 1366 1788
rect 1504 1708 1532 1816
rect 1670 1804 1676 1816
rect 1728 1804 1734 1856
rect 1949 1847 2007 1853
rect 1949 1813 1961 1847
rect 1995 1844 2007 1847
rect 3970 1844 3976 1856
rect 1995 1816 3976 1844
rect 1995 1813 2007 1816
rect 1949 1807 2007 1813
rect 3970 1804 3976 1816
rect 4028 1804 4034 1856
rect 4157 1847 4215 1853
rect 4157 1813 4169 1847
rect 4203 1813 4215 1847
rect 4157 1807 4215 1813
rect 4249 1847 4307 1853
rect 4249 1813 4261 1847
rect 4295 1844 4307 1847
rect 5534 1844 5540 1856
rect 4295 1816 5540 1844
rect 4295 1813 4307 1816
rect 4249 1807 4307 1813
rect 3421 1779 3479 1785
rect 3421 1745 3433 1779
rect 3467 1776 3479 1779
rect 4172 1776 4200 1807
rect 5534 1804 5540 1816
rect 5592 1844 5598 1856
rect 5592 1816 5948 1844
rect 5592 1804 5598 1816
rect 4338 1776 4344 1788
rect 3467 1748 4344 1776
rect 3467 1745 3479 1748
rect 3421 1739 3479 1745
rect 4338 1736 4344 1748
rect 4396 1776 4402 1788
rect 5813 1779 5871 1785
rect 5813 1776 5825 1779
rect 4396 1748 5825 1776
rect 4396 1736 4402 1748
rect 5813 1745 5825 1748
rect 5859 1745 5871 1779
rect 5920 1776 5948 1816
rect 6178 1804 6184 1856
rect 6236 1844 6242 1856
rect 6365 1847 6423 1853
rect 6365 1844 6377 1847
rect 6236 1816 6377 1844
rect 6236 1804 6242 1816
rect 6365 1813 6377 1816
rect 6411 1813 6423 1847
rect 6365 1807 6423 1813
rect 5994 1776 6000 1788
rect 5907 1748 6000 1776
rect 5813 1739 5871 1745
rect 5994 1736 6000 1748
rect 6052 1776 6058 1788
rect 7484 1776 7512 1875
rect 7742 1872 7748 1884
rect 7800 1872 7806 1924
rect 11072 1921 11100 2020
rect 11606 2008 11612 2060
rect 11664 2048 11670 2060
rect 11701 2051 11759 2057
rect 11701 2048 11713 2051
rect 11664 2020 11713 2048
rect 11664 2008 11670 2020
rect 11701 2017 11713 2020
rect 11747 2017 11759 2051
rect 11701 2011 11759 2017
rect 13538 2008 13544 2060
rect 13596 2008 13602 2060
rect 12618 1980 12624 1992
rect 12579 1952 12624 1980
rect 12618 1940 12624 1952
rect 12676 1940 12682 1992
rect 13556 1966 13584 2008
rect 13906 1940 13912 1992
rect 13964 1980 13970 1992
rect 14921 1983 14979 1989
rect 14921 1980 14933 1983
rect 13964 1952 14933 1980
rect 13964 1940 13970 1952
rect 14921 1949 14933 1952
rect 14967 1949 14979 1983
rect 14921 1943 14979 1949
rect 11057 1915 11115 1921
rect 11057 1881 11069 1915
rect 11103 1881 11115 1915
rect 11057 1875 11115 1881
rect 11146 1872 11152 1924
rect 11204 1912 11210 1924
rect 11885 1915 11943 1921
rect 11885 1912 11897 1915
rect 11204 1884 11897 1912
rect 11204 1872 11210 1884
rect 11885 1881 11897 1884
rect 11931 1881 11943 1915
rect 11885 1875 11943 1881
rect 8389 1847 8447 1853
rect 8389 1813 8401 1847
rect 8435 1813 8447 1847
rect 8389 1807 8447 1813
rect 6052 1748 7512 1776
rect 6052 1736 6058 1748
rect 8294 1736 8300 1788
rect 8352 1776 8358 1788
rect 8404 1776 8432 1807
rect 9950 1804 9956 1856
rect 10008 1844 10014 1856
rect 10137 1847 10195 1853
rect 10137 1844 10149 1847
rect 10008 1816 10149 1844
rect 10008 1804 10014 1816
rect 10137 1813 10149 1816
rect 10183 1813 10195 1847
rect 12342 1844 12348 1856
rect 12303 1816 12348 1844
rect 10137 1807 10195 1813
rect 12342 1804 12348 1816
rect 12400 1804 12406 1856
rect 8352 1748 8432 1776
rect 8352 1736 8358 1748
rect 3326 1708 3332 1720
rect 1504 1680 3332 1708
rect 3326 1668 3332 1680
rect 3384 1668 3390 1720
rect 4522 1668 4528 1720
rect 4580 1708 4586 1720
rect 6181 1711 6239 1717
rect 6181 1708 6193 1711
rect 4580 1680 6193 1708
rect 4580 1668 4586 1680
rect 6181 1677 6193 1680
rect 6227 1677 6239 1711
rect 6181 1671 6239 1677
rect 6273 1711 6331 1717
rect 6273 1677 6285 1711
rect 6319 1708 6331 1711
rect 6822 1708 6828 1720
rect 6319 1680 6828 1708
rect 6319 1677 6331 1680
rect 6273 1671 6331 1677
rect 6822 1668 6828 1680
rect 6880 1668 6886 1720
rect 7006 1668 7012 1720
rect 7064 1708 7070 1720
rect 7193 1711 7251 1717
rect 7193 1708 7205 1711
rect 7064 1680 7205 1708
rect 7064 1668 7070 1680
rect 7193 1677 7205 1680
rect 7239 1677 7251 1711
rect 8404 1708 8432 1748
rect 13722 1736 13728 1788
rect 13780 1776 13786 1788
rect 14093 1779 14151 1785
rect 14093 1776 14105 1779
rect 13780 1748 14105 1776
rect 13780 1736 13786 1748
rect 14093 1745 14105 1748
rect 14139 1745 14151 1779
rect 15102 1776 15108 1788
rect 15063 1748 15108 1776
rect 14093 1739 14151 1745
rect 15102 1736 15108 1748
rect 15160 1736 15166 1788
rect 8478 1708 8484 1720
rect 8404 1680 8484 1708
rect 7193 1671 7251 1677
rect 8478 1668 8484 1680
rect 8536 1668 8542 1720
rect 11146 1708 11152 1720
rect 11107 1680 11152 1708
rect 11146 1668 11152 1680
rect 11204 1668 11210 1720
rect 92 1618 15824 1640
rect 92 1566 2606 1618
rect 2658 1566 2670 1618
rect 2722 1566 2734 1618
rect 2786 1566 2798 1618
rect 2850 1566 7878 1618
rect 7930 1566 7942 1618
rect 7994 1566 8006 1618
rect 8058 1566 8070 1618
rect 8122 1566 13150 1618
rect 13202 1566 13214 1618
rect 13266 1566 13278 1618
rect 13330 1566 13342 1618
rect 13394 1566 15824 1618
rect 92 1544 15824 1566
rect 4706 1504 4712 1516
rect 4667 1476 4712 1504
rect 4706 1464 4712 1476
rect 4764 1464 4770 1516
rect 6454 1504 6460 1516
rect 4816 1476 6460 1504
rect 3326 1396 3332 1448
rect 3384 1436 3390 1448
rect 4816 1436 4844 1476
rect 6454 1464 6460 1476
rect 6512 1464 6518 1516
rect 10781 1507 10839 1513
rect 9048 1476 10364 1504
rect 3384 1408 4844 1436
rect 3384 1396 3390 1408
rect 5261 1371 5319 1377
rect 5261 1337 5273 1371
rect 5307 1368 5319 1371
rect 5534 1368 5540 1380
rect 5307 1340 5540 1368
rect 5307 1337 5319 1340
rect 5261 1331 5319 1337
rect 5534 1328 5540 1340
rect 5592 1328 5598 1380
rect 7006 1368 7012 1380
rect 6967 1340 7012 1368
rect 7006 1328 7012 1340
rect 7064 1328 7070 1380
rect 845 1303 903 1309
rect 845 1269 857 1303
rect 891 1300 903 1303
rect 1026 1300 1032 1312
rect 891 1272 1032 1300
rect 891 1269 903 1272
rect 845 1263 903 1269
rect 1026 1260 1032 1272
rect 1084 1260 1090 1312
rect 2314 1300 2320 1312
rect 2275 1272 2320 1300
rect 2314 1260 2320 1272
rect 2372 1260 2378 1312
rect 2792 1272 3556 1300
rect 1489 1235 1547 1241
rect 1489 1201 1501 1235
rect 1535 1232 1547 1235
rect 1946 1232 1952 1244
rect 1535 1204 1952 1232
rect 1535 1201 1547 1204
rect 1489 1195 1547 1201
rect 1946 1192 1952 1204
rect 2004 1232 2010 1244
rect 2792 1232 2820 1272
rect 3528 1244 3556 1272
rect 3970 1260 3976 1312
rect 4028 1300 4034 1312
rect 4249 1303 4307 1309
rect 4249 1300 4261 1303
rect 4028 1272 4261 1300
rect 4028 1260 4034 1272
rect 4249 1269 4261 1272
rect 4295 1269 4307 1303
rect 4249 1263 4307 1269
rect 4338 1260 4344 1312
rect 4396 1300 4402 1312
rect 4433 1303 4491 1309
rect 4433 1300 4445 1303
rect 4396 1272 4445 1300
rect 4396 1260 4402 1272
rect 4433 1269 4445 1272
rect 4479 1269 4491 1303
rect 4433 1263 4491 1269
rect 4522 1260 4528 1312
rect 4580 1300 4586 1312
rect 4801 1303 4859 1309
rect 4580 1272 4625 1300
rect 4580 1260 4586 1272
rect 4801 1269 4813 1303
rect 4847 1300 4859 1303
rect 5626 1300 5632 1312
rect 4847 1272 5632 1300
rect 4847 1269 4859 1272
rect 4801 1263 4859 1269
rect 5626 1260 5632 1272
rect 5684 1260 5690 1312
rect 7285 1303 7343 1309
rect 7285 1269 7297 1303
rect 7331 1300 7343 1303
rect 8294 1300 8300 1312
rect 7331 1272 8300 1300
rect 7331 1269 7343 1272
rect 7285 1263 7343 1269
rect 8294 1260 8300 1272
rect 8352 1300 8358 1312
rect 9048 1309 9076 1476
rect 10336 1436 10364 1476
rect 10781 1473 10793 1507
rect 10827 1504 10839 1507
rect 11698 1504 11704 1516
rect 10827 1476 11704 1504
rect 10827 1473 10839 1476
rect 10781 1467 10839 1473
rect 11698 1464 11704 1476
rect 11756 1464 11762 1516
rect 12069 1439 12127 1445
rect 12069 1436 12081 1439
rect 10336 1408 12081 1436
rect 12069 1405 12081 1408
rect 12115 1436 12127 1439
rect 12434 1436 12440 1448
rect 12115 1408 12440 1436
rect 12115 1405 12127 1408
rect 12069 1399 12127 1405
rect 12434 1396 12440 1408
rect 12492 1396 12498 1448
rect 9309 1371 9367 1377
rect 9309 1337 9321 1371
rect 9355 1368 9367 1371
rect 11238 1368 11244 1380
rect 9355 1340 11244 1368
rect 9355 1337 9367 1340
rect 9309 1331 9367 1337
rect 11238 1328 11244 1340
rect 11296 1328 11302 1380
rect 9033 1303 9091 1309
rect 9033 1300 9045 1303
rect 8352 1272 9045 1300
rect 8352 1260 8358 1272
rect 9033 1269 9045 1272
rect 9079 1269 9091 1303
rect 11422 1300 11428 1312
rect 11383 1272 11428 1300
rect 9033 1263 9091 1269
rect 11422 1260 11428 1272
rect 11480 1260 11486 1312
rect 11882 1300 11888 1312
rect 11843 1272 11888 1300
rect 11882 1260 11888 1272
rect 11940 1260 11946 1312
rect 14277 1303 14335 1309
rect 14277 1269 14289 1303
rect 14323 1300 14335 1303
rect 14826 1300 14832 1312
rect 14323 1272 14832 1300
rect 14323 1269 14335 1272
rect 14277 1263 14335 1269
rect 14826 1260 14832 1272
rect 14884 1260 14890 1312
rect 14921 1303 14979 1309
rect 14921 1269 14933 1303
rect 14967 1269 14979 1303
rect 14921 1263 14979 1269
rect 2004 1204 2820 1232
rect 2004 1192 2010 1204
rect 2958 1192 2964 1244
rect 3016 1232 3022 1244
rect 3237 1235 3295 1241
rect 3237 1232 3249 1235
rect 3016 1204 3249 1232
rect 3016 1192 3022 1204
rect 3237 1201 3249 1204
rect 3283 1201 3295 1235
rect 3237 1195 3295 1201
rect 3421 1235 3479 1241
rect 3421 1201 3433 1235
rect 3467 1201 3479 1235
rect 3421 1195 3479 1201
rect 753 1167 811 1173
rect 753 1133 765 1167
rect 799 1164 811 1167
rect 1118 1164 1124 1176
rect 799 1136 1124 1164
rect 799 1133 811 1136
rect 753 1127 811 1133
rect 1118 1124 1124 1136
rect 1176 1124 1182 1176
rect 1302 1124 1308 1176
rect 1360 1164 1366 1176
rect 3436 1164 3464 1195
rect 3510 1192 3516 1244
rect 3568 1232 3574 1244
rect 5718 1232 5724 1244
rect 3568 1204 5724 1232
rect 3568 1192 3574 1204
rect 5718 1192 5724 1204
rect 5776 1232 5782 1244
rect 5776 1204 5842 1232
rect 5776 1192 5782 1204
rect 9582 1192 9588 1244
rect 9640 1232 9646 1244
rect 9640 1204 9798 1232
rect 9640 1192 9646 1204
rect 14550 1192 14556 1244
rect 14608 1232 14614 1244
rect 14936 1232 14964 1263
rect 14608 1204 14964 1232
rect 14608 1192 14614 1204
rect 11238 1164 11244 1176
rect 1360 1136 3464 1164
rect 11199 1136 11244 1164
rect 1360 1124 1366 1136
rect 11238 1124 11244 1136
rect 11296 1124 11302 1176
rect 14369 1167 14427 1173
rect 14369 1133 14381 1167
rect 14415 1164 14427 1167
rect 14918 1164 14924 1176
rect 14415 1136 14924 1164
rect 14415 1133 14427 1136
rect 14369 1127 14427 1133
rect 14918 1124 14924 1136
rect 14976 1124 14982 1176
rect 15105 1167 15163 1173
rect 15105 1133 15117 1167
rect 15151 1164 15163 1167
rect 15194 1164 15200 1176
rect 15151 1136 15200 1164
rect 15151 1133 15163 1136
rect 15105 1127 15163 1133
rect 15194 1124 15200 1136
rect 15252 1124 15258 1176
rect 92 1074 15824 1096
rect 92 1022 5242 1074
rect 5294 1022 5306 1074
rect 5358 1022 5370 1074
rect 5422 1022 5434 1074
rect 5486 1022 10514 1074
rect 10566 1022 10578 1074
rect 10630 1022 10642 1074
rect 10694 1022 10706 1074
rect 10758 1022 15824 1074
rect 92 1000 15824 1022
rect 4522 920 4528 972
rect 4580 960 4586 972
rect 5905 963 5963 969
rect 5905 960 5917 963
rect 4580 932 5917 960
rect 4580 920 4586 932
rect 5905 929 5917 932
rect 5951 929 5963 963
rect 6822 960 6828 972
rect 6783 932 6828 960
rect 5905 923 5963 929
rect 6822 920 6828 932
rect 6880 920 6886 972
rect 8662 920 8668 972
rect 8720 960 8726 972
rect 9125 963 9183 969
rect 9125 960 9137 963
rect 8720 932 9137 960
rect 8720 920 8726 932
rect 9125 929 9137 932
rect 9171 929 9183 963
rect 9125 923 9183 929
rect 1118 892 1124 904
rect 1079 864 1124 892
rect 1118 852 1124 864
rect 1176 852 1182 904
rect 3513 895 3571 901
rect 3513 861 3525 895
rect 3559 892 3571 895
rect 3786 892 3792 904
rect 3559 864 3792 892
rect 3559 861 3571 864
rect 3513 855 3571 861
rect 3786 852 3792 864
rect 3844 852 3850 904
rect 5074 852 5080 904
rect 5132 892 5138 904
rect 6057 895 6115 901
rect 6057 892 6069 895
rect 5132 864 6069 892
rect 5132 852 5138 864
rect 6057 861 6069 864
rect 6103 861 6115 895
rect 6270 892 6276 904
rect 6231 864 6276 892
rect 6057 855 6115 861
rect 6270 852 6276 864
rect 6328 852 6334 904
rect 11425 895 11483 901
rect 6380 864 10364 892
rect 2130 824 2136 836
rect 2091 796 2136 824
rect 2130 784 2136 796
rect 2188 784 2194 836
rect 5718 824 5724 836
rect 4646 796 5724 824
rect 5718 784 5724 796
rect 5776 784 5782 836
rect 1670 716 1676 768
rect 1728 756 1734 768
rect 3234 756 3240 768
rect 1728 728 3240 756
rect 1728 716 1734 728
rect 3234 716 3240 728
rect 3292 716 3298 768
rect 3510 716 3516 768
rect 3568 756 3574 768
rect 6380 756 6408 864
rect 6917 827 6975 833
rect 6917 793 6929 827
rect 6963 793 6975 827
rect 6917 787 6975 793
rect 7469 827 7527 833
rect 7469 793 7481 827
rect 7515 824 7527 827
rect 8386 824 8392 836
rect 7515 796 8392 824
rect 7515 793 7527 796
rect 7469 787 7527 793
rect 3568 728 6408 756
rect 3568 716 3574 728
rect 934 688 940 700
rect 895 660 940 688
rect 934 648 940 660
rect 992 648 998 700
rect 4614 648 4620 700
rect 4672 688 4678 700
rect 4985 691 5043 697
rect 4985 688 4997 691
rect 4672 660 4997 688
rect 4672 648 4678 660
rect 4985 657 4997 660
rect 5031 657 5043 691
rect 4985 651 5043 657
rect 2225 623 2283 629
rect 2225 589 2237 623
rect 2271 620 2283 623
rect 4890 620 4896 632
rect 2271 592 4896 620
rect 2271 589 2283 592
rect 2225 583 2283 589
rect 4890 580 4896 592
rect 4948 580 4954 632
rect 5534 580 5540 632
rect 5592 620 5598 632
rect 6089 623 6147 629
rect 6089 620 6101 623
rect 5592 592 6101 620
rect 5592 580 5598 592
rect 6089 589 6101 592
rect 6135 620 6147 623
rect 6932 620 6960 787
rect 8386 784 8392 796
rect 8444 784 8450 836
rect 9306 824 9312 836
rect 9267 796 9312 824
rect 9306 784 9312 796
rect 9364 784 9370 836
rect 9401 827 9459 833
rect 9401 793 9413 827
rect 9447 793 9459 827
rect 9401 787 9459 793
rect 9030 716 9036 768
rect 9088 756 9094 768
rect 9416 756 9444 787
rect 9490 784 9496 836
rect 9548 824 9554 836
rect 9677 827 9735 833
rect 9548 796 9593 824
rect 9548 784 9554 796
rect 9677 793 9689 827
rect 9723 824 9735 827
rect 9858 824 9864 836
rect 9723 796 9864 824
rect 9723 793 9735 796
rect 9677 787 9735 793
rect 9858 784 9864 796
rect 9916 784 9922 836
rect 10336 833 10364 864
rect 11425 861 11437 895
rect 11471 892 11483 895
rect 12250 892 12256 904
rect 11471 864 12256 892
rect 11471 861 11483 864
rect 11425 855 11483 861
rect 12250 852 12256 864
rect 12308 852 12314 904
rect 12802 892 12808 904
rect 12763 864 12808 892
rect 12802 852 12808 864
rect 12860 852 12866 904
rect 13998 852 14004 904
rect 14056 892 14062 904
rect 14185 895 14243 901
rect 14185 892 14197 895
rect 14056 864 14197 892
rect 14056 852 14062 864
rect 14185 861 14197 864
rect 14231 861 14243 895
rect 14918 892 14924 904
rect 14879 864 14924 892
rect 14185 855 14243 861
rect 14918 852 14924 864
rect 14976 852 14982 904
rect 10321 827 10379 833
rect 10321 793 10333 827
rect 10367 793 10379 827
rect 10321 787 10379 793
rect 9088 728 9444 756
rect 9088 716 9094 728
rect 7653 691 7711 697
rect 7653 657 7665 691
rect 7699 688 7711 691
rect 8938 688 8944 700
rect 7699 660 8944 688
rect 7699 657 7711 660
rect 7653 651 7711 657
rect 8938 648 8944 660
rect 8996 648 9002 700
rect 10870 648 10876 700
rect 10928 688 10934 700
rect 11241 691 11299 697
rect 11241 688 11253 691
rect 10928 660 11253 688
rect 10928 648 10934 660
rect 11241 657 11253 660
rect 11287 657 11299 691
rect 14366 688 14372 700
rect 14327 660 14372 688
rect 11241 651 11299 657
rect 14366 648 14372 660
rect 14424 648 14430 700
rect 10134 620 10140 632
rect 6135 592 6960 620
rect 10095 592 10140 620
rect 6135 589 6147 592
rect 6089 583 6147 589
rect 10134 580 10140 592
rect 10192 580 10198 632
rect 12894 620 12900 632
rect 12855 592 12900 620
rect 12894 580 12900 592
rect 12952 580 12958 632
rect 14918 580 14924 632
rect 14976 620 14982 632
rect 15013 623 15071 629
rect 15013 620 15025 623
rect 14976 592 15025 620
rect 14976 580 14982 592
rect 15013 589 15025 592
rect 15059 589 15071 623
rect 15013 583 15071 589
rect 92 530 15824 552
rect 92 478 2606 530
rect 2658 478 2670 530
rect 2722 478 2734 530
rect 2786 478 2798 530
rect 2850 478 7878 530
rect 7930 478 7942 530
rect 7994 478 8006 530
rect 8058 478 8070 530
rect 8122 478 13150 530
rect 13202 478 13214 530
rect 13266 478 13278 530
rect 13330 478 13342 530
rect 13394 478 15824 530
rect 92 456 15824 478
rect 2314 376 2320 428
rect 2372 416 2378 428
rect 10134 416 10140 428
rect 2372 388 10140 416
rect 2372 376 2378 388
rect 10134 376 10140 388
rect 10192 376 10198 428
rect 3234 308 3240 360
rect 3292 348 3298 360
rect 4798 348 4804 360
rect 3292 320 4804 348
rect 3292 308 3298 320
rect 4798 308 4804 320
rect 4856 348 4862 360
rect 11238 348 11244 360
rect 4856 320 11244 348
rect 4856 308 4862 320
rect 11238 308 11244 320
rect 11296 308 11302 360
rect 2130 240 2136 292
rect 2188 280 2194 292
rect 11146 280 11152 292
rect 2188 252 11152 280
rect 2188 240 2194 252
rect 11146 240 11152 252
rect 11204 240 11210 292
<< via1 >>
rect 5242 12990 5294 13042
rect 5306 12990 5358 13042
rect 5370 12990 5422 13042
rect 5434 12990 5486 13042
rect 10514 12990 10566 13042
rect 10578 12990 10630 13042
rect 10642 12990 10694 13042
rect 10706 12990 10758 13042
rect 4896 12931 4948 12940
rect 4896 12897 4905 12931
rect 4905 12897 4939 12931
rect 4939 12897 4948 12931
rect 4896 12888 4948 12897
rect 8944 12888 8996 12940
rect 12900 12931 12952 12940
rect 940 12863 992 12872
rect 940 12829 949 12863
rect 949 12829 983 12863
rect 983 12829 992 12863
rect 940 12820 992 12829
rect 2872 12820 2924 12872
rect 3976 12863 4028 12872
rect 3976 12829 3985 12863
rect 3985 12829 4019 12863
rect 4019 12829 4028 12863
rect 3976 12820 4028 12829
rect 6920 12863 6972 12872
rect 6920 12829 6929 12863
rect 6929 12829 6963 12863
rect 6963 12829 6972 12863
rect 12900 12897 12909 12931
rect 12909 12897 12943 12931
rect 12943 12897 12952 12931
rect 12900 12888 12952 12897
rect 14924 12888 14976 12940
rect 6920 12820 6972 12829
rect 10876 12820 10928 12872
rect 14372 12863 14424 12872
rect 14372 12829 14381 12863
rect 14381 12829 14415 12863
rect 14415 12829 14424 12863
rect 14372 12820 14424 12829
rect 1124 12795 1176 12804
rect 1124 12761 1133 12795
rect 1133 12761 1167 12795
rect 1167 12761 1176 12795
rect 1124 12752 1176 12761
rect 1860 12795 1912 12804
rect 1860 12761 1869 12795
rect 1869 12761 1903 12795
rect 1903 12761 1912 12795
rect 1860 12752 1912 12761
rect 3424 12795 3476 12804
rect 3424 12761 3433 12795
rect 3433 12761 3467 12795
rect 3467 12761 3476 12795
rect 3424 12752 3476 12761
rect 3516 12752 3568 12804
rect 4896 12752 4948 12804
rect 7196 12752 7248 12804
rect 8760 12795 8812 12804
rect 8760 12761 8769 12795
rect 8769 12761 8803 12795
rect 8803 12761 8812 12795
rect 8760 12752 8812 12761
rect 8944 12795 8996 12804
rect 8944 12761 8953 12795
rect 8953 12761 8987 12795
rect 8987 12761 8996 12795
rect 8944 12752 8996 12761
rect 9128 12752 9180 12804
rect 11428 12795 11480 12804
rect 11428 12761 11437 12795
rect 11437 12761 11471 12795
rect 11471 12761 11480 12795
rect 11428 12752 11480 12761
rect 12808 12795 12860 12804
rect 12808 12761 12817 12795
rect 12817 12761 12851 12795
rect 12851 12761 12860 12795
rect 12808 12752 12860 12761
rect 14188 12795 14240 12804
rect 14188 12761 14197 12795
rect 14197 12761 14231 12795
rect 14231 12761 14240 12795
rect 14188 12752 14240 12761
rect 14832 12752 14884 12804
rect 7748 12684 7800 12736
rect 12072 12616 12124 12668
rect 1768 12591 1820 12600
rect 1768 12557 1777 12591
rect 1777 12557 1811 12591
rect 1811 12557 1820 12591
rect 1768 12548 1820 12557
rect 9128 12591 9180 12600
rect 9128 12557 9137 12591
rect 9137 12557 9171 12591
rect 9171 12557 9180 12591
rect 9128 12548 9180 12557
rect 2606 12446 2658 12498
rect 2670 12446 2722 12498
rect 2734 12446 2786 12498
rect 2798 12446 2850 12498
rect 7878 12446 7930 12498
rect 7942 12446 7994 12498
rect 8006 12446 8058 12498
rect 8070 12446 8122 12498
rect 13150 12446 13202 12498
rect 13214 12446 13266 12498
rect 13278 12446 13330 12498
rect 13342 12446 13394 12498
rect 940 12344 992 12396
rect 8760 12344 8812 12396
rect 9496 12344 9548 12396
rect 572 12183 624 12192
rect 572 12149 581 12183
rect 581 12149 615 12183
rect 615 12149 624 12183
rect 572 12140 624 12149
rect 6460 12208 6512 12260
rect 4344 12183 4396 12192
rect 848 12115 900 12124
rect 848 12081 857 12115
rect 857 12081 891 12115
rect 891 12081 900 12115
rect 848 12072 900 12081
rect 2504 12072 2556 12124
rect 4344 12149 4353 12183
rect 4353 12149 4387 12183
rect 4387 12149 4396 12183
rect 4344 12140 4396 12149
rect 4528 12183 4580 12192
rect 4528 12149 4537 12183
rect 4537 12149 4571 12183
rect 4571 12149 4580 12183
rect 4528 12140 4580 12149
rect 7196 12183 7248 12192
rect 7196 12149 7205 12183
rect 7205 12149 7239 12183
rect 7239 12149 7248 12183
rect 7196 12140 7248 12149
rect 8208 12140 8260 12192
rect 8944 12208 8996 12260
rect 9404 12208 9456 12260
rect 9864 12208 9916 12260
rect 8852 12183 8904 12192
rect 8852 12149 8861 12183
rect 8861 12149 8895 12183
rect 8895 12149 8904 12183
rect 8852 12140 8904 12149
rect 9588 12140 9640 12192
rect 3240 12072 3292 12124
rect 3516 12115 3568 12124
rect 3516 12081 3525 12115
rect 3525 12081 3559 12115
rect 3559 12081 3568 12115
rect 3516 12072 3568 12081
rect 3700 12115 3752 12124
rect 3700 12081 3709 12115
rect 3709 12081 3743 12115
rect 3743 12081 3752 12115
rect 3700 12072 3752 12081
rect 4804 12072 4856 12124
rect 6920 12072 6972 12124
rect 8944 12115 8996 12124
rect 8944 12081 8979 12115
rect 8979 12081 8996 12115
rect 8944 12072 8996 12081
rect 10876 12072 10928 12124
rect 11152 12115 11204 12124
rect 11152 12081 11161 12115
rect 11161 12081 11195 12115
rect 11195 12081 11204 12115
rect 11152 12072 11204 12081
rect 14280 12072 14332 12124
rect 15108 12115 15160 12124
rect 15108 12081 15117 12115
rect 15117 12081 15151 12115
rect 15151 12081 15160 12115
rect 15108 12072 15160 12081
rect 4160 12004 4212 12056
rect 4712 12004 4764 12056
rect 5540 12004 5592 12056
rect 7288 12047 7340 12056
rect 7288 12013 7297 12047
rect 7297 12013 7331 12047
rect 7331 12013 7340 12047
rect 7288 12004 7340 12013
rect 8668 12004 8720 12056
rect 5242 11902 5294 11954
rect 5306 11902 5358 11954
rect 5370 11902 5422 11954
rect 5434 11902 5486 11954
rect 10514 11902 10566 11954
rect 10578 11902 10630 11954
rect 10642 11902 10694 11954
rect 10706 11902 10758 11954
rect 1860 11800 1912 11852
rect 3976 11800 4028 11852
rect 940 11775 992 11784
rect 940 11741 949 11775
rect 949 11741 983 11775
rect 983 11741 992 11775
rect 940 11732 992 11741
rect 1308 11732 1360 11784
rect 2504 11732 2556 11784
rect 7196 11800 7248 11852
rect 9404 11800 9456 11852
rect 9588 11800 9640 11852
rect 11152 11843 11204 11852
rect 11152 11809 11161 11843
rect 11161 11809 11195 11843
rect 11195 11809 11204 11843
rect 11152 11800 11204 11809
rect 14188 11800 14240 11852
rect 572 11664 624 11716
rect 4712 11707 4764 11716
rect 4712 11673 4721 11707
rect 4721 11673 4755 11707
rect 4755 11673 4764 11707
rect 4712 11664 4764 11673
rect 6460 11732 6512 11784
rect 8392 11732 8444 11784
rect 8668 11775 8720 11784
rect 8668 11741 8677 11775
rect 8677 11741 8711 11775
rect 8711 11741 8720 11775
rect 8668 11732 8720 11741
rect 9956 11732 10008 11784
rect 10876 11732 10928 11784
rect 8300 11664 8352 11716
rect 11152 11664 11204 11716
rect 8392 11639 8444 11648
rect 8392 11605 8401 11639
rect 8401 11605 8435 11639
rect 8435 11605 8444 11639
rect 8392 11596 8444 11605
rect 756 11571 808 11580
rect 756 11537 765 11571
rect 765 11537 799 11571
rect 799 11537 808 11571
rect 756 11528 808 11537
rect 9680 11596 9732 11648
rect 10048 11596 10100 11648
rect 14004 11664 14056 11716
rect 3608 11460 3660 11512
rect 7564 11460 7616 11512
rect 8852 11460 8904 11512
rect 2606 11358 2658 11410
rect 2670 11358 2722 11410
rect 2734 11358 2786 11410
rect 2798 11358 2850 11410
rect 7878 11358 7930 11410
rect 7942 11358 7994 11410
rect 8006 11358 8058 11410
rect 8070 11358 8122 11410
rect 13150 11358 13202 11410
rect 13214 11358 13266 11410
rect 13278 11358 13330 11410
rect 13342 11358 13394 11410
rect 848 11256 900 11308
rect 3608 11256 3660 11308
rect 6920 11299 6972 11308
rect 6920 11265 6929 11299
rect 6929 11265 6963 11299
rect 6963 11265 6972 11299
rect 6920 11256 6972 11265
rect 8300 11256 8352 11308
rect 8576 11256 8628 11308
rect 9956 11256 10008 11308
rect 14280 11299 14332 11308
rect 14280 11265 14289 11299
rect 14289 11265 14323 11299
rect 14323 11265 14332 11299
rect 14280 11256 14332 11265
rect 1860 11095 1912 11104
rect 1860 11061 1869 11095
rect 1869 11061 1903 11095
rect 1903 11061 1912 11095
rect 1860 11052 1912 11061
rect 3424 11188 3476 11240
rect 3700 11120 3752 11172
rect 6184 11120 6236 11172
rect 3240 11095 3292 11104
rect 3240 11061 3249 11095
rect 3249 11061 3283 11095
rect 3283 11061 3292 11095
rect 3240 11052 3292 11061
rect 3516 11095 3568 11104
rect 3516 11061 3525 11095
rect 3525 11061 3559 11095
rect 3559 11061 3568 11095
rect 3976 11095 4028 11104
rect 3516 11052 3568 11061
rect 756 11027 808 11036
rect 756 10993 765 11027
rect 765 10993 799 11027
rect 799 10993 808 11027
rect 756 10984 808 10993
rect 3700 10984 3752 11036
rect 3976 11061 3985 11095
rect 3985 11061 4019 11095
rect 4019 11061 4028 11095
rect 3976 11052 4028 11061
rect 4068 11052 4120 11104
rect 4436 11052 4488 11104
rect 6460 11095 6512 11104
rect 6460 11061 6469 11095
rect 6469 11061 6503 11095
rect 6503 11061 6512 11095
rect 6460 11052 6512 11061
rect 6828 11052 6880 11104
rect 7472 11188 7524 11240
rect 8944 11188 8996 11240
rect 7380 11120 7432 11172
rect 8208 11120 8260 11172
rect 8300 11120 8352 11172
rect 8392 11120 8444 11172
rect 9864 11163 9916 11172
rect 9864 11129 9873 11163
rect 9873 11129 9907 11163
rect 9907 11129 9916 11163
rect 9864 11120 9916 11129
rect 7196 11095 7248 11104
rect 7196 11061 7205 11095
rect 7205 11061 7239 11095
rect 7239 11061 7248 11095
rect 7196 11052 7248 11061
rect 8852 11095 8904 11104
rect 5540 10984 5592 11036
rect 5908 10984 5960 11036
rect 6276 10984 6328 11036
rect 7472 10984 7524 11036
rect 8852 11061 8861 11095
rect 8861 11061 8895 11095
rect 8895 11061 8904 11095
rect 8852 11052 8904 11061
rect 8944 11095 8996 11104
rect 8944 11061 8979 11095
rect 8979 11061 8996 11095
rect 8944 11052 8996 11061
rect 9404 11052 9456 11104
rect 13820 11052 13872 11104
rect 7656 10984 7708 11036
rect 10140 11027 10192 11036
rect 10140 10993 10149 11027
rect 10149 10993 10183 11027
rect 10183 10993 10192 11027
rect 10140 10984 10192 10993
rect 10876 10984 10928 11036
rect 14924 11027 14976 11036
rect 14924 10993 14933 11027
rect 14933 10993 14967 11027
rect 14967 10993 14976 11027
rect 14924 10984 14976 10993
rect 15108 11027 15160 11036
rect 15108 10993 15117 11027
rect 15117 10993 15151 11027
rect 15151 10993 15160 11027
rect 15108 10984 15160 10993
rect 10968 10916 11020 10968
rect 5242 10814 5294 10866
rect 5306 10814 5358 10866
rect 5370 10814 5422 10866
rect 5434 10814 5486 10866
rect 10514 10814 10566 10866
rect 10578 10814 10630 10866
rect 10642 10814 10694 10866
rect 10706 10814 10758 10866
rect 1492 10644 1544 10696
rect 2504 10712 2556 10764
rect 572 10576 624 10628
rect 1216 10551 1268 10560
rect 1216 10517 1225 10551
rect 1225 10517 1259 10551
rect 1259 10517 1268 10551
rect 1216 10508 1268 10517
rect 940 10372 992 10424
rect 3516 10576 3568 10628
rect 4988 10644 5040 10696
rect 5908 10712 5960 10764
rect 7472 10712 7524 10764
rect 9404 10755 9456 10764
rect 6092 10687 6144 10696
rect 6092 10653 6101 10687
rect 6101 10653 6135 10687
rect 6135 10653 6144 10687
rect 6092 10644 6144 10653
rect 4252 10576 4304 10628
rect 4896 10576 4948 10628
rect 6000 10619 6052 10628
rect 6000 10585 6009 10619
rect 6009 10585 6043 10619
rect 6043 10585 6052 10619
rect 6000 10576 6052 10585
rect 6276 10576 6328 10628
rect 6460 10576 6512 10628
rect 6552 10508 6604 10560
rect 7012 10644 7064 10696
rect 9404 10721 9413 10755
rect 9413 10721 9447 10755
rect 9447 10721 9456 10755
rect 9404 10712 9456 10721
rect 9588 10712 9640 10764
rect 11060 10755 11112 10764
rect 11060 10721 11069 10755
rect 11069 10721 11103 10755
rect 11103 10721 11112 10755
rect 11060 10712 11112 10721
rect 11428 10712 11480 10764
rect 8576 10644 8628 10696
rect 9312 10619 9364 10628
rect 9312 10585 9321 10619
rect 9321 10585 9355 10619
rect 9355 10585 9364 10619
rect 9312 10576 9364 10585
rect 9496 10576 9548 10628
rect 9680 10576 9732 10628
rect 9956 10576 10008 10628
rect 10968 10576 11020 10628
rect 11612 10576 11664 10628
rect 12072 10619 12124 10628
rect 12072 10585 12081 10619
rect 12081 10585 12115 10619
rect 12115 10585 12124 10619
rect 12072 10576 12124 10585
rect 6828 10551 6880 10560
rect 6828 10517 6837 10551
rect 6837 10517 6871 10551
rect 6871 10517 6880 10551
rect 7104 10551 7156 10560
rect 6828 10508 6880 10517
rect 7104 10517 7113 10551
rect 7113 10517 7147 10551
rect 7147 10517 7156 10551
rect 7104 10508 7156 10517
rect 7748 10508 7800 10560
rect 11520 10508 11572 10560
rect 11888 10508 11940 10560
rect 15568 10576 15620 10628
rect 3148 10415 3200 10424
rect 3148 10381 3157 10415
rect 3157 10381 3191 10415
rect 3191 10381 3200 10415
rect 3148 10372 3200 10381
rect 4712 10372 4764 10424
rect 4896 10372 4948 10424
rect 6460 10372 6512 10424
rect 8208 10372 8260 10424
rect 10048 10440 10100 10492
rect 12716 10415 12768 10424
rect 12716 10381 12725 10415
rect 12725 10381 12759 10415
rect 12759 10381 12768 10415
rect 12716 10372 12768 10381
rect 15016 10372 15068 10424
rect 2606 10270 2658 10322
rect 2670 10270 2722 10322
rect 2734 10270 2786 10322
rect 2798 10270 2850 10322
rect 7878 10270 7930 10322
rect 7942 10270 7994 10322
rect 8006 10270 8058 10322
rect 8070 10270 8122 10322
rect 13150 10270 13202 10322
rect 13214 10270 13266 10322
rect 13278 10270 13330 10322
rect 13342 10270 13394 10322
rect 1216 10168 1268 10220
rect 1308 10211 1360 10220
rect 1308 10177 1317 10211
rect 1317 10177 1351 10211
rect 1351 10177 1360 10211
rect 1308 10168 1360 10177
rect 1860 10168 1912 10220
rect 2136 10100 2188 10152
rect 3516 10143 3568 10152
rect 3148 10032 3200 10084
rect 3516 10109 3525 10143
rect 3525 10109 3559 10143
rect 3559 10109 3568 10143
rect 3516 10100 3568 10109
rect 4528 10032 4580 10084
rect 4712 10168 4764 10220
rect 6000 10100 6052 10152
rect 6828 10100 6880 10152
rect 6920 10100 6972 10152
rect 7932 10100 7984 10152
rect 8300 10100 8352 10152
rect 3424 9964 3476 10016
rect 6000 10007 6052 10016
rect 6000 9973 6009 10007
rect 6009 9973 6043 10007
rect 6043 9973 6052 10007
rect 6000 9964 6052 9973
rect 1860 9896 1912 9948
rect 2136 9939 2188 9948
rect 2136 9905 2145 9939
rect 2145 9905 2179 9939
rect 2179 9905 2188 9939
rect 2136 9896 2188 9905
rect 3516 9896 3568 9948
rect 5724 9939 5776 9948
rect 1400 9828 1452 9880
rect 2596 9828 2648 9880
rect 4436 9828 4488 9880
rect 5724 9905 5733 9939
rect 5733 9905 5767 9939
rect 5767 9905 5776 9939
rect 5724 9896 5776 9905
rect 6552 9964 6604 10016
rect 9312 9964 9364 10016
rect 5540 9828 5592 9880
rect 7472 9896 7524 9948
rect 8208 9896 8260 9948
rect 10140 10168 10192 10220
rect 14924 10168 14976 10220
rect 12164 10100 12216 10152
rect 11060 10007 11112 10016
rect 6184 9828 6236 9880
rect 7564 9828 7616 9880
rect 7656 9828 7708 9880
rect 9588 9871 9640 9880
rect 9588 9837 9597 9871
rect 9597 9837 9631 9871
rect 9631 9837 9640 9871
rect 9588 9828 9640 9837
rect 9956 9896 10008 9948
rect 11060 9973 11069 10007
rect 11069 9973 11103 10007
rect 11103 9973 11112 10007
rect 11060 9964 11112 9973
rect 11520 10007 11572 10016
rect 11520 9973 11529 10007
rect 11529 9973 11563 10007
rect 11563 9973 11572 10007
rect 11520 9964 11572 9973
rect 12808 10032 12860 10084
rect 14740 9964 14792 10016
rect 11152 9896 11204 9948
rect 14924 9939 14976 9948
rect 14924 9905 14933 9939
rect 14933 9905 14967 9939
rect 14967 9905 14976 9939
rect 14924 9896 14976 9905
rect 15108 9939 15160 9948
rect 15108 9905 15117 9939
rect 15117 9905 15151 9939
rect 15151 9905 15160 9939
rect 15108 9896 15160 9905
rect 11888 9828 11940 9880
rect 12808 9828 12860 9880
rect 5242 9726 5294 9778
rect 5306 9726 5358 9778
rect 5370 9726 5422 9778
rect 5434 9726 5486 9778
rect 10514 9726 10566 9778
rect 10578 9726 10630 9778
rect 10642 9726 10694 9778
rect 10706 9726 10758 9778
rect 1492 9624 1544 9676
rect 940 9599 992 9608
rect 940 9565 949 9599
rect 949 9565 983 9599
rect 983 9565 992 9599
rect 940 9556 992 9565
rect 2596 9624 2648 9676
rect 5724 9624 5776 9676
rect 4712 9556 4764 9608
rect 572 9488 624 9540
rect 1308 9488 1360 9540
rect 4436 9531 4488 9540
rect 4436 9497 4445 9531
rect 4445 9497 4479 9531
rect 4479 9497 4488 9531
rect 4436 9488 4488 9497
rect 7012 9624 7064 9676
rect 7104 9624 7156 9676
rect 6552 9556 6604 9608
rect 14924 9624 14976 9676
rect 756 9463 808 9472
rect 756 9429 765 9463
rect 765 9429 799 9463
rect 799 9429 808 9463
rect 756 9420 808 9429
rect 1768 9463 1820 9472
rect 1768 9429 1777 9463
rect 1777 9429 1811 9463
rect 1811 9429 1820 9463
rect 1768 9420 1820 9429
rect 3240 9463 3292 9472
rect 3240 9429 3249 9463
rect 3249 9429 3283 9463
rect 3283 9429 3292 9463
rect 3240 9420 3292 9429
rect 5908 9420 5960 9472
rect 6920 9488 6972 9540
rect 7380 9531 7432 9540
rect 7380 9497 7389 9531
rect 7389 9497 7423 9531
rect 7423 9497 7432 9531
rect 7380 9488 7432 9497
rect 6644 9420 6696 9472
rect 7104 9352 7156 9404
rect 4528 9284 4580 9336
rect 6920 9284 6972 9336
rect 7932 9488 7984 9540
rect 8392 9488 8444 9540
rect 8668 9488 8720 9540
rect 9128 9531 9180 9540
rect 9128 9497 9137 9531
rect 9137 9497 9171 9531
rect 9171 9497 9180 9531
rect 9128 9488 9180 9497
rect 10140 9531 10192 9540
rect 10140 9497 10149 9531
rect 10149 9497 10183 9531
rect 10183 9497 10192 9531
rect 10140 9488 10192 9497
rect 8208 9420 8260 9472
rect 7564 9352 7616 9404
rect 8576 9420 8628 9472
rect 11520 9531 11572 9540
rect 11520 9497 11529 9531
rect 11529 9497 11563 9531
rect 11563 9497 11572 9531
rect 11796 9531 11848 9540
rect 11520 9488 11572 9497
rect 11796 9497 11805 9531
rect 11805 9497 11839 9531
rect 11839 9497 11848 9531
rect 11796 9488 11848 9497
rect 12256 9531 12308 9540
rect 12256 9497 12265 9531
rect 12265 9497 12299 9531
rect 12299 9497 12308 9531
rect 12256 9488 12308 9497
rect 12440 9531 12492 9540
rect 12440 9497 12442 9531
rect 12442 9497 12476 9531
rect 12476 9497 12492 9531
rect 12440 9488 12492 9497
rect 12624 9488 12676 9540
rect 13636 9488 13688 9540
rect 13912 9488 13964 9540
rect 14648 9531 14700 9540
rect 14648 9497 14657 9531
rect 14657 9497 14691 9531
rect 14691 9497 14700 9531
rect 14648 9488 14700 9497
rect 12072 9420 12124 9472
rect 8392 9352 8444 9404
rect 14464 9352 14516 9404
rect 14832 9352 14884 9404
rect 7656 9284 7708 9336
rect 9036 9327 9088 9336
rect 9036 9293 9045 9327
rect 9045 9293 9079 9327
rect 9079 9293 9088 9327
rect 9036 9284 9088 9293
rect 10048 9327 10100 9336
rect 10048 9293 10057 9327
rect 10057 9293 10091 9327
rect 10091 9293 10100 9327
rect 10048 9284 10100 9293
rect 11428 9284 11480 9336
rect 12256 9284 12308 9336
rect 12532 9284 12584 9336
rect 14096 9327 14148 9336
rect 14096 9293 14105 9327
rect 14105 9293 14139 9327
rect 14139 9293 14148 9327
rect 14096 9284 14148 9293
rect 2606 9182 2658 9234
rect 2670 9182 2722 9234
rect 2734 9182 2786 9234
rect 2798 9182 2850 9234
rect 7878 9182 7930 9234
rect 7942 9182 7994 9234
rect 8006 9182 8058 9234
rect 8070 9182 8122 9234
rect 13150 9182 13202 9234
rect 13214 9182 13266 9234
rect 13278 9182 13330 9234
rect 13342 9182 13394 9234
rect 4344 9080 4396 9132
rect 6460 9080 6512 9132
rect 2044 9012 2096 9064
rect 1308 8944 1360 8996
rect 2504 8944 2556 8996
rect 3516 9012 3568 9064
rect 6920 9012 6972 9064
rect 8668 9012 8720 9064
rect 756 8851 808 8860
rect 756 8817 765 8851
rect 765 8817 799 8851
rect 799 8817 808 8851
rect 756 8808 808 8817
rect 1860 8851 1912 8860
rect 1860 8817 1869 8851
rect 1869 8817 1903 8851
rect 1903 8817 1912 8851
rect 1860 8808 1912 8817
rect 2964 8876 3016 8928
rect 3240 8919 3292 8928
rect 3240 8885 3249 8919
rect 3249 8885 3283 8919
rect 3283 8885 3292 8919
rect 3240 8876 3292 8885
rect 9864 8944 9916 8996
rect 11060 8944 11112 8996
rect 3516 8919 3568 8928
rect 3516 8885 3525 8919
rect 3525 8885 3559 8919
rect 3559 8885 3568 8919
rect 3516 8876 3568 8885
rect 4252 8919 4304 8928
rect 4252 8885 4269 8919
rect 4269 8885 4304 8919
rect 4252 8876 4304 8885
rect 4436 8919 4488 8928
rect 4436 8885 4445 8919
rect 4445 8885 4479 8919
rect 4479 8885 4488 8919
rect 4436 8876 4488 8885
rect 4620 8876 4672 8928
rect 5540 8876 5592 8928
rect 6920 8919 6972 8928
rect 6920 8885 6929 8919
rect 6929 8885 6963 8919
rect 6963 8885 6972 8919
rect 6920 8876 6972 8885
rect 7196 8876 7248 8928
rect 9312 8876 9364 8928
rect 9404 8919 9456 8928
rect 9404 8885 9413 8919
rect 9413 8885 9447 8919
rect 9447 8885 9456 8919
rect 9404 8876 9456 8885
rect 4988 8808 5040 8860
rect 4620 8740 4672 8792
rect 8760 8740 8812 8792
rect 9496 8740 9548 8792
rect 9956 8740 10008 8792
rect 10876 8740 10928 8792
rect 12256 8944 12308 8996
rect 13452 8876 13504 8928
rect 12072 8808 12124 8860
rect 11980 8740 12032 8792
rect 14096 8876 14148 8928
rect 14188 8808 14240 8860
rect 14924 8851 14976 8860
rect 14924 8817 14933 8851
rect 14933 8817 14967 8851
rect 14967 8817 14976 8851
rect 14924 8808 14976 8817
rect 15108 8851 15160 8860
rect 15108 8817 15117 8851
rect 15117 8817 15151 8851
rect 15151 8817 15160 8851
rect 15108 8808 15160 8817
rect 14280 8740 14332 8792
rect 5242 8638 5294 8690
rect 5306 8638 5358 8690
rect 5370 8638 5422 8690
rect 5434 8638 5486 8690
rect 10514 8638 10566 8690
rect 10578 8638 10630 8690
rect 10642 8638 10694 8690
rect 10706 8638 10758 8690
rect 664 8579 716 8588
rect 664 8545 673 8579
rect 673 8545 707 8579
rect 707 8545 716 8579
rect 664 8536 716 8545
rect 5908 8536 5960 8588
rect 9312 8579 9364 8588
rect 1492 8468 1544 8520
rect 1860 8468 1912 8520
rect 4620 8511 4672 8520
rect 4620 8477 4629 8511
rect 4629 8477 4663 8511
rect 4663 8477 4672 8511
rect 4620 8468 4672 8477
rect 5540 8468 5592 8520
rect 7104 8468 7156 8520
rect 2504 8400 2556 8452
rect 4344 8400 4396 8452
rect 4712 8443 4764 8452
rect 4160 8332 4212 8384
rect 4712 8409 4721 8443
rect 4721 8409 4755 8443
rect 4755 8409 4764 8443
rect 4712 8400 4764 8409
rect 4988 8400 5040 8452
rect 9312 8545 9321 8579
rect 9321 8545 9355 8579
rect 9355 8545 9364 8579
rect 9312 8536 9364 8545
rect 11796 8536 11848 8588
rect 11980 8511 12032 8520
rect 9588 8400 9640 8452
rect 7656 8375 7708 8384
rect 3240 8307 3292 8316
rect 3240 8273 3249 8307
rect 3249 8273 3283 8307
rect 3283 8273 3292 8307
rect 3240 8264 3292 8273
rect 3332 8264 3384 8316
rect 7656 8341 7665 8375
rect 7665 8341 7699 8375
rect 7699 8341 7708 8375
rect 7656 8332 7708 8341
rect 9772 8375 9824 8384
rect 9772 8341 9781 8375
rect 9781 8341 9815 8375
rect 9815 8341 9824 8375
rect 9772 8332 9824 8341
rect 10048 8400 10100 8452
rect 10876 8400 10928 8452
rect 11980 8477 11989 8511
rect 11989 8477 12023 8511
rect 12023 8477 12032 8511
rect 11980 8468 12032 8477
rect 13452 8468 13504 8520
rect 11336 8400 11388 8452
rect 12256 8443 12308 8452
rect 12256 8409 12265 8443
rect 12265 8409 12299 8443
rect 12299 8409 12308 8443
rect 12256 8400 12308 8409
rect 12716 8443 12768 8452
rect 12716 8409 12725 8443
rect 12725 8409 12759 8443
rect 12759 8409 12768 8443
rect 12716 8400 12768 8409
rect 11152 8332 11204 8384
rect 8300 8264 8352 8316
rect 9036 8264 9088 8316
rect 9864 8264 9916 8316
rect 11520 8264 11572 8316
rect 12900 8332 12952 8384
rect 6000 8196 6052 8248
rect 7196 8196 7248 8248
rect 9680 8196 9732 8248
rect 13912 8196 13964 8248
rect 2606 8094 2658 8146
rect 2670 8094 2722 8146
rect 2734 8094 2786 8146
rect 2798 8094 2850 8146
rect 7878 8094 7930 8146
rect 7942 8094 7994 8146
rect 8006 8094 8058 8146
rect 8070 8094 8122 8146
rect 13150 8094 13202 8146
rect 13214 8094 13266 8146
rect 13278 8094 13330 8146
rect 13342 8094 13394 8146
rect 1124 7924 1176 7976
rect 4160 7992 4212 8044
rect 5908 7992 5960 8044
rect 7656 7992 7708 8044
rect 4988 7924 5040 7976
rect 8484 7924 8536 7976
rect 5908 7899 5960 7908
rect 5908 7865 5917 7899
rect 5917 7865 5951 7899
rect 5951 7865 5960 7899
rect 5908 7856 5960 7865
rect 7196 7856 7248 7908
rect 9864 7992 9916 8044
rect 10140 7992 10192 8044
rect 11060 8035 11112 8044
rect 11060 8001 11069 8035
rect 11069 8001 11103 8035
rect 11103 8001 11112 8035
rect 11060 7992 11112 8001
rect 11336 7992 11388 8044
rect 11704 7992 11756 8044
rect 12900 7992 12952 8044
rect 11244 7924 11296 7976
rect 12256 7924 12308 7976
rect 8760 7899 8812 7908
rect 664 7831 716 7840
rect 664 7797 673 7831
rect 673 7797 707 7831
rect 707 7797 716 7831
rect 664 7788 716 7797
rect 480 7763 532 7772
rect 480 7729 489 7763
rect 489 7729 523 7763
rect 523 7729 532 7763
rect 480 7720 532 7729
rect 572 7652 624 7704
rect 3424 7831 3476 7840
rect 3424 7797 3433 7831
rect 3433 7797 3467 7831
rect 3467 7797 3476 7831
rect 3424 7788 3476 7797
rect 4068 7831 4120 7840
rect 4068 7797 4077 7831
rect 4077 7797 4111 7831
rect 4111 7797 4120 7831
rect 4068 7788 4120 7797
rect 7472 7831 7524 7840
rect 2964 7720 3016 7772
rect 3148 7720 3200 7772
rect 4712 7720 4764 7772
rect 6644 7720 6696 7772
rect 7472 7797 7481 7831
rect 7481 7797 7515 7831
rect 7515 7797 7524 7831
rect 7472 7788 7524 7797
rect 8760 7865 8769 7899
rect 8769 7865 8803 7899
rect 8803 7865 8812 7899
rect 8760 7856 8812 7865
rect 11980 7856 12032 7908
rect 7380 7720 7432 7772
rect 3332 7652 3384 7704
rect 3792 7652 3844 7704
rect 5724 7652 5776 7704
rect 6828 7652 6880 7704
rect 7840 7652 7892 7704
rect 10048 7720 10100 7772
rect 11060 7720 11112 7772
rect 11336 7831 11388 7840
rect 11336 7797 11345 7831
rect 11345 7797 11379 7831
rect 11379 7797 11388 7831
rect 12532 7831 12584 7840
rect 11336 7788 11388 7797
rect 12532 7797 12541 7831
rect 12541 7797 12575 7831
rect 12575 7797 12584 7831
rect 12532 7788 12584 7797
rect 14372 7856 14424 7908
rect 13912 7831 13964 7840
rect 13912 7797 13938 7831
rect 13938 7797 13964 7831
rect 13912 7788 13964 7797
rect 14096 7788 14148 7840
rect 9496 7652 9548 7704
rect 13728 7695 13780 7704
rect 13728 7661 13737 7695
rect 13737 7661 13771 7695
rect 13771 7661 13780 7695
rect 13728 7652 13780 7661
rect 14096 7652 14148 7704
rect 5242 7550 5294 7602
rect 5306 7550 5358 7602
rect 5370 7550 5422 7602
rect 5434 7550 5486 7602
rect 10514 7550 10566 7602
rect 10578 7550 10630 7602
rect 10642 7550 10694 7602
rect 10706 7550 10758 7602
rect 3148 7448 3200 7500
rect 3976 7448 4028 7500
rect 1492 7380 1544 7432
rect 8576 7448 8628 7500
rect 9404 7448 9456 7500
rect 9956 7448 10008 7500
rect 11152 7448 11204 7500
rect 2504 7312 2556 7364
rect 3516 7312 3568 7364
rect 572 7108 624 7160
rect 664 7108 716 7160
rect 3792 7176 3844 7228
rect 5540 7312 5592 7364
rect 4988 7244 5040 7296
rect 5080 7244 5132 7296
rect 6460 7380 6512 7432
rect 7840 7423 7892 7432
rect 7840 7389 7849 7423
rect 7849 7389 7883 7423
rect 7883 7389 7892 7423
rect 7840 7380 7892 7389
rect 10876 7380 10928 7432
rect 6736 7312 6788 7364
rect 7012 7355 7064 7364
rect 7012 7321 7021 7355
rect 7021 7321 7055 7355
rect 7055 7321 7064 7355
rect 7012 7312 7064 7321
rect 7564 7355 7616 7364
rect 7564 7321 7573 7355
rect 7573 7321 7607 7355
rect 7607 7321 7616 7355
rect 7564 7312 7616 7321
rect 9496 7312 9548 7364
rect 9864 7312 9916 7364
rect 11244 7355 11296 7364
rect 11244 7321 11253 7355
rect 11253 7321 11287 7355
rect 11287 7321 11296 7355
rect 11244 7312 11296 7321
rect 11428 7380 11480 7432
rect 11704 7312 11756 7364
rect 13452 7380 13504 7432
rect 12716 7355 12768 7364
rect 12716 7321 12725 7355
rect 12725 7321 12759 7355
rect 12759 7321 12768 7355
rect 12716 7312 12768 7321
rect 10140 7244 10192 7296
rect 12992 7244 13044 7296
rect 6828 7176 6880 7228
rect 3056 7151 3108 7160
rect 3056 7117 3065 7151
rect 3065 7117 3099 7151
rect 3099 7117 3108 7151
rect 3056 7108 3108 7117
rect 5632 7108 5684 7160
rect 5816 7151 5868 7160
rect 5816 7117 5825 7151
rect 5825 7117 5859 7151
rect 5859 7117 5868 7151
rect 5816 7108 5868 7117
rect 6184 7108 6236 7160
rect 14556 7244 14608 7296
rect 13912 7108 13964 7160
rect 2606 7006 2658 7058
rect 2670 7006 2722 7058
rect 2734 7006 2786 7058
rect 2798 7006 2850 7058
rect 7878 7006 7930 7058
rect 7942 7006 7994 7058
rect 8006 7006 8058 7058
rect 8070 7006 8122 7058
rect 13150 7006 13202 7058
rect 13214 7006 13266 7058
rect 13278 7006 13330 7058
rect 13342 7006 13394 7058
rect 3148 6904 3200 6956
rect 3424 6947 3476 6956
rect 3424 6913 3433 6947
rect 3433 6913 3467 6947
rect 3467 6913 3476 6947
rect 3424 6904 3476 6913
rect 4068 6904 4120 6956
rect 4160 6836 4212 6888
rect 4436 6879 4488 6888
rect 4436 6845 4445 6879
rect 4445 6845 4479 6879
rect 4479 6845 4488 6879
rect 4436 6836 4488 6845
rect 5632 6836 5684 6888
rect 6644 6836 6696 6888
rect 7472 6904 7524 6956
rect 4528 6811 4580 6820
rect 572 6700 624 6752
rect 2320 6743 2372 6752
rect 756 6675 808 6684
rect 756 6641 765 6675
rect 765 6641 799 6675
rect 799 6641 808 6675
rect 756 6632 808 6641
rect 2320 6709 2329 6743
rect 2329 6709 2363 6743
rect 2363 6709 2372 6743
rect 2320 6700 2372 6709
rect 2964 6700 3016 6752
rect 3056 6632 3108 6684
rect 1400 6564 1452 6616
rect 1584 6607 1636 6616
rect 1584 6573 1593 6607
rect 1593 6573 1627 6607
rect 1627 6573 1636 6607
rect 1584 6564 1636 6573
rect 1676 6564 1728 6616
rect 1952 6564 2004 6616
rect 3332 6564 3384 6616
rect 4528 6777 4537 6811
rect 4537 6777 4571 6811
rect 4571 6777 4580 6811
rect 4528 6768 4580 6777
rect 6276 6768 6328 6820
rect 4988 6743 5040 6752
rect 4988 6709 4997 6743
rect 4997 6709 5031 6743
rect 5031 6709 5040 6743
rect 4988 6700 5040 6709
rect 6368 6743 6420 6752
rect 3976 6632 4028 6684
rect 6368 6709 6377 6743
rect 6377 6709 6411 6743
rect 6411 6709 6420 6743
rect 6368 6700 6420 6709
rect 6460 6700 6512 6752
rect 9680 6811 9732 6820
rect 9680 6777 9689 6811
rect 9689 6777 9723 6811
rect 9723 6777 9732 6811
rect 9680 6768 9732 6777
rect 9496 6700 9548 6752
rect 11704 6836 11756 6888
rect 10140 6811 10192 6820
rect 10140 6777 10149 6811
rect 10149 6777 10183 6811
rect 10183 6777 10192 6811
rect 10140 6768 10192 6777
rect 11244 6768 11296 6820
rect 12072 6811 12124 6820
rect 12072 6777 12081 6811
rect 12081 6777 12115 6811
rect 12115 6777 12124 6811
rect 12072 6768 12124 6777
rect 14096 6836 14148 6888
rect 13728 6768 13780 6820
rect 14188 6811 14240 6820
rect 8484 6675 8536 6684
rect 8484 6641 8493 6675
rect 8493 6641 8527 6675
rect 8527 6641 8536 6675
rect 8484 6632 8536 6641
rect 8668 6675 8720 6684
rect 8668 6641 8677 6675
rect 8677 6641 8711 6675
rect 8711 6641 8720 6675
rect 8668 6632 8720 6641
rect 10876 6700 10928 6752
rect 11428 6632 11480 6684
rect 7196 6564 7248 6616
rect 11520 6564 11572 6616
rect 13912 6743 13964 6752
rect 13912 6709 13921 6743
rect 13921 6709 13955 6743
rect 13955 6709 13964 6743
rect 13912 6700 13964 6709
rect 14188 6777 14197 6811
rect 14197 6777 14231 6811
rect 14231 6777 14240 6811
rect 14188 6768 14240 6777
rect 14280 6743 14332 6752
rect 14280 6709 14289 6743
rect 14289 6709 14323 6743
rect 14323 6709 14332 6743
rect 14280 6700 14332 6709
rect 15016 6700 15068 6752
rect 13636 6632 13688 6684
rect 11704 6607 11756 6616
rect 11704 6573 11713 6607
rect 11713 6573 11747 6607
rect 11747 6573 11756 6607
rect 11704 6564 11756 6573
rect 12900 6564 12952 6616
rect 5242 6462 5294 6514
rect 5306 6462 5358 6514
rect 5370 6462 5422 6514
rect 5434 6462 5486 6514
rect 10514 6462 10566 6514
rect 10578 6462 10630 6514
rect 10642 6462 10694 6514
rect 10706 6462 10758 6514
rect 3792 6403 3844 6412
rect 3792 6369 3801 6403
rect 3801 6369 3835 6403
rect 3835 6369 3844 6403
rect 3792 6360 3844 6369
rect 7012 6360 7064 6412
rect 7748 6360 7800 6412
rect 8668 6360 8720 6412
rect 8852 6360 8904 6412
rect 1952 6292 2004 6344
rect 572 6156 624 6208
rect 940 6156 992 6208
rect 6552 6292 6604 6344
rect 6828 6292 6880 6344
rect 3700 6267 3752 6276
rect 3700 6233 3709 6267
rect 3709 6233 3743 6267
rect 3743 6233 3752 6267
rect 3700 6224 3752 6233
rect 4160 6224 4212 6276
rect 4896 6224 4948 6276
rect 5724 6224 5776 6276
rect 6460 6224 6512 6276
rect 9036 6267 9088 6276
rect 3148 6156 3200 6208
rect 3424 6156 3476 6208
rect 4436 6156 4488 6208
rect 8576 6156 8628 6208
rect 9036 6233 9045 6267
rect 9045 6233 9079 6267
rect 9079 6233 9088 6267
rect 9036 6224 9088 6233
rect 9496 6292 9548 6344
rect 11336 6360 11388 6412
rect 12992 6360 13044 6412
rect 14372 6403 14424 6412
rect 14372 6369 14381 6403
rect 14381 6369 14415 6403
rect 14415 6369 14424 6403
rect 14372 6360 14424 6369
rect 12900 6335 12952 6344
rect 10140 6224 10192 6276
rect 11428 6267 11480 6276
rect 11428 6233 11437 6267
rect 11437 6233 11471 6267
rect 11471 6233 11480 6267
rect 11428 6224 11480 6233
rect 11704 6224 11756 6276
rect 12900 6301 12909 6335
rect 12909 6301 12943 6335
rect 12943 6301 12952 6335
rect 12900 6292 12952 6301
rect 12256 6224 12308 6276
rect 13912 6292 13964 6344
rect 15016 6292 15068 6344
rect 2320 6088 2372 6140
rect 5908 6088 5960 6140
rect 11612 6088 11664 6140
rect 1584 6020 1636 6072
rect 4344 6020 4396 6072
rect 4988 6020 5040 6072
rect 5632 6020 5684 6072
rect 11428 6020 11480 6072
rect 12624 6156 12676 6208
rect 13544 6088 13596 6140
rect 15108 6267 15160 6276
rect 15108 6233 15117 6267
rect 15117 6233 15151 6267
rect 15151 6233 15160 6267
rect 15108 6224 15160 6233
rect 14004 6020 14056 6072
rect 2606 5918 2658 5970
rect 2670 5918 2722 5970
rect 2734 5918 2786 5970
rect 2798 5918 2850 5970
rect 7878 5918 7930 5970
rect 7942 5918 7994 5970
rect 8006 5918 8058 5970
rect 8070 5918 8122 5970
rect 13150 5918 13202 5970
rect 13214 5918 13266 5970
rect 13278 5918 13330 5970
rect 13342 5918 13394 5970
rect 1768 5816 1820 5868
rect 3424 5816 3476 5868
rect 1584 5791 1636 5800
rect 1584 5757 1593 5791
rect 1593 5757 1627 5791
rect 1627 5757 1636 5791
rect 1584 5748 1636 5757
rect 3700 5816 3752 5868
rect 6368 5816 6420 5868
rect 8484 5816 8536 5868
rect 1400 5680 1452 5732
rect 3976 5680 4028 5732
rect 6920 5748 6972 5800
rect 7012 5748 7064 5800
rect 11796 5748 11848 5800
rect 12440 5748 12492 5800
rect 6000 5723 6052 5732
rect 6000 5689 6009 5723
rect 6009 5689 6043 5723
rect 6043 5689 6052 5723
rect 6000 5680 6052 5689
rect 2044 5612 2096 5664
rect 2964 5612 3016 5664
rect 4252 5655 4304 5664
rect 4252 5621 4261 5655
rect 4261 5621 4295 5655
rect 4295 5621 4304 5655
rect 4252 5612 4304 5621
rect 4344 5655 4396 5664
rect 4344 5621 4353 5655
rect 4353 5621 4387 5655
rect 4387 5621 4396 5655
rect 4344 5612 4396 5621
rect 4896 5612 4948 5664
rect 5816 5655 5868 5664
rect 5816 5621 5825 5655
rect 5825 5621 5859 5655
rect 5859 5621 5868 5655
rect 5816 5612 5868 5621
rect 5908 5655 5960 5664
rect 5908 5621 5917 5655
rect 5917 5621 5951 5655
rect 5951 5621 5960 5655
rect 6828 5655 6880 5664
rect 5908 5612 5960 5621
rect 6828 5621 6837 5655
rect 6837 5621 6871 5655
rect 6871 5621 6880 5655
rect 6828 5612 6880 5621
rect 6920 5655 6972 5664
rect 6920 5621 6929 5655
rect 6929 5621 6963 5655
rect 6963 5621 6972 5655
rect 6920 5612 6972 5621
rect 8576 5612 8628 5664
rect 8668 5655 8720 5664
rect 8668 5621 8677 5655
rect 8677 5621 8711 5655
rect 8711 5621 8720 5655
rect 9220 5655 9272 5664
rect 8668 5612 8720 5621
rect 9220 5621 9229 5655
rect 9229 5621 9263 5655
rect 9263 5621 9272 5655
rect 9220 5612 9272 5621
rect 3056 5544 3108 5596
rect 3516 5587 3568 5596
rect 3516 5553 3525 5587
rect 3525 5553 3559 5587
rect 3559 5553 3568 5587
rect 3516 5544 3568 5553
rect 6736 5544 6788 5596
rect 3424 5476 3476 5528
rect 9312 5476 9364 5528
rect 9404 5476 9456 5528
rect 9772 5544 9824 5596
rect 9956 5544 10008 5596
rect 9588 5476 9640 5528
rect 12256 5612 12308 5664
rect 14188 5816 14240 5868
rect 13728 5655 13780 5664
rect 13728 5621 13737 5655
rect 13737 5621 13771 5655
rect 13771 5621 13780 5655
rect 13728 5612 13780 5621
rect 11612 5544 11664 5596
rect 15108 5680 15160 5732
rect 14188 5544 14240 5596
rect 15108 5544 15160 5596
rect 10968 5519 11020 5528
rect 10968 5485 10977 5519
rect 10977 5485 11011 5519
rect 11011 5485 11020 5519
rect 10968 5476 11020 5485
rect 11060 5476 11112 5528
rect 15016 5519 15068 5528
rect 15016 5485 15025 5519
rect 15025 5485 15059 5519
rect 15059 5485 15068 5519
rect 15016 5476 15068 5485
rect 5242 5374 5294 5426
rect 5306 5374 5358 5426
rect 5370 5374 5422 5426
rect 5434 5374 5486 5426
rect 10514 5374 10566 5426
rect 10578 5374 10630 5426
rect 10642 5374 10694 5426
rect 10706 5374 10758 5426
rect 2504 5204 2556 5256
rect 1952 5136 2004 5188
rect 572 5111 624 5120
rect 572 5077 581 5111
rect 581 5077 615 5111
rect 615 5077 624 5111
rect 572 5068 624 5077
rect 5632 5272 5684 5324
rect 6000 5272 6052 5324
rect 4436 5204 4488 5256
rect 3976 5179 4028 5188
rect 3976 5145 3985 5179
rect 3985 5145 4019 5179
rect 4019 5145 4028 5179
rect 3976 5136 4028 5145
rect 4160 5136 4212 5188
rect 3516 5111 3568 5120
rect 3516 5077 3525 5111
rect 3525 5077 3559 5111
rect 3559 5077 3568 5111
rect 3516 5068 3568 5077
rect 5908 5136 5960 5188
rect 6276 5272 6328 5324
rect 9404 5315 9456 5324
rect 9404 5281 9413 5315
rect 9413 5281 9447 5315
rect 9447 5281 9456 5315
rect 9404 5272 9456 5281
rect 11244 5272 11296 5324
rect 14188 5272 14240 5324
rect 14740 5272 14792 5324
rect 6920 5204 6972 5256
rect 6276 5179 6328 5188
rect 6276 5145 6285 5179
rect 6285 5145 6319 5179
rect 6319 5145 6328 5179
rect 6276 5136 6328 5145
rect 6736 5136 6788 5188
rect 8944 5204 8996 5256
rect 8484 5179 8536 5188
rect 8484 5145 8493 5179
rect 8493 5145 8527 5179
rect 8527 5145 8536 5179
rect 8484 5136 8536 5145
rect 4620 5000 4672 5052
rect 6368 5068 6420 5120
rect 6644 5068 6696 5120
rect 7104 5111 7156 5120
rect 7104 5077 7113 5111
rect 7113 5077 7147 5111
rect 7147 5077 7156 5111
rect 7104 5068 7156 5077
rect 7380 5111 7432 5120
rect 7380 5077 7389 5111
rect 7389 5077 7423 5111
rect 7423 5077 7432 5111
rect 7380 5068 7432 5077
rect 9036 5136 9088 5188
rect 10968 5136 11020 5188
rect 11796 5136 11848 5188
rect 9128 5068 9180 5120
rect 9864 5068 9916 5120
rect 12440 5204 12492 5256
rect 13452 5204 13504 5256
rect 8852 5000 8904 5052
rect 6184 4932 6236 4984
rect 8760 4932 8812 4984
rect 9220 4932 9272 4984
rect 12348 5068 12400 5120
rect 12532 5111 12584 5120
rect 12532 5077 12541 5111
rect 12541 5077 12575 5111
rect 12575 5077 12584 5111
rect 12532 5068 12584 5077
rect 14832 5204 14884 5256
rect 15292 5204 15344 5256
rect 14740 5179 14792 5188
rect 14740 5145 14752 5179
rect 14752 5145 14786 5179
rect 14786 5145 14792 5179
rect 14740 5136 14792 5145
rect 10140 5000 10192 5052
rect 12348 4932 12400 4984
rect 2606 4830 2658 4882
rect 2670 4830 2722 4882
rect 2734 4830 2786 4882
rect 2798 4830 2850 4882
rect 7878 4830 7930 4882
rect 7942 4830 7994 4882
rect 8006 4830 8058 4882
rect 8070 4830 8122 4882
rect 13150 4830 13202 4882
rect 13214 4830 13266 4882
rect 13278 4830 13330 4882
rect 13342 4830 13394 4882
rect 756 4703 808 4712
rect 756 4669 765 4703
rect 765 4669 799 4703
rect 799 4669 808 4703
rect 756 4660 808 4669
rect 2044 4592 2096 4644
rect 3516 4728 3568 4780
rect 5540 4728 5592 4780
rect 6276 4728 6328 4780
rect 8484 4728 8536 4780
rect 10324 4728 10376 4780
rect 11060 4728 11112 4780
rect 11244 4771 11296 4780
rect 11244 4737 11253 4771
rect 11253 4737 11287 4771
rect 11287 4737 11296 4771
rect 11244 4728 11296 4737
rect 13544 4728 13596 4780
rect 14648 4728 14700 4780
rect 4436 4592 4488 4644
rect 6000 4592 6052 4644
rect 8392 4592 8444 4644
rect 8760 4635 8812 4644
rect 8760 4601 8769 4635
rect 8769 4601 8803 4635
rect 8803 4601 8812 4635
rect 8760 4592 8812 4601
rect 13636 4660 13688 4712
rect 940 4567 992 4576
rect 940 4533 949 4567
rect 949 4533 983 4567
rect 983 4533 992 4567
rect 940 4524 992 4533
rect 3148 4524 3200 4576
rect 3976 4524 4028 4576
rect 6092 4524 6144 4576
rect 10876 4592 10928 4644
rect 11796 4567 11848 4576
rect 1400 4456 1452 4508
rect 4436 4456 4488 4508
rect 5724 4456 5776 4508
rect 7196 4456 7248 4508
rect 1216 4388 1268 4440
rect 1676 4388 1728 4440
rect 3608 4431 3660 4440
rect 3608 4397 3617 4431
rect 3617 4397 3651 4431
rect 3651 4397 3660 4431
rect 3608 4388 3660 4397
rect 4712 4388 4764 4440
rect 6736 4388 6788 4440
rect 9036 4499 9088 4508
rect 9036 4465 9045 4499
rect 9045 4465 9079 4499
rect 9079 4465 9088 4499
rect 9036 4456 9088 4465
rect 9680 4456 9732 4508
rect 11152 4499 11204 4508
rect 10324 4388 10376 4440
rect 10416 4388 10468 4440
rect 10876 4388 10928 4440
rect 11152 4465 11161 4499
rect 11161 4465 11195 4499
rect 11195 4465 11204 4499
rect 11152 4456 11204 4465
rect 11796 4533 11805 4567
rect 11805 4533 11839 4567
rect 11839 4533 11848 4567
rect 11796 4524 11848 4533
rect 12348 4524 12400 4576
rect 11704 4456 11756 4508
rect 12624 4567 12676 4576
rect 12624 4533 12633 4567
rect 12633 4533 12667 4567
rect 12667 4533 12676 4567
rect 12624 4524 12676 4533
rect 14740 4567 14792 4576
rect 14740 4533 14749 4567
rect 14749 4533 14783 4567
rect 14783 4533 14792 4567
rect 14740 4524 14792 4533
rect 14832 4524 14884 4576
rect 15016 4567 15068 4576
rect 15016 4533 15025 4567
rect 15025 4533 15059 4567
rect 15059 4533 15068 4567
rect 15016 4524 15068 4533
rect 12716 4456 12768 4508
rect 14188 4456 14240 4508
rect 14464 4388 14516 4440
rect 14832 4388 14884 4440
rect 5242 4286 5294 4338
rect 5306 4286 5358 4338
rect 5370 4286 5422 4338
rect 5434 4286 5486 4338
rect 10514 4286 10566 4338
rect 10578 4286 10630 4338
rect 10642 4286 10694 4338
rect 10706 4286 10758 4338
rect 1952 4184 2004 4236
rect 3148 4227 3200 4236
rect 3148 4193 3157 4227
rect 3157 4193 3191 4227
rect 3191 4193 3200 4227
rect 3148 4184 3200 4193
rect 3608 4184 3660 4236
rect 4620 4184 4672 4236
rect 4712 4184 4764 4236
rect 7104 4184 7156 4236
rect 3424 4048 3476 4100
rect 5908 4116 5960 4168
rect 9036 4184 9088 4236
rect 8484 4116 8536 4168
rect 8668 4116 8720 4168
rect 11796 4184 11848 4236
rect 9772 4159 9824 4168
rect 9772 4125 9781 4159
rect 9781 4125 9815 4159
rect 9815 4125 9824 4159
rect 12624 4184 12676 4236
rect 14188 4184 14240 4236
rect 9772 4116 9824 4125
rect 13452 4116 13504 4168
rect 14648 4116 14700 4168
rect 572 3980 624 4032
rect 756 3980 808 4032
rect 1124 4023 1176 4032
rect 1124 3989 1133 4023
rect 1133 3989 1167 4023
rect 1167 3989 1176 4023
rect 1124 3980 1176 3989
rect 2136 3980 2188 4032
rect 3976 3980 4028 4032
rect 4896 4048 4948 4100
rect 6092 4048 6144 4100
rect 6368 4048 6420 4100
rect 6276 3980 6328 4032
rect 9128 4048 9180 4100
rect 9312 4048 9364 4100
rect 9680 4091 9732 4100
rect 9680 4057 9689 4091
rect 9689 4057 9723 4091
rect 9723 4057 9732 4091
rect 9680 4048 9732 4057
rect 10140 4048 10192 4100
rect 8944 3980 8996 4032
rect 10968 3980 11020 4032
rect 11612 4048 11664 4100
rect 12072 4091 12124 4100
rect 12072 4057 12081 4091
rect 12081 4057 12115 4091
rect 12115 4057 12124 4091
rect 12072 4048 12124 4057
rect 12532 4091 12584 4100
rect 12532 4057 12541 4091
rect 12541 4057 12575 4091
rect 12575 4057 12584 4091
rect 12532 4048 12584 4057
rect 12348 3980 12400 4032
rect 14004 3980 14056 4032
rect 15476 3980 15528 4032
rect 7380 3912 7432 3964
rect 11060 3912 11112 3964
rect 3148 3844 3200 3896
rect 5908 3844 5960 3896
rect 6184 3887 6236 3896
rect 6184 3853 6193 3887
rect 6193 3853 6227 3887
rect 6227 3853 6236 3887
rect 6184 3844 6236 3853
rect 10968 3844 11020 3896
rect 12256 3844 12308 3896
rect 2606 3742 2658 3794
rect 2670 3742 2722 3794
rect 2734 3742 2786 3794
rect 2798 3742 2850 3794
rect 7878 3742 7930 3794
rect 7942 3742 7994 3794
rect 8006 3742 8058 3794
rect 8070 3742 8122 3794
rect 13150 3742 13202 3794
rect 13214 3742 13266 3794
rect 13278 3742 13330 3794
rect 13342 3742 13394 3794
rect 848 3683 900 3692
rect 848 3649 857 3683
rect 857 3649 891 3683
rect 891 3649 900 3683
rect 848 3640 900 3649
rect 2044 3640 2096 3692
rect 4160 3640 4212 3692
rect 5080 3640 5132 3692
rect 5908 3640 5960 3692
rect 3148 3504 3200 3556
rect 4068 3572 4120 3624
rect 11336 3640 11388 3692
rect 12072 3640 12124 3692
rect 7840 3572 7892 3624
rect 8944 3572 8996 3624
rect 9312 3572 9364 3624
rect 11244 3572 11296 3624
rect 2228 3436 2280 3488
rect 4896 3504 4948 3556
rect 4988 3504 5040 3556
rect 5816 3504 5868 3556
rect 6276 3504 6328 3556
rect 4252 3436 4304 3488
rect 5632 3436 5684 3488
rect 5724 3436 5776 3488
rect 6644 3436 6696 3488
rect 8392 3504 8444 3556
rect 12440 3572 12492 3624
rect 12624 3572 12676 3624
rect 13820 3615 13872 3624
rect 13820 3581 13829 3615
rect 13829 3581 13863 3615
rect 13863 3581 13872 3615
rect 13820 3572 13872 3581
rect 7196 3479 7248 3488
rect 7196 3445 7205 3479
rect 7205 3445 7239 3479
rect 7239 3445 7248 3479
rect 7196 3436 7248 3445
rect 9312 3436 9364 3488
rect 9864 3479 9916 3488
rect 4344 3368 4396 3420
rect 5264 3368 5316 3420
rect 5908 3368 5960 3420
rect 4252 3300 4304 3352
rect 8484 3368 8536 3420
rect 8668 3411 8720 3420
rect 8668 3377 8677 3411
rect 8677 3377 8711 3411
rect 8711 3377 8720 3411
rect 8668 3368 8720 3377
rect 7748 3300 7800 3352
rect 9128 3368 9180 3420
rect 9864 3445 9873 3479
rect 9873 3445 9907 3479
rect 9907 3445 9916 3479
rect 9864 3436 9916 3445
rect 10416 3479 10468 3488
rect 10416 3445 10425 3479
rect 10425 3445 10459 3479
rect 10459 3445 10468 3479
rect 10416 3436 10468 3445
rect 11060 3479 11112 3488
rect 11060 3445 11069 3479
rect 11069 3445 11103 3479
rect 11103 3445 11112 3479
rect 11060 3436 11112 3445
rect 11612 3436 11664 3488
rect 13636 3504 13688 3556
rect 12532 3479 12584 3488
rect 12532 3445 12541 3479
rect 12541 3445 12575 3479
rect 12575 3445 12584 3479
rect 12532 3436 12584 3445
rect 9956 3368 10008 3420
rect 11428 3368 11480 3420
rect 11796 3368 11848 3420
rect 13728 3368 13780 3420
rect 14188 3411 14240 3420
rect 14188 3377 14197 3411
rect 14197 3377 14231 3411
rect 14231 3377 14240 3411
rect 14188 3368 14240 3377
rect 8944 3300 8996 3352
rect 9588 3300 9640 3352
rect 10140 3300 10192 3352
rect 12532 3300 12584 3352
rect 12716 3300 12768 3352
rect 15016 3436 15068 3488
rect 5242 3198 5294 3250
rect 5306 3198 5358 3250
rect 5370 3198 5422 3250
rect 5434 3198 5486 3250
rect 10514 3198 10566 3250
rect 10578 3198 10630 3250
rect 10642 3198 10694 3250
rect 10706 3198 10758 3250
rect 2964 3096 3016 3148
rect 4252 3139 4304 3148
rect 4252 3105 4261 3139
rect 4261 3105 4295 3139
rect 4295 3105 4304 3139
rect 4252 3096 4304 3105
rect 5816 3139 5868 3148
rect 5816 3105 5825 3139
rect 5825 3105 5859 3139
rect 5859 3105 5868 3139
rect 5816 3096 5868 3105
rect 5908 3096 5960 3148
rect 1216 3071 1268 3080
rect 1216 3037 1225 3071
rect 1225 3037 1259 3071
rect 1259 3037 1268 3071
rect 1216 3028 1268 3037
rect 1952 3028 2004 3080
rect 5632 3028 5684 3080
rect 3148 3003 3200 3012
rect 3148 2969 3157 3003
rect 3157 2969 3191 3003
rect 3191 2969 3200 3003
rect 3148 2960 3200 2969
rect 756 2892 808 2944
rect 1584 2892 1636 2944
rect 4620 2960 4672 3012
rect 6000 3003 6052 3012
rect 6000 2969 6009 3003
rect 6009 2969 6043 3003
rect 6043 2969 6052 3003
rect 6000 2960 6052 2969
rect 6184 3003 6236 3012
rect 6184 2969 6193 3003
rect 6193 2969 6227 3003
rect 6227 2969 6236 3003
rect 6184 2960 6236 2969
rect 6828 2960 6880 3012
rect 8852 3096 8904 3148
rect 9404 3096 9456 3148
rect 9588 3096 9640 3148
rect 11152 3096 11204 3148
rect 11612 3096 11664 3148
rect 12900 3096 12952 3148
rect 14188 3139 14240 3148
rect 14188 3105 14197 3139
rect 14197 3105 14231 3139
rect 14231 3105 14240 3139
rect 14188 3096 14240 3105
rect 7840 3071 7892 3080
rect 7840 3037 7849 3071
rect 7849 3037 7883 3071
rect 7883 3037 7892 3071
rect 7840 3028 7892 3037
rect 8576 3028 8628 3080
rect 8760 3028 8812 3080
rect 9220 3028 9272 3080
rect 10876 3028 10928 3080
rect 12256 3028 12308 3080
rect 13452 3028 13504 3080
rect 15292 3028 15344 3080
rect 11244 3003 11296 3012
rect 6276 2892 6328 2944
rect 6920 2892 6972 2944
rect 11244 2969 11253 3003
rect 11253 2969 11287 3003
rect 11287 2969 11296 3003
rect 11244 2960 11296 2969
rect 11428 3003 11480 3012
rect 11428 2969 11437 3003
rect 11437 2969 11471 3003
rect 11471 2969 11480 3003
rect 11428 2960 11480 2969
rect 8668 2935 8720 2944
rect 8668 2901 8677 2935
rect 8677 2901 8711 2935
rect 8711 2901 8720 2935
rect 8668 2892 8720 2901
rect 9864 2892 9916 2944
rect 10968 2892 11020 2944
rect 11704 2935 11756 2944
rect 11704 2901 11713 2935
rect 11713 2901 11747 2935
rect 11747 2901 11756 2935
rect 11704 2892 11756 2901
rect 6644 2824 6696 2876
rect 2228 2756 2280 2808
rect 5908 2756 5960 2808
rect 9772 2824 9824 2876
rect 12440 2935 12492 2944
rect 12440 2901 12449 2935
rect 12449 2901 12483 2935
rect 12483 2901 12492 2935
rect 12440 2892 12492 2901
rect 15108 2867 15160 2876
rect 15108 2833 15117 2867
rect 15117 2833 15151 2867
rect 15151 2833 15160 2867
rect 15108 2824 15160 2833
rect 9680 2756 9732 2808
rect 10876 2756 10928 2808
rect 11060 2799 11112 2808
rect 11060 2765 11069 2799
rect 11069 2765 11103 2799
rect 11103 2765 11112 2799
rect 11060 2756 11112 2765
rect 11152 2756 11204 2808
rect 11336 2756 11388 2808
rect 2606 2654 2658 2706
rect 2670 2654 2722 2706
rect 2734 2654 2786 2706
rect 2798 2654 2850 2706
rect 7878 2654 7930 2706
rect 7942 2654 7994 2706
rect 8006 2654 8058 2706
rect 8070 2654 8122 2706
rect 13150 2654 13202 2706
rect 13214 2654 13266 2706
rect 13278 2654 13330 2706
rect 13342 2654 13394 2706
rect 1124 2552 1176 2604
rect 4712 2552 4764 2604
rect 5724 2552 5776 2604
rect 9772 2552 9824 2604
rect 9956 2552 10008 2604
rect 1676 2391 1728 2400
rect 1676 2357 1685 2391
rect 1685 2357 1719 2391
rect 1719 2357 1728 2391
rect 1676 2348 1728 2357
rect 2228 2348 2280 2400
rect 848 2323 900 2332
rect 848 2289 857 2323
rect 857 2289 891 2323
rect 891 2289 900 2323
rect 848 2280 900 2289
rect 1216 2280 1268 2332
rect 5632 2416 5684 2468
rect 6736 2416 6788 2468
rect 7196 2416 7248 2468
rect 4160 2391 4212 2400
rect 4160 2357 4169 2391
rect 4169 2357 4203 2391
rect 4203 2357 4212 2391
rect 4160 2348 4212 2357
rect 4712 2391 4764 2400
rect 4712 2357 4721 2391
rect 4721 2357 4755 2391
rect 4755 2357 4764 2391
rect 4712 2348 4764 2357
rect 3792 2255 3844 2264
rect 3792 2221 3801 2255
rect 3801 2221 3835 2255
rect 3835 2221 3844 2255
rect 3792 2212 3844 2221
rect 4528 2280 4580 2332
rect 5264 2280 5316 2332
rect 5724 2280 5776 2332
rect 6276 2280 6328 2332
rect 4436 2212 4488 2264
rect 4896 2212 4948 2264
rect 7288 2348 7340 2400
rect 11060 2416 11112 2468
rect 6920 2280 6972 2332
rect 9496 2280 9548 2332
rect 8484 2212 8536 2264
rect 11244 2348 11296 2400
rect 12532 2552 12584 2604
rect 14004 2595 14056 2604
rect 14004 2561 14013 2595
rect 14013 2561 14047 2595
rect 14047 2561 14056 2595
rect 14004 2552 14056 2561
rect 14924 2552 14976 2604
rect 11704 2416 11756 2468
rect 12624 2391 12676 2400
rect 12624 2357 12633 2391
rect 12633 2357 12667 2391
rect 12667 2357 12676 2391
rect 12624 2348 12676 2357
rect 12900 2348 12952 2400
rect 13728 2391 13780 2400
rect 13728 2357 13737 2391
rect 13737 2357 13771 2391
rect 13771 2357 13780 2391
rect 13728 2348 13780 2357
rect 15016 2348 15068 2400
rect 10968 2280 11020 2332
rect 11704 2323 11756 2332
rect 11704 2289 11739 2323
rect 11739 2289 11756 2323
rect 11704 2280 11756 2289
rect 11244 2255 11296 2264
rect 11244 2221 11253 2255
rect 11253 2221 11287 2255
rect 11287 2221 11296 2255
rect 11244 2212 11296 2221
rect 12624 2212 12676 2264
rect 5242 2110 5294 2162
rect 5306 2110 5358 2162
rect 5370 2110 5422 2162
rect 5434 2110 5486 2162
rect 10514 2110 10566 2162
rect 10578 2110 10630 2162
rect 10642 2110 10694 2162
rect 10706 2110 10758 2162
rect 5080 2008 5132 2060
rect 6644 2051 6696 2060
rect 6644 2017 6653 2051
rect 6653 2017 6687 2051
rect 6687 2017 6696 2051
rect 6644 2008 6696 2017
rect 7288 2008 7340 2060
rect 3516 1940 3568 1992
rect 4160 1940 4212 1992
rect 4712 1983 4764 1992
rect 4712 1949 4721 1983
rect 4721 1949 4755 1983
rect 4755 1949 4764 1983
rect 4712 1940 4764 1949
rect 1216 1915 1268 1924
rect 1216 1881 1225 1915
rect 1225 1881 1259 1915
rect 1259 1881 1268 1915
rect 1216 1872 1268 1881
rect 4620 1915 4672 1924
rect 4620 1881 4629 1915
rect 4629 1881 4663 1915
rect 4663 1881 4672 1915
rect 6276 1940 6328 1992
rect 6828 1940 6880 1992
rect 8944 1940 8996 1992
rect 9680 1940 9732 1992
rect 4620 1872 4672 1881
rect 5908 1872 5960 1924
rect 6736 1872 6788 1924
rect 7748 1915 7800 1924
rect 1676 1847 1728 1856
rect 1308 1736 1360 1788
rect 1676 1813 1685 1847
rect 1685 1813 1719 1847
rect 1719 1813 1728 1847
rect 1676 1804 1728 1813
rect 3976 1804 4028 1856
rect 5540 1804 5592 1856
rect 4344 1736 4396 1788
rect 6184 1804 6236 1856
rect 6000 1736 6052 1788
rect 7748 1881 7757 1915
rect 7757 1881 7791 1915
rect 7791 1881 7800 1915
rect 7748 1872 7800 1881
rect 11612 2008 11664 2060
rect 13544 2008 13596 2060
rect 12624 1983 12676 1992
rect 12624 1949 12633 1983
rect 12633 1949 12667 1983
rect 12667 1949 12676 1983
rect 12624 1940 12676 1949
rect 13912 1940 13964 1992
rect 11152 1872 11204 1924
rect 8300 1736 8352 1788
rect 9956 1804 10008 1856
rect 12348 1847 12400 1856
rect 12348 1813 12357 1847
rect 12357 1813 12391 1847
rect 12391 1813 12400 1847
rect 12348 1804 12400 1813
rect 3332 1668 3384 1720
rect 4528 1668 4580 1720
rect 6828 1668 6880 1720
rect 7012 1668 7064 1720
rect 13728 1736 13780 1788
rect 15108 1779 15160 1788
rect 15108 1745 15117 1779
rect 15117 1745 15151 1779
rect 15151 1745 15160 1779
rect 15108 1736 15160 1745
rect 8484 1668 8536 1720
rect 11152 1711 11204 1720
rect 11152 1677 11161 1711
rect 11161 1677 11195 1711
rect 11195 1677 11204 1711
rect 11152 1668 11204 1677
rect 2606 1566 2658 1618
rect 2670 1566 2722 1618
rect 2734 1566 2786 1618
rect 2798 1566 2850 1618
rect 7878 1566 7930 1618
rect 7942 1566 7994 1618
rect 8006 1566 8058 1618
rect 8070 1566 8122 1618
rect 13150 1566 13202 1618
rect 13214 1566 13266 1618
rect 13278 1566 13330 1618
rect 13342 1566 13394 1618
rect 4712 1507 4764 1516
rect 4712 1473 4721 1507
rect 4721 1473 4755 1507
rect 4755 1473 4764 1507
rect 4712 1464 4764 1473
rect 3332 1396 3384 1448
rect 6460 1464 6512 1516
rect 5540 1328 5592 1380
rect 7012 1371 7064 1380
rect 7012 1337 7021 1371
rect 7021 1337 7055 1371
rect 7055 1337 7064 1371
rect 7012 1328 7064 1337
rect 1032 1260 1084 1312
rect 2320 1303 2372 1312
rect 2320 1269 2329 1303
rect 2329 1269 2363 1303
rect 2363 1269 2372 1303
rect 2320 1260 2372 1269
rect 1952 1192 2004 1244
rect 3976 1260 4028 1312
rect 4344 1260 4396 1312
rect 4528 1303 4580 1312
rect 4528 1269 4537 1303
rect 4537 1269 4571 1303
rect 4571 1269 4580 1303
rect 4528 1260 4580 1269
rect 5632 1260 5684 1312
rect 8300 1260 8352 1312
rect 11704 1464 11756 1516
rect 12440 1396 12492 1448
rect 11244 1328 11296 1380
rect 11428 1303 11480 1312
rect 11428 1269 11437 1303
rect 11437 1269 11471 1303
rect 11471 1269 11480 1303
rect 11428 1260 11480 1269
rect 11888 1303 11940 1312
rect 11888 1269 11897 1303
rect 11897 1269 11931 1303
rect 11931 1269 11940 1303
rect 11888 1260 11940 1269
rect 14832 1260 14884 1312
rect 2964 1192 3016 1244
rect 1124 1124 1176 1176
rect 1308 1124 1360 1176
rect 3516 1192 3568 1244
rect 5724 1192 5776 1244
rect 9588 1192 9640 1244
rect 14556 1192 14608 1244
rect 11244 1167 11296 1176
rect 11244 1133 11253 1167
rect 11253 1133 11287 1167
rect 11287 1133 11296 1167
rect 11244 1124 11296 1133
rect 14924 1124 14976 1176
rect 15200 1124 15252 1176
rect 5242 1022 5294 1074
rect 5306 1022 5358 1074
rect 5370 1022 5422 1074
rect 5434 1022 5486 1074
rect 10514 1022 10566 1074
rect 10578 1022 10630 1074
rect 10642 1022 10694 1074
rect 10706 1022 10758 1074
rect 4528 920 4580 972
rect 6828 963 6880 972
rect 6828 929 6837 963
rect 6837 929 6871 963
rect 6871 929 6880 963
rect 6828 920 6880 929
rect 8668 920 8720 972
rect 1124 895 1176 904
rect 1124 861 1133 895
rect 1133 861 1167 895
rect 1167 861 1176 895
rect 1124 852 1176 861
rect 3792 852 3844 904
rect 5080 852 5132 904
rect 6276 895 6328 904
rect 6276 861 6285 895
rect 6285 861 6319 895
rect 6319 861 6328 895
rect 6276 852 6328 861
rect 2136 827 2188 836
rect 2136 793 2145 827
rect 2145 793 2179 827
rect 2179 793 2188 827
rect 2136 784 2188 793
rect 5724 784 5776 836
rect 1676 716 1728 768
rect 3240 759 3292 768
rect 3240 725 3249 759
rect 3249 725 3283 759
rect 3283 725 3292 759
rect 3240 716 3292 725
rect 3516 716 3568 768
rect 940 691 992 700
rect 940 657 949 691
rect 949 657 983 691
rect 983 657 992 691
rect 940 648 992 657
rect 4620 648 4672 700
rect 4896 580 4948 632
rect 5540 580 5592 632
rect 8392 784 8444 836
rect 9312 827 9364 836
rect 9312 793 9321 827
rect 9321 793 9355 827
rect 9355 793 9364 827
rect 9312 784 9364 793
rect 9036 716 9088 768
rect 9496 827 9548 836
rect 9496 793 9505 827
rect 9505 793 9539 827
rect 9539 793 9548 827
rect 9496 784 9548 793
rect 9864 784 9916 836
rect 12256 852 12308 904
rect 12808 895 12860 904
rect 12808 861 12817 895
rect 12817 861 12851 895
rect 12851 861 12860 895
rect 12808 852 12860 861
rect 14004 852 14056 904
rect 14924 895 14976 904
rect 14924 861 14933 895
rect 14933 861 14967 895
rect 14967 861 14976 895
rect 14924 852 14976 861
rect 8944 648 8996 700
rect 10876 648 10928 700
rect 14372 691 14424 700
rect 14372 657 14381 691
rect 14381 657 14415 691
rect 14415 657 14424 691
rect 14372 648 14424 657
rect 10140 623 10192 632
rect 10140 589 10149 623
rect 10149 589 10183 623
rect 10183 589 10192 623
rect 10140 580 10192 589
rect 12900 623 12952 632
rect 12900 589 12909 623
rect 12909 589 12943 623
rect 12943 589 12952 623
rect 12900 580 12952 589
rect 14924 580 14976 632
rect 2606 478 2658 530
rect 2670 478 2722 530
rect 2734 478 2786 530
rect 2798 478 2850 530
rect 7878 478 7930 530
rect 7942 478 7994 530
rect 8006 478 8058 530
rect 8070 478 8122 530
rect 13150 478 13202 530
rect 13214 478 13266 530
rect 13278 478 13330 530
rect 13342 478 13394 530
rect 2320 376 2372 428
rect 10140 376 10192 428
rect 3240 308 3292 360
rect 4804 308 4856 360
rect 11244 308 11296 360
rect 2136 240 2188 292
rect 11152 240 11204 292
<< metal2 >>
rect 938 13760 994 13960
rect 2870 13760 2926 13960
rect 4894 13760 4950 13960
rect 6918 13760 6974 13960
rect 8942 13760 8998 13960
rect 10874 13760 10930 13960
rect 12898 13760 12954 13960
rect 14922 13760 14978 13960
rect 952 12878 980 13760
rect 2884 12878 2912 13760
rect 3974 13384 4030 13393
rect 3974 13319 4030 13328
rect 3988 12878 4016 13319
rect 4908 12946 4936 13760
rect 5216 13044 5512 13064
rect 5272 13042 5296 13044
rect 5352 13042 5376 13044
rect 5432 13042 5456 13044
rect 5294 12990 5296 13042
rect 5358 12990 5370 13042
rect 5432 12990 5434 13042
rect 5272 12988 5296 12990
rect 5352 12988 5376 12990
rect 5432 12988 5456 12990
rect 5216 12968 5512 12988
rect 4896 12940 4948 12946
rect 4896 12882 4948 12888
rect 6932 12878 6960 13760
rect 8956 12946 8984 13760
rect 10488 13044 10784 13064
rect 10544 13042 10568 13044
rect 10624 13042 10648 13044
rect 10704 13042 10728 13044
rect 10566 12990 10568 13042
rect 10630 12990 10642 13042
rect 10704 12990 10706 13042
rect 10544 12988 10568 12990
rect 10624 12988 10648 12990
rect 10704 12988 10728 12990
rect 10488 12968 10784 12988
rect 8944 12940 8996 12946
rect 8944 12882 8996 12888
rect 10888 12878 10916 13760
rect 12912 12946 12940 13760
rect 14370 13384 14426 13393
rect 14370 13319 14426 13328
rect 12900 12940 12952 12946
rect 12900 12882 12952 12888
rect 14384 12878 14412 13319
rect 14936 12946 14964 13760
rect 14924 12940 14976 12946
rect 14924 12882 14976 12888
rect 940 12872 992 12878
rect 940 12814 992 12820
rect 2872 12872 2924 12878
rect 2872 12814 2924 12820
rect 3976 12872 4028 12878
rect 3976 12814 4028 12820
rect 6920 12872 6972 12878
rect 6920 12814 6972 12820
rect 10876 12872 10928 12878
rect 10876 12814 10928 12820
rect 14372 12872 14424 12878
rect 14372 12814 14424 12820
rect 1124 12804 1176 12810
rect 1124 12746 1176 12752
rect 1860 12804 1912 12810
rect 1860 12746 1912 12752
rect 3424 12804 3476 12810
rect 3424 12746 3476 12752
rect 3516 12804 3568 12810
rect 3516 12746 3568 12752
rect 4896 12804 4948 12810
rect 4896 12746 4948 12752
rect 7196 12804 7248 12810
rect 7196 12746 7248 12752
rect 8760 12804 8812 12810
rect 8760 12746 8812 12752
rect 8944 12804 8996 12810
rect 8944 12746 8996 12752
rect 9128 12804 9180 12810
rect 9128 12746 9180 12752
rect 11428 12804 11480 12810
rect 11428 12746 11480 12752
rect 12808 12804 12860 12810
rect 12808 12746 12860 12752
rect 14188 12804 14240 12810
rect 14188 12746 14240 12752
rect 14832 12804 14884 12810
rect 14832 12746 14884 12752
rect 940 12396 992 12402
rect 940 12338 992 12344
rect 572 12192 624 12198
rect 572 12134 624 12140
rect 584 11722 612 12134
rect 848 12124 900 12130
rect 848 12066 900 12072
rect 572 11716 624 11722
rect 572 11658 624 11664
rect 584 10634 612 11658
rect 756 11580 808 11586
rect 756 11522 808 11528
rect 768 11353 796 11522
rect 754 11344 810 11353
rect 860 11314 888 12066
rect 952 11790 980 12338
rect 940 11784 992 11790
rect 940 11726 992 11732
rect 754 11279 810 11288
rect 848 11308 900 11314
rect 848 11250 900 11256
rect 756 11036 808 11042
rect 756 10978 808 10984
rect 572 10628 624 10634
rect 572 10570 624 10576
rect 584 9546 612 10570
rect 768 10401 796 10978
rect 940 10424 992 10430
rect 754 10392 810 10401
rect 940 10366 992 10372
rect 754 10327 810 10336
rect 952 9614 980 10366
rect 940 9608 992 9614
rect 940 9550 992 9556
rect 572 9540 624 9546
rect 572 9482 624 9488
rect 756 9472 808 9478
rect 754 9440 756 9449
rect 808 9440 810 9449
rect 754 9375 810 9384
rect 756 8860 808 8866
rect 756 8802 808 8808
rect 664 8588 716 8594
rect 664 8530 716 8536
rect 676 7846 704 8530
rect 768 8361 796 8802
rect 754 8352 810 8361
rect 754 8287 810 8296
rect 1136 7982 1164 12746
rect 1768 12600 1820 12606
rect 1768 12542 1820 12548
rect 1780 12441 1808 12542
rect 1766 12432 1822 12441
rect 1766 12367 1822 12376
rect 1872 11858 1900 12746
rect 2580 12500 2876 12520
rect 2636 12498 2660 12500
rect 2716 12498 2740 12500
rect 2796 12498 2820 12500
rect 2658 12446 2660 12498
rect 2722 12446 2734 12498
rect 2796 12446 2798 12498
rect 2636 12444 2660 12446
rect 2716 12444 2740 12446
rect 2796 12444 2820 12446
rect 2580 12424 2876 12444
rect 3436 12394 3464 12746
rect 3344 12366 3464 12394
rect 2504 12124 2556 12130
rect 2504 12066 2556 12072
rect 3240 12124 3292 12130
rect 3240 12066 3292 12072
rect 1860 11852 1912 11858
rect 1860 11794 1912 11800
rect 2516 11790 2544 12066
rect 1308 11784 1360 11790
rect 1308 11726 1360 11732
rect 2504 11784 2556 11790
rect 2504 11726 2556 11732
rect 1216 10560 1268 10566
rect 1216 10502 1268 10508
rect 1228 10226 1256 10502
rect 1320 10226 1348 11726
rect 1860 11104 1912 11110
rect 1860 11046 1912 11052
rect 1492 10696 1544 10702
rect 1492 10638 1544 10644
rect 1216 10220 1268 10226
rect 1216 10162 1268 10168
rect 1308 10220 1360 10226
rect 1308 10162 1360 10168
rect 1400 9880 1452 9886
rect 1400 9822 1452 9828
rect 1308 9540 1360 9546
rect 1308 9482 1360 9488
rect 1320 9002 1348 9482
rect 1308 8996 1360 9002
rect 1308 8938 1360 8944
rect 1124 7976 1176 7982
rect 1124 7918 1176 7924
rect 664 7840 716 7846
rect 664 7782 716 7788
rect 480 7772 532 7778
rect 480 7714 532 7720
rect 492 7409 520 7714
rect 572 7704 624 7710
rect 572 7646 624 7652
rect 478 7400 534 7409
rect 478 7335 534 7344
rect 584 7166 612 7646
rect 572 7160 624 7166
rect 572 7102 624 7108
rect 664 7160 716 7166
rect 664 7102 716 7108
rect 584 6758 612 7102
rect 572 6752 624 6758
rect 572 6694 624 6700
rect 676 6298 704 7102
rect 1136 6874 1164 7918
rect 1044 6846 1164 6874
rect 1412 6874 1440 9822
rect 1504 9682 1532 10638
rect 1872 10226 1900 11046
rect 2516 10770 2544 11726
rect 2580 11412 2876 11432
rect 2636 11410 2660 11412
rect 2716 11410 2740 11412
rect 2796 11410 2820 11412
rect 2658 11358 2660 11410
rect 2722 11358 2734 11410
rect 2796 11358 2798 11410
rect 2636 11356 2660 11358
rect 2716 11356 2740 11358
rect 2796 11356 2820 11358
rect 2580 11336 2876 11356
rect 3252 11110 3280 12066
rect 3240 11104 3292 11110
rect 3240 11046 3292 11052
rect 2504 10764 2556 10770
rect 2504 10706 2556 10712
rect 3148 10424 3200 10430
rect 3148 10366 3200 10372
rect 2580 10324 2876 10344
rect 2636 10322 2660 10324
rect 2716 10322 2740 10324
rect 2796 10322 2820 10324
rect 2658 10270 2660 10322
rect 2722 10270 2734 10322
rect 2796 10270 2798 10322
rect 2636 10268 2660 10270
rect 2716 10268 2740 10270
rect 2796 10268 2820 10270
rect 2580 10248 2876 10268
rect 1860 10220 1912 10226
rect 1860 10162 1912 10168
rect 1872 9954 1900 10162
rect 2136 10152 2188 10158
rect 2136 10094 2188 10100
rect 2148 9954 2176 10094
rect 3160 10090 3188 10366
rect 3148 10084 3200 10090
rect 3148 10026 3200 10032
rect 1860 9948 1912 9954
rect 1860 9890 1912 9896
rect 2136 9948 2188 9954
rect 2136 9890 2188 9896
rect 2596 9880 2648 9886
rect 2596 9822 2648 9828
rect 2608 9682 2636 9822
rect 1492 9676 1544 9682
rect 1492 9618 1544 9624
rect 2596 9676 2648 9682
rect 2596 9618 2648 9624
rect 1504 8526 1532 9618
rect 1768 9472 1820 9478
rect 1768 9414 1820 9420
rect 3240 9472 3292 9478
rect 3240 9414 3292 9420
rect 1492 8520 1544 8526
rect 1492 8462 1544 8468
rect 1504 7438 1532 8462
rect 1492 7432 1544 7438
rect 1492 7374 1544 7380
rect 1504 7250 1532 7374
rect 1504 7222 1716 7250
rect 1412 6846 1624 6874
rect 756 6684 808 6690
rect 756 6626 808 6632
rect 768 6457 796 6626
rect 754 6448 810 6457
rect 754 6383 810 6392
rect 584 6270 704 6298
rect 584 6214 612 6270
rect 572 6208 624 6214
rect 572 6150 624 6156
rect 940 6208 992 6214
rect 940 6150 992 6156
rect 584 5126 612 6150
rect 754 5360 810 5369
rect 754 5295 810 5304
rect 572 5120 624 5126
rect 572 5062 624 5068
rect 584 4038 612 5062
rect 768 4718 796 5295
rect 756 4712 808 4718
rect 756 4654 808 4660
rect 952 4582 980 6150
rect 940 4576 992 4582
rect 940 4518 992 4524
rect 846 4408 902 4417
rect 846 4343 902 4352
rect 572 4032 624 4038
rect 572 3974 624 3980
rect 756 4032 808 4038
rect 756 3974 808 3980
rect 768 2950 796 3974
rect 860 3698 888 4343
rect 848 3692 900 3698
rect 848 3634 900 3640
rect 756 2944 808 2950
rect 756 2886 808 2892
rect 846 2368 902 2377
rect 846 2303 848 2312
rect 900 2303 902 2312
rect 848 2274 900 2280
rect 1044 1318 1072 6846
rect 1596 6622 1624 6846
rect 1688 6622 1716 7222
rect 1400 6616 1452 6622
rect 1400 6558 1452 6564
rect 1584 6616 1636 6622
rect 1584 6558 1636 6564
rect 1676 6616 1728 6622
rect 1676 6558 1728 6564
rect 1412 5738 1440 6558
rect 1584 6072 1636 6078
rect 1584 6014 1636 6020
rect 1596 5806 1624 6014
rect 1780 5874 1808 9414
rect 2580 9236 2876 9256
rect 2636 9234 2660 9236
rect 2716 9234 2740 9236
rect 2796 9234 2820 9236
rect 2658 9182 2660 9234
rect 2722 9182 2734 9234
rect 2796 9182 2798 9234
rect 2636 9180 2660 9182
rect 2716 9180 2740 9182
rect 2796 9180 2820 9182
rect 2580 9160 2876 9180
rect 2044 9064 2096 9070
rect 2044 9006 2096 9012
rect 1860 8860 1912 8866
rect 1860 8802 1912 8808
rect 1872 8526 1900 8802
rect 1860 8520 1912 8526
rect 1860 8462 1912 8468
rect 1952 6616 2004 6622
rect 1952 6558 2004 6564
rect 1964 6350 1992 6558
rect 1952 6344 2004 6350
rect 1952 6286 2004 6292
rect 1768 5868 1820 5874
rect 1768 5810 1820 5816
rect 1584 5800 1636 5806
rect 1584 5742 1636 5748
rect 1400 5732 1452 5738
rect 1400 5674 1452 5680
rect 1412 4514 1440 5674
rect 1964 5194 1992 6286
rect 2056 5670 2084 9006
rect 2504 8996 2556 9002
rect 2504 8938 2556 8944
rect 2516 8458 2544 8938
rect 3252 8934 3280 9414
rect 2964 8928 3016 8934
rect 2964 8870 3016 8876
rect 3240 8928 3292 8934
rect 3240 8870 3292 8876
rect 2504 8452 2556 8458
rect 2504 8394 2556 8400
rect 2580 8148 2876 8168
rect 2636 8146 2660 8148
rect 2716 8146 2740 8148
rect 2796 8146 2820 8148
rect 2658 8094 2660 8146
rect 2722 8094 2734 8146
rect 2796 8094 2798 8146
rect 2636 8092 2660 8094
rect 2716 8092 2740 8094
rect 2796 8092 2820 8094
rect 2580 8072 2876 8092
rect 2976 7778 3004 8870
rect 3344 8746 3372 12366
rect 3528 12130 3556 12746
rect 4908 12394 4936 12746
rect 4816 12366 4936 12394
rect 4344 12192 4396 12198
rect 4344 12134 4396 12140
rect 4528 12192 4580 12198
rect 4528 12134 4580 12140
rect 3516 12124 3568 12130
rect 3516 12066 3568 12072
rect 3700 12124 3752 12130
rect 3700 12066 3752 12072
rect 3608 11512 3660 11518
rect 3608 11454 3660 11460
rect 3620 11314 3648 11454
rect 3608 11308 3660 11314
rect 3608 11250 3660 11256
rect 3424 11240 3476 11246
rect 3424 11182 3476 11188
rect 3436 10022 3464 11182
rect 3712 11178 3740 12066
rect 4160 12056 4212 12062
rect 4160 11998 4212 12004
rect 3976 11852 4028 11858
rect 3976 11794 4028 11800
rect 3700 11172 3752 11178
rect 3700 11114 3752 11120
rect 3516 11104 3568 11110
rect 3516 11046 3568 11052
rect 3528 10634 3556 11046
rect 3712 11042 3740 11114
rect 3988 11110 4016 11794
rect 3976 11104 4028 11110
rect 4068 11104 4120 11110
rect 3976 11046 4028 11052
rect 4066 11072 4068 11081
rect 4120 11072 4122 11081
rect 3700 11036 3752 11042
rect 4066 11007 4122 11016
rect 3700 10978 3752 10984
rect 3516 10628 3568 10634
rect 3516 10570 3568 10576
rect 3528 10158 3556 10570
rect 3516 10152 3568 10158
rect 3516 10094 3568 10100
rect 3424 10016 3476 10022
rect 3424 9958 3476 9964
rect 3516 9948 3568 9954
rect 3516 9890 3568 9896
rect 3528 9070 3556 9890
rect 3516 9064 3568 9070
rect 3516 9006 3568 9012
rect 3528 8934 3556 9006
rect 3516 8928 3568 8934
rect 3516 8870 3568 8876
rect 3252 8718 3372 8746
rect 3252 8322 3280 8718
rect 4172 8390 4200 11998
rect 4252 10628 4304 10634
rect 4252 10570 4304 10576
rect 4264 8934 4292 10570
rect 4356 9138 4384 12134
rect 4436 11104 4488 11110
rect 4436 11046 4488 11052
rect 4448 10673 4476 11046
rect 4434 10664 4490 10673
rect 4434 10599 4490 10608
rect 4540 10090 4568 12134
rect 4816 12130 4844 12366
rect 6460 12260 6512 12266
rect 6460 12202 6512 12208
rect 4804 12124 4856 12130
rect 4804 12066 4856 12072
rect 4712 12056 4764 12062
rect 4712 11998 4764 12004
rect 4724 11722 4752 11998
rect 4712 11716 4764 11722
rect 4712 11658 4764 11664
rect 4724 11081 4752 11658
rect 4710 11072 4766 11081
rect 4710 11007 4766 11016
rect 4712 10424 4764 10430
rect 4712 10366 4764 10372
rect 4724 10226 4752 10366
rect 4712 10220 4764 10226
rect 4712 10162 4764 10168
rect 4528 10084 4580 10090
rect 4528 10026 4580 10032
rect 4436 9880 4488 9886
rect 4436 9822 4488 9828
rect 4448 9546 4476 9822
rect 4436 9540 4488 9546
rect 4436 9482 4488 9488
rect 4448 9449 4476 9482
rect 4434 9440 4490 9449
rect 4434 9375 4490 9384
rect 4344 9132 4396 9138
rect 4344 9074 4396 9080
rect 4448 8934 4476 9375
rect 4540 9342 4568 10026
rect 4712 9608 4764 9614
rect 4712 9550 4764 9556
rect 4528 9336 4580 9342
rect 4528 9278 4580 9284
rect 4252 8928 4304 8934
rect 4252 8870 4304 8876
rect 4436 8928 4488 8934
rect 4436 8870 4488 8876
rect 4620 8928 4672 8934
rect 4724 8916 4752 9550
rect 4672 8888 4752 8916
rect 4620 8870 4672 8876
rect 4264 8440 4292 8870
rect 4620 8792 4672 8798
rect 4620 8734 4672 8740
rect 4632 8526 4660 8734
rect 4620 8520 4672 8526
rect 4620 8462 4672 8468
rect 4724 8458 4752 8888
rect 4344 8452 4396 8458
rect 4264 8412 4344 8440
rect 4344 8394 4396 8400
rect 4712 8452 4764 8458
rect 4712 8394 4764 8400
rect 4160 8384 4212 8390
rect 4160 8326 4212 8332
rect 3240 8316 3292 8322
rect 3240 8258 3292 8264
rect 3332 8316 3384 8322
rect 3332 8258 3384 8264
rect 2964 7772 3016 7778
rect 2964 7714 3016 7720
rect 3148 7772 3200 7778
rect 3148 7714 3200 7720
rect 3160 7506 3188 7714
rect 3148 7500 3200 7506
rect 3148 7442 3200 7448
rect 2504 7364 2556 7370
rect 2504 7306 2556 7312
rect 2320 6752 2372 6758
rect 2320 6694 2372 6700
rect 2332 6146 2360 6694
rect 2320 6140 2372 6146
rect 2320 6082 2372 6088
rect 2044 5664 2096 5670
rect 2044 5606 2096 5612
rect 2516 5262 2544 7306
rect 3056 7160 3108 7166
rect 3056 7102 3108 7108
rect 2580 7060 2876 7080
rect 2636 7058 2660 7060
rect 2716 7058 2740 7060
rect 2796 7058 2820 7060
rect 2658 7006 2660 7058
rect 2722 7006 2734 7058
rect 2796 7006 2798 7058
rect 2636 7004 2660 7006
rect 2716 7004 2740 7006
rect 2796 7004 2820 7006
rect 2580 6984 2876 7004
rect 2964 6752 3016 6758
rect 2964 6694 3016 6700
rect 2580 5972 2876 5992
rect 2636 5970 2660 5972
rect 2716 5970 2740 5972
rect 2796 5970 2820 5972
rect 2658 5918 2660 5970
rect 2722 5918 2734 5970
rect 2796 5918 2798 5970
rect 2636 5916 2660 5918
rect 2716 5916 2740 5918
rect 2796 5916 2820 5918
rect 2580 5896 2876 5916
rect 2976 5670 3004 6694
rect 3068 6690 3096 7102
rect 3148 6956 3200 6962
rect 3148 6898 3200 6904
rect 3056 6684 3108 6690
rect 3056 6626 3108 6632
rect 2964 5664 3016 5670
rect 2964 5606 3016 5612
rect 2504 5256 2556 5262
rect 2504 5198 2556 5204
rect 1952 5188 2004 5194
rect 1952 5130 2004 5136
rect 1400 4508 1452 4514
rect 1400 4450 1452 4456
rect 1216 4440 1268 4446
rect 1216 4382 1268 4388
rect 1676 4440 1728 4446
rect 1676 4382 1728 4388
rect 1124 4032 1176 4038
rect 1124 3974 1176 3980
rect 1136 2610 1164 3974
rect 1228 3086 1256 4382
rect 1216 3080 1268 3086
rect 1216 3022 1268 3028
rect 1584 2944 1636 2950
rect 1584 2886 1636 2892
rect 1124 2604 1176 2610
rect 1124 2546 1176 2552
rect 1216 2332 1268 2338
rect 1216 2274 1268 2280
rect 1228 1930 1256 2274
rect 1596 2218 1624 2886
rect 1688 2406 1716 4382
rect 1964 4242 1992 5130
rect 2580 4884 2876 4904
rect 2636 4882 2660 4884
rect 2716 4882 2740 4884
rect 2796 4882 2820 4884
rect 2658 4830 2660 4882
rect 2722 4830 2734 4882
rect 2796 4830 2798 4882
rect 2636 4828 2660 4830
rect 2716 4828 2740 4830
rect 2796 4828 2820 4830
rect 2580 4808 2876 4828
rect 2044 4644 2096 4650
rect 2044 4586 2096 4592
rect 1952 4236 2004 4242
rect 1952 4178 2004 4184
rect 1964 3086 1992 4178
rect 2056 3986 2084 4586
rect 2136 4032 2188 4038
rect 2056 3980 2136 3986
rect 2056 3974 2188 3980
rect 2056 3958 2176 3974
rect 2056 3698 2084 3958
rect 2580 3796 2876 3816
rect 2636 3794 2660 3796
rect 2716 3794 2740 3796
rect 2796 3794 2820 3796
rect 2658 3742 2660 3794
rect 2722 3742 2734 3794
rect 2796 3742 2798 3794
rect 2636 3740 2660 3742
rect 2716 3740 2740 3742
rect 2796 3740 2820 3742
rect 2580 3720 2876 3740
rect 2044 3692 2096 3698
rect 2044 3634 2096 3640
rect 2228 3488 2280 3494
rect 2228 3430 2280 3436
rect 1952 3080 2004 3086
rect 1952 3022 2004 3028
rect 1676 2400 1728 2406
rect 1676 2342 1728 2348
rect 1596 2190 1716 2218
rect 1216 1924 1268 1930
rect 1216 1866 1268 1872
rect 1688 1862 1716 2190
rect 1676 1856 1728 1862
rect 1676 1798 1728 1804
rect 1308 1788 1360 1794
rect 1308 1730 1360 1736
rect 1032 1312 1084 1318
rect 1032 1254 1084 1260
rect 1320 1182 1348 1730
rect 1124 1176 1176 1182
rect 1124 1118 1176 1124
rect 1308 1176 1360 1182
rect 1308 1118 1360 1124
rect 1136 910 1164 1118
rect 1124 904 1176 910
rect 1124 846 1176 852
rect 1688 774 1716 1798
rect 1964 1250 1992 3022
rect 2240 2814 2268 3430
rect 2976 3154 3004 5606
rect 3068 5602 3096 6626
rect 3160 6214 3188 6898
rect 3148 6208 3200 6214
rect 3148 6150 3200 6156
rect 3056 5596 3108 5602
rect 3056 5538 3108 5544
rect 3148 4576 3200 4582
rect 3148 4518 3200 4524
rect 3160 4242 3188 4518
rect 3148 4236 3200 4242
rect 3148 4178 3200 4184
rect 3148 3896 3200 3902
rect 3148 3838 3200 3844
rect 3160 3562 3188 3838
rect 3148 3556 3200 3562
rect 3148 3498 3200 3504
rect 2964 3148 3016 3154
rect 2964 3090 3016 3096
rect 3160 3018 3188 3498
rect 3148 3012 3200 3018
rect 3148 2954 3200 2960
rect 2228 2808 2280 2814
rect 2228 2750 2280 2756
rect 2240 2406 2268 2750
rect 3252 2734 3280 8258
rect 3344 7710 3372 8258
rect 4160 8044 4212 8050
rect 4160 7986 4212 7992
rect 3424 7840 3476 7846
rect 3424 7782 3476 7788
rect 4068 7840 4120 7846
rect 4068 7782 4120 7788
rect 3332 7704 3384 7710
rect 3332 7646 3384 7652
rect 3436 6962 3464 7782
rect 3792 7704 3844 7710
rect 3792 7646 3844 7652
rect 3516 7364 3568 7370
rect 3516 7306 3568 7312
rect 3424 6956 3476 6962
rect 3424 6898 3476 6904
rect 3332 6616 3384 6622
rect 3528 6570 3556 7306
rect 3804 7234 3832 7646
rect 3976 7500 4028 7506
rect 3976 7442 4028 7448
rect 3792 7228 3844 7234
rect 3792 7170 3844 7176
rect 3384 6564 3556 6570
rect 3332 6558 3556 6564
rect 3344 6542 3556 6558
rect 3424 6208 3476 6214
rect 3424 6150 3476 6156
rect 3436 5874 3464 6150
rect 3424 5868 3476 5874
rect 3424 5810 3476 5816
rect 3528 5602 3556 6542
rect 3804 6418 3832 7170
rect 3988 6690 4016 7442
rect 4080 6962 4108 7782
rect 4068 6956 4120 6962
rect 4068 6898 4120 6904
rect 4172 6894 4200 7986
rect 4724 7778 4752 8394
rect 4712 7772 4764 7778
rect 4712 7714 4764 7720
rect 4160 6888 4212 6894
rect 4160 6830 4212 6836
rect 4436 6888 4488 6894
rect 4436 6830 4488 6836
rect 4526 6856 4582 6865
rect 3976 6684 4028 6690
rect 3976 6626 4028 6632
rect 3792 6412 3844 6418
rect 3792 6354 3844 6360
rect 3700 6276 3752 6282
rect 3700 6218 3752 6224
rect 3712 5874 3740 6218
rect 3700 5868 3752 5874
rect 3700 5810 3752 5816
rect 3988 5738 4016 6626
rect 4160 6276 4212 6282
rect 4160 6218 4212 6224
rect 3976 5732 4028 5738
rect 3976 5674 4028 5680
rect 3516 5596 3568 5602
rect 3516 5538 3568 5544
rect 3424 5528 3476 5534
rect 3424 5470 3476 5476
rect 3436 4106 3464 5470
rect 3988 5194 4016 5674
rect 4172 5194 4200 6218
rect 4448 6214 4476 6830
rect 4526 6791 4528 6800
rect 4580 6791 4582 6800
rect 4528 6762 4580 6768
rect 4436 6208 4488 6214
rect 4436 6150 4488 6156
rect 4344 6072 4396 6078
rect 4344 6014 4396 6020
rect 4356 5670 4384 6014
rect 4252 5664 4304 5670
rect 4252 5606 4304 5612
rect 4344 5664 4396 5670
rect 4344 5606 4396 5612
rect 3976 5188 4028 5194
rect 3976 5130 4028 5136
rect 4160 5188 4212 5194
rect 4160 5130 4212 5136
rect 3516 5120 3568 5126
rect 3516 5062 3568 5068
rect 3528 4786 3556 5062
rect 3516 4780 3568 4786
rect 3516 4722 3568 4728
rect 3988 4582 4016 5130
rect 3976 4576 4028 4582
rect 3976 4518 4028 4524
rect 3608 4440 3660 4446
rect 3608 4382 3660 4388
rect 3620 4242 3648 4382
rect 3608 4236 3660 4242
rect 3608 4178 3660 4184
rect 3424 4100 3476 4106
rect 3424 4042 3476 4048
rect 3988 4038 4016 4518
rect 3976 4032 4028 4038
rect 3976 3974 4028 3980
rect 4172 3698 4200 5130
rect 4160 3692 4212 3698
rect 4160 3634 4212 3640
rect 4068 3624 4120 3630
rect 4068 3566 4120 3572
rect 4080 3465 4108 3566
rect 4264 3494 4292 5606
rect 4252 3488 4304 3494
rect 4066 3456 4122 3465
rect 4252 3430 4304 3436
rect 4356 3426 4384 5606
rect 4448 5262 4476 6150
rect 4436 5256 4488 5262
rect 4436 5198 4488 5204
rect 4448 4650 4476 5198
rect 4620 5052 4672 5058
rect 4620 4994 4672 5000
rect 4436 4644 4488 4650
rect 4436 4586 4488 4592
rect 4436 4508 4488 4514
rect 4436 4450 4488 4456
rect 4066 3391 4122 3400
rect 4344 3420 4396 3426
rect 4344 3362 4396 3368
rect 4252 3352 4304 3358
rect 4252 3294 4304 3300
rect 4264 3154 4292 3294
rect 4252 3148 4304 3154
rect 4252 3090 4304 3096
rect 2580 2708 2876 2728
rect 2636 2706 2660 2708
rect 2716 2706 2740 2708
rect 2796 2706 2820 2708
rect 3252 2706 3372 2734
rect 2658 2654 2660 2706
rect 2722 2654 2734 2706
rect 2796 2654 2798 2706
rect 2636 2652 2660 2654
rect 2716 2652 2740 2654
rect 2796 2652 2820 2654
rect 2580 2632 2876 2652
rect 2228 2400 2280 2406
rect 2228 2342 2280 2348
rect 3344 1726 3372 2706
rect 4160 2400 4212 2406
rect 4160 2342 4212 2348
rect 3792 2264 3844 2270
rect 3792 2206 3844 2212
rect 3516 1992 3568 1998
rect 3516 1934 3568 1940
rect 3332 1720 3384 1726
rect 3332 1662 3384 1668
rect 2580 1620 2876 1640
rect 2636 1618 2660 1620
rect 2716 1618 2740 1620
rect 2796 1618 2820 1620
rect 2658 1566 2660 1618
rect 2722 1566 2734 1618
rect 2796 1566 2798 1618
rect 2636 1564 2660 1566
rect 2716 1564 2740 1566
rect 2796 1564 2820 1566
rect 2580 1544 2876 1564
rect 3332 1448 3384 1454
rect 3330 1416 3332 1425
rect 3384 1416 3386 1425
rect 3330 1351 3386 1360
rect 2320 1312 2372 1318
rect 2320 1254 2372 1260
rect 1952 1244 2004 1250
rect 1952 1186 2004 1192
rect 2136 836 2188 842
rect 2136 778 2188 784
rect 1676 768 1728 774
rect 1676 710 1728 716
rect 940 700 992 706
rect 940 642 992 648
rect 952 160 980 642
rect 2148 298 2176 778
rect 2332 434 2360 1254
rect 3528 1250 3556 1934
rect 2964 1244 3016 1250
rect 2964 1186 3016 1192
rect 3516 1244 3568 1250
rect 3516 1186 3568 1192
rect 2580 532 2876 552
rect 2636 530 2660 532
rect 2716 530 2740 532
rect 2796 530 2820 532
rect 2658 478 2660 530
rect 2722 478 2734 530
rect 2796 478 2798 530
rect 2636 476 2660 478
rect 2716 476 2740 478
rect 2796 476 2820 478
rect 2580 456 2876 476
rect 2320 428 2372 434
rect 2320 370 2372 376
rect 2976 314 3004 1186
rect 3804 910 3832 2206
rect 4172 1998 4200 2342
rect 4448 2270 4476 4450
rect 4632 4242 4660 4994
rect 4712 4440 4764 4446
rect 4712 4382 4764 4388
rect 4724 4242 4752 4382
rect 4620 4236 4672 4242
rect 4620 4178 4672 4184
rect 4712 4236 4764 4242
rect 4712 4178 4764 4184
rect 4620 3012 4672 3018
rect 4620 2954 4672 2960
rect 4528 2332 4580 2338
rect 4528 2274 4580 2280
rect 4436 2264 4488 2270
rect 4436 2206 4488 2212
rect 4160 1992 4212 1998
rect 4160 1934 4212 1940
rect 3976 1856 4028 1862
rect 3976 1798 4028 1804
rect 3988 1318 4016 1798
rect 4344 1788 4396 1794
rect 4344 1730 4396 1736
rect 4356 1318 4384 1730
rect 4540 1726 4568 2274
rect 4632 1930 4660 2954
rect 4724 2610 4752 4178
rect 4816 2734 4844 12066
rect 5540 12056 5592 12062
rect 5540 11998 5592 12004
rect 5216 11956 5512 11976
rect 5272 11954 5296 11956
rect 5352 11954 5376 11956
rect 5432 11954 5456 11956
rect 5294 11902 5296 11954
rect 5358 11902 5370 11954
rect 5432 11902 5434 11954
rect 5272 11900 5296 11902
rect 5352 11900 5376 11902
rect 5432 11900 5456 11902
rect 5216 11880 5512 11900
rect 5552 11042 5580 11998
rect 6472 11790 6500 12202
rect 7208 12198 7236 12746
rect 7748 12736 7800 12742
rect 7748 12678 7800 12684
rect 7196 12192 7248 12198
rect 7196 12134 7248 12140
rect 6920 12124 6972 12130
rect 6920 12066 6972 12072
rect 6460 11784 6512 11790
rect 6460 11726 6512 11732
rect 6184 11172 6236 11178
rect 6236 11132 6316 11160
rect 6184 11114 6236 11120
rect 6288 11042 6316 11132
rect 6472 11110 6500 11726
rect 6932 11314 6960 12066
rect 7208 11858 7236 12134
rect 7288 12056 7340 12062
rect 7288 11998 7340 12004
rect 7196 11852 7248 11858
rect 7196 11794 7248 11800
rect 6920 11308 6972 11314
rect 6920 11250 6972 11256
rect 6460 11104 6512 11110
rect 6460 11046 6512 11052
rect 6828 11104 6880 11110
rect 6828 11046 6880 11052
rect 7196 11104 7248 11110
rect 7196 11046 7248 11052
rect 5540 11036 5592 11042
rect 5540 10978 5592 10984
rect 5908 11036 5960 11042
rect 5908 10978 5960 10984
rect 6276 11036 6328 11042
rect 6276 10978 6328 10984
rect 5216 10868 5512 10888
rect 5272 10866 5296 10868
rect 5352 10866 5376 10868
rect 5432 10866 5456 10868
rect 5294 10814 5296 10866
rect 5358 10814 5370 10866
rect 5432 10814 5434 10866
rect 5272 10812 5296 10814
rect 5352 10812 5376 10814
rect 5432 10812 5456 10814
rect 5216 10792 5512 10812
rect 4988 10696 5040 10702
rect 4988 10638 5040 10644
rect 4896 10628 4948 10634
rect 4896 10570 4948 10576
rect 4908 10430 4936 10570
rect 4896 10424 4948 10430
rect 4896 10366 4948 10372
rect 5000 8866 5028 10638
rect 5552 9886 5580 10978
rect 5920 10770 5948 10978
rect 5908 10764 5960 10770
rect 5908 10706 5960 10712
rect 6092 10696 6144 10702
rect 6144 10644 6224 10650
rect 6092 10638 6224 10644
rect 6000 10628 6052 10634
rect 6104 10622 6224 10638
rect 6288 10634 6316 10978
rect 6000 10570 6052 10576
rect 6012 10265 6040 10570
rect 5998 10256 6054 10265
rect 5998 10191 6054 10200
rect 6000 10152 6052 10158
rect 6000 10094 6052 10100
rect 6012 10022 6040 10094
rect 6000 10016 6052 10022
rect 6000 9958 6052 9964
rect 5724 9948 5776 9954
rect 5724 9890 5776 9896
rect 5540 9880 5592 9886
rect 5540 9822 5592 9828
rect 5216 9780 5512 9800
rect 5272 9778 5296 9780
rect 5352 9778 5376 9780
rect 5432 9778 5456 9780
rect 5294 9726 5296 9778
rect 5358 9726 5370 9778
rect 5432 9726 5434 9778
rect 5272 9724 5296 9726
rect 5352 9724 5376 9726
rect 5432 9724 5456 9726
rect 5216 9704 5512 9724
rect 5552 8934 5580 9822
rect 5736 9682 5764 9890
rect 6196 9886 6224 10622
rect 6276 10628 6328 10634
rect 6276 10570 6328 10576
rect 6460 10628 6512 10634
rect 6460 10570 6512 10576
rect 6472 10430 6500 10570
rect 6840 10566 6868 11046
rect 7012 10696 7064 10702
rect 7012 10638 7064 10644
rect 6552 10560 6604 10566
rect 6552 10502 6604 10508
rect 6828 10560 6880 10566
rect 6828 10502 6880 10508
rect 6460 10424 6512 10430
rect 6460 10366 6512 10372
rect 6274 10256 6330 10265
rect 6274 10191 6330 10200
rect 6184 9880 6236 9886
rect 6184 9822 6236 9828
rect 5724 9676 5776 9682
rect 6196 9634 6224 9822
rect 5724 9618 5776 9624
rect 5920 9606 6224 9634
rect 5920 9478 5948 9606
rect 5908 9472 5960 9478
rect 5908 9414 5960 9420
rect 5540 8928 5592 8934
rect 5540 8870 5592 8876
rect 4988 8860 5040 8866
rect 4988 8802 5040 8808
rect 5000 8458 5028 8802
rect 5216 8692 5512 8712
rect 5272 8690 5296 8692
rect 5352 8690 5376 8692
rect 5432 8690 5456 8692
rect 5294 8638 5296 8690
rect 5358 8638 5370 8690
rect 5432 8638 5434 8690
rect 5272 8636 5296 8638
rect 5352 8636 5376 8638
rect 5432 8636 5456 8638
rect 5216 8616 5512 8636
rect 5552 8526 5580 8870
rect 5908 8588 5960 8594
rect 5908 8530 5960 8536
rect 5540 8520 5592 8526
rect 5540 8462 5592 8468
rect 4988 8452 5040 8458
rect 4988 8394 5040 8400
rect 5000 7982 5028 8394
rect 5920 8050 5948 8530
rect 6000 8248 6052 8254
rect 6000 8190 6052 8196
rect 5908 8044 5960 8050
rect 5908 7986 5960 7992
rect 4988 7976 5040 7982
rect 4988 7918 5040 7924
rect 5920 7914 5948 7986
rect 5908 7908 5960 7914
rect 5908 7850 5960 7856
rect 5724 7704 5776 7710
rect 5724 7646 5776 7652
rect 5216 7604 5512 7624
rect 5272 7602 5296 7604
rect 5352 7602 5376 7604
rect 5432 7602 5456 7604
rect 5294 7550 5296 7602
rect 5358 7550 5370 7602
rect 5432 7550 5434 7602
rect 5272 7548 5296 7550
rect 5352 7548 5376 7550
rect 5432 7548 5456 7550
rect 5216 7528 5512 7548
rect 5540 7364 5592 7370
rect 5540 7306 5592 7312
rect 4988 7296 5040 7302
rect 4988 7238 5040 7244
rect 5080 7296 5132 7302
rect 5080 7238 5132 7244
rect 5000 6758 5028 7238
rect 4988 6752 5040 6758
rect 4988 6694 5040 6700
rect 4896 6276 4948 6282
rect 4896 6218 4948 6224
rect 4908 5670 4936 6218
rect 5000 6078 5028 6694
rect 4988 6072 5040 6078
rect 4988 6014 5040 6020
rect 4896 5664 4948 5670
rect 4896 5606 4948 5612
rect 4908 4106 4936 5606
rect 4896 4100 4948 4106
rect 4896 4042 4948 4048
rect 4908 3562 4936 4042
rect 5092 3850 5120 7238
rect 5216 6516 5512 6536
rect 5272 6514 5296 6516
rect 5352 6514 5376 6516
rect 5432 6514 5456 6516
rect 5294 6462 5296 6514
rect 5358 6462 5370 6514
rect 5432 6462 5434 6514
rect 5272 6460 5296 6462
rect 5352 6460 5376 6462
rect 5432 6460 5456 6462
rect 5216 6440 5512 6460
rect 5216 5428 5512 5448
rect 5272 5426 5296 5428
rect 5352 5426 5376 5428
rect 5432 5426 5456 5428
rect 5294 5374 5296 5426
rect 5358 5374 5370 5426
rect 5432 5374 5434 5426
rect 5272 5372 5296 5374
rect 5352 5372 5376 5374
rect 5432 5372 5456 5374
rect 5216 5352 5512 5372
rect 5552 4786 5580 7306
rect 5632 7160 5684 7166
rect 5632 7102 5684 7108
rect 5644 6894 5672 7102
rect 5632 6888 5684 6894
rect 5632 6830 5684 6836
rect 5630 6720 5686 6729
rect 5630 6655 5686 6664
rect 5644 6078 5672 6655
rect 5736 6282 5764 7646
rect 5816 7160 5868 7166
rect 5816 7102 5868 7108
rect 5724 6276 5776 6282
rect 5724 6218 5776 6224
rect 5632 6072 5684 6078
rect 5632 6014 5684 6020
rect 5644 5330 5672 6014
rect 5632 5324 5684 5330
rect 5632 5266 5684 5272
rect 5540 4780 5592 4786
rect 5540 4722 5592 4728
rect 5736 4514 5764 6218
rect 5828 5670 5856 7102
rect 6012 6865 6040 8190
rect 6288 7420 6316 10191
rect 6472 9138 6500 10366
rect 6564 10022 6592 10502
rect 6840 10158 6868 10502
rect 6828 10152 6880 10158
rect 6828 10094 6880 10100
rect 6920 10152 6972 10158
rect 6920 10094 6972 10100
rect 6552 10016 6604 10022
rect 6552 9958 6604 9964
rect 6552 9608 6604 9614
rect 6552 9550 6604 9556
rect 6460 9132 6512 9138
rect 6460 9074 6512 9080
rect 6460 7432 6512 7438
rect 6288 7392 6460 7420
rect 6184 7160 6236 7166
rect 6184 7102 6236 7108
rect 5998 6856 6054 6865
rect 5998 6791 6054 6800
rect 5908 6140 5960 6146
rect 5908 6082 5960 6088
rect 5920 5670 5948 6082
rect 6000 5732 6052 5738
rect 6000 5674 6052 5680
rect 5816 5664 5868 5670
rect 5816 5606 5868 5612
rect 5908 5664 5960 5670
rect 5908 5606 5960 5612
rect 6012 5330 6040 5674
rect 6000 5324 6052 5330
rect 6000 5266 6052 5272
rect 5908 5188 5960 5194
rect 5908 5130 5960 5136
rect 5724 4508 5776 4514
rect 5724 4450 5776 4456
rect 5216 4340 5512 4360
rect 5272 4338 5296 4340
rect 5352 4338 5376 4340
rect 5432 4338 5456 4340
rect 5294 4286 5296 4338
rect 5358 4286 5370 4338
rect 5432 4286 5434 4338
rect 5272 4284 5296 4286
rect 5352 4284 5376 4286
rect 5432 4284 5456 4286
rect 5216 4264 5512 4284
rect 5920 4174 5948 5130
rect 6012 4650 6040 5266
rect 6196 4990 6224 7102
rect 6288 6826 6316 7392
rect 6460 7374 6512 7380
rect 6276 6820 6328 6826
rect 6276 6762 6328 6768
rect 6288 5330 6316 6762
rect 6368 6752 6420 6758
rect 6460 6752 6512 6758
rect 6368 6694 6420 6700
rect 6458 6720 6460 6729
rect 6512 6720 6514 6729
rect 6380 5874 6408 6694
rect 6458 6655 6514 6664
rect 6564 6350 6592 9550
rect 6644 9472 6696 9478
rect 6642 9440 6644 9449
rect 6696 9440 6698 9449
rect 6642 9375 6698 9384
rect 6840 8882 6868 10094
rect 6932 9546 6960 10094
rect 7024 9682 7052 10638
rect 7104 10560 7156 10566
rect 7104 10502 7156 10508
rect 7116 9682 7144 10502
rect 7012 9676 7064 9682
rect 7012 9618 7064 9624
rect 7104 9676 7156 9682
rect 7104 9618 7156 9624
rect 7024 9585 7052 9618
rect 7010 9576 7066 9585
rect 6920 9540 6972 9546
rect 7010 9511 7066 9520
rect 6920 9482 6972 9488
rect 7102 9440 7158 9449
rect 7102 9375 7104 9384
rect 7156 9375 7158 9384
rect 7104 9346 7156 9352
rect 6920 9336 6972 9342
rect 6920 9278 6972 9284
rect 6932 9070 6960 9278
rect 6920 9064 6972 9070
rect 6920 9006 6972 9012
rect 7208 8934 7236 11046
rect 6920 8928 6972 8934
rect 6840 8876 6920 8882
rect 6840 8870 6972 8876
rect 7196 8928 7248 8934
rect 7196 8870 7248 8876
rect 6840 8854 6960 8870
rect 7104 8520 7156 8526
rect 6840 8468 7104 8474
rect 6840 8462 7156 8468
rect 6840 8446 7144 8462
rect 6644 7772 6696 7778
rect 6644 7714 6696 7720
rect 6656 7522 6684 7714
rect 6840 7710 6868 8446
rect 7196 8248 7248 8254
rect 7196 8190 7248 8196
rect 7208 7914 7236 8190
rect 7196 7908 7248 7914
rect 7196 7850 7248 7856
rect 6828 7704 6880 7710
rect 6828 7646 6880 7652
rect 6656 7494 6960 7522
rect 6736 7364 6788 7370
rect 6736 7306 6788 7312
rect 6644 6888 6696 6894
rect 6642 6856 6644 6865
rect 6696 6856 6698 6865
rect 6642 6791 6698 6800
rect 6748 6604 6776 7306
rect 6828 7228 6880 7234
rect 6828 7170 6880 7176
rect 6656 6576 6776 6604
rect 6552 6344 6604 6350
rect 6552 6286 6604 6292
rect 6460 6276 6512 6282
rect 6460 6218 6512 6224
rect 6368 5868 6420 5874
rect 6368 5810 6420 5816
rect 6276 5324 6328 5330
rect 6276 5266 6328 5272
rect 6276 5188 6328 5194
rect 6276 5130 6328 5136
rect 6184 4984 6236 4990
rect 6184 4926 6236 4932
rect 6000 4644 6052 4650
rect 6000 4586 6052 4592
rect 6092 4576 6144 4582
rect 6092 4518 6144 4524
rect 5908 4168 5960 4174
rect 5908 4110 5960 4116
rect 6104 4106 6132 4518
rect 6092 4100 6144 4106
rect 6092 4042 6144 4048
rect 6196 3902 6224 4926
rect 6288 4786 6316 5130
rect 6368 5120 6420 5126
rect 6368 5062 6420 5068
rect 6276 4780 6328 4786
rect 6276 4722 6328 4728
rect 6288 4038 6316 4722
rect 6380 4106 6408 5062
rect 6368 4100 6420 4106
rect 6368 4042 6420 4048
rect 6276 4032 6328 4038
rect 6276 3974 6328 3980
rect 5908 3896 5960 3902
rect 5092 3822 5304 3850
rect 5908 3838 5960 3844
rect 6184 3896 6236 3902
rect 6184 3838 6236 3844
rect 5080 3692 5132 3698
rect 5080 3634 5132 3640
rect 4896 3556 4948 3562
rect 4896 3498 4948 3504
rect 4988 3556 5040 3562
rect 4988 3498 5040 3504
rect 5000 2734 5028 3498
rect 5092 3034 5120 3634
rect 5276 3426 5304 3822
rect 5920 3698 5948 3838
rect 5908 3692 5960 3698
rect 5908 3634 5960 3640
rect 6288 3562 6316 3974
rect 5816 3556 5868 3562
rect 5816 3498 5868 3504
rect 6276 3556 6328 3562
rect 6276 3498 6328 3504
rect 5632 3488 5684 3494
rect 5632 3430 5684 3436
rect 5724 3488 5776 3494
rect 5724 3430 5776 3436
rect 5264 3420 5316 3426
rect 5264 3362 5316 3368
rect 5216 3252 5512 3272
rect 5272 3250 5296 3252
rect 5352 3250 5376 3252
rect 5432 3250 5456 3252
rect 5294 3198 5296 3250
rect 5358 3198 5370 3250
rect 5432 3198 5434 3250
rect 5272 3196 5296 3198
rect 5352 3196 5376 3198
rect 5432 3196 5456 3198
rect 5216 3176 5512 3196
rect 5644 3086 5672 3430
rect 5632 3080 5684 3086
rect 5092 3006 5304 3034
rect 5632 3022 5684 3028
rect 4816 2706 4936 2734
rect 5000 2706 5120 2734
rect 4712 2604 4764 2610
rect 4712 2546 4764 2552
rect 4712 2400 4764 2406
rect 4764 2360 4844 2388
rect 4712 2342 4764 2348
rect 4712 1992 4764 1998
rect 4712 1934 4764 1940
rect 4620 1924 4672 1930
rect 4620 1866 4672 1872
rect 4528 1720 4580 1726
rect 4528 1662 4580 1668
rect 4540 1402 4568 1662
rect 4724 1522 4752 1934
rect 4712 1516 4764 1522
rect 4712 1458 4764 1464
rect 4540 1374 4660 1402
rect 3976 1312 4028 1318
rect 3976 1254 4028 1260
rect 4344 1312 4396 1318
rect 4344 1254 4396 1260
rect 4528 1312 4580 1318
rect 4528 1254 4580 1260
rect 4540 978 4568 1254
rect 4528 972 4580 978
rect 4528 914 4580 920
rect 3792 904 3844 910
rect 3792 846 3844 852
rect 3240 768 3292 774
rect 3516 768 3568 774
rect 3240 710 3292 716
rect 3514 736 3516 745
rect 3568 736 3570 745
rect 3252 366 3280 710
rect 4632 706 4660 1374
rect 3514 671 3570 680
rect 4620 700 4672 706
rect 4620 642 4672 648
rect 4816 366 4844 2360
rect 4908 2270 4936 2706
rect 4896 2264 4948 2270
rect 4896 2206 4948 2212
rect 5092 2066 5120 2706
rect 5276 2338 5304 3006
rect 5736 2610 5764 3430
rect 5828 3154 5856 3498
rect 5908 3420 5960 3426
rect 5908 3362 5960 3368
rect 5920 3154 5948 3362
rect 5816 3148 5868 3154
rect 5816 3090 5868 3096
rect 5908 3148 5960 3154
rect 5908 3090 5960 3096
rect 6000 3012 6052 3018
rect 6000 2954 6052 2960
rect 6184 3012 6236 3018
rect 6184 2954 6236 2960
rect 5908 2808 5960 2814
rect 5908 2750 5960 2756
rect 5724 2604 5776 2610
rect 5724 2546 5776 2552
rect 5632 2468 5684 2474
rect 5632 2410 5684 2416
rect 5264 2332 5316 2338
rect 5264 2274 5316 2280
rect 5216 2164 5512 2184
rect 5272 2162 5296 2164
rect 5352 2162 5376 2164
rect 5432 2162 5456 2164
rect 5294 2110 5296 2162
rect 5358 2110 5370 2162
rect 5432 2110 5434 2162
rect 5272 2108 5296 2110
rect 5352 2108 5376 2110
rect 5432 2108 5456 2110
rect 5216 2088 5512 2108
rect 5080 2060 5132 2066
rect 5080 2002 5132 2008
rect 5092 910 5120 2002
rect 5540 1856 5592 1862
rect 5540 1798 5592 1804
rect 5552 1386 5580 1798
rect 5540 1380 5592 1386
rect 5540 1322 5592 1328
rect 5216 1076 5512 1096
rect 5272 1074 5296 1076
rect 5352 1074 5376 1076
rect 5432 1074 5456 1076
rect 5294 1022 5296 1074
rect 5358 1022 5370 1074
rect 5432 1022 5434 1074
rect 5272 1020 5296 1022
rect 5352 1020 5376 1022
rect 5432 1020 5456 1022
rect 5216 1000 5512 1020
rect 5080 904 5132 910
rect 5080 846 5132 852
rect 5552 638 5580 1322
rect 5644 1318 5672 2410
rect 5724 2332 5776 2338
rect 5724 2274 5776 2280
rect 5632 1312 5684 1318
rect 5632 1254 5684 1260
rect 5736 1250 5764 2274
rect 5920 1930 5948 2750
rect 5908 1924 5960 1930
rect 5908 1866 5960 1872
rect 6012 1794 6040 2954
rect 6196 1862 6224 2954
rect 6276 2944 6328 2950
rect 6276 2886 6328 2892
rect 6288 2338 6316 2886
rect 6276 2332 6328 2338
rect 6276 2274 6328 2280
rect 6288 1998 6316 2274
rect 6276 1992 6328 1998
rect 6276 1934 6328 1940
rect 6184 1856 6236 1862
rect 6184 1798 6236 1804
rect 6000 1788 6052 1794
rect 6000 1730 6052 1736
rect 5724 1244 5776 1250
rect 5724 1186 5776 1192
rect 5736 842 5764 1186
rect 6288 910 6316 1934
rect 6472 1522 6500 6218
rect 6656 5126 6684 6576
rect 6840 6350 6868 7170
rect 6828 6344 6880 6350
rect 6828 6286 6880 6292
rect 6840 5670 6868 6286
rect 6932 5806 6960 7494
rect 7012 7364 7064 7370
rect 7012 7306 7064 7312
rect 7024 6418 7052 7306
rect 7208 6622 7236 7850
rect 7196 6616 7248 6622
rect 7196 6558 7248 6564
rect 7012 6412 7064 6418
rect 7012 6354 7064 6360
rect 7024 5806 7052 6354
rect 6920 5800 6972 5806
rect 6920 5742 6972 5748
rect 7012 5800 7064 5806
rect 7012 5742 7064 5748
rect 6828 5664 6880 5670
rect 6828 5606 6880 5612
rect 6920 5664 6972 5670
rect 6920 5606 6972 5612
rect 6736 5596 6788 5602
rect 6736 5538 6788 5544
rect 6748 5194 6776 5538
rect 6932 5262 6960 5606
rect 6920 5256 6972 5262
rect 6920 5198 6972 5204
rect 6736 5188 6788 5194
rect 6736 5130 6788 5136
rect 6644 5120 6696 5126
rect 6644 5062 6696 5068
rect 6748 4530 6776 5130
rect 6656 4502 6776 4530
rect 6656 3494 6684 4502
rect 6736 4440 6788 4446
rect 6736 4382 6788 4388
rect 6644 3488 6696 3494
rect 6644 3430 6696 3436
rect 6644 2876 6696 2882
rect 6644 2818 6696 2824
rect 6656 2066 6684 2818
rect 6748 2474 6776 4382
rect 6828 3012 6880 3018
rect 6828 2954 6880 2960
rect 6736 2468 6788 2474
rect 6736 2410 6788 2416
rect 6644 2060 6696 2066
rect 6644 2002 6696 2008
rect 6748 1930 6776 2410
rect 6840 1998 6868 2954
rect 6932 2950 6960 5198
rect 7104 5120 7156 5126
rect 7104 5062 7156 5068
rect 7116 4242 7144 5062
rect 7196 4508 7248 4514
rect 7196 4450 7248 4456
rect 7104 4236 7156 4242
rect 7104 4178 7156 4184
rect 7208 3494 7236 4450
rect 7196 3488 7248 3494
rect 7196 3430 7248 3436
rect 6920 2944 6972 2950
rect 6920 2886 6972 2892
rect 7300 2734 7328 11998
rect 7564 11512 7616 11518
rect 7564 11454 7616 11460
rect 7472 11240 7524 11246
rect 7472 11182 7524 11188
rect 7380 11172 7432 11178
rect 7380 11114 7432 11120
rect 7392 9546 7420 11114
rect 7484 11042 7512 11182
rect 7472 11036 7524 11042
rect 7472 10978 7524 10984
rect 7472 10764 7524 10770
rect 7472 10706 7524 10712
rect 7484 9954 7512 10706
rect 7472 9948 7524 9954
rect 7472 9890 7524 9896
rect 7576 9886 7604 11454
rect 7654 11072 7710 11081
rect 7654 11007 7656 11016
rect 7708 11007 7710 11016
rect 7656 10978 7708 10984
rect 7760 10566 7788 12678
rect 7852 12500 8148 12520
rect 7908 12498 7932 12500
rect 7988 12498 8012 12500
rect 8068 12498 8092 12500
rect 7930 12446 7932 12498
rect 7994 12446 8006 12498
rect 8068 12446 8070 12498
rect 7908 12444 7932 12446
rect 7988 12444 8012 12446
rect 8068 12444 8092 12446
rect 7852 12424 8148 12444
rect 8772 12402 8800 12746
rect 8760 12396 8812 12402
rect 8760 12338 8812 12344
rect 8956 12266 8984 12746
rect 9140 12606 9168 12746
rect 9128 12600 9180 12606
rect 9128 12542 9180 12548
rect 8944 12260 8996 12266
rect 8944 12202 8996 12208
rect 8208 12192 8260 12198
rect 8208 12134 8260 12140
rect 8852 12192 8904 12198
rect 8852 12134 8904 12140
rect 7852 11412 8148 11432
rect 7908 11410 7932 11412
rect 7988 11410 8012 11412
rect 8068 11410 8092 11412
rect 7930 11358 7932 11410
rect 7994 11358 8006 11410
rect 8068 11358 8070 11410
rect 7908 11356 7932 11358
rect 7988 11356 8012 11358
rect 8068 11356 8092 11358
rect 7852 11336 8148 11356
rect 8220 11178 8248 12134
rect 8668 12056 8720 12062
rect 8668 11998 8720 12004
rect 8680 11790 8708 11998
rect 8392 11784 8444 11790
rect 8668 11784 8720 11790
rect 8444 11744 8616 11772
rect 8392 11726 8444 11732
rect 8300 11716 8352 11722
rect 8300 11658 8352 11664
rect 8312 11314 8340 11658
rect 8392 11648 8444 11654
rect 8392 11590 8444 11596
rect 8300 11308 8352 11314
rect 8300 11250 8352 11256
rect 8404 11178 8432 11590
rect 8588 11314 8616 11744
rect 8668 11726 8720 11732
rect 8864 11518 8892 12134
rect 8944 12124 8996 12130
rect 8944 12066 8996 12072
rect 8852 11512 8904 11518
rect 8852 11454 8904 11460
rect 8576 11308 8628 11314
rect 8576 11250 8628 11256
rect 8208 11172 8260 11178
rect 8208 11114 8260 11120
rect 8300 11172 8352 11178
rect 8300 11114 8352 11120
rect 8392 11172 8444 11178
rect 8392 11114 8444 11120
rect 7748 10560 7800 10566
rect 7748 10502 7800 10508
rect 7564 9880 7616 9886
rect 7564 9822 7616 9828
rect 7656 9880 7708 9886
rect 7656 9822 7708 9828
rect 7576 9634 7604 9822
rect 7484 9606 7604 9634
rect 7380 9540 7432 9546
rect 7484 9528 7512 9606
rect 7484 9500 7604 9528
rect 7380 9482 7432 9488
rect 7392 7778 7420 9482
rect 7576 9410 7604 9500
rect 7564 9404 7616 9410
rect 7564 9346 7616 9352
rect 7668 9342 7696 9822
rect 7760 9634 7788 10502
rect 8208 10424 8260 10430
rect 8208 10366 8260 10372
rect 7852 10324 8148 10344
rect 7908 10322 7932 10324
rect 7988 10322 8012 10324
rect 8068 10322 8092 10324
rect 7930 10270 7932 10322
rect 7994 10270 8006 10322
rect 8068 10270 8070 10322
rect 7908 10268 7932 10270
rect 7988 10268 8012 10270
rect 8068 10268 8092 10270
rect 7852 10248 8148 10268
rect 7932 10152 7984 10158
rect 7932 10094 7984 10100
rect 7760 9606 7880 9634
rect 7852 9460 7880 9606
rect 7944 9546 7972 10094
rect 8220 9954 8248 10366
rect 8312 10158 8340 11114
rect 8588 10702 8616 11250
rect 8864 11110 8892 11454
rect 8956 11246 8984 12066
rect 8944 11240 8996 11246
rect 8944 11182 8996 11188
rect 8956 11110 8984 11182
rect 8852 11104 8904 11110
rect 8852 11046 8904 11052
rect 8944 11104 8996 11110
rect 8944 11046 8996 11052
rect 8576 10696 8628 10702
rect 8576 10638 8628 10644
rect 8300 10152 8352 10158
rect 8300 10094 8352 10100
rect 8208 9948 8260 9954
rect 8208 9890 8260 9896
rect 8220 9585 8248 9890
rect 8206 9576 8262 9585
rect 7932 9540 7984 9546
rect 9140 9546 9168 12542
rect 9496 12396 9548 12402
rect 9496 12338 9548 12344
rect 9404 12260 9456 12266
rect 9404 12202 9456 12208
rect 9416 11858 9444 12202
rect 9404 11852 9456 11858
rect 9404 11794 9456 11800
rect 9416 11110 9444 11794
rect 9404 11104 9456 11110
rect 9404 11046 9456 11052
rect 9416 10770 9444 11046
rect 9404 10764 9456 10770
rect 9404 10706 9456 10712
rect 9310 10664 9366 10673
rect 9508 10634 9536 12338
rect 9864 12260 9916 12266
rect 9864 12202 9916 12208
rect 9588 12192 9640 12198
rect 9588 12134 9640 12140
rect 9600 11858 9628 12134
rect 9588 11852 9640 11858
rect 9588 11794 9640 11800
rect 9600 10770 9628 11794
rect 9680 11648 9732 11654
rect 9680 11590 9732 11596
rect 9588 10764 9640 10770
rect 9588 10706 9640 10712
rect 9310 10599 9312 10608
rect 9364 10599 9366 10608
rect 9496 10628 9548 10634
rect 9312 10570 9364 10576
rect 9496 10570 9548 10576
rect 9324 10022 9352 10570
rect 9312 10016 9364 10022
rect 9312 9958 9364 9964
rect 9600 9886 9628 10706
rect 9692 10634 9720 11590
rect 9876 11178 9904 12202
rect 10876 12124 10928 12130
rect 10876 12066 10928 12072
rect 11152 12124 11204 12130
rect 11152 12066 11204 12072
rect 10488 11956 10784 11976
rect 10544 11954 10568 11956
rect 10624 11954 10648 11956
rect 10704 11954 10728 11956
rect 10566 11902 10568 11954
rect 10630 11902 10642 11954
rect 10704 11902 10706 11954
rect 10544 11900 10568 11902
rect 10624 11900 10648 11902
rect 10704 11900 10728 11902
rect 10488 11880 10784 11900
rect 10888 11790 10916 12066
rect 11164 11858 11192 12066
rect 11152 11852 11204 11858
rect 11152 11794 11204 11800
rect 9956 11784 10008 11790
rect 9956 11726 10008 11732
rect 10876 11784 10928 11790
rect 10876 11726 10928 11732
rect 9968 11314 9996 11726
rect 10048 11648 10100 11654
rect 10048 11590 10100 11596
rect 9956 11308 10008 11314
rect 9956 11250 10008 11256
rect 9864 11172 9916 11178
rect 9864 11114 9916 11120
rect 9680 10628 9732 10634
rect 9680 10570 9732 10576
rect 9588 9880 9640 9886
rect 9588 9822 9640 9828
rect 8206 9511 8262 9520
rect 8392 9540 8444 9546
rect 7932 9482 7984 9488
rect 8220 9478 8248 9511
rect 8668 9540 8720 9546
rect 8444 9500 8524 9528
rect 8392 9482 8444 9488
rect 7760 9432 7880 9460
rect 8208 9472 8260 9478
rect 7656 9336 7708 9342
rect 7656 9278 7708 9284
rect 7656 8384 7708 8390
rect 7656 8326 7708 8332
rect 7668 8050 7696 8326
rect 7656 8044 7708 8050
rect 7656 7986 7708 7992
rect 7472 7840 7524 7846
rect 7472 7782 7524 7788
rect 7380 7772 7432 7778
rect 7380 7714 7432 7720
rect 7484 6962 7512 7782
rect 7564 7364 7616 7370
rect 7668 7352 7696 7986
rect 7616 7324 7696 7352
rect 7564 7306 7616 7312
rect 7472 6956 7524 6962
rect 7472 6898 7524 6904
rect 7760 6418 7788 9432
rect 8208 9414 8260 9420
rect 8390 9440 8446 9449
rect 8390 9375 8392 9384
rect 8444 9375 8446 9384
rect 8392 9346 8444 9352
rect 7852 9236 8148 9256
rect 7908 9234 7932 9236
rect 7988 9234 8012 9236
rect 8068 9234 8092 9236
rect 7930 9182 7932 9234
rect 7994 9182 8006 9234
rect 8068 9182 8070 9234
rect 7908 9180 7932 9182
rect 7988 9180 8012 9182
rect 8068 9180 8092 9182
rect 7852 9160 8148 9180
rect 8300 8316 8352 8322
rect 8300 8258 8352 8264
rect 7852 8148 8148 8168
rect 7908 8146 7932 8148
rect 7988 8146 8012 8148
rect 8068 8146 8092 8148
rect 7930 8094 7932 8146
rect 7994 8094 8006 8146
rect 8068 8094 8070 8146
rect 7908 8092 7932 8094
rect 7988 8092 8012 8094
rect 8068 8092 8092 8094
rect 7852 8072 8148 8092
rect 7840 7704 7892 7710
rect 7840 7646 7892 7652
rect 7852 7438 7880 7646
rect 7840 7432 7892 7438
rect 7840 7374 7892 7380
rect 7852 7060 8148 7080
rect 7908 7058 7932 7060
rect 7988 7058 8012 7060
rect 8068 7058 8092 7060
rect 7930 7006 7932 7058
rect 7994 7006 8006 7058
rect 8068 7006 8070 7058
rect 7908 7004 7932 7006
rect 7988 7004 8012 7006
rect 8068 7004 8092 7006
rect 7852 6984 8148 7004
rect 7748 6412 7800 6418
rect 7748 6354 7800 6360
rect 7852 5972 8148 5992
rect 7908 5970 7932 5972
rect 7988 5970 8012 5972
rect 8068 5970 8092 5972
rect 7930 5918 7932 5970
rect 7994 5918 8006 5970
rect 8068 5918 8070 5970
rect 7908 5916 7932 5918
rect 7988 5916 8012 5918
rect 8068 5916 8092 5918
rect 7852 5896 8148 5916
rect 7380 5120 7432 5126
rect 7380 5062 7432 5068
rect 7392 3970 7420 5062
rect 7852 4884 8148 4904
rect 7908 4882 7932 4884
rect 7988 4882 8012 4884
rect 8068 4882 8092 4884
rect 7930 4830 7932 4882
rect 7994 4830 8006 4882
rect 8068 4830 8070 4882
rect 7908 4828 7932 4830
rect 7988 4828 8012 4830
rect 8068 4828 8092 4830
rect 7852 4808 8148 4828
rect 7380 3964 7432 3970
rect 7380 3906 7432 3912
rect 7852 3796 8148 3816
rect 7908 3794 7932 3796
rect 7988 3794 8012 3796
rect 8068 3794 8092 3796
rect 7930 3742 7932 3794
rect 7994 3742 8006 3794
rect 8068 3742 8070 3794
rect 7908 3740 7932 3742
rect 7988 3740 8012 3742
rect 8068 3740 8092 3742
rect 7852 3720 8148 3740
rect 7840 3624 7892 3630
rect 7840 3566 7892 3572
rect 7748 3352 7800 3358
rect 7748 3294 7800 3300
rect 7208 2706 7328 2734
rect 7208 2474 7236 2706
rect 7196 2468 7248 2474
rect 7196 2410 7248 2416
rect 7288 2400 7340 2406
rect 7288 2342 7340 2348
rect 6920 2332 6972 2338
rect 6920 2274 6972 2280
rect 6828 1992 6880 1998
rect 6828 1934 6880 1940
rect 6736 1924 6788 1930
rect 6736 1866 6788 1872
rect 6840 1726 6868 1934
rect 6828 1720 6880 1726
rect 6828 1662 6880 1668
rect 6460 1516 6512 1522
rect 6460 1458 6512 1464
rect 6840 978 6868 1662
rect 6828 972 6880 978
rect 6828 914 6880 920
rect 6276 904 6328 910
rect 6276 846 6328 852
rect 5724 836 5776 842
rect 5724 778 5776 784
rect 4896 632 4948 638
rect 4896 574 4948 580
rect 5540 632 5592 638
rect 5540 574 5592 580
rect 2136 292 2188 298
rect 2136 234 2188 240
rect 2884 286 3004 314
rect 3240 360 3292 366
rect 3240 302 3292 308
rect 4804 360 4856 366
rect 4804 302 4856 308
rect 2884 160 2912 286
rect 4908 160 4936 574
rect 6932 160 6960 2274
rect 7300 2066 7328 2342
rect 7288 2060 7340 2066
rect 7288 2002 7340 2008
rect 7760 1930 7788 3294
rect 7852 3086 7880 3566
rect 8312 3442 8340 8258
rect 8496 7982 8524 9500
rect 8668 9482 8720 9488
rect 9128 9540 9180 9546
rect 9128 9482 9180 9488
rect 8576 9472 8628 9478
rect 8576 9414 8628 9420
rect 8484 7976 8536 7982
rect 8484 7918 8536 7924
rect 8588 7506 8616 9414
rect 8680 9070 8708 9482
rect 9036 9336 9088 9342
rect 9036 9278 9088 9284
rect 8668 9064 8720 9070
rect 8668 9006 8720 9012
rect 8760 8792 8812 8798
rect 8760 8734 8812 8740
rect 8772 7914 8800 8734
rect 9048 8322 9076 9278
rect 9876 9002 9904 11114
rect 9956 10628 10008 10634
rect 9956 10570 10008 10576
rect 9968 9954 9996 10570
rect 10060 10498 10088 11590
rect 10888 11042 10916 11726
rect 11152 11716 11204 11722
rect 11152 11658 11204 11664
rect 10140 11036 10192 11042
rect 10140 10978 10192 10984
rect 10876 11036 10928 11042
rect 10876 10978 10928 10984
rect 10048 10492 10100 10498
rect 10048 10434 10100 10440
rect 10152 10226 10180 10978
rect 10488 10868 10784 10888
rect 10544 10866 10568 10868
rect 10624 10866 10648 10868
rect 10704 10866 10728 10868
rect 10566 10814 10568 10866
rect 10630 10814 10642 10866
rect 10704 10814 10706 10866
rect 10544 10812 10568 10814
rect 10624 10812 10648 10814
rect 10704 10812 10728 10814
rect 10488 10792 10784 10812
rect 10140 10220 10192 10226
rect 10140 10162 10192 10168
rect 9956 9948 10008 9954
rect 9956 9890 10008 9896
rect 10488 9780 10784 9800
rect 10544 9778 10568 9780
rect 10624 9778 10648 9780
rect 10704 9778 10728 9780
rect 10566 9726 10568 9778
rect 10630 9726 10642 9778
rect 10704 9726 10706 9778
rect 10544 9724 10568 9726
rect 10624 9724 10648 9726
rect 10704 9724 10728 9726
rect 10488 9704 10784 9724
rect 10140 9540 10192 9546
rect 10140 9482 10192 9488
rect 10048 9336 10100 9342
rect 10048 9278 10100 9284
rect 9864 8996 9916 9002
rect 9864 8938 9916 8944
rect 9312 8928 9364 8934
rect 9312 8870 9364 8876
rect 9404 8928 9456 8934
rect 9404 8870 9456 8876
rect 9324 8594 9352 8870
rect 9312 8588 9364 8594
rect 9312 8530 9364 8536
rect 9036 8316 9088 8322
rect 9036 8258 9088 8264
rect 8760 7908 8812 7914
rect 8760 7850 8812 7856
rect 9416 7506 9444 8870
rect 9496 8792 9548 8798
rect 9496 8734 9548 8740
rect 9508 7710 9536 8734
rect 9588 8452 9640 8458
rect 9588 8394 9640 8400
rect 9496 7704 9548 7710
rect 9496 7646 9548 7652
rect 8576 7500 8628 7506
rect 8576 7442 8628 7448
rect 9404 7500 9456 7506
rect 9404 7442 9456 7448
rect 9508 7370 9536 7646
rect 9496 7364 9548 7370
rect 9496 7306 9548 7312
rect 9496 6752 9548 6758
rect 9600 6740 9628 8394
rect 9772 8384 9824 8390
rect 9772 8326 9824 8332
rect 9680 8248 9732 8254
rect 9680 8190 9732 8196
rect 9692 6826 9720 8190
rect 9680 6820 9732 6826
rect 9680 6762 9732 6768
rect 9548 6712 9628 6740
rect 9496 6694 9548 6700
rect 8484 6684 8536 6690
rect 8484 6626 8536 6632
rect 8668 6684 8720 6690
rect 8668 6626 8720 6632
rect 8496 5874 8524 6626
rect 8680 6418 8708 6626
rect 8668 6412 8720 6418
rect 8668 6354 8720 6360
rect 8852 6412 8904 6418
rect 8852 6354 8904 6360
rect 8576 6208 8628 6214
rect 8576 6150 8628 6156
rect 8484 5868 8536 5874
rect 8484 5810 8536 5816
rect 8496 5346 8524 5810
rect 8588 5670 8616 6150
rect 8576 5664 8628 5670
rect 8576 5606 8628 5612
rect 8668 5664 8720 5670
rect 8668 5606 8720 5612
rect 8404 5318 8524 5346
rect 8404 4650 8432 5318
rect 8484 5188 8536 5194
rect 8484 5130 8536 5136
rect 8496 4786 8524 5130
rect 8484 4780 8536 4786
rect 8484 4722 8536 4728
rect 8392 4644 8444 4650
rect 8392 4586 8444 4592
rect 8404 3562 8432 4586
rect 8484 4168 8536 4174
rect 8484 4110 8536 4116
rect 8392 3556 8444 3562
rect 8392 3498 8444 3504
rect 8312 3414 8432 3442
rect 8496 3426 8524 4110
rect 8588 3442 8616 5606
rect 8680 4174 8708 5606
rect 8864 5058 8892 6354
rect 9508 6350 9536 6694
rect 9496 6344 9548 6350
rect 9496 6286 9548 6292
rect 9036 6276 9088 6282
rect 9036 6218 9088 6224
rect 8944 5256 8996 5262
rect 8944 5198 8996 5204
rect 8852 5052 8904 5058
rect 8852 4994 8904 5000
rect 8760 4984 8812 4990
rect 8760 4926 8812 4932
rect 8772 4650 8800 4926
rect 8760 4644 8812 4650
rect 8760 4586 8812 4592
rect 8668 4168 8720 4174
rect 8668 4110 8720 4116
rect 8588 3426 8708 3442
rect 7840 3080 7892 3086
rect 7840 3022 7892 3028
rect 7852 2708 8148 2728
rect 7908 2706 7932 2708
rect 7988 2706 8012 2708
rect 8068 2706 8092 2708
rect 7930 2654 7932 2706
rect 7994 2654 8006 2706
rect 8068 2654 8070 2706
rect 7908 2652 7932 2654
rect 7988 2652 8012 2654
rect 8068 2652 8092 2654
rect 7852 2632 8148 2652
rect 7748 1924 7800 1930
rect 7748 1866 7800 1872
rect 8300 1788 8352 1794
rect 8300 1730 8352 1736
rect 7012 1720 7064 1726
rect 7012 1662 7064 1668
rect 7024 1386 7052 1662
rect 7852 1620 8148 1640
rect 7908 1618 7932 1620
rect 7988 1618 8012 1620
rect 8068 1618 8092 1620
rect 7930 1566 7932 1618
rect 7994 1566 8006 1618
rect 8068 1566 8070 1618
rect 7908 1564 7932 1566
rect 7988 1564 8012 1566
rect 8068 1564 8092 1566
rect 7852 1544 8148 1564
rect 7012 1380 7064 1386
rect 7012 1322 7064 1328
rect 8312 1318 8340 1730
rect 8300 1312 8352 1318
rect 8300 1254 8352 1260
rect 8404 842 8432 3414
rect 8484 3420 8536 3426
rect 8588 3420 8720 3426
rect 8588 3414 8668 3420
rect 8484 3362 8536 3368
rect 8668 3362 8720 3368
rect 8772 3086 8800 4586
rect 8864 3154 8892 4994
rect 8956 4038 8984 5198
rect 9048 5194 9076 6218
rect 9220 5664 9272 5670
rect 9220 5606 9272 5612
rect 9036 5188 9088 5194
rect 9036 5130 9088 5136
rect 9128 5120 9180 5126
rect 9128 5062 9180 5068
rect 9036 4508 9088 4514
rect 9036 4450 9088 4456
rect 9048 4242 9076 4450
rect 9036 4236 9088 4242
rect 9036 4178 9088 4184
rect 9140 4106 9168 5062
rect 9232 4990 9260 5606
rect 9324 5590 9628 5618
rect 9784 5602 9812 8326
rect 9876 8322 9904 8938
rect 9956 8792 10008 8798
rect 9956 8734 10008 8740
rect 9864 8316 9916 8322
rect 9864 8258 9916 8264
rect 9876 8050 9904 8258
rect 9864 8044 9916 8050
rect 9864 7986 9916 7992
rect 9876 7370 9904 7986
rect 9968 7658 9996 8734
rect 10060 8458 10088 9278
rect 10048 8452 10100 8458
rect 10048 8394 10100 8400
rect 10152 8050 10180 9482
rect 10888 8798 10916 10978
rect 10968 10968 11020 10974
rect 10968 10910 11020 10916
rect 10980 10634 11008 10910
rect 11060 10764 11112 10770
rect 11060 10706 11112 10712
rect 10968 10628 11020 10634
rect 10968 10570 11020 10576
rect 11072 10022 11100 10706
rect 11060 10016 11112 10022
rect 11060 9958 11112 9964
rect 11164 9954 11192 11658
rect 11440 10770 11468 12746
rect 12072 12668 12124 12674
rect 12072 12610 12124 12616
rect 11428 10764 11480 10770
rect 11428 10706 11480 10712
rect 12084 10634 12112 12610
rect 11612 10628 11664 10634
rect 11612 10570 11664 10576
rect 12072 10628 12124 10634
rect 12072 10570 12124 10576
rect 11520 10560 11572 10566
rect 11520 10502 11572 10508
rect 11532 10022 11560 10502
rect 11520 10016 11572 10022
rect 11520 9958 11572 9964
rect 11152 9948 11204 9954
rect 11152 9890 11204 9896
rect 11520 9540 11572 9546
rect 11520 9482 11572 9488
rect 11428 9336 11480 9342
rect 11428 9278 11480 9284
rect 11060 8996 11112 9002
rect 11060 8938 11112 8944
rect 10876 8792 10928 8798
rect 10876 8734 10928 8740
rect 10488 8692 10784 8712
rect 10544 8690 10568 8692
rect 10624 8690 10648 8692
rect 10704 8690 10728 8692
rect 10566 8638 10568 8690
rect 10630 8638 10642 8690
rect 10704 8638 10706 8690
rect 10544 8636 10568 8638
rect 10624 8636 10648 8638
rect 10704 8636 10728 8638
rect 10488 8616 10784 8636
rect 10876 8452 10928 8458
rect 10876 8394 10928 8400
rect 10140 8044 10192 8050
rect 10140 7986 10192 7992
rect 10048 7772 10100 7778
rect 10048 7714 10100 7720
rect 10060 7658 10088 7714
rect 9968 7630 10088 7658
rect 9968 7506 9996 7630
rect 9956 7500 10008 7506
rect 9956 7442 10008 7448
rect 9864 7364 9916 7370
rect 9864 7306 9916 7312
rect 9968 5602 9996 7442
rect 10152 7302 10180 7986
rect 10488 7604 10784 7624
rect 10544 7602 10568 7604
rect 10624 7602 10648 7604
rect 10704 7602 10728 7604
rect 10566 7550 10568 7602
rect 10630 7550 10642 7602
rect 10704 7550 10706 7602
rect 10544 7548 10568 7550
rect 10624 7548 10648 7550
rect 10704 7548 10728 7550
rect 10488 7528 10784 7548
rect 10888 7438 10916 8394
rect 11072 8050 11100 8938
rect 11336 8452 11388 8458
rect 11336 8394 11388 8400
rect 11152 8384 11204 8390
rect 11152 8326 11204 8332
rect 11060 8044 11112 8050
rect 11060 7986 11112 7992
rect 11060 7772 11112 7778
rect 11060 7714 11112 7720
rect 10876 7432 10928 7438
rect 10876 7374 10928 7380
rect 10140 7296 10192 7302
rect 10140 7238 10192 7244
rect 10152 6826 10180 7238
rect 10140 6820 10192 6826
rect 10140 6762 10192 6768
rect 10888 6758 10916 7374
rect 10876 6752 10928 6758
rect 10876 6694 10928 6700
rect 10488 6516 10784 6536
rect 10544 6514 10568 6516
rect 10624 6514 10648 6516
rect 10704 6514 10728 6516
rect 10566 6462 10568 6514
rect 10630 6462 10642 6514
rect 10704 6462 10706 6514
rect 10544 6460 10568 6462
rect 10624 6460 10648 6462
rect 10704 6460 10728 6462
rect 10488 6440 10784 6460
rect 10140 6276 10192 6282
rect 10140 6218 10192 6224
rect 9324 5534 9352 5590
rect 9600 5534 9628 5590
rect 9772 5596 9824 5602
rect 9772 5538 9824 5544
rect 9956 5596 10008 5602
rect 9956 5538 10008 5544
rect 9312 5528 9364 5534
rect 9312 5470 9364 5476
rect 9404 5528 9456 5534
rect 9404 5470 9456 5476
rect 9588 5528 9640 5534
rect 9968 5482 9996 5538
rect 9588 5470 9640 5476
rect 9416 5330 9444 5470
rect 9692 5454 9996 5482
rect 9404 5324 9456 5330
rect 9404 5266 9456 5272
rect 9220 4984 9272 4990
rect 9220 4926 9272 4932
rect 9692 4514 9720 5454
rect 9862 5224 9918 5233
rect 9862 5159 9918 5168
rect 9876 5126 9904 5159
rect 9864 5120 9916 5126
rect 9864 5062 9916 5068
rect 10152 5058 10180 6218
rect 10488 5428 10784 5448
rect 10544 5426 10568 5428
rect 10624 5426 10648 5428
rect 10704 5426 10728 5428
rect 10566 5374 10568 5426
rect 10630 5374 10642 5426
rect 10704 5374 10706 5426
rect 10544 5372 10568 5374
rect 10624 5372 10648 5374
rect 10704 5372 10728 5374
rect 10488 5352 10784 5372
rect 10140 5052 10192 5058
rect 10140 4994 10192 5000
rect 9680 4508 9732 4514
rect 9680 4450 9732 4456
rect 9692 4224 9720 4450
rect 9600 4196 9720 4224
rect 9128 4100 9180 4106
rect 9128 4042 9180 4048
rect 9312 4100 9364 4106
rect 9600 4088 9628 4196
rect 9772 4168 9824 4174
rect 9772 4110 9824 4116
rect 9312 4042 9364 4048
rect 9416 4060 9628 4088
rect 9680 4100 9732 4106
rect 8944 4032 8996 4038
rect 8944 3974 8996 3980
rect 8956 3630 8984 3974
rect 9324 3630 9352 4042
rect 8944 3624 8996 3630
rect 9312 3624 9364 3630
rect 8996 3584 9076 3612
rect 8944 3566 8996 3572
rect 8944 3352 8996 3358
rect 8944 3294 8996 3300
rect 8852 3148 8904 3154
rect 8852 3090 8904 3096
rect 8576 3080 8628 3086
rect 8576 3022 8628 3028
rect 8760 3080 8812 3086
rect 8760 3022 8812 3028
rect 8588 2734 8616 3022
rect 8668 2944 8720 2950
rect 8668 2886 8720 2892
rect 8496 2706 8616 2734
rect 8496 2270 8524 2706
rect 8484 2264 8536 2270
rect 8484 2206 8536 2212
rect 8496 1726 8524 2206
rect 8484 1720 8536 1726
rect 8484 1662 8536 1668
rect 8680 978 8708 2886
rect 8956 1998 8984 3294
rect 8944 1992 8996 1998
rect 8944 1934 8996 1940
rect 8668 972 8720 978
rect 8668 914 8720 920
rect 8392 836 8444 842
rect 8392 778 8444 784
rect 9048 774 9076 3584
rect 9312 3566 9364 3572
rect 9324 3494 9352 3566
rect 9312 3488 9364 3494
rect 9126 3456 9182 3465
rect 9312 3430 9364 3436
rect 9126 3391 9128 3400
rect 9180 3391 9182 3400
rect 9128 3362 9180 3368
rect 9220 3080 9272 3086
rect 9218 3048 9220 3057
rect 9272 3048 9274 3057
rect 9218 2983 9274 2992
rect 9324 842 9352 3430
rect 9416 3340 9444 4060
rect 9680 4042 9732 4048
rect 9692 3476 9720 4042
rect 9600 3465 9720 3476
rect 9586 3456 9720 3465
rect 9642 3448 9720 3456
rect 9586 3391 9642 3400
rect 9588 3352 9640 3358
rect 9416 3312 9536 3340
rect 9404 3148 9456 3154
rect 9404 3090 9456 3096
rect 9312 836 9364 842
rect 9416 824 9444 3090
rect 9508 3057 9536 3312
rect 9588 3294 9640 3300
rect 9600 3154 9628 3294
rect 9588 3148 9640 3154
rect 9588 3090 9640 3096
rect 9494 3048 9550 3057
rect 9494 2983 9550 2992
rect 9508 2338 9536 2983
rect 9692 2814 9720 3448
rect 9784 2882 9812 4110
rect 10152 4106 10180 4994
rect 10324 4780 10376 4786
rect 10324 4722 10376 4728
rect 10336 4446 10364 4722
rect 10888 4650 10916 6694
rect 11072 5534 11100 7714
rect 11164 7506 11192 8326
rect 11348 8050 11376 8394
rect 11336 8044 11388 8050
rect 11336 7986 11388 7992
rect 11244 7976 11296 7982
rect 11244 7918 11296 7924
rect 11152 7500 11204 7506
rect 11152 7442 11204 7448
rect 11256 7370 11284 7918
rect 11336 7840 11388 7846
rect 11336 7782 11388 7788
rect 11244 7364 11296 7370
rect 11244 7306 11296 7312
rect 11256 6826 11284 7306
rect 11244 6820 11296 6826
rect 11244 6762 11296 6768
rect 11348 6418 11376 7782
rect 11440 7438 11468 9278
rect 11532 8322 11560 9482
rect 11520 8316 11572 8322
rect 11520 8258 11572 8264
rect 11428 7432 11480 7438
rect 11428 7374 11480 7380
rect 11440 6690 11468 7374
rect 11428 6684 11480 6690
rect 11428 6626 11480 6632
rect 11532 6622 11560 8258
rect 11520 6616 11572 6622
rect 11520 6558 11572 6564
rect 11624 6434 11652 10570
rect 11888 10560 11940 10566
rect 11888 10502 11940 10508
rect 11900 9886 11928 10502
rect 12716 10424 12768 10430
rect 12716 10366 12768 10372
rect 12164 10152 12216 10158
rect 12164 10094 12216 10100
rect 11888 9880 11940 9886
rect 11888 9822 11940 9828
rect 11796 9540 11848 9546
rect 11796 9482 11848 9488
rect 11808 8594 11836 9482
rect 11796 8588 11848 8594
rect 11796 8530 11848 8536
rect 11704 8044 11756 8050
rect 11704 7986 11756 7992
rect 11716 7370 11744 7986
rect 11704 7364 11756 7370
rect 11704 7306 11756 7312
rect 11716 6894 11744 7306
rect 11704 6888 11756 6894
rect 11704 6830 11756 6836
rect 11704 6616 11756 6622
rect 11704 6558 11756 6564
rect 11336 6412 11388 6418
rect 11336 6354 11388 6360
rect 11532 6406 11652 6434
rect 11428 6276 11480 6282
rect 11428 6218 11480 6224
rect 11440 6078 11468 6218
rect 11428 6072 11480 6078
rect 11428 6014 11480 6020
rect 10968 5528 11020 5534
rect 10968 5470 11020 5476
rect 11060 5528 11112 5534
rect 11060 5470 11112 5476
rect 10980 5194 11008 5470
rect 10968 5188 11020 5194
rect 10968 5130 11020 5136
rect 10876 4644 10928 4650
rect 10876 4586 10928 4592
rect 10980 4530 11008 5130
rect 11072 4786 11100 5470
rect 11244 5324 11296 5330
rect 11244 5266 11296 5272
rect 11256 4786 11284 5266
rect 11060 4780 11112 4786
rect 11060 4722 11112 4728
rect 11244 4780 11296 4786
rect 11244 4722 11296 4728
rect 10888 4502 11008 4530
rect 11152 4508 11204 4514
rect 10888 4446 10916 4502
rect 11152 4450 11204 4456
rect 10324 4440 10376 4446
rect 10324 4382 10376 4388
rect 10416 4440 10468 4446
rect 10416 4382 10468 4388
rect 10876 4440 10928 4446
rect 10876 4382 10928 4388
rect 10140 4100 10192 4106
rect 10140 4042 10192 4048
rect 9864 3488 9916 3494
rect 9864 3430 9916 3436
rect 9876 2950 9904 3430
rect 9956 3420 10008 3426
rect 9956 3362 10008 3368
rect 9864 2944 9916 2950
rect 9864 2886 9916 2892
rect 9772 2876 9824 2882
rect 9772 2818 9824 2824
rect 9680 2808 9732 2814
rect 9680 2750 9732 2756
rect 9784 2610 9812 2818
rect 9772 2604 9824 2610
rect 9772 2546 9824 2552
rect 9496 2332 9548 2338
rect 9496 2274 9548 2280
rect 9508 1980 9536 2274
rect 9680 1992 9732 1998
rect 9508 1952 9680 1980
rect 9600 1250 9628 1952
rect 9680 1934 9732 1940
rect 9588 1244 9640 1250
rect 9588 1186 9640 1192
rect 9876 842 9904 2886
rect 9968 2610 9996 3362
rect 10152 3358 10180 4042
rect 10428 3494 10456 4382
rect 10488 4340 10784 4360
rect 10544 4338 10568 4340
rect 10624 4338 10648 4340
rect 10704 4338 10728 4340
rect 10566 4286 10568 4338
rect 10630 4286 10642 4338
rect 10704 4286 10706 4338
rect 10544 4284 10568 4286
rect 10624 4284 10648 4286
rect 10704 4284 10728 4286
rect 10488 4264 10784 4284
rect 10968 4032 11020 4038
rect 10968 3974 11020 3980
rect 10980 3902 11008 3974
rect 11060 3964 11112 3970
rect 11060 3906 11112 3912
rect 10968 3896 11020 3902
rect 10968 3838 11020 3844
rect 10416 3488 10468 3494
rect 10416 3430 10468 3436
rect 10140 3352 10192 3358
rect 10140 3294 10192 3300
rect 10488 3252 10784 3272
rect 10544 3250 10568 3252
rect 10624 3250 10648 3252
rect 10704 3250 10728 3252
rect 10566 3198 10568 3250
rect 10630 3198 10642 3250
rect 10704 3198 10706 3250
rect 10544 3196 10568 3198
rect 10624 3196 10648 3198
rect 10704 3196 10728 3198
rect 10488 3176 10784 3196
rect 10876 3080 10928 3086
rect 10876 3022 10928 3028
rect 10888 2814 10916 3022
rect 10980 2950 11008 3838
rect 11072 3494 11100 3906
rect 11060 3488 11112 3494
rect 11060 3430 11112 3436
rect 11164 3154 11192 4450
rect 11336 3692 11388 3698
rect 11336 3634 11388 3640
rect 11244 3624 11296 3630
rect 11244 3566 11296 3572
rect 11152 3148 11204 3154
rect 11152 3090 11204 3096
rect 11256 3018 11284 3566
rect 11244 3012 11296 3018
rect 11244 2954 11296 2960
rect 10968 2944 11020 2950
rect 10968 2886 11020 2892
rect 10876 2808 10928 2814
rect 11060 2808 11112 2814
rect 10928 2756 11008 2762
rect 10876 2750 11008 2756
rect 11060 2750 11112 2756
rect 11152 2808 11204 2814
rect 11152 2750 11204 2756
rect 10888 2734 11008 2750
rect 9956 2604 10008 2610
rect 9956 2546 10008 2552
rect 9968 1862 9996 2546
rect 10980 2338 11008 2734
rect 11072 2474 11100 2750
rect 11060 2468 11112 2474
rect 11060 2410 11112 2416
rect 10968 2332 11020 2338
rect 10968 2274 11020 2280
rect 10488 2164 10784 2184
rect 10544 2162 10568 2164
rect 10624 2162 10648 2164
rect 10704 2162 10728 2164
rect 10566 2110 10568 2162
rect 10630 2110 10642 2162
rect 10704 2110 10706 2162
rect 10544 2108 10568 2110
rect 10624 2108 10648 2110
rect 10704 2108 10728 2110
rect 10488 2088 10784 2108
rect 11164 1930 11192 2750
rect 11256 2406 11284 2954
rect 11348 2814 11376 3634
rect 11428 3420 11480 3426
rect 11428 3362 11480 3368
rect 11440 3018 11468 3362
rect 11428 3012 11480 3018
rect 11428 2954 11480 2960
rect 11336 2808 11388 2814
rect 11336 2750 11388 2756
rect 11532 2734 11560 6406
rect 11716 6282 11744 6558
rect 11704 6276 11756 6282
rect 11704 6218 11756 6224
rect 11612 6140 11664 6146
rect 11612 6082 11664 6088
rect 11624 5602 11652 6082
rect 11796 5800 11848 5806
rect 11796 5742 11848 5748
rect 11612 5596 11664 5602
rect 11612 5538 11664 5544
rect 11624 4106 11652 5538
rect 11808 5233 11836 5742
rect 11794 5224 11850 5233
rect 11794 5159 11796 5168
rect 11848 5159 11850 5168
rect 11796 5130 11848 5136
rect 11808 5099 11836 5130
rect 11796 4576 11848 4582
rect 11796 4518 11848 4524
rect 11704 4508 11756 4514
rect 11704 4450 11756 4456
rect 11612 4100 11664 4106
rect 11612 4042 11664 4048
rect 11624 3494 11652 4042
rect 11612 3488 11664 3494
rect 11612 3430 11664 3436
rect 11624 3154 11652 3430
rect 11612 3148 11664 3154
rect 11612 3090 11664 3096
rect 11716 3034 11744 4450
rect 11808 4242 11836 4518
rect 11796 4236 11848 4242
rect 11796 4178 11848 4184
rect 11796 3420 11848 3426
rect 11796 3362 11848 3368
rect 11440 2706 11560 2734
rect 11624 3006 11744 3034
rect 11244 2400 11296 2406
rect 11244 2342 11296 2348
rect 11244 2264 11296 2270
rect 11244 2206 11296 2212
rect 11152 1924 11204 1930
rect 11152 1866 11204 1872
rect 9956 1856 10008 1862
rect 9956 1798 10008 1804
rect 11152 1720 11204 1726
rect 11152 1662 11204 1668
rect 10488 1076 10784 1096
rect 10544 1074 10568 1076
rect 10624 1074 10648 1076
rect 10704 1074 10728 1076
rect 10566 1022 10568 1074
rect 10630 1022 10642 1074
rect 10704 1022 10706 1074
rect 10544 1020 10568 1022
rect 10624 1020 10648 1022
rect 10704 1020 10728 1022
rect 10488 1000 10784 1020
rect 9496 836 9548 842
rect 9416 796 9496 824
rect 9312 778 9364 784
rect 9496 778 9548 784
rect 9864 836 9916 842
rect 9864 778 9916 784
rect 9036 768 9088 774
rect 9036 710 9088 716
rect 8944 700 8996 706
rect 8944 642 8996 648
rect 10876 700 10928 706
rect 10876 642 10928 648
rect 7852 532 8148 552
rect 7908 530 7932 532
rect 7988 530 8012 532
rect 8068 530 8092 532
rect 7930 478 7932 530
rect 7994 478 8006 530
rect 8068 478 8070 530
rect 7908 476 7932 478
rect 7988 476 8012 478
rect 8068 476 8092 478
rect 7852 456 8148 476
rect 8956 160 8984 642
rect 10140 632 10192 638
rect 10140 574 10192 580
rect 10152 434 10180 574
rect 10140 428 10192 434
rect 10140 370 10192 376
rect 10888 160 10916 642
rect 11164 298 11192 1662
rect 11256 1386 11284 2206
rect 11244 1380 11296 1386
rect 11244 1322 11296 1328
rect 11440 1318 11468 2706
rect 11624 2066 11652 3006
rect 11704 2944 11756 2950
rect 11704 2886 11756 2892
rect 11716 2474 11744 2886
rect 11704 2468 11756 2474
rect 11704 2410 11756 2416
rect 11808 2354 11836 3362
rect 11716 2338 11836 2354
rect 11704 2332 11836 2338
rect 11756 2326 11836 2332
rect 11704 2274 11756 2280
rect 11612 2060 11664 2066
rect 11612 2002 11664 2008
rect 11716 1522 11744 2274
rect 11704 1516 11756 1522
rect 11704 1458 11756 1464
rect 11900 1318 11928 9822
rect 12072 9472 12124 9478
rect 12072 9414 12124 9420
rect 12084 8866 12112 9414
rect 12072 8860 12124 8866
rect 12072 8802 12124 8808
rect 11980 8792 12032 8798
rect 11980 8734 12032 8740
rect 11992 8526 12020 8734
rect 11980 8520 12032 8526
rect 11980 8462 12032 8468
rect 11992 7914 12020 8462
rect 11980 7908 12032 7914
rect 11980 7850 12032 7856
rect 12084 6826 12112 8802
rect 12072 6820 12124 6826
rect 12072 6762 12124 6768
rect 12072 4100 12124 4106
rect 12072 4042 12124 4048
rect 12084 3698 12112 4042
rect 12072 3692 12124 3698
rect 12072 3634 12124 3640
rect 12176 2734 12204 10094
rect 12256 9540 12308 9546
rect 12440 9540 12492 9546
rect 12308 9500 12388 9528
rect 12256 9482 12308 9488
rect 12256 9336 12308 9342
rect 12256 9278 12308 9284
rect 12268 9002 12296 9278
rect 12256 8996 12308 9002
rect 12256 8938 12308 8944
rect 12268 8458 12296 8938
rect 12256 8452 12308 8458
rect 12256 8394 12308 8400
rect 12268 7982 12296 8394
rect 12256 7976 12308 7982
rect 12256 7918 12308 7924
rect 12256 6276 12308 6282
rect 12256 6218 12308 6224
rect 12268 5670 12296 6218
rect 12256 5664 12308 5670
rect 12256 5606 12308 5612
rect 12360 5126 12388 9500
rect 12440 9482 12492 9488
rect 12624 9540 12676 9546
rect 12624 9482 12676 9488
rect 12452 5806 12480 9482
rect 12532 9336 12584 9342
rect 12532 9278 12584 9284
rect 12544 7846 12572 9278
rect 12532 7840 12584 7846
rect 12532 7782 12584 7788
rect 12636 6214 12664 9482
rect 12728 8458 12756 10366
rect 12820 10090 12848 12746
rect 13124 12500 13420 12520
rect 13180 12498 13204 12500
rect 13260 12498 13284 12500
rect 13340 12498 13364 12500
rect 13202 12446 13204 12498
rect 13266 12446 13278 12498
rect 13340 12446 13342 12498
rect 13180 12444 13204 12446
rect 13260 12444 13284 12446
rect 13340 12444 13364 12446
rect 13124 12424 13420 12444
rect 14200 11858 14228 12746
rect 14280 12124 14332 12130
rect 14280 12066 14332 12072
rect 14188 11852 14240 11858
rect 14188 11794 14240 11800
rect 14004 11716 14056 11722
rect 14004 11658 14056 11664
rect 13124 11412 13420 11432
rect 13180 11410 13204 11412
rect 13260 11410 13284 11412
rect 13340 11410 13364 11412
rect 13202 11358 13204 11410
rect 13266 11358 13278 11410
rect 13340 11358 13342 11410
rect 13180 11356 13204 11358
rect 13260 11356 13284 11358
rect 13340 11356 13364 11358
rect 13124 11336 13420 11356
rect 13820 11104 13872 11110
rect 13820 11046 13872 11052
rect 13124 10324 13420 10344
rect 13180 10322 13204 10324
rect 13260 10322 13284 10324
rect 13340 10322 13364 10324
rect 13202 10270 13204 10322
rect 13266 10270 13278 10322
rect 13340 10270 13342 10322
rect 13180 10268 13204 10270
rect 13260 10268 13284 10270
rect 13340 10268 13364 10270
rect 13124 10248 13420 10268
rect 12808 10084 12860 10090
rect 12808 10026 12860 10032
rect 12808 9880 12860 9886
rect 12808 9822 12860 9828
rect 12716 8452 12768 8458
rect 12716 8394 12768 8400
rect 12728 7370 12756 8394
rect 12716 7364 12768 7370
rect 12716 7306 12768 7312
rect 12624 6208 12676 6214
rect 12624 6150 12676 6156
rect 12440 5800 12492 5806
rect 12440 5742 12492 5748
rect 12440 5256 12492 5262
rect 12440 5198 12492 5204
rect 12348 5120 12400 5126
rect 12348 5062 12400 5068
rect 12348 4984 12400 4990
rect 12348 4926 12400 4932
rect 12360 4582 12388 4926
rect 12348 4576 12400 4582
rect 12348 4518 12400 4524
rect 12348 4032 12400 4038
rect 12348 3974 12400 3980
rect 12256 3896 12308 3902
rect 12256 3838 12308 3844
rect 12268 3086 12296 3838
rect 12360 3442 12388 3974
rect 12452 3630 12480 5198
rect 12532 5120 12584 5126
rect 12532 5062 12584 5068
rect 12544 4106 12572 5062
rect 12624 4576 12676 4582
rect 12624 4518 12676 4524
rect 12636 4242 12664 4518
rect 12716 4508 12768 4514
rect 12716 4450 12768 4456
rect 12624 4236 12676 4242
rect 12624 4178 12676 4184
rect 12532 4100 12584 4106
rect 12532 4042 12584 4048
rect 12728 3952 12756 4450
rect 12544 3924 12756 3952
rect 12440 3624 12492 3630
rect 12440 3566 12492 3572
rect 12544 3494 12572 3924
rect 12624 3624 12676 3630
rect 12624 3566 12676 3572
rect 12532 3488 12584 3494
rect 12360 3414 12480 3442
rect 12532 3430 12584 3436
rect 12256 3080 12308 3086
rect 12256 3022 12308 3028
rect 12452 2950 12480 3414
rect 12532 3352 12584 3358
rect 12532 3294 12584 3300
rect 12440 2944 12492 2950
rect 12440 2886 12492 2892
rect 12176 2706 12296 2734
rect 11428 1312 11480 1318
rect 11428 1254 11480 1260
rect 11888 1312 11940 1318
rect 11888 1254 11940 1260
rect 11244 1176 11296 1182
rect 11244 1118 11296 1124
rect 11256 366 11284 1118
rect 12268 910 12296 2706
rect 12348 1856 12400 1862
rect 12452 1810 12480 2886
rect 12544 2610 12572 3294
rect 12532 2604 12584 2610
rect 12532 2546 12584 2552
rect 12636 2406 12664 3566
rect 12728 3358 12756 3924
rect 12716 3352 12768 3358
rect 12716 3294 12768 3300
rect 12624 2400 12676 2406
rect 12624 2342 12676 2348
rect 12624 2264 12676 2270
rect 12624 2206 12676 2212
rect 12636 1998 12664 2206
rect 12624 1992 12676 1998
rect 12624 1934 12676 1940
rect 12400 1804 12480 1810
rect 12348 1798 12480 1804
rect 12360 1782 12480 1798
rect 12452 1454 12480 1782
rect 12440 1448 12492 1454
rect 12440 1390 12492 1396
rect 12820 910 12848 9822
rect 13636 9540 13688 9546
rect 13636 9482 13688 9488
rect 13124 9236 13420 9256
rect 13180 9234 13204 9236
rect 13260 9234 13284 9236
rect 13340 9234 13364 9236
rect 13202 9182 13204 9234
rect 13266 9182 13278 9234
rect 13340 9182 13342 9234
rect 13180 9180 13204 9182
rect 13260 9180 13284 9182
rect 13340 9180 13364 9182
rect 13124 9160 13420 9180
rect 13452 8928 13504 8934
rect 13452 8870 13504 8876
rect 13464 8526 13492 8870
rect 13452 8520 13504 8526
rect 13452 8462 13504 8468
rect 12900 8384 12952 8390
rect 12900 8326 12952 8332
rect 12912 8050 12940 8326
rect 13124 8148 13420 8168
rect 13180 8146 13204 8148
rect 13260 8146 13284 8148
rect 13340 8146 13364 8148
rect 13202 8094 13204 8146
rect 13266 8094 13278 8146
rect 13340 8094 13342 8146
rect 13180 8092 13204 8094
rect 13260 8092 13284 8094
rect 13340 8092 13364 8094
rect 13124 8072 13420 8092
rect 12900 8044 12952 8050
rect 12900 7986 12952 7992
rect 13464 7438 13492 8462
rect 13452 7432 13504 7438
rect 13452 7374 13504 7380
rect 12992 7296 13044 7302
rect 12992 7238 13044 7244
rect 12900 6616 12952 6622
rect 12900 6558 12952 6564
rect 12912 6350 12940 6558
rect 13004 6418 13032 7238
rect 13124 7060 13420 7080
rect 13180 7058 13204 7060
rect 13260 7058 13284 7060
rect 13340 7058 13364 7060
rect 13202 7006 13204 7058
rect 13266 7006 13278 7058
rect 13340 7006 13342 7058
rect 13180 7004 13204 7006
rect 13260 7004 13284 7006
rect 13340 7004 13364 7006
rect 13124 6984 13420 7004
rect 12992 6412 13044 6418
rect 12992 6354 13044 6360
rect 12900 6344 12952 6350
rect 12900 6286 12952 6292
rect 13124 5972 13420 5992
rect 13180 5970 13204 5972
rect 13260 5970 13284 5972
rect 13340 5970 13364 5972
rect 13202 5918 13204 5970
rect 13266 5918 13278 5970
rect 13340 5918 13342 5970
rect 13180 5916 13204 5918
rect 13260 5916 13284 5918
rect 13340 5916 13364 5918
rect 13124 5896 13420 5916
rect 13464 5262 13492 7374
rect 13648 6690 13676 9482
rect 13728 7704 13780 7710
rect 13728 7646 13780 7652
rect 13740 6826 13768 7646
rect 13728 6820 13780 6826
rect 13728 6762 13780 6768
rect 13636 6684 13688 6690
rect 13636 6626 13688 6632
rect 13544 6140 13596 6146
rect 13544 6082 13596 6088
rect 13452 5256 13504 5262
rect 13452 5198 13504 5204
rect 13124 4884 13420 4904
rect 13180 4882 13204 4884
rect 13260 4882 13284 4884
rect 13340 4882 13364 4884
rect 13202 4830 13204 4882
rect 13266 4830 13278 4882
rect 13340 4830 13342 4882
rect 13180 4828 13204 4830
rect 13260 4828 13284 4830
rect 13340 4828 13364 4830
rect 13124 4808 13420 4828
rect 13464 4174 13492 5198
rect 13556 4786 13584 6082
rect 13740 5670 13768 6762
rect 13728 5664 13780 5670
rect 13728 5606 13780 5612
rect 13544 4780 13596 4786
rect 13544 4722 13596 4728
rect 13636 4712 13688 4718
rect 13636 4654 13688 4660
rect 13452 4168 13504 4174
rect 13452 4110 13504 4116
rect 13124 3796 13420 3816
rect 13180 3794 13204 3796
rect 13260 3794 13284 3796
rect 13340 3794 13364 3796
rect 13202 3742 13204 3794
rect 13266 3742 13278 3794
rect 13340 3742 13342 3794
rect 13180 3740 13204 3742
rect 13260 3740 13284 3742
rect 13340 3740 13364 3742
rect 13124 3720 13420 3740
rect 12900 3148 12952 3154
rect 12900 3090 12952 3096
rect 12912 2406 12940 3090
rect 13464 3086 13492 4110
rect 13648 3562 13676 4654
rect 13832 3630 13860 11046
rect 13912 9540 13964 9546
rect 13912 9482 13964 9488
rect 13924 8254 13952 9482
rect 13912 8248 13964 8254
rect 13912 8190 13964 8196
rect 13924 7846 13952 8190
rect 13912 7840 13964 7846
rect 13912 7782 13964 7788
rect 13912 7160 13964 7166
rect 13912 7102 13964 7108
rect 13924 6758 13952 7102
rect 13912 6752 13964 6758
rect 13912 6694 13964 6700
rect 13924 6350 13952 6694
rect 13912 6344 13964 6350
rect 13912 6286 13964 6292
rect 14016 6162 14044 11658
rect 14292 11314 14320 12066
rect 14280 11308 14332 11314
rect 14280 11250 14332 11256
rect 14740 10016 14792 10022
rect 14740 9958 14792 9964
rect 14648 9540 14700 9546
rect 14648 9482 14700 9488
rect 14464 9404 14516 9410
rect 14464 9346 14516 9352
rect 14096 9336 14148 9342
rect 14096 9278 14148 9284
rect 14108 8934 14136 9278
rect 14096 8928 14148 8934
rect 14096 8870 14148 8876
rect 14108 7846 14136 8870
rect 14188 8860 14240 8866
rect 14188 8802 14240 8808
rect 14096 7840 14148 7846
rect 14096 7782 14148 7788
rect 14096 7704 14148 7710
rect 14096 7646 14148 7652
rect 14108 6894 14136 7646
rect 14096 6888 14148 6894
rect 14096 6830 14148 6836
rect 14200 6826 14228 8802
rect 14280 8792 14332 8798
rect 14280 8734 14332 8740
rect 14188 6820 14240 6826
rect 14188 6762 14240 6768
rect 14016 6134 14136 6162
rect 14004 6072 14056 6078
rect 14004 6014 14056 6020
rect 14016 4038 14044 6014
rect 14004 4032 14056 4038
rect 14004 3974 14056 3980
rect 13820 3624 13872 3630
rect 13820 3566 13872 3572
rect 13636 3556 13688 3562
rect 13636 3498 13688 3504
rect 13728 3420 13780 3426
rect 13728 3362 13780 3368
rect 13452 3080 13504 3086
rect 13504 3040 13584 3068
rect 13452 3022 13504 3028
rect 13124 2708 13420 2728
rect 13180 2706 13204 2708
rect 13260 2706 13284 2708
rect 13340 2706 13364 2708
rect 13202 2654 13204 2706
rect 13266 2654 13278 2706
rect 13340 2654 13342 2706
rect 13180 2652 13204 2654
rect 13260 2652 13284 2654
rect 13340 2652 13364 2654
rect 13124 2632 13420 2652
rect 12900 2400 12952 2406
rect 12900 2342 12952 2348
rect 13556 2066 13584 3040
rect 13740 2406 13768 3362
rect 13832 2734 13860 3566
rect 14108 2734 14136 6134
rect 14200 5874 14228 6762
rect 14292 6758 14320 8734
rect 14372 7908 14424 7914
rect 14372 7850 14424 7856
rect 14280 6752 14332 6758
rect 14280 6694 14332 6700
rect 14384 6418 14412 7850
rect 14372 6412 14424 6418
rect 14372 6354 14424 6360
rect 14188 5868 14240 5874
rect 14188 5810 14240 5816
rect 14188 5596 14240 5602
rect 14188 5538 14240 5544
rect 14200 5330 14228 5538
rect 14188 5324 14240 5330
rect 14188 5266 14240 5272
rect 14188 4508 14240 4514
rect 14188 4450 14240 4456
rect 14200 4242 14228 4450
rect 14476 4446 14504 9346
rect 14556 7296 14608 7302
rect 14556 7238 14608 7244
rect 14464 4440 14516 4446
rect 14464 4382 14516 4388
rect 14188 4236 14240 4242
rect 14188 4178 14240 4184
rect 14188 3420 14240 3426
rect 14188 3362 14240 3368
rect 14200 3154 14228 3362
rect 14188 3148 14240 3154
rect 14188 3090 14240 3096
rect 13832 2706 13952 2734
rect 13728 2400 13780 2406
rect 13728 2342 13780 2348
rect 13544 2060 13596 2066
rect 13544 2002 13596 2008
rect 13740 1794 13768 2342
rect 13924 1998 13952 2706
rect 14016 2706 14136 2734
rect 14016 2610 14044 2706
rect 14004 2604 14056 2610
rect 14004 2546 14056 2552
rect 13912 1992 13964 1998
rect 13912 1934 13964 1940
rect 13728 1788 13780 1794
rect 13728 1730 13780 1736
rect 13124 1620 13420 1640
rect 13180 1618 13204 1620
rect 13260 1618 13284 1620
rect 13340 1618 13364 1620
rect 13202 1566 13204 1618
rect 13266 1566 13278 1618
rect 13340 1566 13342 1618
rect 13180 1564 13204 1566
rect 13260 1564 13284 1566
rect 13340 1564 13364 1566
rect 13124 1544 13420 1564
rect 14016 910 14044 2546
rect 14568 1250 14596 7238
rect 14660 4786 14688 9482
rect 14752 5330 14780 9958
rect 14844 9410 14872 12746
rect 15106 12160 15162 12169
rect 15106 12095 15108 12104
rect 15160 12095 15162 12104
rect 15108 12066 15160 12072
rect 15106 11072 15162 11081
rect 14924 11036 14976 11042
rect 15106 11007 15108 11016
rect 14924 10978 14976 10984
rect 15160 11007 15162 11016
rect 15108 10978 15160 10984
rect 14936 10226 14964 10978
rect 15568 10628 15620 10634
rect 15568 10570 15620 10576
rect 15016 10424 15068 10430
rect 15016 10366 15068 10372
rect 14924 10220 14976 10226
rect 14924 10162 14976 10168
rect 14924 9948 14976 9954
rect 14924 9890 14976 9896
rect 14936 9682 14964 9890
rect 14924 9676 14976 9682
rect 14924 9618 14976 9624
rect 14832 9404 14884 9410
rect 14832 9346 14884 9352
rect 14924 8860 14976 8866
rect 14924 8802 14976 8808
rect 14740 5324 14792 5330
rect 14740 5266 14792 5272
rect 14832 5256 14884 5262
rect 14832 5198 14884 5204
rect 14740 5188 14792 5194
rect 14740 5130 14792 5136
rect 14648 4780 14700 4786
rect 14648 4722 14700 4728
rect 14660 4174 14688 4722
rect 14752 4582 14780 5130
rect 14844 4582 14872 5198
rect 14740 4576 14792 4582
rect 14740 4518 14792 4524
rect 14832 4576 14884 4582
rect 14832 4518 14884 4524
rect 14832 4440 14884 4446
rect 14832 4382 14884 4388
rect 14648 4168 14700 4174
rect 14648 4110 14700 4116
rect 14844 1318 14872 4382
rect 14936 2610 14964 8802
rect 15028 6758 15056 10366
rect 15108 9948 15160 9954
rect 15108 9890 15160 9896
rect 15120 9857 15148 9890
rect 15106 9848 15162 9857
rect 15106 9783 15162 9792
rect 15108 8860 15160 8866
rect 15108 8802 15160 8808
rect 15120 8769 15148 8802
rect 15106 8760 15162 8769
rect 15106 8695 15162 8704
rect 15580 7545 15608 10570
rect 15566 7536 15622 7545
rect 15566 7471 15622 7480
rect 15016 6752 15068 6758
rect 15016 6694 15068 6700
rect 15028 6350 15056 6694
rect 15016 6344 15068 6350
rect 15016 6286 15068 6292
rect 15198 6312 15254 6321
rect 15108 6276 15160 6282
rect 15198 6247 15254 6256
rect 15108 6218 15160 6224
rect 15120 5738 15148 6218
rect 15108 5732 15160 5738
rect 15108 5674 15160 5680
rect 15108 5596 15160 5602
rect 15108 5538 15160 5544
rect 15016 5528 15068 5534
rect 15016 5470 15068 5476
rect 15028 5233 15056 5470
rect 15014 5224 15070 5233
rect 15014 5159 15070 5168
rect 15016 4576 15068 4582
rect 15016 4518 15068 4524
rect 15028 3494 15056 4518
rect 15016 3488 15068 3494
rect 15016 3430 15068 3436
rect 15120 3306 15148 5538
rect 15028 3278 15148 3306
rect 14924 2604 14976 2610
rect 14924 2546 14976 2552
rect 15028 2406 15056 3278
rect 15106 2912 15162 2921
rect 15106 2847 15108 2856
rect 15160 2847 15162 2856
rect 15108 2818 15160 2824
rect 15016 2400 15068 2406
rect 15016 2342 15068 2348
rect 15108 1788 15160 1794
rect 15108 1730 15160 1736
rect 15120 1697 15148 1730
rect 15106 1688 15162 1697
rect 15106 1623 15162 1632
rect 14832 1312 14884 1318
rect 14832 1254 14884 1260
rect 14556 1244 14608 1250
rect 14556 1186 14608 1192
rect 15212 1182 15240 6247
rect 15292 5256 15344 5262
rect 15292 5198 15344 5204
rect 15304 3086 15332 5198
rect 15476 4032 15528 4038
rect 15474 4000 15476 4009
rect 15528 4000 15530 4009
rect 15474 3935 15530 3944
rect 15292 3080 15344 3086
rect 15292 3022 15344 3028
rect 14924 1176 14976 1182
rect 14924 1118 14976 1124
rect 15200 1176 15252 1182
rect 15200 1118 15252 1124
rect 14936 910 14964 1118
rect 12256 904 12308 910
rect 12256 846 12308 852
rect 12808 904 12860 910
rect 12808 846 12860 852
rect 14004 904 14056 910
rect 14004 846 14056 852
rect 14924 904 14976 910
rect 14924 846 14976 852
rect 14372 700 14424 706
rect 14372 642 14424 648
rect 12900 632 12952 638
rect 14384 609 14412 642
rect 14924 632 14976 638
rect 12900 574 12952 580
rect 14370 600 14426 609
rect 11244 360 11296 366
rect 11244 302 11296 308
rect 11152 292 11204 298
rect 11152 234 11204 240
rect 12912 160 12940 574
rect 13124 532 13420 552
rect 14924 574 14976 580
rect 14370 535 14426 544
rect 13180 530 13204 532
rect 13260 530 13284 532
rect 13340 530 13364 532
rect 13202 478 13204 530
rect 13266 478 13278 530
rect 13340 478 13342 530
rect 13180 476 13204 478
rect 13260 476 13284 478
rect 13340 476 13364 478
rect 13124 456 13420 476
rect 14936 160 14964 574
rect 938 -40 994 160
rect 2870 -40 2926 160
rect 4894 -40 4950 160
rect 6918 -40 6974 160
rect 8942 -40 8998 160
rect 10874 -40 10930 160
rect 12898 -40 12954 160
rect 14922 -40 14978 160
<< via2 >>
rect 3974 13328 4030 13384
rect 5216 13042 5272 13044
rect 5296 13042 5352 13044
rect 5376 13042 5432 13044
rect 5456 13042 5512 13044
rect 5216 12990 5242 13042
rect 5242 12990 5272 13042
rect 5296 12990 5306 13042
rect 5306 12990 5352 13042
rect 5376 12990 5422 13042
rect 5422 12990 5432 13042
rect 5456 12990 5486 13042
rect 5486 12990 5512 13042
rect 5216 12988 5272 12990
rect 5296 12988 5352 12990
rect 5376 12988 5432 12990
rect 5456 12988 5512 12990
rect 10488 13042 10544 13044
rect 10568 13042 10624 13044
rect 10648 13042 10704 13044
rect 10728 13042 10784 13044
rect 10488 12990 10514 13042
rect 10514 12990 10544 13042
rect 10568 12990 10578 13042
rect 10578 12990 10624 13042
rect 10648 12990 10694 13042
rect 10694 12990 10704 13042
rect 10728 12990 10758 13042
rect 10758 12990 10784 13042
rect 10488 12988 10544 12990
rect 10568 12988 10624 12990
rect 10648 12988 10704 12990
rect 10728 12988 10784 12990
rect 14370 13328 14426 13384
rect 754 11288 810 11344
rect 754 10336 810 10392
rect 754 9420 756 9440
rect 756 9420 808 9440
rect 808 9420 810 9440
rect 754 9384 810 9420
rect 754 8296 810 8352
rect 1766 12376 1822 12432
rect 2580 12498 2636 12500
rect 2660 12498 2716 12500
rect 2740 12498 2796 12500
rect 2820 12498 2876 12500
rect 2580 12446 2606 12498
rect 2606 12446 2636 12498
rect 2660 12446 2670 12498
rect 2670 12446 2716 12498
rect 2740 12446 2786 12498
rect 2786 12446 2796 12498
rect 2820 12446 2850 12498
rect 2850 12446 2876 12498
rect 2580 12444 2636 12446
rect 2660 12444 2716 12446
rect 2740 12444 2796 12446
rect 2820 12444 2876 12446
rect 478 7344 534 7400
rect 2580 11410 2636 11412
rect 2660 11410 2716 11412
rect 2740 11410 2796 11412
rect 2820 11410 2876 11412
rect 2580 11358 2606 11410
rect 2606 11358 2636 11410
rect 2660 11358 2670 11410
rect 2670 11358 2716 11410
rect 2740 11358 2786 11410
rect 2786 11358 2796 11410
rect 2820 11358 2850 11410
rect 2850 11358 2876 11410
rect 2580 11356 2636 11358
rect 2660 11356 2716 11358
rect 2740 11356 2796 11358
rect 2820 11356 2876 11358
rect 2580 10322 2636 10324
rect 2660 10322 2716 10324
rect 2740 10322 2796 10324
rect 2820 10322 2876 10324
rect 2580 10270 2606 10322
rect 2606 10270 2636 10322
rect 2660 10270 2670 10322
rect 2670 10270 2716 10322
rect 2740 10270 2786 10322
rect 2786 10270 2796 10322
rect 2820 10270 2850 10322
rect 2850 10270 2876 10322
rect 2580 10268 2636 10270
rect 2660 10268 2716 10270
rect 2740 10268 2796 10270
rect 2820 10268 2876 10270
rect 754 6392 810 6448
rect 754 5304 810 5360
rect 846 4352 902 4408
rect 846 2332 902 2368
rect 846 2312 848 2332
rect 848 2312 900 2332
rect 900 2312 902 2332
rect 2580 9234 2636 9236
rect 2660 9234 2716 9236
rect 2740 9234 2796 9236
rect 2820 9234 2876 9236
rect 2580 9182 2606 9234
rect 2606 9182 2636 9234
rect 2660 9182 2670 9234
rect 2670 9182 2716 9234
rect 2740 9182 2786 9234
rect 2786 9182 2796 9234
rect 2820 9182 2850 9234
rect 2850 9182 2876 9234
rect 2580 9180 2636 9182
rect 2660 9180 2716 9182
rect 2740 9180 2796 9182
rect 2820 9180 2876 9182
rect 2580 8146 2636 8148
rect 2660 8146 2716 8148
rect 2740 8146 2796 8148
rect 2820 8146 2876 8148
rect 2580 8094 2606 8146
rect 2606 8094 2636 8146
rect 2660 8094 2670 8146
rect 2670 8094 2716 8146
rect 2740 8094 2786 8146
rect 2786 8094 2796 8146
rect 2820 8094 2850 8146
rect 2850 8094 2876 8146
rect 2580 8092 2636 8094
rect 2660 8092 2716 8094
rect 2740 8092 2796 8094
rect 2820 8092 2876 8094
rect 4066 11052 4068 11072
rect 4068 11052 4120 11072
rect 4120 11052 4122 11072
rect 4066 11016 4122 11052
rect 4434 10608 4490 10664
rect 4710 11016 4766 11072
rect 4434 9384 4490 9440
rect 2580 7058 2636 7060
rect 2660 7058 2716 7060
rect 2740 7058 2796 7060
rect 2820 7058 2876 7060
rect 2580 7006 2606 7058
rect 2606 7006 2636 7058
rect 2660 7006 2670 7058
rect 2670 7006 2716 7058
rect 2740 7006 2786 7058
rect 2786 7006 2796 7058
rect 2820 7006 2850 7058
rect 2850 7006 2876 7058
rect 2580 7004 2636 7006
rect 2660 7004 2716 7006
rect 2740 7004 2796 7006
rect 2820 7004 2876 7006
rect 2580 5970 2636 5972
rect 2660 5970 2716 5972
rect 2740 5970 2796 5972
rect 2820 5970 2876 5972
rect 2580 5918 2606 5970
rect 2606 5918 2636 5970
rect 2660 5918 2670 5970
rect 2670 5918 2716 5970
rect 2740 5918 2786 5970
rect 2786 5918 2796 5970
rect 2820 5918 2850 5970
rect 2850 5918 2876 5970
rect 2580 5916 2636 5918
rect 2660 5916 2716 5918
rect 2740 5916 2796 5918
rect 2820 5916 2876 5918
rect 2580 4882 2636 4884
rect 2660 4882 2716 4884
rect 2740 4882 2796 4884
rect 2820 4882 2876 4884
rect 2580 4830 2606 4882
rect 2606 4830 2636 4882
rect 2660 4830 2670 4882
rect 2670 4830 2716 4882
rect 2740 4830 2786 4882
rect 2786 4830 2796 4882
rect 2820 4830 2850 4882
rect 2850 4830 2876 4882
rect 2580 4828 2636 4830
rect 2660 4828 2716 4830
rect 2740 4828 2796 4830
rect 2820 4828 2876 4830
rect 2580 3794 2636 3796
rect 2660 3794 2716 3796
rect 2740 3794 2796 3796
rect 2820 3794 2876 3796
rect 2580 3742 2606 3794
rect 2606 3742 2636 3794
rect 2660 3742 2670 3794
rect 2670 3742 2716 3794
rect 2740 3742 2786 3794
rect 2786 3742 2796 3794
rect 2820 3742 2850 3794
rect 2850 3742 2876 3794
rect 2580 3740 2636 3742
rect 2660 3740 2716 3742
rect 2740 3740 2796 3742
rect 2820 3740 2876 3742
rect 4526 6820 4582 6856
rect 4526 6800 4528 6820
rect 4528 6800 4580 6820
rect 4580 6800 4582 6820
rect 4066 3400 4122 3456
rect 2580 2706 2636 2708
rect 2660 2706 2716 2708
rect 2740 2706 2796 2708
rect 2820 2706 2876 2708
rect 2580 2654 2606 2706
rect 2606 2654 2636 2706
rect 2660 2654 2670 2706
rect 2670 2654 2716 2706
rect 2740 2654 2786 2706
rect 2786 2654 2796 2706
rect 2820 2654 2850 2706
rect 2850 2654 2876 2706
rect 2580 2652 2636 2654
rect 2660 2652 2716 2654
rect 2740 2652 2796 2654
rect 2820 2652 2876 2654
rect 2580 1618 2636 1620
rect 2660 1618 2716 1620
rect 2740 1618 2796 1620
rect 2820 1618 2876 1620
rect 2580 1566 2606 1618
rect 2606 1566 2636 1618
rect 2660 1566 2670 1618
rect 2670 1566 2716 1618
rect 2740 1566 2786 1618
rect 2786 1566 2796 1618
rect 2820 1566 2850 1618
rect 2850 1566 2876 1618
rect 2580 1564 2636 1566
rect 2660 1564 2716 1566
rect 2740 1564 2796 1566
rect 2820 1564 2876 1566
rect 3330 1396 3332 1416
rect 3332 1396 3384 1416
rect 3384 1396 3386 1416
rect 3330 1360 3386 1396
rect 2580 530 2636 532
rect 2660 530 2716 532
rect 2740 530 2796 532
rect 2820 530 2876 532
rect 2580 478 2606 530
rect 2606 478 2636 530
rect 2660 478 2670 530
rect 2670 478 2716 530
rect 2740 478 2786 530
rect 2786 478 2796 530
rect 2820 478 2850 530
rect 2850 478 2876 530
rect 2580 476 2636 478
rect 2660 476 2716 478
rect 2740 476 2796 478
rect 2820 476 2876 478
rect 5216 11954 5272 11956
rect 5296 11954 5352 11956
rect 5376 11954 5432 11956
rect 5456 11954 5512 11956
rect 5216 11902 5242 11954
rect 5242 11902 5272 11954
rect 5296 11902 5306 11954
rect 5306 11902 5352 11954
rect 5376 11902 5422 11954
rect 5422 11902 5432 11954
rect 5456 11902 5486 11954
rect 5486 11902 5512 11954
rect 5216 11900 5272 11902
rect 5296 11900 5352 11902
rect 5376 11900 5432 11902
rect 5456 11900 5512 11902
rect 5216 10866 5272 10868
rect 5296 10866 5352 10868
rect 5376 10866 5432 10868
rect 5456 10866 5512 10868
rect 5216 10814 5242 10866
rect 5242 10814 5272 10866
rect 5296 10814 5306 10866
rect 5306 10814 5352 10866
rect 5376 10814 5422 10866
rect 5422 10814 5432 10866
rect 5456 10814 5486 10866
rect 5486 10814 5512 10866
rect 5216 10812 5272 10814
rect 5296 10812 5352 10814
rect 5376 10812 5432 10814
rect 5456 10812 5512 10814
rect 5998 10200 6054 10256
rect 5216 9778 5272 9780
rect 5296 9778 5352 9780
rect 5376 9778 5432 9780
rect 5456 9778 5512 9780
rect 5216 9726 5242 9778
rect 5242 9726 5272 9778
rect 5296 9726 5306 9778
rect 5306 9726 5352 9778
rect 5376 9726 5422 9778
rect 5422 9726 5432 9778
rect 5456 9726 5486 9778
rect 5486 9726 5512 9778
rect 5216 9724 5272 9726
rect 5296 9724 5352 9726
rect 5376 9724 5432 9726
rect 5456 9724 5512 9726
rect 6274 10200 6330 10256
rect 5216 8690 5272 8692
rect 5296 8690 5352 8692
rect 5376 8690 5432 8692
rect 5456 8690 5512 8692
rect 5216 8638 5242 8690
rect 5242 8638 5272 8690
rect 5296 8638 5306 8690
rect 5306 8638 5352 8690
rect 5376 8638 5422 8690
rect 5422 8638 5432 8690
rect 5456 8638 5486 8690
rect 5486 8638 5512 8690
rect 5216 8636 5272 8638
rect 5296 8636 5352 8638
rect 5376 8636 5432 8638
rect 5456 8636 5512 8638
rect 5216 7602 5272 7604
rect 5296 7602 5352 7604
rect 5376 7602 5432 7604
rect 5456 7602 5512 7604
rect 5216 7550 5242 7602
rect 5242 7550 5272 7602
rect 5296 7550 5306 7602
rect 5306 7550 5352 7602
rect 5376 7550 5422 7602
rect 5422 7550 5432 7602
rect 5456 7550 5486 7602
rect 5486 7550 5512 7602
rect 5216 7548 5272 7550
rect 5296 7548 5352 7550
rect 5376 7548 5432 7550
rect 5456 7548 5512 7550
rect 5216 6514 5272 6516
rect 5296 6514 5352 6516
rect 5376 6514 5432 6516
rect 5456 6514 5512 6516
rect 5216 6462 5242 6514
rect 5242 6462 5272 6514
rect 5296 6462 5306 6514
rect 5306 6462 5352 6514
rect 5376 6462 5422 6514
rect 5422 6462 5432 6514
rect 5456 6462 5486 6514
rect 5486 6462 5512 6514
rect 5216 6460 5272 6462
rect 5296 6460 5352 6462
rect 5376 6460 5432 6462
rect 5456 6460 5512 6462
rect 5216 5426 5272 5428
rect 5296 5426 5352 5428
rect 5376 5426 5432 5428
rect 5456 5426 5512 5428
rect 5216 5374 5242 5426
rect 5242 5374 5272 5426
rect 5296 5374 5306 5426
rect 5306 5374 5352 5426
rect 5376 5374 5422 5426
rect 5422 5374 5432 5426
rect 5456 5374 5486 5426
rect 5486 5374 5512 5426
rect 5216 5372 5272 5374
rect 5296 5372 5352 5374
rect 5376 5372 5432 5374
rect 5456 5372 5512 5374
rect 5630 6664 5686 6720
rect 5998 6800 6054 6856
rect 5216 4338 5272 4340
rect 5296 4338 5352 4340
rect 5376 4338 5432 4340
rect 5456 4338 5512 4340
rect 5216 4286 5242 4338
rect 5242 4286 5272 4338
rect 5296 4286 5306 4338
rect 5306 4286 5352 4338
rect 5376 4286 5422 4338
rect 5422 4286 5432 4338
rect 5456 4286 5486 4338
rect 5486 4286 5512 4338
rect 5216 4284 5272 4286
rect 5296 4284 5352 4286
rect 5376 4284 5432 4286
rect 5456 4284 5512 4286
rect 6458 6700 6460 6720
rect 6460 6700 6512 6720
rect 6512 6700 6514 6720
rect 6458 6664 6514 6700
rect 6642 9420 6644 9440
rect 6644 9420 6696 9440
rect 6696 9420 6698 9440
rect 6642 9384 6698 9420
rect 7010 9520 7066 9576
rect 7102 9404 7158 9440
rect 7102 9384 7104 9404
rect 7104 9384 7156 9404
rect 7156 9384 7158 9404
rect 6642 6836 6644 6856
rect 6644 6836 6696 6856
rect 6696 6836 6698 6856
rect 6642 6800 6698 6836
rect 5216 3250 5272 3252
rect 5296 3250 5352 3252
rect 5376 3250 5432 3252
rect 5456 3250 5512 3252
rect 5216 3198 5242 3250
rect 5242 3198 5272 3250
rect 5296 3198 5306 3250
rect 5306 3198 5352 3250
rect 5376 3198 5422 3250
rect 5422 3198 5432 3250
rect 5456 3198 5486 3250
rect 5486 3198 5512 3250
rect 5216 3196 5272 3198
rect 5296 3196 5352 3198
rect 5376 3196 5432 3198
rect 5456 3196 5512 3198
rect 3514 716 3516 736
rect 3516 716 3568 736
rect 3568 716 3570 736
rect 3514 680 3570 716
rect 5216 2162 5272 2164
rect 5296 2162 5352 2164
rect 5376 2162 5432 2164
rect 5456 2162 5512 2164
rect 5216 2110 5242 2162
rect 5242 2110 5272 2162
rect 5296 2110 5306 2162
rect 5306 2110 5352 2162
rect 5376 2110 5422 2162
rect 5422 2110 5432 2162
rect 5456 2110 5486 2162
rect 5486 2110 5512 2162
rect 5216 2108 5272 2110
rect 5296 2108 5352 2110
rect 5376 2108 5432 2110
rect 5456 2108 5512 2110
rect 5216 1074 5272 1076
rect 5296 1074 5352 1076
rect 5376 1074 5432 1076
rect 5456 1074 5512 1076
rect 5216 1022 5242 1074
rect 5242 1022 5272 1074
rect 5296 1022 5306 1074
rect 5306 1022 5352 1074
rect 5376 1022 5422 1074
rect 5422 1022 5432 1074
rect 5456 1022 5486 1074
rect 5486 1022 5512 1074
rect 5216 1020 5272 1022
rect 5296 1020 5352 1022
rect 5376 1020 5432 1022
rect 5456 1020 5512 1022
rect 7654 11036 7710 11072
rect 7654 11016 7656 11036
rect 7656 11016 7708 11036
rect 7708 11016 7710 11036
rect 7852 12498 7908 12500
rect 7932 12498 7988 12500
rect 8012 12498 8068 12500
rect 8092 12498 8148 12500
rect 7852 12446 7878 12498
rect 7878 12446 7908 12498
rect 7932 12446 7942 12498
rect 7942 12446 7988 12498
rect 8012 12446 8058 12498
rect 8058 12446 8068 12498
rect 8092 12446 8122 12498
rect 8122 12446 8148 12498
rect 7852 12444 7908 12446
rect 7932 12444 7988 12446
rect 8012 12444 8068 12446
rect 8092 12444 8148 12446
rect 7852 11410 7908 11412
rect 7932 11410 7988 11412
rect 8012 11410 8068 11412
rect 8092 11410 8148 11412
rect 7852 11358 7878 11410
rect 7878 11358 7908 11410
rect 7932 11358 7942 11410
rect 7942 11358 7988 11410
rect 8012 11358 8058 11410
rect 8058 11358 8068 11410
rect 8092 11358 8122 11410
rect 8122 11358 8148 11410
rect 7852 11356 7908 11358
rect 7932 11356 7988 11358
rect 8012 11356 8068 11358
rect 8092 11356 8148 11358
rect 7852 10322 7908 10324
rect 7932 10322 7988 10324
rect 8012 10322 8068 10324
rect 8092 10322 8148 10324
rect 7852 10270 7878 10322
rect 7878 10270 7908 10322
rect 7932 10270 7942 10322
rect 7942 10270 7988 10322
rect 8012 10270 8058 10322
rect 8058 10270 8068 10322
rect 8092 10270 8122 10322
rect 8122 10270 8148 10322
rect 7852 10268 7908 10270
rect 7932 10268 7988 10270
rect 8012 10268 8068 10270
rect 8092 10268 8148 10270
rect 8206 9520 8262 9576
rect 9310 10628 9366 10664
rect 9310 10608 9312 10628
rect 9312 10608 9364 10628
rect 9364 10608 9366 10628
rect 10488 11954 10544 11956
rect 10568 11954 10624 11956
rect 10648 11954 10704 11956
rect 10728 11954 10784 11956
rect 10488 11902 10514 11954
rect 10514 11902 10544 11954
rect 10568 11902 10578 11954
rect 10578 11902 10624 11954
rect 10648 11902 10694 11954
rect 10694 11902 10704 11954
rect 10728 11902 10758 11954
rect 10758 11902 10784 11954
rect 10488 11900 10544 11902
rect 10568 11900 10624 11902
rect 10648 11900 10704 11902
rect 10728 11900 10784 11902
rect 8390 9404 8446 9440
rect 8390 9384 8392 9404
rect 8392 9384 8444 9404
rect 8444 9384 8446 9404
rect 7852 9234 7908 9236
rect 7932 9234 7988 9236
rect 8012 9234 8068 9236
rect 8092 9234 8148 9236
rect 7852 9182 7878 9234
rect 7878 9182 7908 9234
rect 7932 9182 7942 9234
rect 7942 9182 7988 9234
rect 8012 9182 8058 9234
rect 8058 9182 8068 9234
rect 8092 9182 8122 9234
rect 8122 9182 8148 9234
rect 7852 9180 7908 9182
rect 7932 9180 7988 9182
rect 8012 9180 8068 9182
rect 8092 9180 8148 9182
rect 7852 8146 7908 8148
rect 7932 8146 7988 8148
rect 8012 8146 8068 8148
rect 8092 8146 8148 8148
rect 7852 8094 7878 8146
rect 7878 8094 7908 8146
rect 7932 8094 7942 8146
rect 7942 8094 7988 8146
rect 8012 8094 8058 8146
rect 8058 8094 8068 8146
rect 8092 8094 8122 8146
rect 8122 8094 8148 8146
rect 7852 8092 7908 8094
rect 7932 8092 7988 8094
rect 8012 8092 8068 8094
rect 8092 8092 8148 8094
rect 7852 7058 7908 7060
rect 7932 7058 7988 7060
rect 8012 7058 8068 7060
rect 8092 7058 8148 7060
rect 7852 7006 7878 7058
rect 7878 7006 7908 7058
rect 7932 7006 7942 7058
rect 7942 7006 7988 7058
rect 8012 7006 8058 7058
rect 8058 7006 8068 7058
rect 8092 7006 8122 7058
rect 8122 7006 8148 7058
rect 7852 7004 7908 7006
rect 7932 7004 7988 7006
rect 8012 7004 8068 7006
rect 8092 7004 8148 7006
rect 7852 5970 7908 5972
rect 7932 5970 7988 5972
rect 8012 5970 8068 5972
rect 8092 5970 8148 5972
rect 7852 5918 7878 5970
rect 7878 5918 7908 5970
rect 7932 5918 7942 5970
rect 7942 5918 7988 5970
rect 8012 5918 8058 5970
rect 8058 5918 8068 5970
rect 8092 5918 8122 5970
rect 8122 5918 8148 5970
rect 7852 5916 7908 5918
rect 7932 5916 7988 5918
rect 8012 5916 8068 5918
rect 8092 5916 8148 5918
rect 7852 4882 7908 4884
rect 7932 4882 7988 4884
rect 8012 4882 8068 4884
rect 8092 4882 8148 4884
rect 7852 4830 7878 4882
rect 7878 4830 7908 4882
rect 7932 4830 7942 4882
rect 7942 4830 7988 4882
rect 8012 4830 8058 4882
rect 8058 4830 8068 4882
rect 8092 4830 8122 4882
rect 8122 4830 8148 4882
rect 7852 4828 7908 4830
rect 7932 4828 7988 4830
rect 8012 4828 8068 4830
rect 8092 4828 8148 4830
rect 7852 3794 7908 3796
rect 7932 3794 7988 3796
rect 8012 3794 8068 3796
rect 8092 3794 8148 3796
rect 7852 3742 7878 3794
rect 7878 3742 7908 3794
rect 7932 3742 7942 3794
rect 7942 3742 7988 3794
rect 8012 3742 8058 3794
rect 8058 3742 8068 3794
rect 8092 3742 8122 3794
rect 8122 3742 8148 3794
rect 7852 3740 7908 3742
rect 7932 3740 7988 3742
rect 8012 3740 8068 3742
rect 8092 3740 8148 3742
rect 10488 10866 10544 10868
rect 10568 10866 10624 10868
rect 10648 10866 10704 10868
rect 10728 10866 10784 10868
rect 10488 10814 10514 10866
rect 10514 10814 10544 10866
rect 10568 10814 10578 10866
rect 10578 10814 10624 10866
rect 10648 10814 10694 10866
rect 10694 10814 10704 10866
rect 10728 10814 10758 10866
rect 10758 10814 10784 10866
rect 10488 10812 10544 10814
rect 10568 10812 10624 10814
rect 10648 10812 10704 10814
rect 10728 10812 10784 10814
rect 10488 9778 10544 9780
rect 10568 9778 10624 9780
rect 10648 9778 10704 9780
rect 10728 9778 10784 9780
rect 10488 9726 10514 9778
rect 10514 9726 10544 9778
rect 10568 9726 10578 9778
rect 10578 9726 10624 9778
rect 10648 9726 10694 9778
rect 10694 9726 10704 9778
rect 10728 9726 10758 9778
rect 10758 9726 10784 9778
rect 10488 9724 10544 9726
rect 10568 9724 10624 9726
rect 10648 9724 10704 9726
rect 10728 9724 10784 9726
rect 7852 2706 7908 2708
rect 7932 2706 7988 2708
rect 8012 2706 8068 2708
rect 8092 2706 8148 2708
rect 7852 2654 7878 2706
rect 7878 2654 7908 2706
rect 7932 2654 7942 2706
rect 7942 2654 7988 2706
rect 8012 2654 8058 2706
rect 8058 2654 8068 2706
rect 8092 2654 8122 2706
rect 8122 2654 8148 2706
rect 7852 2652 7908 2654
rect 7932 2652 7988 2654
rect 8012 2652 8068 2654
rect 8092 2652 8148 2654
rect 7852 1618 7908 1620
rect 7932 1618 7988 1620
rect 8012 1618 8068 1620
rect 8092 1618 8148 1620
rect 7852 1566 7878 1618
rect 7878 1566 7908 1618
rect 7932 1566 7942 1618
rect 7942 1566 7988 1618
rect 8012 1566 8058 1618
rect 8058 1566 8068 1618
rect 8092 1566 8122 1618
rect 8122 1566 8148 1618
rect 7852 1564 7908 1566
rect 7932 1564 7988 1566
rect 8012 1564 8068 1566
rect 8092 1564 8148 1566
rect 10488 8690 10544 8692
rect 10568 8690 10624 8692
rect 10648 8690 10704 8692
rect 10728 8690 10784 8692
rect 10488 8638 10514 8690
rect 10514 8638 10544 8690
rect 10568 8638 10578 8690
rect 10578 8638 10624 8690
rect 10648 8638 10694 8690
rect 10694 8638 10704 8690
rect 10728 8638 10758 8690
rect 10758 8638 10784 8690
rect 10488 8636 10544 8638
rect 10568 8636 10624 8638
rect 10648 8636 10704 8638
rect 10728 8636 10784 8638
rect 10488 7602 10544 7604
rect 10568 7602 10624 7604
rect 10648 7602 10704 7604
rect 10728 7602 10784 7604
rect 10488 7550 10514 7602
rect 10514 7550 10544 7602
rect 10568 7550 10578 7602
rect 10578 7550 10624 7602
rect 10648 7550 10694 7602
rect 10694 7550 10704 7602
rect 10728 7550 10758 7602
rect 10758 7550 10784 7602
rect 10488 7548 10544 7550
rect 10568 7548 10624 7550
rect 10648 7548 10704 7550
rect 10728 7548 10784 7550
rect 10488 6514 10544 6516
rect 10568 6514 10624 6516
rect 10648 6514 10704 6516
rect 10728 6514 10784 6516
rect 10488 6462 10514 6514
rect 10514 6462 10544 6514
rect 10568 6462 10578 6514
rect 10578 6462 10624 6514
rect 10648 6462 10694 6514
rect 10694 6462 10704 6514
rect 10728 6462 10758 6514
rect 10758 6462 10784 6514
rect 10488 6460 10544 6462
rect 10568 6460 10624 6462
rect 10648 6460 10704 6462
rect 10728 6460 10784 6462
rect 9862 5168 9918 5224
rect 10488 5426 10544 5428
rect 10568 5426 10624 5428
rect 10648 5426 10704 5428
rect 10728 5426 10784 5428
rect 10488 5374 10514 5426
rect 10514 5374 10544 5426
rect 10568 5374 10578 5426
rect 10578 5374 10624 5426
rect 10648 5374 10694 5426
rect 10694 5374 10704 5426
rect 10728 5374 10758 5426
rect 10758 5374 10784 5426
rect 10488 5372 10544 5374
rect 10568 5372 10624 5374
rect 10648 5372 10704 5374
rect 10728 5372 10784 5374
rect 9126 3420 9182 3456
rect 9126 3400 9128 3420
rect 9128 3400 9180 3420
rect 9180 3400 9182 3420
rect 9218 3028 9220 3048
rect 9220 3028 9272 3048
rect 9272 3028 9274 3048
rect 9218 2992 9274 3028
rect 9586 3400 9642 3456
rect 9494 2992 9550 3048
rect 10488 4338 10544 4340
rect 10568 4338 10624 4340
rect 10648 4338 10704 4340
rect 10728 4338 10784 4340
rect 10488 4286 10514 4338
rect 10514 4286 10544 4338
rect 10568 4286 10578 4338
rect 10578 4286 10624 4338
rect 10648 4286 10694 4338
rect 10694 4286 10704 4338
rect 10728 4286 10758 4338
rect 10758 4286 10784 4338
rect 10488 4284 10544 4286
rect 10568 4284 10624 4286
rect 10648 4284 10704 4286
rect 10728 4284 10784 4286
rect 10488 3250 10544 3252
rect 10568 3250 10624 3252
rect 10648 3250 10704 3252
rect 10728 3250 10784 3252
rect 10488 3198 10514 3250
rect 10514 3198 10544 3250
rect 10568 3198 10578 3250
rect 10578 3198 10624 3250
rect 10648 3198 10694 3250
rect 10694 3198 10704 3250
rect 10728 3198 10758 3250
rect 10758 3198 10784 3250
rect 10488 3196 10544 3198
rect 10568 3196 10624 3198
rect 10648 3196 10704 3198
rect 10728 3196 10784 3198
rect 10488 2162 10544 2164
rect 10568 2162 10624 2164
rect 10648 2162 10704 2164
rect 10728 2162 10784 2164
rect 10488 2110 10514 2162
rect 10514 2110 10544 2162
rect 10568 2110 10578 2162
rect 10578 2110 10624 2162
rect 10648 2110 10694 2162
rect 10694 2110 10704 2162
rect 10728 2110 10758 2162
rect 10758 2110 10784 2162
rect 10488 2108 10544 2110
rect 10568 2108 10624 2110
rect 10648 2108 10704 2110
rect 10728 2108 10784 2110
rect 11794 5188 11850 5224
rect 11794 5168 11796 5188
rect 11796 5168 11848 5188
rect 11848 5168 11850 5188
rect 10488 1074 10544 1076
rect 10568 1074 10624 1076
rect 10648 1074 10704 1076
rect 10728 1074 10784 1076
rect 10488 1022 10514 1074
rect 10514 1022 10544 1074
rect 10568 1022 10578 1074
rect 10578 1022 10624 1074
rect 10648 1022 10694 1074
rect 10694 1022 10704 1074
rect 10728 1022 10758 1074
rect 10758 1022 10784 1074
rect 10488 1020 10544 1022
rect 10568 1020 10624 1022
rect 10648 1020 10704 1022
rect 10728 1020 10784 1022
rect 7852 530 7908 532
rect 7932 530 7988 532
rect 8012 530 8068 532
rect 8092 530 8148 532
rect 7852 478 7878 530
rect 7878 478 7908 530
rect 7932 478 7942 530
rect 7942 478 7988 530
rect 8012 478 8058 530
rect 8058 478 8068 530
rect 8092 478 8122 530
rect 8122 478 8148 530
rect 7852 476 7908 478
rect 7932 476 7988 478
rect 8012 476 8068 478
rect 8092 476 8148 478
rect 13124 12498 13180 12500
rect 13204 12498 13260 12500
rect 13284 12498 13340 12500
rect 13364 12498 13420 12500
rect 13124 12446 13150 12498
rect 13150 12446 13180 12498
rect 13204 12446 13214 12498
rect 13214 12446 13260 12498
rect 13284 12446 13330 12498
rect 13330 12446 13340 12498
rect 13364 12446 13394 12498
rect 13394 12446 13420 12498
rect 13124 12444 13180 12446
rect 13204 12444 13260 12446
rect 13284 12444 13340 12446
rect 13364 12444 13420 12446
rect 13124 11410 13180 11412
rect 13204 11410 13260 11412
rect 13284 11410 13340 11412
rect 13364 11410 13420 11412
rect 13124 11358 13150 11410
rect 13150 11358 13180 11410
rect 13204 11358 13214 11410
rect 13214 11358 13260 11410
rect 13284 11358 13330 11410
rect 13330 11358 13340 11410
rect 13364 11358 13394 11410
rect 13394 11358 13420 11410
rect 13124 11356 13180 11358
rect 13204 11356 13260 11358
rect 13284 11356 13340 11358
rect 13364 11356 13420 11358
rect 13124 10322 13180 10324
rect 13204 10322 13260 10324
rect 13284 10322 13340 10324
rect 13364 10322 13420 10324
rect 13124 10270 13150 10322
rect 13150 10270 13180 10322
rect 13204 10270 13214 10322
rect 13214 10270 13260 10322
rect 13284 10270 13330 10322
rect 13330 10270 13340 10322
rect 13364 10270 13394 10322
rect 13394 10270 13420 10322
rect 13124 10268 13180 10270
rect 13204 10268 13260 10270
rect 13284 10268 13340 10270
rect 13364 10268 13420 10270
rect 13124 9234 13180 9236
rect 13204 9234 13260 9236
rect 13284 9234 13340 9236
rect 13364 9234 13420 9236
rect 13124 9182 13150 9234
rect 13150 9182 13180 9234
rect 13204 9182 13214 9234
rect 13214 9182 13260 9234
rect 13284 9182 13330 9234
rect 13330 9182 13340 9234
rect 13364 9182 13394 9234
rect 13394 9182 13420 9234
rect 13124 9180 13180 9182
rect 13204 9180 13260 9182
rect 13284 9180 13340 9182
rect 13364 9180 13420 9182
rect 13124 8146 13180 8148
rect 13204 8146 13260 8148
rect 13284 8146 13340 8148
rect 13364 8146 13420 8148
rect 13124 8094 13150 8146
rect 13150 8094 13180 8146
rect 13204 8094 13214 8146
rect 13214 8094 13260 8146
rect 13284 8094 13330 8146
rect 13330 8094 13340 8146
rect 13364 8094 13394 8146
rect 13394 8094 13420 8146
rect 13124 8092 13180 8094
rect 13204 8092 13260 8094
rect 13284 8092 13340 8094
rect 13364 8092 13420 8094
rect 13124 7058 13180 7060
rect 13204 7058 13260 7060
rect 13284 7058 13340 7060
rect 13364 7058 13420 7060
rect 13124 7006 13150 7058
rect 13150 7006 13180 7058
rect 13204 7006 13214 7058
rect 13214 7006 13260 7058
rect 13284 7006 13330 7058
rect 13330 7006 13340 7058
rect 13364 7006 13394 7058
rect 13394 7006 13420 7058
rect 13124 7004 13180 7006
rect 13204 7004 13260 7006
rect 13284 7004 13340 7006
rect 13364 7004 13420 7006
rect 13124 5970 13180 5972
rect 13204 5970 13260 5972
rect 13284 5970 13340 5972
rect 13364 5970 13420 5972
rect 13124 5918 13150 5970
rect 13150 5918 13180 5970
rect 13204 5918 13214 5970
rect 13214 5918 13260 5970
rect 13284 5918 13330 5970
rect 13330 5918 13340 5970
rect 13364 5918 13394 5970
rect 13394 5918 13420 5970
rect 13124 5916 13180 5918
rect 13204 5916 13260 5918
rect 13284 5916 13340 5918
rect 13364 5916 13420 5918
rect 13124 4882 13180 4884
rect 13204 4882 13260 4884
rect 13284 4882 13340 4884
rect 13364 4882 13420 4884
rect 13124 4830 13150 4882
rect 13150 4830 13180 4882
rect 13204 4830 13214 4882
rect 13214 4830 13260 4882
rect 13284 4830 13330 4882
rect 13330 4830 13340 4882
rect 13364 4830 13394 4882
rect 13394 4830 13420 4882
rect 13124 4828 13180 4830
rect 13204 4828 13260 4830
rect 13284 4828 13340 4830
rect 13364 4828 13420 4830
rect 13124 3794 13180 3796
rect 13204 3794 13260 3796
rect 13284 3794 13340 3796
rect 13364 3794 13420 3796
rect 13124 3742 13150 3794
rect 13150 3742 13180 3794
rect 13204 3742 13214 3794
rect 13214 3742 13260 3794
rect 13284 3742 13330 3794
rect 13330 3742 13340 3794
rect 13364 3742 13394 3794
rect 13394 3742 13420 3794
rect 13124 3740 13180 3742
rect 13204 3740 13260 3742
rect 13284 3740 13340 3742
rect 13364 3740 13420 3742
rect 13124 2706 13180 2708
rect 13204 2706 13260 2708
rect 13284 2706 13340 2708
rect 13364 2706 13420 2708
rect 13124 2654 13150 2706
rect 13150 2654 13180 2706
rect 13204 2654 13214 2706
rect 13214 2654 13260 2706
rect 13284 2654 13330 2706
rect 13330 2654 13340 2706
rect 13364 2654 13394 2706
rect 13394 2654 13420 2706
rect 13124 2652 13180 2654
rect 13204 2652 13260 2654
rect 13284 2652 13340 2654
rect 13364 2652 13420 2654
rect 13124 1618 13180 1620
rect 13204 1618 13260 1620
rect 13284 1618 13340 1620
rect 13364 1618 13420 1620
rect 13124 1566 13150 1618
rect 13150 1566 13180 1618
rect 13204 1566 13214 1618
rect 13214 1566 13260 1618
rect 13284 1566 13330 1618
rect 13330 1566 13340 1618
rect 13364 1566 13394 1618
rect 13394 1566 13420 1618
rect 13124 1564 13180 1566
rect 13204 1564 13260 1566
rect 13284 1564 13340 1566
rect 13364 1564 13420 1566
rect 15106 12124 15162 12160
rect 15106 12104 15108 12124
rect 15108 12104 15160 12124
rect 15160 12104 15162 12124
rect 15106 11036 15162 11072
rect 15106 11016 15108 11036
rect 15108 11016 15160 11036
rect 15160 11016 15162 11036
rect 15106 9792 15162 9848
rect 15106 8704 15162 8760
rect 15566 7480 15622 7536
rect 15198 6256 15254 6312
rect 15014 5168 15070 5224
rect 15106 2876 15162 2912
rect 15106 2856 15108 2876
rect 15108 2856 15160 2876
rect 15160 2856 15162 2876
rect 15106 1632 15162 1688
rect 15474 3980 15476 4000
rect 15476 3980 15528 4000
rect 15528 3980 15530 4000
rect 15474 3944 15530 3980
rect 14370 544 14426 600
rect 13124 530 13180 532
rect 13204 530 13260 532
rect 13284 530 13340 532
rect 13364 530 13420 532
rect 13124 478 13150 530
rect 13150 478 13180 530
rect 13204 478 13214 530
rect 13214 478 13260 530
rect 13284 478 13330 530
rect 13330 478 13340 530
rect 13364 478 13394 530
rect 13394 478 13420 530
rect 13124 476 13180 478
rect 13204 476 13260 478
rect 13284 476 13340 478
rect 13364 476 13420 478
<< metal3 >>
rect 3969 13386 4035 13389
rect 0 13384 4035 13386
rect 0 13328 3974 13384
rect 4030 13328 4035 13384
rect 0 13326 4035 13328
rect 3969 13323 4035 13326
rect 14365 13386 14431 13389
rect 14365 13384 16000 13386
rect 14365 13328 14370 13384
rect 14426 13328 16000 13384
rect 14365 13326 16000 13328
rect 14365 13323 14431 13326
rect 5204 13048 5524 13049
rect 5204 12984 5212 13048
rect 5276 12984 5292 13048
rect 5356 12984 5372 13048
rect 5436 12984 5452 13048
rect 5516 12984 5524 13048
rect 5204 12983 5524 12984
rect 10476 13048 10796 13049
rect 10476 12984 10484 13048
rect 10548 12984 10564 13048
rect 10628 12984 10644 13048
rect 10708 12984 10724 13048
rect 10788 12984 10796 13048
rect 10476 12983 10796 12984
rect 2568 12504 2888 12505
rect 2568 12440 2576 12504
rect 2640 12440 2656 12504
rect 2720 12440 2736 12504
rect 2800 12440 2816 12504
rect 2880 12440 2888 12504
rect 2568 12439 2888 12440
rect 7840 12504 8160 12505
rect 7840 12440 7848 12504
rect 7912 12440 7928 12504
rect 7992 12440 8008 12504
rect 8072 12440 8088 12504
rect 8152 12440 8160 12504
rect 7840 12439 8160 12440
rect 13112 12504 13432 12505
rect 13112 12440 13120 12504
rect 13184 12440 13200 12504
rect 13264 12440 13280 12504
rect 13344 12440 13360 12504
rect 13424 12440 13432 12504
rect 13112 12439 13432 12440
rect 1761 12434 1827 12437
rect 0 12432 1827 12434
rect 0 12376 1766 12432
rect 1822 12376 1827 12432
rect 0 12374 1827 12376
rect 1761 12371 1827 12374
rect 15101 12162 15167 12165
rect 15101 12160 16000 12162
rect 15101 12104 15106 12160
rect 15162 12104 16000 12160
rect 15101 12102 16000 12104
rect 15101 12099 15167 12102
rect 5204 11960 5524 11961
rect 5204 11896 5212 11960
rect 5276 11896 5292 11960
rect 5356 11896 5372 11960
rect 5436 11896 5452 11960
rect 5516 11896 5524 11960
rect 5204 11895 5524 11896
rect 10476 11960 10796 11961
rect 10476 11896 10484 11960
rect 10548 11896 10564 11960
rect 10628 11896 10644 11960
rect 10708 11896 10724 11960
rect 10788 11896 10796 11960
rect 10476 11895 10796 11896
rect 2568 11416 2888 11417
rect 2568 11352 2576 11416
rect 2640 11352 2656 11416
rect 2720 11352 2736 11416
rect 2800 11352 2816 11416
rect 2880 11352 2888 11416
rect 2568 11351 2888 11352
rect 7840 11416 8160 11417
rect 7840 11352 7848 11416
rect 7912 11352 7928 11416
rect 7992 11352 8008 11416
rect 8072 11352 8088 11416
rect 8152 11352 8160 11416
rect 7840 11351 8160 11352
rect 13112 11416 13432 11417
rect 13112 11352 13120 11416
rect 13184 11352 13200 11416
rect 13264 11352 13280 11416
rect 13344 11352 13360 11416
rect 13424 11352 13432 11416
rect 13112 11351 13432 11352
rect 749 11346 815 11349
rect 0 11344 815 11346
rect 0 11288 754 11344
rect 810 11288 815 11344
rect 0 11286 815 11288
rect 749 11283 815 11286
rect 4061 11074 4127 11077
rect 4705 11074 4771 11077
rect 7649 11074 7715 11077
rect 4061 11072 7715 11074
rect 4061 11016 4066 11072
rect 4122 11016 4710 11072
rect 4766 11016 7654 11072
rect 7710 11016 7715 11072
rect 4061 11014 7715 11016
rect 4061 11011 4127 11014
rect 4705 11011 4771 11014
rect 7649 11011 7715 11014
rect 15101 11074 15167 11077
rect 15101 11072 16000 11074
rect 15101 11016 15106 11072
rect 15162 11016 16000 11072
rect 15101 11014 16000 11016
rect 15101 11011 15167 11014
rect 5204 10872 5524 10873
rect 5204 10808 5212 10872
rect 5276 10808 5292 10872
rect 5356 10808 5372 10872
rect 5436 10808 5452 10872
rect 5516 10808 5524 10872
rect 5204 10807 5524 10808
rect 10476 10872 10796 10873
rect 10476 10808 10484 10872
rect 10548 10808 10564 10872
rect 10628 10808 10644 10872
rect 10708 10808 10724 10872
rect 10788 10808 10796 10872
rect 10476 10807 10796 10808
rect 4429 10666 4495 10669
rect 9305 10666 9371 10669
rect 4429 10664 9371 10666
rect 4429 10608 4434 10664
rect 4490 10608 9310 10664
rect 9366 10608 9371 10664
rect 4429 10606 9371 10608
rect 4429 10603 4495 10606
rect 9305 10603 9371 10606
rect 749 10394 815 10397
rect 0 10392 815 10394
rect 0 10336 754 10392
rect 810 10336 815 10392
rect 0 10334 815 10336
rect 749 10331 815 10334
rect 2568 10328 2888 10329
rect 2568 10264 2576 10328
rect 2640 10264 2656 10328
rect 2720 10264 2736 10328
rect 2800 10264 2816 10328
rect 2880 10264 2888 10328
rect 2568 10263 2888 10264
rect 7840 10328 8160 10329
rect 7840 10264 7848 10328
rect 7912 10264 7928 10328
rect 7992 10264 8008 10328
rect 8072 10264 8088 10328
rect 8152 10264 8160 10328
rect 7840 10263 8160 10264
rect 13112 10328 13432 10329
rect 13112 10264 13120 10328
rect 13184 10264 13200 10328
rect 13264 10264 13280 10328
rect 13344 10264 13360 10328
rect 13424 10264 13432 10328
rect 13112 10263 13432 10264
rect 5993 10258 6059 10261
rect 6269 10258 6335 10261
rect 5993 10256 6335 10258
rect 5993 10200 5998 10256
rect 6054 10200 6274 10256
rect 6330 10200 6335 10256
rect 5993 10198 6335 10200
rect 5993 10195 6059 10198
rect 6269 10195 6335 10198
rect 15101 9850 15167 9853
rect 15101 9848 16000 9850
rect 15101 9792 15106 9848
rect 15162 9792 16000 9848
rect 15101 9790 16000 9792
rect 15101 9787 15167 9790
rect 5204 9784 5524 9785
rect 5204 9720 5212 9784
rect 5276 9720 5292 9784
rect 5356 9720 5372 9784
rect 5436 9720 5452 9784
rect 5516 9720 5524 9784
rect 5204 9719 5524 9720
rect 10476 9784 10796 9785
rect 10476 9720 10484 9784
rect 10548 9720 10564 9784
rect 10628 9720 10644 9784
rect 10708 9720 10724 9784
rect 10788 9720 10796 9784
rect 10476 9719 10796 9720
rect 7005 9578 7071 9581
rect 8201 9578 8267 9581
rect 7005 9576 8267 9578
rect 7005 9520 7010 9576
rect 7066 9520 8206 9576
rect 8262 9520 8267 9576
rect 7005 9518 8267 9520
rect 7005 9515 7071 9518
rect 8201 9515 8267 9518
rect 749 9442 815 9445
rect 0 9440 815 9442
rect 0 9384 754 9440
rect 810 9384 815 9440
rect 0 9382 815 9384
rect 749 9379 815 9382
rect 4429 9442 4495 9445
rect 6637 9442 6703 9445
rect 4429 9440 6703 9442
rect 4429 9384 4434 9440
rect 4490 9384 6642 9440
rect 6698 9384 6703 9440
rect 4429 9382 6703 9384
rect 4429 9379 4495 9382
rect 6637 9379 6703 9382
rect 7097 9442 7163 9445
rect 8385 9442 8451 9445
rect 7097 9440 8451 9442
rect 7097 9384 7102 9440
rect 7158 9384 8390 9440
rect 8446 9384 8451 9440
rect 7097 9382 8451 9384
rect 7097 9379 7163 9382
rect 8385 9379 8451 9382
rect 2568 9240 2888 9241
rect 2568 9176 2576 9240
rect 2640 9176 2656 9240
rect 2720 9176 2736 9240
rect 2800 9176 2816 9240
rect 2880 9176 2888 9240
rect 2568 9175 2888 9176
rect 7840 9240 8160 9241
rect 7840 9176 7848 9240
rect 7912 9176 7928 9240
rect 7992 9176 8008 9240
rect 8072 9176 8088 9240
rect 8152 9176 8160 9240
rect 7840 9175 8160 9176
rect 13112 9240 13432 9241
rect 13112 9176 13120 9240
rect 13184 9176 13200 9240
rect 13264 9176 13280 9240
rect 13344 9176 13360 9240
rect 13424 9176 13432 9240
rect 13112 9175 13432 9176
rect 15101 8762 15167 8765
rect 15101 8760 16000 8762
rect 15101 8704 15106 8760
rect 15162 8704 16000 8760
rect 15101 8702 16000 8704
rect 15101 8699 15167 8702
rect 5204 8696 5524 8697
rect 5204 8632 5212 8696
rect 5276 8632 5292 8696
rect 5356 8632 5372 8696
rect 5436 8632 5452 8696
rect 5516 8632 5524 8696
rect 5204 8631 5524 8632
rect 10476 8696 10796 8697
rect 10476 8632 10484 8696
rect 10548 8632 10564 8696
rect 10628 8632 10644 8696
rect 10708 8632 10724 8696
rect 10788 8632 10796 8696
rect 10476 8631 10796 8632
rect 749 8354 815 8357
rect 0 8352 815 8354
rect 0 8296 754 8352
rect 810 8296 815 8352
rect 0 8294 815 8296
rect 749 8291 815 8294
rect 2568 8152 2888 8153
rect 2568 8088 2576 8152
rect 2640 8088 2656 8152
rect 2720 8088 2736 8152
rect 2800 8088 2816 8152
rect 2880 8088 2888 8152
rect 2568 8087 2888 8088
rect 7840 8152 8160 8153
rect 7840 8088 7848 8152
rect 7912 8088 7928 8152
rect 7992 8088 8008 8152
rect 8072 8088 8088 8152
rect 8152 8088 8160 8152
rect 7840 8087 8160 8088
rect 13112 8152 13432 8153
rect 13112 8088 13120 8152
rect 13184 8088 13200 8152
rect 13264 8088 13280 8152
rect 13344 8088 13360 8152
rect 13424 8088 13432 8152
rect 13112 8087 13432 8088
rect 5204 7608 5524 7609
rect 5204 7544 5212 7608
rect 5276 7544 5292 7608
rect 5356 7544 5372 7608
rect 5436 7544 5452 7608
rect 5516 7544 5524 7608
rect 5204 7543 5524 7544
rect 10476 7608 10796 7609
rect 10476 7544 10484 7608
rect 10548 7544 10564 7608
rect 10628 7544 10644 7608
rect 10708 7544 10724 7608
rect 10788 7544 10796 7608
rect 10476 7543 10796 7544
rect 15561 7538 15627 7541
rect 15561 7536 16000 7538
rect 15561 7480 15566 7536
rect 15622 7480 16000 7536
rect 15561 7478 16000 7480
rect 15561 7475 15627 7478
rect 473 7402 539 7405
rect 0 7400 539 7402
rect 0 7344 478 7400
rect 534 7344 539 7400
rect 0 7342 539 7344
rect 473 7339 539 7342
rect 2568 7064 2888 7065
rect 2568 7000 2576 7064
rect 2640 7000 2656 7064
rect 2720 7000 2736 7064
rect 2800 7000 2816 7064
rect 2880 7000 2888 7064
rect 2568 6999 2888 7000
rect 7840 7064 8160 7065
rect 7840 7000 7848 7064
rect 7912 7000 7928 7064
rect 7992 7000 8008 7064
rect 8072 7000 8088 7064
rect 8152 7000 8160 7064
rect 7840 6999 8160 7000
rect 13112 7064 13432 7065
rect 13112 7000 13120 7064
rect 13184 7000 13200 7064
rect 13264 7000 13280 7064
rect 13344 7000 13360 7064
rect 13424 7000 13432 7064
rect 13112 6999 13432 7000
rect 4521 6858 4587 6861
rect 5993 6858 6059 6861
rect 6637 6858 6703 6861
rect 4521 6856 6703 6858
rect 4521 6800 4526 6856
rect 4582 6800 5998 6856
rect 6054 6800 6642 6856
rect 6698 6800 6703 6856
rect 4521 6798 6703 6800
rect 4521 6795 4587 6798
rect 5993 6795 6059 6798
rect 6637 6795 6703 6798
rect 5625 6722 5691 6725
rect 6453 6722 6519 6725
rect 5625 6720 6519 6722
rect 5625 6664 5630 6720
rect 5686 6664 6458 6720
rect 6514 6664 6519 6720
rect 5625 6662 6519 6664
rect 5625 6659 5691 6662
rect 6453 6659 6519 6662
rect 5204 6520 5524 6521
rect 5204 6456 5212 6520
rect 5276 6456 5292 6520
rect 5356 6456 5372 6520
rect 5436 6456 5452 6520
rect 5516 6456 5524 6520
rect 5204 6455 5524 6456
rect 10476 6520 10796 6521
rect 10476 6456 10484 6520
rect 10548 6456 10564 6520
rect 10628 6456 10644 6520
rect 10708 6456 10724 6520
rect 10788 6456 10796 6520
rect 10476 6455 10796 6456
rect 749 6450 815 6453
rect 0 6448 815 6450
rect 0 6392 754 6448
rect 810 6392 815 6448
rect 0 6390 815 6392
rect 749 6387 815 6390
rect 15193 6314 15259 6317
rect 15193 6312 16000 6314
rect 15193 6256 15198 6312
rect 15254 6256 16000 6312
rect 15193 6254 16000 6256
rect 15193 6251 15259 6254
rect 2568 5976 2888 5977
rect 2568 5912 2576 5976
rect 2640 5912 2656 5976
rect 2720 5912 2736 5976
rect 2800 5912 2816 5976
rect 2880 5912 2888 5976
rect 2568 5911 2888 5912
rect 7840 5976 8160 5977
rect 7840 5912 7848 5976
rect 7912 5912 7928 5976
rect 7992 5912 8008 5976
rect 8072 5912 8088 5976
rect 8152 5912 8160 5976
rect 7840 5911 8160 5912
rect 13112 5976 13432 5977
rect 13112 5912 13120 5976
rect 13184 5912 13200 5976
rect 13264 5912 13280 5976
rect 13344 5912 13360 5976
rect 13424 5912 13432 5976
rect 13112 5911 13432 5912
rect 5204 5432 5524 5433
rect 5204 5368 5212 5432
rect 5276 5368 5292 5432
rect 5356 5368 5372 5432
rect 5436 5368 5452 5432
rect 5516 5368 5524 5432
rect 5204 5367 5524 5368
rect 10476 5432 10796 5433
rect 10476 5368 10484 5432
rect 10548 5368 10564 5432
rect 10628 5368 10644 5432
rect 10708 5368 10724 5432
rect 10788 5368 10796 5432
rect 10476 5367 10796 5368
rect 749 5362 815 5365
rect 0 5360 815 5362
rect 0 5304 754 5360
rect 810 5304 815 5360
rect 0 5302 815 5304
rect 749 5299 815 5302
rect 9857 5226 9923 5229
rect 11789 5226 11855 5229
rect 9857 5224 11855 5226
rect 9857 5168 9862 5224
rect 9918 5168 11794 5224
rect 11850 5168 11855 5224
rect 9857 5166 11855 5168
rect 9857 5163 9923 5166
rect 11789 5163 11855 5166
rect 15009 5226 15075 5229
rect 15009 5224 16000 5226
rect 15009 5168 15014 5224
rect 15070 5168 16000 5224
rect 15009 5166 16000 5168
rect 15009 5163 15075 5166
rect 2568 4888 2888 4889
rect 2568 4824 2576 4888
rect 2640 4824 2656 4888
rect 2720 4824 2736 4888
rect 2800 4824 2816 4888
rect 2880 4824 2888 4888
rect 2568 4823 2888 4824
rect 7840 4888 8160 4889
rect 7840 4824 7848 4888
rect 7912 4824 7928 4888
rect 7992 4824 8008 4888
rect 8072 4824 8088 4888
rect 8152 4824 8160 4888
rect 7840 4823 8160 4824
rect 13112 4888 13432 4889
rect 13112 4824 13120 4888
rect 13184 4824 13200 4888
rect 13264 4824 13280 4888
rect 13344 4824 13360 4888
rect 13424 4824 13432 4888
rect 13112 4823 13432 4824
rect 841 4410 907 4413
rect 0 4408 907 4410
rect 0 4352 846 4408
rect 902 4352 907 4408
rect 0 4350 907 4352
rect 841 4347 907 4350
rect 5204 4344 5524 4345
rect 5204 4280 5212 4344
rect 5276 4280 5292 4344
rect 5356 4280 5372 4344
rect 5436 4280 5452 4344
rect 5516 4280 5524 4344
rect 5204 4279 5524 4280
rect 10476 4344 10796 4345
rect 10476 4280 10484 4344
rect 10548 4280 10564 4344
rect 10628 4280 10644 4344
rect 10708 4280 10724 4344
rect 10788 4280 10796 4344
rect 10476 4279 10796 4280
rect 15469 4002 15535 4005
rect 15469 4000 16000 4002
rect 15469 3944 15474 4000
rect 15530 3944 16000 4000
rect 15469 3942 16000 3944
rect 15469 3939 15535 3942
rect 2568 3800 2888 3801
rect 2568 3736 2576 3800
rect 2640 3736 2656 3800
rect 2720 3736 2736 3800
rect 2800 3736 2816 3800
rect 2880 3736 2888 3800
rect 2568 3735 2888 3736
rect 7840 3800 8160 3801
rect 7840 3736 7848 3800
rect 7912 3736 7928 3800
rect 7992 3736 8008 3800
rect 8072 3736 8088 3800
rect 8152 3736 8160 3800
rect 7840 3735 8160 3736
rect 13112 3800 13432 3801
rect 13112 3736 13120 3800
rect 13184 3736 13200 3800
rect 13264 3736 13280 3800
rect 13344 3736 13360 3800
rect 13424 3736 13432 3800
rect 13112 3735 13432 3736
rect 4061 3458 4127 3461
rect 0 3456 4127 3458
rect 0 3400 4066 3456
rect 4122 3400 4127 3456
rect 0 3398 4127 3400
rect 4061 3395 4127 3398
rect 9121 3458 9187 3461
rect 9581 3458 9647 3461
rect 9121 3456 9647 3458
rect 9121 3400 9126 3456
rect 9182 3400 9586 3456
rect 9642 3400 9647 3456
rect 9121 3398 9647 3400
rect 9121 3395 9187 3398
rect 9581 3395 9647 3398
rect 5204 3256 5524 3257
rect 5204 3192 5212 3256
rect 5276 3192 5292 3256
rect 5356 3192 5372 3256
rect 5436 3192 5452 3256
rect 5516 3192 5524 3256
rect 5204 3191 5524 3192
rect 10476 3256 10796 3257
rect 10476 3192 10484 3256
rect 10548 3192 10564 3256
rect 10628 3192 10644 3256
rect 10708 3192 10724 3256
rect 10788 3192 10796 3256
rect 10476 3191 10796 3192
rect 9213 3050 9279 3053
rect 9489 3050 9555 3053
rect 9213 3048 9555 3050
rect 9213 2992 9218 3048
rect 9274 2992 9494 3048
rect 9550 2992 9555 3048
rect 9213 2990 9555 2992
rect 9213 2987 9279 2990
rect 9489 2987 9555 2990
rect 15101 2914 15167 2917
rect 15101 2912 16000 2914
rect 15101 2856 15106 2912
rect 15162 2856 16000 2912
rect 15101 2854 16000 2856
rect 15101 2851 15167 2854
rect 2568 2712 2888 2713
rect 2568 2648 2576 2712
rect 2640 2648 2656 2712
rect 2720 2648 2736 2712
rect 2800 2648 2816 2712
rect 2880 2648 2888 2712
rect 2568 2647 2888 2648
rect 7840 2712 8160 2713
rect 7840 2648 7848 2712
rect 7912 2648 7928 2712
rect 7992 2648 8008 2712
rect 8072 2648 8088 2712
rect 8152 2648 8160 2712
rect 7840 2647 8160 2648
rect 13112 2712 13432 2713
rect 13112 2648 13120 2712
rect 13184 2648 13200 2712
rect 13264 2648 13280 2712
rect 13344 2648 13360 2712
rect 13424 2648 13432 2712
rect 13112 2647 13432 2648
rect 841 2370 907 2373
rect 0 2368 907 2370
rect 0 2312 846 2368
rect 902 2312 907 2368
rect 0 2310 907 2312
rect 841 2307 907 2310
rect 5204 2168 5524 2169
rect 5204 2104 5212 2168
rect 5276 2104 5292 2168
rect 5356 2104 5372 2168
rect 5436 2104 5452 2168
rect 5516 2104 5524 2168
rect 5204 2103 5524 2104
rect 10476 2168 10796 2169
rect 10476 2104 10484 2168
rect 10548 2104 10564 2168
rect 10628 2104 10644 2168
rect 10708 2104 10724 2168
rect 10788 2104 10796 2168
rect 10476 2103 10796 2104
rect 15101 1690 15167 1693
rect 15101 1688 16000 1690
rect 15101 1632 15106 1688
rect 15162 1632 16000 1688
rect 15101 1630 16000 1632
rect 15101 1627 15167 1630
rect 2568 1624 2888 1625
rect 2568 1560 2576 1624
rect 2640 1560 2656 1624
rect 2720 1560 2736 1624
rect 2800 1560 2816 1624
rect 2880 1560 2888 1624
rect 2568 1559 2888 1560
rect 7840 1624 8160 1625
rect 7840 1560 7848 1624
rect 7912 1560 7928 1624
rect 7992 1560 8008 1624
rect 8072 1560 8088 1624
rect 8152 1560 8160 1624
rect 7840 1559 8160 1560
rect 13112 1624 13432 1625
rect 13112 1560 13120 1624
rect 13184 1560 13200 1624
rect 13264 1560 13280 1624
rect 13344 1560 13360 1624
rect 13424 1560 13432 1624
rect 13112 1559 13432 1560
rect 3325 1418 3391 1421
rect 0 1416 3391 1418
rect 0 1360 3330 1416
rect 3386 1360 3391 1416
rect 0 1358 3391 1360
rect 3325 1355 3391 1358
rect 5204 1080 5524 1081
rect 5204 1016 5212 1080
rect 5276 1016 5292 1080
rect 5356 1016 5372 1080
rect 5436 1016 5452 1080
rect 5516 1016 5524 1080
rect 5204 1015 5524 1016
rect 10476 1080 10796 1081
rect 10476 1016 10484 1080
rect 10548 1016 10564 1080
rect 10628 1016 10644 1080
rect 10708 1016 10724 1080
rect 10788 1016 10796 1080
rect 10476 1015 10796 1016
rect 3509 738 3575 741
rect 2270 736 3575 738
rect 2270 680 3514 736
rect 3570 680 3575 736
rect 2270 678 3575 680
rect 2270 466 2330 678
rect 3509 675 3575 678
rect 14365 602 14431 605
rect 14365 600 16000 602
rect 14365 544 14370 600
rect 14426 544 16000 600
rect 14365 542 16000 544
rect 14365 539 14431 542
rect 2568 536 2888 537
rect 2568 472 2576 536
rect 2640 472 2656 536
rect 2720 472 2736 536
rect 2800 472 2816 536
rect 2880 472 2888 536
rect 2568 471 2888 472
rect 7840 536 8160 537
rect 7840 472 7848 536
rect 7912 472 7928 536
rect 7992 472 8008 536
rect 8072 472 8088 536
rect 8152 472 8160 536
rect 7840 471 8160 472
rect 13112 536 13432 537
rect 13112 472 13120 536
rect 13184 472 13200 536
rect 13264 472 13280 536
rect 13344 472 13360 536
rect 13424 472 13432 536
rect 13112 471 13432 472
rect 0 406 2330 466
<< via3 >>
rect 5212 13044 5276 13048
rect 5212 12988 5216 13044
rect 5216 12988 5272 13044
rect 5272 12988 5276 13044
rect 5212 12984 5276 12988
rect 5292 13044 5356 13048
rect 5292 12988 5296 13044
rect 5296 12988 5352 13044
rect 5352 12988 5356 13044
rect 5292 12984 5356 12988
rect 5372 13044 5436 13048
rect 5372 12988 5376 13044
rect 5376 12988 5432 13044
rect 5432 12988 5436 13044
rect 5372 12984 5436 12988
rect 5452 13044 5516 13048
rect 5452 12988 5456 13044
rect 5456 12988 5512 13044
rect 5512 12988 5516 13044
rect 5452 12984 5516 12988
rect 10484 13044 10548 13048
rect 10484 12988 10488 13044
rect 10488 12988 10544 13044
rect 10544 12988 10548 13044
rect 10484 12984 10548 12988
rect 10564 13044 10628 13048
rect 10564 12988 10568 13044
rect 10568 12988 10624 13044
rect 10624 12988 10628 13044
rect 10564 12984 10628 12988
rect 10644 13044 10708 13048
rect 10644 12988 10648 13044
rect 10648 12988 10704 13044
rect 10704 12988 10708 13044
rect 10644 12984 10708 12988
rect 10724 13044 10788 13048
rect 10724 12988 10728 13044
rect 10728 12988 10784 13044
rect 10784 12988 10788 13044
rect 10724 12984 10788 12988
rect 2576 12500 2640 12504
rect 2576 12444 2580 12500
rect 2580 12444 2636 12500
rect 2636 12444 2640 12500
rect 2576 12440 2640 12444
rect 2656 12500 2720 12504
rect 2656 12444 2660 12500
rect 2660 12444 2716 12500
rect 2716 12444 2720 12500
rect 2656 12440 2720 12444
rect 2736 12500 2800 12504
rect 2736 12444 2740 12500
rect 2740 12444 2796 12500
rect 2796 12444 2800 12500
rect 2736 12440 2800 12444
rect 2816 12500 2880 12504
rect 2816 12444 2820 12500
rect 2820 12444 2876 12500
rect 2876 12444 2880 12500
rect 2816 12440 2880 12444
rect 7848 12500 7912 12504
rect 7848 12444 7852 12500
rect 7852 12444 7908 12500
rect 7908 12444 7912 12500
rect 7848 12440 7912 12444
rect 7928 12500 7992 12504
rect 7928 12444 7932 12500
rect 7932 12444 7988 12500
rect 7988 12444 7992 12500
rect 7928 12440 7992 12444
rect 8008 12500 8072 12504
rect 8008 12444 8012 12500
rect 8012 12444 8068 12500
rect 8068 12444 8072 12500
rect 8008 12440 8072 12444
rect 8088 12500 8152 12504
rect 8088 12444 8092 12500
rect 8092 12444 8148 12500
rect 8148 12444 8152 12500
rect 8088 12440 8152 12444
rect 13120 12500 13184 12504
rect 13120 12444 13124 12500
rect 13124 12444 13180 12500
rect 13180 12444 13184 12500
rect 13120 12440 13184 12444
rect 13200 12500 13264 12504
rect 13200 12444 13204 12500
rect 13204 12444 13260 12500
rect 13260 12444 13264 12500
rect 13200 12440 13264 12444
rect 13280 12500 13344 12504
rect 13280 12444 13284 12500
rect 13284 12444 13340 12500
rect 13340 12444 13344 12500
rect 13280 12440 13344 12444
rect 13360 12500 13424 12504
rect 13360 12444 13364 12500
rect 13364 12444 13420 12500
rect 13420 12444 13424 12500
rect 13360 12440 13424 12444
rect 5212 11956 5276 11960
rect 5212 11900 5216 11956
rect 5216 11900 5272 11956
rect 5272 11900 5276 11956
rect 5212 11896 5276 11900
rect 5292 11956 5356 11960
rect 5292 11900 5296 11956
rect 5296 11900 5352 11956
rect 5352 11900 5356 11956
rect 5292 11896 5356 11900
rect 5372 11956 5436 11960
rect 5372 11900 5376 11956
rect 5376 11900 5432 11956
rect 5432 11900 5436 11956
rect 5372 11896 5436 11900
rect 5452 11956 5516 11960
rect 5452 11900 5456 11956
rect 5456 11900 5512 11956
rect 5512 11900 5516 11956
rect 5452 11896 5516 11900
rect 10484 11956 10548 11960
rect 10484 11900 10488 11956
rect 10488 11900 10544 11956
rect 10544 11900 10548 11956
rect 10484 11896 10548 11900
rect 10564 11956 10628 11960
rect 10564 11900 10568 11956
rect 10568 11900 10624 11956
rect 10624 11900 10628 11956
rect 10564 11896 10628 11900
rect 10644 11956 10708 11960
rect 10644 11900 10648 11956
rect 10648 11900 10704 11956
rect 10704 11900 10708 11956
rect 10644 11896 10708 11900
rect 10724 11956 10788 11960
rect 10724 11900 10728 11956
rect 10728 11900 10784 11956
rect 10784 11900 10788 11956
rect 10724 11896 10788 11900
rect 2576 11412 2640 11416
rect 2576 11356 2580 11412
rect 2580 11356 2636 11412
rect 2636 11356 2640 11412
rect 2576 11352 2640 11356
rect 2656 11412 2720 11416
rect 2656 11356 2660 11412
rect 2660 11356 2716 11412
rect 2716 11356 2720 11412
rect 2656 11352 2720 11356
rect 2736 11412 2800 11416
rect 2736 11356 2740 11412
rect 2740 11356 2796 11412
rect 2796 11356 2800 11412
rect 2736 11352 2800 11356
rect 2816 11412 2880 11416
rect 2816 11356 2820 11412
rect 2820 11356 2876 11412
rect 2876 11356 2880 11412
rect 2816 11352 2880 11356
rect 7848 11412 7912 11416
rect 7848 11356 7852 11412
rect 7852 11356 7908 11412
rect 7908 11356 7912 11412
rect 7848 11352 7912 11356
rect 7928 11412 7992 11416
rect 7928 11356 7932 11412
rect 7932 11356 7988 11412
rect 7988 11356 7992 11412
rect 7928 11352 7992 11356
rect 8008 11412 8072 11416
rect 8008 11356 8012 11412
rect 8012 11356 8068 11412
rect 8068 11356 8072 11412
rect 8008 11352 8072 11356
rect 8088 11412 8152 11416
rect 8088 11356 8092 11412
rect 8092 11356 8148 11412
rect 8148 11356 8152 11412
rect 8088 11352 8152 11356
rect 13120 11412 13184 11416
rect 13120 11356 13124 11412
rect 13124 11356 13180 11412
rect 13180 11356 13184 11412
rect 13120 11352 13184 11356
rect 13200 11412 13264 11416
rect 13200 11356 13204 11412
rect 13204 11356 13260 11412
rect 13260 11356 13264 11412
rect 13200 11352 13264 11356
rect 13280 11412 13344 11416
rect 13280 11356 13284 11412
rect 13284 11356 13340 11412
rect 13340 11356 13344 11412
rect 13280 11352 13344 11356
rect 13360 11412 13424 11416
rect 13360 11356 13364 11412
rect 13364 11356 13420 11412
rect 13420 11356 13424 11412
rect 13360 11352 13424 11356
rect 5212 10868 5276 10872
rect 5212 10812 5216 10868
rect 5216 10812 5272 10868
rect 5272 10812 5276 10868
rect 5212 10808 5276 10812
rect 5292 10868 5356 10872
rect 5292 10812 5296 10868
rect 5296 10812 5352 10868
rect 5352 10812 5356 10868
rect 5292 10808 5356 10812
rect 5372 10868 5436 10872
rect 5372 10812 5376 10868
rect 5376 10812 5432 10868
rect 5432 10812 5436 10868
rect 5372 10808 5436 10812
rect 5452 10868 5516 10872
rect 5452 10812 5456 10868
rect 5456 10812 5512 10868
rect 5512 10812 5516 10868
rect 5452 10808 5516 10812
rect 10484 10868 10548 10872
rect 10484 10812 10488 10868
rect 10488 10812 10544 10868
rect 10544 10812 10548 10868
rect 10484 10808 10548 10812
rect 10564 10868 10628 10872
rect 10564 10812 10568 10868
rect 10568 10812 10624 10868
rect 10624 10812 10628 10868
rect 10564 10808 10628 10812
rect 10644 10868 10708 10872
rect 10644 10812 10648 10868
rect 10648 10812 10704 10868
rect 10704 10812 10708 10868
rect 10644 10808 10708 10812
rect 10724 10868 10788 10872
rect 10724 10812 10728 10868
rect 10728 10812 10784 10868
rect 10784 10812 10788 10868
rect 10724 10808 10788 10812
rect 2576 10324 2640 10328
rect 2576 10268 2580 10324
rect 2580 10268 2636 10324
rect 2636 10268 2640 10324
rect 2576 10264 2640 10268
rect 2656 10324 2720 10328
rect 2656 10268 2660 10324
rect 2660 10268 2716 10324
rect 2716 10268 2720 10324
rect 2656 10264 2720 10268
rect 2736 10324 2800 10328
rect 2736 10268 2740 10324
rect 2740 10268 2796 10324
rect 2796 10268 2800 10324
rect 2736 10264 2800 10268
rect 2816 10324 2880 10328
rect 2816 10268 2820 10324
rect 2820 10268 2876 10324
rect 2876 10268 2880 10324
rect 2816 10264 2880 10268
rect 7848 10324 7912 10328
rect 7848 10268 7852 10324
rect 7852 10268 7908 10324
rect 7908 10268 7912 10324
rect 7848 10264 7912 10268
rect 7928 10324 7992 10328
rect 7928 10268 7932 10324
rect 7932 10268 7988 10324
rect 7988 10268 7992 10324
rect 7928 10264 7992 10268
rect 8008 10324 8072 10328
rect 8008 10268 8012 10324
rect 8012 10268 8068 10324
rect 8068 10268 8072 10324
rect 8008 10264 8072 10268
rect 8088 10324 8152 10328
rect 8088 10268 8092 10324
rect 8092 10268 8148 10324
rect 8148 10268 8152 10324
rect 8088 10264 8152 10268
rect 13120 10324 13184 10328
rect 13120 10268 13124 10324
rect 13124 10268 13180 10324
rect 13180 10268 13184 10324
rect 13120 10264 13184 10268
rect 13200 10324 13264 10328
rect 13200 10268 13204 10324
rect 13204 10268 13260 10324
rect 13260 10268 13264 10324
rect 13200 10264 13264 10268
rect 13280 10324 13344 10328
rect 13280 10268 13284 10324
rect 13284 10268 13340 10324
rect 13340 10268 13344 10324
rect 13280 10264 13344 10268
rect 13360 10324 13424 10328
rect 13360 10268 13364 10324
rect 13364 10268 13420 10324
rect 13420 10268 13424 10324
rect 13360 10264 13424 10268
rect 5212 9780 5276 9784
rect 5212 9724 5216 9780
rect 5216 9724 5272 9780
rect 5272 9724 5276 9780
rect 5212 9720 5276 9724
rect 5292 9780 5356 9784
rect 5292 9724 5296 9780
rect 5296 9724 5352 9780
rect 5352 9724 5356 9780
rect 5292 9720 5356 9724
rect 5372 9780 5436 9784
rect 5372 9724 5376 9780
rect 5376 9724 5432 9780
rect 5432 9724 5436 9780
rect 5372 9720 5436 9724
rect 5452 9780 5516 9784
rect 5452 9724 5456 9780
rect 5456 9724 5512 9780
rect 5512 9724 5516 9780
rect 5452 9720 5516 9724
rect 10484 9780 10548 9784
rect 10484 9724 10488 9780
rect 10488 9724 10544 9780
rect 10544 9724 10548 9780
rect 10484 9720 10548 9724
rect 10564 9780 10628 9784
rect 10564 9724 10568 9780
rect 10568 9724 10624 9780
rect 10624 9724 10628 9780
rect 10564 9720 10628 9724
rect 10644 9780 10708 9784
rect 10644 9724 10648 9780
rect 10648 9724 10704 9780
rect 10704 9724 10708 9780
rect 10644 9720 10708 9724
rect 10724 9780 10788 9784
rect 10724 9724 10728 9780
rect 10728 9724 10784 9780
rect 10784 9724 10788 9780
rect 10724 9720 10788 9724
rect 2576 9236 2640 9240
rect 2576 9180 2580 9236
rect 2580 9180 2636 9236
rect 2636 9180 2640 9236
rect 2576 9176 2640 9180
rect 2656 9236 2720 9240
rect 2656 9180 2660 9236
rect 2660 9180 2716 9236
rect 2716 9180 2720 9236
rect 2656 9176 2720 9180
rect 2736 9236 2800 9240
rect 2736 9180 2740 9236
rect 2740 9180 2796 9236
rect 2796 9180 2800 9236
rect 2736 9176 2800 9180
rect 2816 9236 2880 9240
rect 2816 9180 2820 9236
rect 2820 9180 2876 9236
rect 2876 9180 2880 9236
rect 2816 9176 2880 9180
rect 7848 9236 7912 9240
rect 7848 9180 7852 9236
rect 7852 9180 7908 9236
rect 7908 9180 7912 9236
rect 7848 9176 7912 9180
rect 7928 9236 7992 9240
rect 7928 9180 7932 9236
rect 7932 9180 7988 9236
rect 7988 9180 7992 9236
rect 7928 9176 7992 9180
rect 8008 9236 8072 9240
rect 8008 9180 8012 9236
rect 8012 9180 8068 9236
rect 8068 9180 8072 9236
rect 8008 9176 8072 9180
rect 8088 9236 8152 9240
rect 8088 9180 8092 9236
rect 8092 9180 8148 9236
rect 8148 9180 8152 9236
rect 8088 9176 8152 9180
rect 13120 9236 13184 9240
rect 13120 9180 13124 9236
rect 13124 9180 13180 9236
rect 13180 9180 13184 9236
rect 13120 9176 13184 9180
rect 13200 9236 13264 9240
rect 13200 9180 13204 9236
rect 13204 9180 13260 9236
rect 13260 9180 13264 9236
rect 13200 9176 13264 9180
rect 13280 9236 13344 9240
rect 13280 9180 13284 9236
rect 13284 9180 13340 9236
rect 13340 9180 13344 9236
rect 13280 9176 13344 9180
rect 13360 9236 13424 9240
rect 13360 9180 13364 9236
rect 13364 9180 13420 9236
rect 13420 9180 13424 9236
rect 13360 9176 13424 9180
rect 5212 8692 5276 8696
rect 5212 8636 5216 8692
rect 5216 8636 5272 8692
rect 5272 8636 5276 8692
rect 5212 8632 5276 8636
rect 5292 8692 5356 8696
rect 5292 8636 5296 8692
rect 5296 8636 5352 8692
rect 5352 8636 5356 8692
rect 5292 8632 5356 8636
rect 5372 8692 5436 8696
rect 5372 8636 5376 8692
rect 5376 8636 5432 8692
rect 5432 8636 5436 8692
rect 5372 8632 5436 8636
rect 5452 8692 5516 8696
rect 5452 8636 5456 8692
rect 5456 8636 5512 8692
rect 5512 8636 5516 8692
rect 5452 8632 5516 8636
rect 10484 8692 10548 8696
rect 10484 8636 10488 8692
rect 10488 8636 10544 8692
rect 10544 8636 10548 8692
rect 10484 8632 10548 8636
rect 10564 8692 10628 8696
rect 10564 8636 10568 8692
rect 10568 8636 10624 8692
rect 10624 8636 10628 8692
rect 10564 8632 10628 8636
rect 10644 8692 10708 8696
rect 10644 8636 10648 8692
rect 10648 8636 10704 8692
rect 10704 8636 10708 8692
rect 10644 8632 10708 8636
rect 10724 8692 10788 8696
rect 10724 8636 10728 8692
rect 10728 8636 10784 8692
rect 10784 8636 10788 8692
rect 10724 8632 10788 8636
rect 2576 8148 2640 8152
rect 2576 8092 2580 8148
rect 2580 8092 2636 8148
rect 2636 8092 2640 8148
rect 2576 8088 2640 8092
rect 2656 8148 2720 8152
rect 2656 8092 2660 8148
rect 2660 8092 2716 8148
rect 2716 8092 2720 8148
rect 2656 8088 2720 8092
rect 2736 8148 2800 8152
rect 2736 8092 2740 8148
rect 2740 8092 2796 8148
rect 2796 8092 2800 8148
rect 2736 8088 2800 8092
rect 2816 8148 2880 8152
rect 2816 8092 2820 8148
rect 2820 8092 2876 8148
rect 2876 8092 2880 8148
rect 2816 8088 2880 8092
rect 7848 8148 7912 8152
rect 7848 8092 7852 8148
rect 7852 8092 7908 8148
rect 7908 8092 7912 8148
rect 7848 8088 7912 8092
rect 7928 8148 7992 8152
rect 7928 8092 7932 8148
rect 7932 8092 7988 8148
rect 7988 8092 7992 8148
rect 7928 8088 7992 8092
rect 8008 8148 8072 8152
rect 8008 8092 8012 8148
rect 8012 8092 8068 8148
rect 8068 8092 8072 8148
rect 8008 8088 8072 8092
rect 8088 8148 8152 8152
rect 8088 8092 8092 8148
rect 8092 8092 8148 8148
rect 8148 8092 8152 8148
rect 8088 8088 8152 8092
rect 13120 8148 13184 8152
rect 13120 8092 13124 8148
rect 13124 8092 13180 8148
rect 13180 8092 13184 8148
rect 13120 8088 13184 8092
rect 13200 8148 13264 8152
rect 13200 8092 13204 8148
rect 13204 8092 13260 8148
rect 13260 8092 13264 8148
rect 13200 8088 13264 8092
rect 13280 8148 13344 8152
rect 13280 8092 13284 8148
rect 13284 8092 13340 8148
rect 13340 8092 13344 8148
rect 13280 8088 13344 8092
rect 13360 8148 13424 8152
rect 13360 8092 13364 8148
rect 13364 8092 13420 8148
rect 13420 8092 13424 8148
rect 13360 8088 13424 8092
rect 5212 7604 5276 7608
rect 5212 7548 5216 7604
rect 5216 7548 5272 7604
rect 5272 7548 5276 7604
rect 5212 7544 5276 7548
rect 5292 7604 5356 7608
rect 5292 7548 5296 7604
rect 5296 7548 5352 7604
rect 5352 7548 5356 7604
rect 5292 7544 5356 7548
rect 5372 7604 5436 7608
rect 5372 7548 5376 7604
rect 5376 7548 5432 7604
rect 5432 7548 5436 7604
rect 5372 7544 5436 7548
rect 5452 7604 5516 7608
rect 5452 7548 5456 7604
rect 5456 7548 5512 7604
rect 5512 7548 5516 7604
rect 5452 7544 5516 7548
rect 10484 7604 10548 7608
rect 10484 7548 10488 7604
rect 10488 7548 10544 7604
rect 10544 7548 10548 7604
rect 10484 7544 10548 7548
rect 10564 7604 10628 7608
rect 10564 7548 10568 7604
rect 10568 7548 10624 7604
rect 10624 7548 10628 7604
rect 10564 7544 10628 7548
rect 10644 7604 10708 7608
rect 10644 7548 10648 7604
rect 10648 7548 10704 7604
rect 10704 7548 10708 7604
rect 10644 7544 10708 7548
rect 10724 7604 10788 7608
rect 10724 7548 10728 7604
rect 10728 7548 10784 7604
rect 10784 7548 10788 7604
rect 10724 7544 10788 7548
rect 2576 7060 2640 7064
rect 2576 7004 2580 7060
rect 2580 7004 2636 7060
rect 2636 7004 2640 7060
rect 2576 7000 2640 7004
rect 2656 7060 2720 7064
rect 2656 7004 2660 7060
rect 2660 7004 2716 7060
rect 2716 7004 2720 7060
rect 2656 7000 2720 7004
rect 2736 7060 2800 7064
rect 2736 7004 2740 7060
rect 2740 7004 2796 7060
rect 2796 7004 2800 7060
rect 2736 7000 2800 7004
rect 2816 7060 2880 7064
rect 2816 7004 2820 7060
rect 2820 7004 2876 7060
rect 2876 7004 2880 7060
rect 2816 7000 2880 7004
rect 7848 7060 7912 7064
rect 7848 7004 7852 7060
rect 7852 7004 7908 7060
rect 7908 7004 7912 7060
rect 7848 7000 7912 7004
rect 7928 7060 7992 7064
rect 7928 7004 7932 7060
rect 7932 7004 7988 7060
rect 7988 7004 7992 7060
rect 7928 7000 7992 7004
rect 8008 7060 8072 7064
rect 8008 7004 8012 7060
rect 8012 7004 8068 7060
rect 8068 7004 8072 7060
rect 8008 7000 8072 7004
rect 8088 7060 8152 7064
rect 8088 7004 8092 7060
rect 8092 7004 8148 7060
rect 8148 7004 8152 7060
rect 8088 7000 8152 7004
rect 13120 7060 13184 7064
rect 13120 7004 13124 7060
rect 13124 7004 13180 7060
rect 13180 7004 13184 7060
rect 13120 7000 13184 7004
rect 13200 7060 13264 7064
rect 13200 7004 13204 7060
rect 13204 7004 13260 7060
rect 13260 7004 13264 7060
rect 13200 7000 13264 7004
rect 13280 7060 13344 7064
rect 13280 7004 13284 7060
rect 13284 7004 13340 7060
rect 13340 7004 13344 7060
rect 13280 7000 13344 7004
rect 13360 7060 13424 7064
rect 13360 7004 13364 7060
rect 13364 7004 13420 7060
rect 13420 7004 13424 7060
rect 13360 7000 13424 7004
rect 5212 6516 5276 6520
rect 5212 6460 5216 6516
rect 5216 6460 5272 6516
rect 5272 6460 5276 6516
rect 5212 6456 5276 6460
rect 5292 6516 5356 6520
rect 5292 6460 5296 6516
rect 5296 6460 5352 6516
rect 5352 6460 5356 6516
rect 5292 6456 5356 6460
rect 5372 6516 5436 6520
rect 5372 6460 5376 6516
rect 5376 6460 5432 6516
rect 5432 6460 5436 6516
rect 5372 6456 5436 6460
rect 5452 6516 5516 6520
rect 5452 6460 5456 6516
rect 5456 6460 5512 6516
rect 5512 6460 5516 6516
rect 5452 6456 5516 6460
rect 10484 6516 10548 6520
rect 10484 6460 10488 6516
rect 10488 6460 10544 6516
rect 10544 6460 10548 6516
rect 10484 6456 10548 6460
rect 10564 6516 10628 6520
rect 10564 6460 10568 6516
rect 10568 6460 10624 6516
rect 10624 6460 10628 6516
rect 10564 6456 10628 6460
rect 10644 6516 10708 6520
rect 10644 6460 10648 6516
rect 10648 6460 10704 6516
rect 10704 6460 10708 6516
rect 10644 6456 10708 6460
rect 10724 6516 10788 6520
rect 10724 6460 10728 6516
rect 10728 6460 10784 6516
rect 10784 6460 10788 6516
rect 10724 6456 10788 6460
rect 2576 5972 2640 5976
rect 2576 5916 2580 5972
rect 2580 5916 2636 5972
rect 2636 5916 2640 5972
rect 2576 5912 2640 5916
rect 2656 5972 2720 5976
rect 2656 5916 2660 5972
rect 2660 5916 2716 5972
rect 2716 5916 2720 5972
rect 2656 5912 2720 5916
rect 2736 5972 2800 5976
rect 2736 5916 2740 5972
rect 2740 5916 2796 5972
rect 2796 5916 2800 5972
rect 2736 5912 2800 5916
rect 2816 5972 2880 5976
rect 2816 5916 2820 5972
rect 2820 5916 2876 5972
rect 2876 5916 2880 5972
rect 2816 5912 2880 5916
rect 7848 5972 7912 5976
rect 7848 5916 7852 5972
rect 7852 5916 7908 5972
rect 7908 5916 7912 5972
rect 7848 5912 7912 5916
rect 7928 5972 7992 5976
rect 7928 5916 7932 5972
rect 7932 5916 7988 5972
rect 7988 5916 7992 5972
rect 7928 5912 7992 5916
rect 8008 5972 8072 5976
rect 8008 5916 8012 5972
rect 8012 5916 8068 5972
rect 8068 5916 8072 5972
rect 8008 5912 8072 5916
rect 8088 5972 8152 5976
rect 8088 5916 8092 5972
rect 8092 5916 8148 5972
rect 8148 5916 8152 5972
rect 8088 5912 8152 5916
rect 13120 5972 13184 5976
rect 13120 5916 13124 5972
rect 13124 5916 13180 5972
rect 13180 5916 13184 5972
rect 13120 5912 13184 5916
rect 13200 5972 13264 5976
rect 13200 5916 13204 5972
rect 13204 5916 13260 5972
rect 13260 5916 13264 5972
rect 13200 5912 13264 5916
rect 13280 5972 13344 5976
rect 13280 5916 13284 5972
rect 13284 5916 13340 5972
rect 13340 5916 13344 5972
rect 13280 5912 13344 5916
rect 13360 5972 13424 5976
rect 13360 5916 13364 5972
rect 13364 5916 13420 5972
rect 13420 5916 13424 5972
rect 13360 5912 13424 5916
rect 5212 5428 5276 5432
rect 5212 5372 5216 5428
rect 5216 5372 5272 5428
rect 5272 5372 5276 5428
rect 5212 5368 5276 5372
rect 5292 5428 5356 5432
rect 5292 5372 5296 5428
rect 5296 5372 5352 5428
rect 5352 5372 5356 5428
rect 5292 5368 5356 5372
rect 5372 5428 5436 5432
rect 5372 5372 5376 5428
rect 5376 5372 5432 5428
rect 5432 5372 5436 5428
rect 5372 5368 5436 5372
rect 5452 5428 5516 5432
rect 5452 5372 5456 5428
rect 5456 5372 5512 5428
rect 5512 5372 5516 5428
rect 5452 5368 5516 5372
rect 10484 5428 10548 5432
rect 10484 5372 10488 5428
rect 10488 5372 10544 5428
rect 10544 5372 10548 5428
rect 10484 5368 10548 5372
rect 10564 5428 10628 5432
rect 10564 5372 10568 5428
rect 10568 5372 10624 5428
rect 10624 5372 10628 5428
rect 10564 5368 10628 5372
rect 10644 5428 10708 5432
rect 10644 5372 10648 5428
rect 10648 5372 10704 5428
rect 10704 5372 10708 5428
rect 10644 5368 10708 5372
rect 10724 5428 10788 5432
rect 10724 5372 10728 5428
rect 10728 5372 10784 5428
rect 10784 5372 10788 5428
rect 10724 5368 10788 5372
rect 2576 4884 2640 4888
rect 2576 4828 2580 4884
rect 2580 4828 2636 4884
rect 2636 4828 2640 4884
rect 2576 4824 2640 4828
rect 2656 4884 2720 4888
rect 2656 4828 2660 4884
rect 2660 4828 2716 4884
rect 2716 4828 2720 4884
rect 2656 4824 2720 4828
rect 2736 4884 2800 4888
rect 2736 4828 2740 4884
rect 2740 4828 2796 4884
rect 2796 4828 2800 4884
rect 2736 4824 2800 4828
rect 2816 4884 2880 4888
rect 2816 4828 2820 4884
rect 2820 4828 2876 4884
rect 2876 4828 2880 4884
rect 2816 4824 2880 4828
rect 7848 4884 7912 4888
rect 7848 4828 7852 4884
rect 7852 4828 7908 4884
rect 7908 4828 7912 4884
rect 7848 4824 7912 4828
rect 7928 4884 7992 4888
rect 7928 4828 7932 4884
rect 7932 4828 7988 4884
rect 7988 4828 7992 4884
rect 7928 4824 7992 4828
rect 8008 4884 8072 4888
rect 8008 4828 8012 4884
rect 8012 4828 8068 4884
rect 8068 4828 8072 4884
rect 8008 4824 8072 4828
rect 8088 4884 8152 4888
rect 8088 4828 8092 4884
rect 8092 4828 8148 4884
rect 8148 4828 8152 4884
rect 8088 4824 8152 4828
rect 13120 4884 13184 4888
rect 13120 4828 13124 4884
rect 13124 4828 13180 4884
rect 13180 4828 13184 4884
rect 13120 4824 13184 4828
rect 13200 4884 13264 4888
rect 13200 4828 13204 4884
rect 13204 4828 13260 4884
rect 13260 4828 13264 4884
rect 13200 4824 13264 4828
rect 13280 4884 13344 4888
rect 13280 4828 13284 4884
rect 13284 4828 13340 4884
rect 13340 4828 13344 4884
rect 13280 4824 13344 4828
rect 13360 4884 13424 4888
rect 13360 4828 13364 4884
rect 13364 4828 13420 4884
rect 13420 4828 13424 4884
rect 13360 4824 13424 4828
rect 5212 4340 5276 4344
rect 5212 4284 5216 4340
rect 5216 4284 5272 4340
rect 5272 4284 5276 4340
rect 5212 4280 5276 4284
rect 5292 4340 5356 4344
rect 5292 4284 5296 4340
rect 5296 4284 5352 4340
rect 5352 4284 5356 4340
rect 5292 4280 5356 4284
rect 5372 4340 5436 4344
rect 5372 4284 5376 4340
rect 5376 4284 5432 4340
rect 5432 4284 5436 4340
rect 5372 4280 5436 4284
rect 5452 4340 5516 4344
rect 5452 4284 5456 4340
rect 5456 4284 5512 4340
rect 5512 4284 5516 4340
rect 5452 4280 5516 4284
rect 10484 4340 10548 4344
rect 10484 4284 10488 4340
rect 10488 4284 10544 4340
rect 10544 4284 10548 4340
rect 10484 4280 10548 4284
rect 10564 4340 10628 4344
rect 10564 4284 10568 4340
rect 10568 4284 10624 4340
rect 10624 4284 10628 4340
rect 10564 4280 10628 4284
rect 10644 4340 10708 4344
rect 10644 4284 10648 4340
rect 10648 4284 10704 4340
rect 10704 4284 10708 4340
rect 10644 4280 10708 4284
rect 10724 4340 10788 4344
rect 10724 4284 10728 4340
rect 10728 4284 10784 4340
rect 10784 4284 10788 4340
rect 10724 4280 10788 4284
rect 2576 3796 2640 3800
rect 2576 3740 2580 3796
rect 2580 3740 2636 3796
rect 2636 3740 2640 3796
rect 2576 3736 2640 3740
rect 2656 3796 2720 3800
rect 2656 3740 2660 3796
rect 2660 3740 2716 3796
rect 2716 3740 2720 3796
rect 2656 3736 2720 3740
rect 2736 3796 2800 3800
rect 2736 3740 2740 3796
rect 2740 3740 2796 3796
rect 2796 3740 2800 3796
rect 2736 3736 2800 3740
rect 2816 3796 2880 3800
rect 2816 3740 2820 3796
rect 2820 3740 2876 3796
rect 2876 3740 2880 3796
rect 2816 3736 2880 3740
rect 7848 3796 7912 3800
rect 7848 3740 7852 3796
rect 7852 3740 7908 3796
rect 7908 3740 7912 3796
rect 7848 3736 7912 3740
rect 7928 3796 7992 3800
rect 7928 3740 7932 3796
rect 7932 3740 7988 3796
rect 7988 3740 7992 3796
rect 7928 3736 7992 3740
rect 8008 3796 8072 3800
rect 8008 3740 8012 3796
rect 8012 3740 8068 3796
rect 8068 3740 8072 3796
rect 8008 3736 8072 3740
rect 8088 3796 8152 3800
rect 8088 3740 8092 3796
rect 8092 3740 8148 3796
rect 8148 3740 8152 3796
rect 8088 3736 8152 3740
rect 13120 3796 13184 3800
rect 13120 3740 13124 3796
rect 13124 3740 13180 3796
rect 13180 3740 13184 3796
rect 13120 3736 13184 3740
rect 13200 3796 13264 3800
rect 13200 3740 13204 3796
rect 13204 3740 13260 3796
rect 13260 3740 13264 3796
rect 13200 3736 13264 3740
rect 13280 3796 13344 3800
rect 13280 3740 13284 3796
rect 13284 3740 13340 3796
rect 13340 3740 13344 3796
rect 13280 3736 13344 3740
rect 13360 3796 13424 3800
rect 13360 3740 13364 3796
rect 13364 3740 13420 3796
rect 13420 3740 13424 3796
rect 13360 3736 13424 3740
rect 5212 3252 5276 3256
rect 5212 3196 5216 3252
rect 5216 3196 5272 3252
rect 5272 3196 5276 3252
rect 5212 3192 5276 3196
rect 5292 3252 5356 3256
rect 5292 3196 5296 3252
rect 5296 3196 5352 3252
rect 5352 3196 5356 3252
rect 5292 3192 5356 3196
rect 5372 3252 5436 3256
rect 5372 3196 5376 3252
rect 5376 3196 5432 3252
rect 5432 3196 5436 3252
rect 5372 3192 5436 3196
rect 5452 3252 5516 3256
rect 5452 3196 5456 3252
rect 5456 3196 5512 3252
rect 5512 3196 5516 3252
rect 5452 3192 5516 3196
rect 10484 3252 10548 3256
rect 10484 3196 10488 3252
rect 10488 3196 10544 3252
rect 10544 3196 10548 3252
rect 10484 3192 10548 3196
rect 10564 3252 10628 3256
rect 10564 3196 10568 3252
rect 10568 3196 10624 3252
rect 10624 3196 10628 3252
rect 10564 3192 10628 3196
rect 10644 3252 10708 3256
rect 10644 3196 10648 3252
rect 10648 3196 10704 3252
rect 10704 3196 10708 3252
rect 10644 3192 10708 3196
rect 10724 3252 10788 3256
rect 10724 3196 10728 3252
rect 10728 3196 10784 3252
rect 10784 3196 10788 3252
rect 10724 3192 10788 3196
rect 2576 2708 2640 2712
rect 2576 2652 2580 2708
rect 2580 2652 2636 2708
rect 2636 2652 2640 2708
rect 2576 2648 2640 2652
rect 2656 2708 2720 2712
rect 2656 2652 2660 2708
rect 2660 2652 2716 2708
rect 2716 2652 2720 2708
rect 2656 2648 2720 2652
rect 2736 2708 2800 2712
rect 2736 2652 2740 2708
rect 2740 2652 2796 2708
rect 2796 2652 2800 2708
rect 2736 2648 2800 2652
rect 2816 2708 2880 2712
rect 2816 2652 2820 2708
rect 2820 2652 2876 2708
rect 2876 2652 2880 2708
rect 2816 2648 2880 2652
rect 7848 2708 7912 2712
rect 7848 2652 7852 2708
rect 7852 2652 7908 2708
rect 7908 2652 7912 2708
rect 7848 2648 7912 2652
rect 7928 2708 7992 2712
rect 7928 2652 7932 2708
rect 7932 2652 7988 2708
rect 7988 2652 7992 2708
rect 7928 2648 7992 2652
rect 8008 2708 8072 2712
rect 8008 2652 8012 2708
rect 8012 2652 8068 2708
rect 8068 2652 8072 2708
rect 8008 2648 8072 2652
rect 8088 2708 8152 2712
rect 8088 2652 8092 2708
rect 8092 2652 8148 2708
rect 8148 2652 8152 2708
rect 8088 2648 8152 2652
rect 13120 2708 13184 2712
rect 13120 2652 13124 2708
rect 13124 2652 13180 2708
rect 13180 2652 13184 2708
rect 13120 2648 13184 2652
rect 13200 2708 13264 2712
rect 13200 2652 13204 2708
rect 13204 2652 13260 2708
rect 13260 2652 13264 2708
rect 13200 2648 13264 2652
rect 13280 2708 13344 2712
rect 13280 2652 13284 2708
rect 13284 2652 13340 2708
rect 13340 2652 13344 2708
rect 13280 2648 13344 2652
rect 13360 2708 13424 2712
rect 13360 2652 13364 2708
rect 13364 2652 13420 2708
rect 13420 2652 13424 2708
rect 13360 2648 13424 2652
rect 5212 2164 5276 2168
rect 5212 2108 5216 2164
rect 5216 2108 5272 2164
rect 5272 2108 5276 2164
rect 5212 2104 5276 2108
rect 5292 2164 5356 2168
rect 5292 2108 5296 2164
rect 5296 2108 5352 2164
rect 5352 2108 5356 2164
rect 5292 2104 5356 2108
rect 5372 2164 5436 2168
rect 5372 2108 5376 2164
rect 5376 2108 5432 2164
rect 5432 2108 5436 2164
rect 5372 2104 5436 2108
rect 5452 2164 5516 2168
rect 5452 2108 5456 2164
rect 5456 2108 5512 2164
rect 5512 2108 5516 2164
rect 5452 2104 5516 2108
rect 10484 2164 10548 2168
rect 10484 2108 10488 2164
rect 10488 2108 10544 2164
rect 10544 2108 10548 2164
rect 10484 2104 10548 2108
rect 10564 2164 10628 2168
rect 10564 2108 10568 2164
rect 10568 2108 10624 2164
rect 10624 2108 10628 2164
rect 10564 2104 10628 2108
rect 10644 2164 10708 2168
rect 10644 2108 10648 2164
rect 10648 2108 10704 2164
rect 10704 2108 10708 2164
rect 10644 2104 10708 2108
rect 10724 2164 10788 2168
rect 10724 2108 10728 2164
rect 10728 2108 10784 2164
rect 10784 2108 10788 2164
rect 10724 2104 10788 2108
rect 2576 1620 2640 1624
rect 2576 1564 2580 1620
rect 2580 1564 2636 1620
rect 2636 1564 2640 1620
rect 2576 1560 2640 1564
rect 2656 1620 2720 1624
rect 2656 1564 2660 1620
rect 2660 1564 2716 1620
rect 2716 1564 2720 1620
rect 2656 1560 2720 1564
rect 2736 1620 2800 1624
rect 2736 1564 2740 1620
rect 2740 1564 2796 1620
rect 2796 1564 2800 1620
rect 2736 1560 2800 1564
rect 2816 1620 2880 1624
rect 2816 1564 2820 1620
rect 2820 1564 2876 1620
rect 2876 1564 2880 1620
rect 2816 1560 2880 1564
rect 7848 1620 7912 1624
rect 7848 1564 7852 1620
rect 7852 1564 7908 1620
rect 7908 1564 7912 1620
rect 7848 1560 7912 1564
rect 7928 1620 7992 1624
rect 7928 1564 7932 1620
rect 7932 1564 7988 1620
rect 7988 1564 7992 1620
rect 7928 1560 7992 1564
rect 8008 1620 8072 1624
rect 8008 1564 8012 1620
rect 8012 1564 8068 1620
rect 8068 1564 8072 1620
rect 8008 1560 8072 1564
rect 8088 1620 8152 1624
rect 8088 1564 8092 1620
rect 8092 1564 8148 1620
rect 8148 1564 8152 1620
rect 8088 1560 8152 1564
rect 13120 1620 13184 1624
rect 13120 1564 13124 1620
rect 13124 1564 13180 1620
rect 13180 1564 13184 1620
rect 13120 1560 13184 1564
rect 13200 1620 13264 1624
rect 13200 1564 13204 1620
rect 13204 1564 13260 1620
rect 13260 1564 13264 1620
rect 13200 1560 13264 1564
rect 13280 1620 13344 1624
rect 13280 1564 13284 1620
rect 13284 1564 13340 1620
rect 13340 1564 13344 1620
rect 13280 1560 13344 1564
rect 13360 1620 13424 1624
rect 13360 1564 13364 1620
rect 13364 1564 13420 1620
rect 13420 1564 13424 1620
rect 13360 1560 13424 1564
rect 5212 1076 5276 1080
rect 5212 1020 5216 1076
rect 5216 1020 5272 1076
rect 5272 1020 5276 1076
rect 5212 1016 5276 1020
rect 5292 1076 5356 1080
rect 5292 1020 5296 1076
rect 5296 1020 5352 1076
rect 5352 1020 5356 1076
rect 5292 1016 5356 1020
rect 5372 1076 5436 1080
rect 5372 1020 5376 1076
rect 5376 1020 5432 1076
rect 5432 1020 5436 1076
rect 5372 1016 5436 1020
rect 5452 1076 5516 1080
rect 5452 1020 5456 1076
rect 5456 1020 5512 1076
rect 5512 1020 5516 1076
rect 5452 1016 5516 1020
rect 10484 1076 10548 1080
rect 10484 1020 10488 1076
rect 10488 1020 10544 1076
rect 10544 1020 10548 1076
rect 10484 1016 10548 1020
rect 10564 1076 10628 1080
rect 10564 1020 10568 1076
rect 10568 1020 10624 1076
rect 10624 1020 10628 1076
rect 10564 1016 10628 1020
rect 10644 1076 10708 1080
rect 10644 1020 10648 1076
rect 10648 1020 10704 1076
rect 10704 1020 10708 1076
rect 10644 1016 10708 1020
rect 10724 1076 10788 1080
rect 10724 1020 10728 1076
rect 10728 1020 10784 1076
rect 10784 1020 10788 1076
rect 10724 1016 10788 1020
rect 2576 532 2640 536
rect 2576 476 2580 532
rect 2580 476 2636 532
rect 2636 476 2640 532
rect 2576 472 2640 476
rect 2656 532 2720 536
rect 2656 476 2660 532
rect 2660 476 2716 532
rect 2716 476 2720 532
rect 2656 472 2720 476
rect 2736 532 2800 536
rect 2736 476 2740 532
rect 2740 476 2796 532
rect 2796 476 2800 532
rect 2736 472 2800 476
rect 2816 532 2880 536
rect 2816 476 2820 532
rect 2820 476 2876 532
rect 2876 476 2880 532
rect 2816 472 2880 476
rect 7848 532 7912 536
rect 7848 476 7852 532
rect 7852 476 7908 532
rect 7908 476 7912 532
rect 7848 472 7912 476
rect 7928 532 7992 536
rect 7928 476 7932 532
rect 7932 476 7988 532
rect 7988 476 7992 532
rect 7928 472 7992 476
rect 8008 532 8072 536
rect 8008 476 8012 532
rect 8012 476 8068 532
rect 8068 476 8072 532
rect 8008 472 8072 476
rect 8088 532 8152 536
rect 8088 476 8092 532
rect 8092 476 8148 532
rect 8148 476 8152 532
rect 8088 472 8152 476
rect 13120 532 13184 536
rect 13120 476 13124 532
rect 13124 476 13180 532
rect 13180 476 13184 532
rect 13120 472 13184 476
rect 13200 532 13264 536
rect 13200 476 13204 532
rect 13204 476 13260 532
rect 13260 476 13264 532
rect 13200 472 13264 476
rect 13280 532 13344 536
rect 13280 476 13284 532
rect 13284 476 13340 532
rect 13340 476 13344 532
rect 13280 472 13344 476
rect 13360 532 13424 536
rect 13360 476 13364 532
rect 13364 476 13420 532
rect 13420 476 13424 532
rect 13360 472 13424 476
<< metal4 >>
rect 2568 12504 2888 13064
rect 2568 12440 2576 12504
rect 2640 12440 2656 12504
rect 2720 12440 2736 12504
rect 2800 12440 2816 12504
rect 2880 12440 2888 12504
rect 2568 11416 2888 12440
rect 2568 11352 2576 11416
rect 2640 11352 2656 11416
rect 2720 11352 2736 11416
rect 2800 11352 2816 11416
rect 2880 11352 2888 11416
rect 2568 11334 2888 11352
rect 2568 11098 2610 11334
rect 2846 11098 2888 11334
rect 2568 10328 2888 11098
rect 2568 10264 2576 10328
rect 2640 10264 2656 10328
rect 2720 10264 2736 10328
rect 2800 10264 2816 10328
rect 2880 10264 2888 10328
rect 2568 9240 2888 10264
rect 2568 9176 2576 9240
rect 2640 9176 2656 9240
rect 2720 9176 2736 9240
rect 2800 9176 2816 9240
rect 2880 9176 2888 9240
rect 2568 8152 2888 9176
rect 2568 8088 2576 8152
rect 2640 8088 2656 8152
rect 2720 8088 2736 8152
rect 2800 8088 2816 8152
rect 2880 8088 2888 8152
rect 2568 7064 2888 8088
rect 2568 7000 2576 7064
rect 2640 7030 2656 7064
rect 2720 7030 2736 7064
rect 2800 7030 2816 7064
rect 2880 7000 2888 7064
rect 2568 6794 2610 7000
rect 2846 6794 2888 7000
rect 2568 5976 2888 6794
rect 2568 5912 2576 5976
rect 2640 5912 2656 5976
rect 2720 5912 2736 5976
rect 2800 5912 2816 5976
rect 2880 5912 2888 5976
rect 2568 4888 2888 5912
rect 2568 4824 2576 4888
rect 2640 4824 2656 4888
rect 2720 4824 2736 4888
rect 2800 4824 2816 4888
rect 2880 4824 2888 4888
rect 2568 3800 2888 4824
rect 2568 3736 2576 3800
rect 2640 3736 2656 3800
rect 2720 3736 2736 3800
rect 2800 3736 2816 3800
rect 2880 3736 2888 3800
rect 2568 2726 2888 3736
rect 2568 2712 2610 2726
rect 2846 2712 2888 2726
rect 2568 2648 2576 2712
rect 2880 2648 2888 2712
rect 2568 2490 2610 2648
rect 2846 2490 2888 2648
rect 2568 1624 2888 2490
rect 2568 1560 2576 1624
rect 2640 1560 2656 1624
rect 2720 1560 2736 1624
rect 2800 1560 2816 1624
rect 2880 1560 2888 1624
rect 2568 536 2888 1560
rect 2568 472 2576 536
rect 2640 472 2656 536
rect 2720 472 2736 536
rect 2800 472 2816 536
rect 2880 472 2888 536
rect 2568 456 2888 472
rect 5204 13048 5524 13064
rect 5204 12984 5212 13048
rect 5276 12984 5292 13048
rect 5356 12984 5372 13048
rect 5436 12984 5452 13048
rect 5516 12984 5524 13048
rect 5204 11960 5524 12984
rect 5204 11896 5212 11960
rect 5276 11896 5292 11960
rect 5356 11896 5372 11960
rect 5436 11896 5452 11960
rect 5516 11896 5524 11960
rect 5204 10872 5524 11896
rect 5204 10808 5212 10872
rect 5276 10808 5292 10872
rect 5356 10808 5372 10872
rect 5436 10808 5452 10872
rect 5516 10808 5524 10872
rect 5204 9784 5524 10808
rect 5204 9720 5212 9784
rect 5276 9720 5292 9784
rect 5356 9720 5372 9784
rect 5436 9720 5452 9784
rect 5516 9720 5524 9784
rect 5204 9182 5524 9720
rect 5204 8946 5246 9182
rect 5482 8946 5524 9182
rect 5204 8696 5524 8946
rect 5204 8632 5212 8696
rect 5276 8632 5292 8696
rect 5356 8632 5372 8696
rect 5436 8632 5452 8696
rect 5516 8632 5524 8696
rect 5204 7608 5524 8632
rect 5204 7544 5212 7608
rect 5276 7544 5292 7608
rect 5356 7544 5372 7608
rect 5436 7544 5452 7608
rect 5516 7544 5524 7608
rect 5204 6520 5524 7544
rect 5204 6456 5212 6520
rect 5276 6456 5292 6520
rect 5356 6456 5372 6520
rect 5436 6456 5452 6520
rect 5516 6456 5524 6520
rect 5204 5432 5524 6456
rect 5204 5368 5212 5432
rect 5276 5368 5292 5432
rect 5356 5368 5372 5432
rect 5436 5368 5452 5432
rect 5516 5368 5524 5432
rect 5204 4878 5524 5368
rect 5204 4642 5246 4878
rect 5482 4642 5524 4878
rect 5204 4344 5524 4642
rect 5204 4280 5212 4344
rect 5276 4280 5292 4344
rect 5356 4280 5372 4344
rect 5436 4280 5452 4344
rect 5516 4280 5524 4344
rect 5204 3256 5524 4280
rect 5204 3192 5212 3256
rect 5276 3192 5292 3256
rect 5356 3192 5372 3256
rect 5436 3192 5452 3256
rect 5516 3192 5524 3256
rect 5204 2168 5524 3192
rect 5204 2104 5212 2168
rect 5276 2104 5292 2168
rect 5356 2104 5372 2168
rect 5436 2104 5452 2168
rect 5516 2104 5524 2168
rect 5204 1080 5524 2104
rect 5204 1016 5212 1080
rect 5276 1016 5292 1080
rect 5356 1016 5372 1080
rect 5436 1016 5452 1080
rect 5516 1016 5524 1080
rect 5204 456 5524 1016
rect 7840 12504 8160 13064
rect 7840 12440 7848 12504
rect 7912 12440 7928 12504
rect 7992 12440 8008 12504
rect 8072 12440 8088 12504
rect 8152 12440 8160 12504
rect 7840 11416 8160 12440
rect 7840 11352 7848 11416
rect 7912 11352 7928 11416
rect 7992 11352 8008 11416
rect 8072 11352 8088 11416
rect 8152 11352 8160 11416
rect 7840 11334 8160 11352
rect 7840 11098 7882 11334
rect 8118 11098 8160 11334
rect 7840 10328 8160 11098
rect 7840 10264 7848 10328
rect 7912 10264 7928 10328
rect 7992 10264 8008 10328
rect 8072 10264 8088 10328
rect 8152 10264 8160 10328
rect 7840 9240 8160 10264
rect 7840 9176 7848 9240
rect 7912 9176 7928 9240
rect 7992 9176 8008 9240
rect 8072 9176 8088 9240
rect 8152 9176 8160 9240
rect 7840 8152 8160 9176
rect 7840 8088 7848 8152
rect 7912 8088 7928 8152
rect 7992 8088 8008 8152
rect 8072 8088 8088 8152
rect 8152 8088 8160 8152
rect 7840 7064 8160 8088
rect 7840 7000 7848 7064
rect 7912 7030 7928 7064
rect 7992 7030 8008 7064
rect 8072 7030 8088 7064
rect 8152 7000 8160 7064
rect 7840 6794 7882 7000
rect 8118 6794 8160 7000
rect 7840 5976 8160 6794
rect 7840 5912 7848 5976
rect 7912 5912 7928 5976
rect 7992 5912 8008 5976
rect 8072 5912 8088 5976
rect 8152 5912 8160 5976
rect 7840 4888 8160 5912
rect 7840 4824 7848 4888
rect 7912 4824 7928 4888
rect 7992 4824 8008 4888
rect 8072 4824 8088 4888
rect 8152 4824 8160 4888
rect 7840 3800 8160 4824
rect 7840 3736 7848 3800
rect 7912 3736 7928 3800
rect 7992 3736 8008 3800
rect 8072 3736 8088 3800
rect 8152 3736 8160 3800
rect 7840 2726 8160 3736
rect 7840 2712 7882 2726
rect 8118 2712 8160 2726
rect 7840 2648 7848 2712
rect 8152 2648 8160 2712
rect 7840 2490 7882 2648
rect 8118 2490 8160 2648
rect 7840 1624 8160 2490
rect 7840 1560 7848 1624
rect 7912 1560 7928 1624
rect 7992 1560 8008 1624
rect 8072 1560 8088 1624
rect 8152 1560 8160 1624
rect 7840 536 8160 1560
rect 7840 472 7848 536
rect 7912 472 7928 536
rect 7992 472 8008 536
rect 8072 472 8088 536
rect 8152 472 8160 536
rect 7840 456 8160 472
rect 10476 13048 10796 13064
rect 10476 12984 10484 13048
rect 10548 12984 10564 13048
rect 10628 12984 10644 13048
rect 10708 12984 10724 13048
rect 10788 12984 10796 13048
rect 10476 11960 10796 12984
rect 10476 11896 10484 11960
rect 10548 11896 10564 11960
rect 10628 11896 10644 11960
rect 10708 11896 10724 11960
rect 10788 11896 10796 11960
rect 10476 10872 10796 11896
rect 10476 10808 10484 10872
rect 10548 10808 10564 10872
rect 10628 10808 10644 10872
rect 10708 10808 10724 10872
rect 10788 10808 10796 10872
rect 10476 9784 10796 10808
rect 10476 9720 10484 9784
rect 10548 9720 10564 9784
rect 10628 9720 10644 9784
rect 10708 9720 10724 9784
rect 10788 9720 10796 9784
rect 10476 9182 10796 9720
rect 10476 8946 10518 9182
rect 10754 8946 10796 9182
rect 10476 8696 10796 8946
rect 10476 8632 10484 8696
rect 10548 8632 10564 8696
rect 10628 8632 10644 8696
rect 10708 8632 10724 8696
rect 10788 8632 10796 8696
rect 10476 7608 10796 8632
rect 10476 7544 10484 7608
rect 10548 7544 10564 7608
rect 10628 7544 10644 7608
rect 10708 7544 10724 7608
rect 10788 7544 10796 7608
rect 10476 6520 10796 7544
rect 10476 6456 10484 6520
rect 10548 6456 10564 6520
rect 10628 6456 10644 6520
rect 10708 6456 10724 6520
rect 10788 6456 10796 6520
rect 10476 5432 10796 6456
rect 10476 5368 10484 5432
rect 10548 5368 10564 5432
rect 10628 5368 10644 5432
rect 10708 5368 10724 5432
rect 10788 5368 10796 5432
rect 10476 4878 10796 5368
rect 10476 4642 10518 4878
rect 10754 4642 10796 4878
rect 10476 4344 10796 4642
rect 10476 4280 10484 4344
rect 10548 4280 10564 4344
rect 10628 4280 10644 4344
rect 10708 4280 10724 4344
rect 10788 4280 10796 4344
rect 10476 3256 10796 4280
rect 10476 3192 10484 3256
rect 10548 3192 10564 3256
rect 10628 3192 10644 3256
rect 10708 3192 10724 3256
rect 10788 3192 10796 3256
rect 10476 2168 10796 3192
rect 10476 2104 10484 2168
rect 10548 2104 10564 2168
rect 10628 2104 10644 2168
rect 10708 2104 10724 2168
rect 10788 2104 10796 2168
rect 10476 1080 10796 2104
rect 10476 1016 10484 1080
rect 10548 1016 10564 1080
rect 10628 1016 10644 1080
rect 10708 1016 10724 1080
rect 10788 1016 10796 1080
rect 10476 456 10796 1016
rect 13112 12504 13432 13064
rect 13112 12440 13120 12504
rect 13184 12440 13200 12504
rect 13264 12440 13280 12504
rect 13344 12440 13360 12504
rect 13424 12440 13432 12504
rect 13112 11416 13432 12440
rect 13112 11352 13120 11416
rect 13184 11352 13200 11416
rect 13264 11352 13280 11416
rect 13344 11352 13360 11416
rect 13424 11352 13432 11416
rect 13112 11334 13432 11352
rect 13112 11098 13154 11334
rect 13390 11098 13432 11334
rect 13112 10328 13432 11098
rect 13112 10264 13120 10328
rect 13184 10264 13200 10328
rect 13264 10264 13280 10328
rect 13344 10264 13360 10328
rect 13424 10264 13432 10328
rect 13112 9240 13432 10264
rect 13112 9176 13120 9240
rect 13184 9176 13200 9240
rect 13264 9176 13280 9240
rect 13344 9176 13360 9240
rect 13424 9176 13432 9240
rect 13112 8152 13432 9176
rect 13112 8088 13120 8152
rect 13184 8088 13200 8152
rect 13264 8088 13280 8152
rect 13344 8088 13360 8152
rect 13424 8088 13432 8152
rect 13112 7064 13432 8088
rect 13112 7000 13120 7064
rect 13184 7030 13200 7064
rect 13264 7030 13280 7064
rect 13344 7030 13360 7064
rect 13424 7000 13432 7064
rect 13112 6794 13154 7000
rect 13390 6794 13432 7000
rect 13112 5976 13432 6794
rect 13112 5912 13120 5976
rect 13184 5912 13200 5976
rect 13264 5912 13280 5976
rect 13344 5912 13360 5976
rect 13424 5912 13432 5976
rect 13112 4888 13432 5912
rect 13112 4824 13120 4888
rect 13184 4824 13200 4888
rect 13264 4824 13280 4888
rect 13344 4824 13360 4888
rect 13424 4824 13432 4888
rect 13112 3800 13432 4824
rect 13112 3736 13120 3800
rect 13184 3736 13200 3800
rect 13264 3736 13280 3800
rect 13344 3736 13360 3800
rect 13424 3736 13432 3800
rect 13112 2726 13432 3736
rect 13112 2712 13154 2726
rect 13390 2712 13432 2726
rect 13112 2648 13120 2712
rect 13424 2648 13432 2712
rect 13112 2490 13154 2648
rect 13390 2490 13432 2648
rect 13112 1624 13432 2490
rect 13112 1560 13120 1624
rect 13184 1560 13200 1624
rect 13264 1560 13280 1624
rect 13344 1560 13360 1624
rect 13424 1560 13432 1624
rect 13112 536 13432 1560
rect 13112 472 13120 536
rect 13184 472 13200 536
rect 13264 472 13280 536
rect 13344 472 13360 536
rect 13424 472 13432 536
rect 13112 456 13432 472
<< via4 >>
rect 2610 11098 2846 11334
rect 2610 7000 2640 7030
rect 2640 7000 2656 7030
rect 2656 7000 2720 7030
rect 2720 7000 2736 7030
rect 2736 7000 2800 7030
rect 2800 7000 2816 7030
rect 2816 7000 2846 7030
rect 2610 6794 2846 7000
rect 2610 2712 2846 2726
rect 2610 2648 2640 2712
rect 2640 2648 2656 2712
rect 2656 2648 2720 2712
rect 2720 2648 2736 2712
rect 2736 2648 2800 2712
rect 2800 2648 2816 2712
rect 2816 2648 2846 2712
rect 2610 2490 2846 2648
rect 5246 8946 5482 9182
rect 5246 4642 5482 4878
rect 7882 11098 8118 11334
rect 7882 7000 7912 7030
rect 7912 7000 7928 7030
rect 7928 7000 7992 7030
rect 7992 7000 8008 7030
rect 8008 7000 8072 7030
rect 8072 7000 8088 7030
rect 8088 7000 8118 7030
rect 7882 6794 8118 7000
rect 7882 2712 8118 2726
rect 7882 2648 7912 2712
rect 7912 2648 7928 2712
rect 7928 2648 7992 2712
rect 7992 2648 8008 2712
rect 8008 2648 8072 2712
rect 8072 2648 8088 2712
rect 8088 2648 8118 2712
rect 7882 2490 8118 2648
rect 10518 8946 10754 9182
rect 10518 4642 10754 4878
rect 13154 11098 13390 11334
rect 13154 7000 13184 7030
rect 13184 7000 13200 7030
rect 13200 7000 13264 7030
rect 13264 7000 13280 7030
rect 13280 7000 13344 7030
rect 13344 7000 13360 7030
rect 13360 7000 13390 7030
rect 13154 6794 13390 7000
rect 13154 2712 13390 2726
rect 13154 2648 13184 2712
rect 13184 2648 13200 2712
rect 13200 2648 13264 2712
rect 13264 2648 13280 2712
rect 13280 2648 13344 2712
rect 13344 2648 13360 2712
rect 13360 2648 13390 2712
rect 13154 2490 13390 2648
<< metal5 >>
rect 92 11334 15824 11376
rect 92 11098 2610 11334
rect 2846 11098 7882 11334
rect 8118 11098 13154 11334
rect 13390 11098 15824 11334
rect 92 11056 15824 11098
rect 92 9182 15824 9224
rect 92 8946 5246 9182
rect 5482 8946 10518 9182
rect 10754 8946 15824 9182
rect 92 8904 15824 8946
rect 92 7030 15824 7072
rect 92 6794 2610 7030
rect 2846 6794 7882 7030
rect 8118 6794 13154 7030
rect 13390 6794 15824 7030
rect 92 6752 15824 6794
rect 92 4878 15824 4920
rect 92 4642 5246 4878
rect 5482 4642 10518 4878
rect 10754 4642 15824 4878
rect 92 4600 15824 4642
rect 92 2726 15824 2768
rect 92 2490 2610 2726
rect 2846 2490 7882 2726
rect 8118 2490 13154 2726
rect 13390 2490 15824 2726
rect 92 2448 15824 2490
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1696364841
transform -1 0 3220 0 -1 7536
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1696364841
transform -1 0 6256 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1696364841
transform 1 0 3128 0 -1 3184
box -38 -88 314 552
use sky130_fd_sc_hd__and3_1  _143_
timestamp 1696364841
transform 1 0 3220 0 1 6528
box -38 -88 498 552
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1696364841
transform 1 0 4048 0 1 7616
box -38 -88 314 552
use sky130_fd_sc_hd__nand2_1  _145_
timestamp 1696364841
transform 1 0 2116 0 1 6528
box -38 -88 314 552
use sky130_fd_sc_hd__and3_2  _146_
timestamp 1696364841
transform 1 0 3312 0 1 5440
box -38 -88 590 552
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1696364841
transform 1 0 11868 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1696364841
transform 1 0 4140 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1696364841
transform 1 0 2024 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__or3_4  _150_
timestamp 1696364841
transform 1 0 3956 0 -1 5360
box -38 -88 866 552
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1696364841
transform 1 0 4692 0 -1 3184
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1696364841
transform -1 0 6992 0 -1 1008
box -38 -88 314 552
use sky130_fd_sc_hd__or4b_4  _153_
timestamp 1696364841
transform 1 0 5796 0 -1 2096
box -38 -88 1050 552
use sky130_fd_sc_hd__buf_1  _154_
timestamp 1696364841
transform 1 0 4048 0 -1 3184
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1696364841
transform -1 0 8740 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _156_
timestamp 1696364841
transform 1 0 8464 0 1 6528
box -38 -88 498 552
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1696364841
transform 1 0 9660 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1696364841
transform 1 0 13984 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1696364841
transform -1 0 14536 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1696364841
transform -1 0 15088 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1696364841
transform -1 0 12880 0 1 6528
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1696364841
transform -1 0 15088 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__o22a_1  _163_
timestamp 1696364841
transform 1 0 13708 0 1 7616
box -38 -88 682 552
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1696364841
transform 1 0 13708 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__o22a_1  _165_
timestamp 1696364841
transform 1 0 13708 0 1 8704
box -38 -88 682 552
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1696364841
transform -1 0 11316 0 -1 8624
box -38 -88 314 552
use sky130_fd_sc_hd__a22o_1  _167_
timestamp 1696364841
transform -1 0 12328 0 -1 8624
box -38 -88 682 552
use sky130_fd_sc_hd__a2bb2oi_1  _168_
timestamp 1696364841
transform -1 0 12144 0 1 6528
box -38 -88 682 552
use sky130_fd_sc_hd__nor2_1  _169_
timestamp 1696364841
transform -1 0 11684 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__a2bb2o_1  _170_
timestamp 1696364841
transform 1 0 11040 0 1 7616
box -38 -88 774 552
use sky130_fd_sc_hd__o22a_1  _171_
timestamp 1696364841
transform 1 0 13708 0 1 6528
box -38 -88 682 552
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1696364841
transform -1 0 13156 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__a2bb2o_1  _173_
timestamp 1696364841
transform -1 0 12880 0 1 7616
box -38 -88 774 552
use sky130_fd_sc_hd__a22o_1  _174_
timestamp 1696364841
transform 1 0 12696 0 -1 6448
box -38 -88 682 552
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1696364841
transform -1 0 2392 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1696364841
transform 1 0 1472 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1696364841
transform 1 0 1288 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__or3_4  _178_
timestamp 1696364841
transform 1 0 4232 0 1 5440
box -38 -88 866 552
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1696364841
transform -1 0 6348 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__or3_1  _180_
timestamp 1696364841
transform 1 0 4508 0 -1 6448
box -38 -88 498 552
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1696364841
transform -1 0 7176 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__o211a_1  _182_
timestamp 1696364841
transform 1 0 4048 0 -1 4272
box -38 -88 774 552
use sky130_fd_sc_hd__o221ai_4  _183_
timestamp 1696364841
transform -1 0 5980 0 1 6528
box -38 -88 1970 552
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1696364841
transform 1 0 3220 0 1 4352
box -38 -88 866 552
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1696364841
transform -1 0 1748 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__o21a_1  _186_
timestamp 1696364841
transform 1 0 3036 0 -1 5360
box -38 -88 590 552
use sky130_fd_sc_hd__buf_1  _187_
timestamp 1696364841
transform 1 0 3404 0 1 7616
box -38 -88 314 552
use sky130_fd_sc_hd__mux2_1  _188_
timestamp 1696364841
transform 1 0 3312 0 -1 6448
box -38 -88 866 552
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1696364841
transform -1 0 7176 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1696364841
transform 1 0 7544 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1696364841
transform -1 0 2392 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__or2_1  _192_
timestamp 1696364841
transform 1 0 7360 0 -1 4272
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1696364841
transform 1 0 11040 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__buf_1  _194_
timestamp 1696364841
transform 1 0 11040 0 -1 4272
box -38 -88 314 552
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1696364841
transform -1 0 9752 0 -1 1008
box -38 -88 682 552
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1696364841
transform 1 0 12052 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _197_
timestamp 1696364841
transform -1 0 8832 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__a32o_1  _198_
timestamp 1696364841
transform 1 0 9200 0 1 3264
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _199_
timestamp 1696364841
transform 1 0 11224 0 1 2176
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _200_
timestamp 1696364841
transform 1 0 11040 0 -1 3184
box -38 -88 774 552
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1696364841
transform 1 0 10304 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__a32o_1  _202_
timestamp 1696364841
transform 1 0 9384 0 -1 4272
box -38 -88 774 552
use sky130_fd_sc_hd__a31o_1  _203_
timestamp 1696364841
transform 1 0 6624 0 1 4352
box -38 -88 682 552
use sky130_fd_sc_hd__a31oi_2  _204_
timestamp 1696364841
transform 1 0 4048 0 -1 2096
box -38 -88 958 552
use sky130_fd_sc_hd__o21a_1  _205_
timestamp 1696364841
transform 1 0 3772 0 1 2176
box -38 -88 590 552
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1696364841
transform -1 0 1288 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__and3_1  _207_
timestamp 1696364841
transform -1 0 6348 0 -1 1008
box -38 -88 498 552
use sky130_fd_sc_hd__o22a_1  _208_
timestamp 1696364841
transform 1 0 4232 0 1 1088
box -38 -88 682 552
use sky130_fd_sc_hd__a22o_1  _209_
timestamp 1696364841
transform -1 0 6440 0 -1 3184
box -38 -88 682 552
use sky130_fd_sc_hd__o22ai_1  _210_
timestamp 1696364841
transform -1 0 5612 0 1 3264
box -38 -88 498 552
use sky130_fd_sc_hd__a22o_1  _211_
timestamp 1696364841
transform -1 0 7820 0 -1 2096
box -38 -88 682 552
use sky130_fd_sc_hd__buf_1  _212_
timestamp 1696364841
transform 1 0 3956 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1696364841
transform 1 0 7360 0 1 8704
box -38 -88 314 552
use sky130_fd_sc_hd__a22o_1  _214_
timestamp 1696364841
transform -1 0 6440 0 -1 10800
box -38 -88 682 552
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1696364841
transform 1 0 12512 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  _216_
timestamp 1696364841
transform 1 0 6440 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  _217_
timestamp 1696364841
transform 1 0 4600 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__a32o_1  _218_
timestamp 1696364841
transform 1 0 6900 0 1 10880
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _219_
timestamp 1696364841
transform 1 0 8464 0 1 10880
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _220_
timestamp 1696364841
transform 1 0 8464 0 1 11968
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _221_
timestamp 1696364841
transform 1 0 7176 0 -1 9712
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _222_
timestamp 1696364841
transform 1 0 5796 0 -1 9712
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _223_
timestamp 1696364841
transform -1 0 4784 0 1 8704
box -38 -88 774 552
use sky130_fd_sc_hd__a32o_1  _224_
timestamp 1696364841
transform -1 0 4968 0 -1 8624
box -38 -88 774 552
use sky130_fd_sc_hd__and2_1  _225_
timestamp 1696364841
transform -1 0 7268 0 1 3264
box -38 -88 498 552
use sky130_fd_sc_hd__o21a_1  _226_
timestamp 1696364841
transform 1 0 3128 0 -1 4272
box -38 -88 590 552
use sky130_fd_sc_hd__nand2_1  _227_
timestamp 1696364841
transform -1 0 8372 0 -1 8624
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1696364841
transform -1 0 1748 0 1 6528
box -38 -88 314 552
use sky130_fd_sc_hd__a2bb2o_1  _229_
timestamp 1696364841
transform 1 0 1472 0 1 4352
box -38 -88 774 552
use sky130_fd_sc_hd__clkbuf_2  _230_
timestamp 1696364841
transform 1 0 2024 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__o2111a_1  _231_
timestamp 1696364841
transform 1 0 3588 0 -1 7536
box -38 -88 866 552
use sky130_fd_sc_hd__clkbuf_2  _232_
timestamp 1696364841
transform 1 0 3220 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__a21oi_1  _233_
timestamp 1696364841
transform 1 0 3220 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1696364841
transform -1 0 2116 0 1 10880
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 1696364841
transform 1 0 3956 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _236_
timestamp 1696364841
transform -1 0 1380 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _237_
timestamp 1696364841
transform -1 0 9660 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _238_
timestamp 1696364841
transform -1 0 11316 0 -1 11888
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _239_
timestamp 1696364841
transform -1 0 9844 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _240_
timestamp 1696364841
transform 1 0 10212 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _241_
timestamp 1696364841
transform 1 0 3128 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _242_
timestamp 1696364841
transform -1 0 736 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _243_
timestamp 1696364841
transform 1 0 3220 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1696364841
transform -1 0 920 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _245_
timestamp 1696364841
transform 1 0 1840 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _246_
timestamp 1696364841
transform 1 0 4324 0 1 11968
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _247_
timestamp 1696364841
transform 1 0 2024 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _248_
timestamp 1696364841
transform 1 0 8280 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1696364841
transform -1 0 9476 0 1 8704
box -38 -88 314 552
use sky130_fd_sc_hd__o22a_1  _250_
timestamp 1696364841
transform 1 0 6624 0 1 5440
box -38 -88 682 552
use sky130_fd_sc_hd__o211a_1  _251_
timestamp 1696364841
transform -1 0 7084 0 1 6528
box -38 -88 774 552
use sky130_fd_sc_hd__o21ai_1  _252_
timestamp 1696364841
transform -1 0 7636 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1696364841
transform -1 0 10212 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1696364841
transform 1 0 11776 0 1 4352
box -38 -88 314 552
use sky130_fd_sc_hd__or3_2  _255_
timestamp 1696364841
transform 1 0 5980 0 -1 4272
box -38 -88 590 552
use sky130_fd_sc_hd__a31o_1  _256_
timestamp 1696364841
transform -1 0 7636 0 -1 5360
box -38 -88 682 552
use sky130_fd_sc_hd__o21ba_1  _257_
timestamp 1696364841
transform -1 0 9016 0 -1 5360
box -38 -88 774 552
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1696364841
transform 1 0 9384 0 -1 5360
box -38 -88 866 552
use sky130_fd_sc_hd__a21oi_1  _259_
timestamp 1696364841
transform -1 0 12880 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_2  _260_
timestamp 1696364841
transform 1 0 8832 0 -1 6448
box -38 -88 498 552
use sky130_fd_sc_hd__nor2_1  _261_
timestamp 1696364841
transform -1 0 12880 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _262_
timestamp 1696364841
transform 1 0 14628 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _263_
timestamp 1696364841
transform -1 0 12144 0 -1 4272
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _264_
timestamp 1696364841
transform -1 0 12880 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _265_
timestamp 1696364841
transform 1 0 14904 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__a21oi_1  _266_
timestamp 1696364841
transform 1 0 14720 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__nor2_1  _267_
timestamp 1696364841
transform -1 0 12144 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _268_
timestamp 1696364841
transform -1 0 1656 0 1 7616
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1696364841
transform -1 0 920 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _270_
timestamp 1696364841
transform 1 0 2852 0 -1 8624
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1696364841
transform -1 0 644 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _272_
timestamp 1696364841
transform 1 0 4232 0 -1 9712
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1696364841
transform 1 0 14260 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _274_
timestamp 1696364841
transform 1 0 8464 0 1 9792
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1696364841
transform 1 0 12604 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1696364841
transform -1 0 11500 0 -1 10800
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1696364841
transform -1 0 11132 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__or2_1  _278_
timestamp 1696364841
transform 1 0 8740 0 -1 12976
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1696364841
transform -1 0 9200 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__or2_1  _280_
timestamp 1696364841
transform 1 0 4508 0 -1 11888
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1696364841
transform 1 0 7176 0 1 11968
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _282_
timestamp 1696364841
transform 1 0 3496 0 1 11968
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1696364841
transform 1 0 11040 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _284_
timestamp 1696364841
transform 1 0 14720 0 -1 5360
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1696364841
transform -1 0 14444 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__nand2_1  _286_
timestamp 1696364841
transform -1 0 12512 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _287_
timestamp 1696364841
transform 1 0 13892 0 1 4352
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1696364841
transform 1 0 14628 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _289_
timestamp 1696364841
transform -1 0 14260 0 1 3264
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1696364841
transform 1 0 14168 0 1 10880
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _291_
timestamp 1696364841
transform 1 0 13708 0 1 2176
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1696364841
transform 1 0 14260 0 -1 11888
box -38 -88 314 552
use sky130_fd_sc_hd__or2_2  _293_
timestamp 1696364841
transform 1 0 10948 0 1 4352
box -38 -88 498 552
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1696364841
transform 1 0 14904 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__o2111a_1  _295_
timestamp 1696364841
transform 1 0 5796 0 -1 5360
box -38 -88 866 552
use sky130_fd_sc_hd__o221ai_1  _296_
timestamp 1696364841
transform 1 0 5796 0 -1 7536
box -38 -88 682 552
use sky130_fd_sc_hd__nor2_2  _297_
timestamp 1696364841
transform 1 0 9752 0 -1 7536
box -38 -88 498 552
use sky130_fd_sc_hd__and3_1  _298_
timestamp 1696364841
transform -1 0 3772 0 1 3264
box -38 -88 498 552
use sky130_fd_sc_hd__o22a_1  _299_
timestamp 1696364841
transform 1 0 11224 0 -1 9712
box -38 -88 682 552
use sky130_fd_sc_hd__a221oi_2  _300_
timestamp 1696364841
transform 1 0 9568 0 1 6528
box -38 -88 1142 552
use sky130_fd_sc_hd__o221a_1  _301_
timestamp 1696364841
transform -1 0 11868 0 -1 7536
box -38 -88 866 552
use sky130_fd_sc_hd__o32a_1  _302_
timestamp 1696364841
transform 1 0 9292 0 -1 8624
box -38 -88 774 552
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1696364841
transform -1 0 8832 0 1 8704
box -38 -88 314 552
use sky130_fd_sc_hd__mux2_2  _304_
timestamp 1696364841
transform 1 0 5244 0 1 7616
box -38 -88 866 552
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 1696364841
transform 1 0 8188 0 -1 4272
box -38 -88 866 552
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1696364841
transform 1 0 11040 0 -1 5360
box -38 -88 866 552
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1696364841
transform 1 0 5428 0 1 5440
box -38 -88 866 552
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1696364841
transform 1 0 4968 0 1 4352
box -38 -88 866 552
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1696364841
transform 1 0 12512 0 -1 5360
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1696364841
transform 1 0 12512 0 -1 4272
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _311_
timestamp 1696364841
transform 1 0 12420 0 -1 3184
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 1696364841
transform 1 0 12328 0 -1 2096
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1696364841
transform 1 0 9200 0 1 5440
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1696364841
transform 1 0 7544 0 -1 7536
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1696364841
transform -1 0 2300 0 -1 7536
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1696364841
transform -1 0 2484 0 -1 8624
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1696364841
transform 1 0 1472 0 -1 9712
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1696364841
transform 1 0 920 0 -1 10800
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1696364841
transform 1 0 9844 0 1 10880
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1696364841
transform -1 0 11500 0 1 11968
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1696364841
transform 1 0 1748 0 -1 11888
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1696364841
transform 1 0 552 0 1 11968
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1696364841
transform 1 0 920 0 -1 3184
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_2  _324_
timestamp 1696364841
transform -1 0 7728 0 -1 8624
box -38 -88 1970 552
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1696364841
transform -1 0 6992 0 1 8704
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1696364841
transform -1 0 6072 0 1 9792
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1696364841
transform 1 0 6808 0 -1 10800
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1696364841
transform 1 0 8372 0 -1 11888
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1696364841
transform 1 0 6164 0 -1 11888
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1696364841
transform -1 0 6808 0 1 11968
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 1696364841
transform -1 0 6532 0 1 10880
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_4  _332_
timestamp 1696364841
transform -1 0 7360 0 1 1088
box -38 -88 2154 552
use sky130_fd_sc_hd__dfrtp_4  _333_
timestamp 1696364841
transform 1 0 4692 0 1 2176
box -38 -88 2154 552
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1696364841
transform 1 0 1656 0 -1 2096
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1696364841
transform 1 0 3220 0 -1 1008
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1696364841
transform 1 0 8740 0 1 4352
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1696364841
transform -1 0 10856 0 1 2176
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1696364841
transform 1 0 9016 0 1 1088
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1696364841
transform 1 0 8372 0 -1 2096
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1696364841
transform 1 0 8372 0 -1 3184
box -38 -88 1878 552
use sky130_fd_sc_hd__dfrtp_4  _341_
timestamp 1696364841
transform 1 0 644 0 -1 6448
box -38 -88 2154 552
use sky130_fd_sc_hd__dfrtp_4  _342_
timestamp 1696364841
transform 1 0 552 0 -1 5360
box -38 -88 2154 552
use sky130_fd_sc_hd__dfrtp_1  _343_
timestamp 1696364841
transform 1 0 828 0 -1 4272
box -38 -88 1878 552
use sky130_fd_sc_hd__dfstp_1  _344_
timestamp 1696364841
transform 1 0 12696 0 -1 7536
box -38 -88 1970 552
use sky130_fd_sc_hd__dfstp_1  _345_
timestamp 1696364841
transform 1 0 12696 0 -1 8624
box -38 -88 1970 552
use sky130_fd_sc_hd__dfstp_1  _346_
timestamp 1696364841
transform 1 0 10396 0 1 8704
box -38 -88 1970 552
use sky130_fd_sc_hd__dfrtp_1  _347_
timestamp 1696364841
transform 1 0 8464 0 1 7616
box -38 -88 1878 552
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1696364841
transform 1 0 6624 0 -1 6448
box -38 -88 1878 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1696364841
transform -1 0 6164 0 -1 12976
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1696364841
transform -1 0 11776 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1696364841
transform 1 0 11224 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1696364841
transform 1 0 11868 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1696364841
transform -1 0 12144 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1696364841
transform -1 0 12788 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 1696364841
transform 1 0 368 0 -1 1008
box -38 -88 590 552
use sky130_fd_sc_hd__decap_8  FILLER_0_13
timestamp 1696364841
transform 1 0 1288 0 -1 1008
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_0_25
timestamp 1696364841
transform 1 0 2392 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1696364841
transform 1 0 2852 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1696364841
transform 1 0 5060 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1696364841
transform 1 0 5520 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1696364841
transform 1 0 6348 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1696364841
transform 1 0 6992 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1696364841
transform 1 0 7728 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_0_88
timestamp 1696364841
transform 1 0 8188 0 -1 1008
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 1696364841
transform 1 0 8924 0 -1 1008
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1696364841
transform 1 0 9752 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1696364841
transform 1 0 10396 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1696364841
transform 1 0 10856 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1696364841
transform 1 0 11592 0 -1 1008
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1696364841
transform 1 0 13064 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_0_146
timestamp 1696364841
transform 1 0 13524 0 -1 1008
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1696364841
transform 1 0 14444 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1696364841
transform 1 0 15180 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1696364841
transform 1 0 368 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1696364841
transform 1 0 920 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1696364841
transform 1 0 2392 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1696364841
transform 1 0 2852 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_1_38
timestamp 1696364841
transform 1 0 3588 0 1 1088
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 1696364841
transform 1 0 4140 0 1 1088
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1696364841
transform 1 0 4876 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_1_79
timestamp 1696364841
transform 1 0 7360 0 1 1088
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1696364841
transform 1 0 7912 0 1 1088
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_1_87
timestamp 1696364841
transform 1 0 8096 0 1 1088
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_1_95
timestamp 1696364841
transform 1 0 8832 0 1 1088
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1696364841
transform 1 0 10856 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1696364841
transform 1 0 11500 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_12  FILLER_1_131
timestamp 1696364841
transform 1 0 12144 0 1 1088
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_8  FILLER_1_144
timestamp 1696364841
transform 1 0 13340 0 1 1088
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1696364841
transform 1 0 14076 0 1 1088
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1696364841
transform 1 0 14536 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1696364841
transform 1 0 15180 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1696364841
transform 1 0 644 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1696364841
transform 1 0 1288 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_2_37
timestamp 1696364841
transform 1 0 3496 0 -1 2096
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1696364841
transform 1 0 4968 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1696364841
transform 1 0 5428 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1696364841
transform 1 0 6808 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_2_84
timestamp 1696364841
transform 1 0 7820 0 -1 2096
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1696364841
transform 1 0 10212 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1696364841
transform 1 0 10672 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1696364841
transform 1 0 11316 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1696364841
transform 1 0 11960 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1696364841
transform 1 0 14168 0 -1 2096
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_2_159
timestamp 1696364841
transform 1 0 14720 0 -1 2096
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1696364841
transform 1 0 15180 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1696364841
transform 1 0 368 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1696364841
transform 1 0 1104 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1696364841
transform 1 0 1748 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1696364841
transform 1 0 2392 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_3_30
timestamp 1696364841
transform 1 0 2852 0 1 2176
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1696364841
transform 1 0 3588 0 1 2176
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1696364841
transform 1 0 4324 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_73
timestamp 1696364841
transform 1 0 6808 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1696364841
transform 1 0 7544 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_3_85
timestamp 1696364841
transform 1 0 7912 0 1 2176
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_3_87
timestamp 1696364841
transform 1 0 8096 0 1 2176
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1696364841
transform 1 0 8832 0 1 2176
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1696364841
transform 1 0 10856 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_3_129
timestamp 1696364841
transform 1 0 11960 0 1 2176
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1696364841
transform 1 0 12512 0 1 2176
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1696364841
transform 1 0 12880 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 1696364841
transform 1 0 13340 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_3_153
timestamp 1696364841
transform 1 0 14168 0 1 2176
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1696364841
transform 1 0 15180 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1696364841
transform 1 0 368 0 -1 3184
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1696364841
transform 1 0 2760 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_4_36
timestamp 1696364841
transform 1 0 3404 0 -1 3184
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1696364841
transform 1 0 3956 0 -1 3184
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1696364841
transform 1 0 4324 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1696364841
transform 1 0 4968 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1696364841
transform 1 0 5428 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1696364841
transform 1 0 6440 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_77
timestamp 1696364841
transform 1 0 7176 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1696364841
transform 1 0 7912 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1696364841
transform 1 0 8280 0 -1 3184
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1696364841
transform 1 0 10212 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1696364841
transform 1 0 10672 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_4_127
timestamp 1696364841
transform 1 0 11776 0 -1 3184
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_4_133
timestamp 1696364841
transform 1 0 12328 0 -1 3184
box -38 -88 130 552
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1696364841
transform 1 0 14260 0 -1 3184
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1696364841
transform 1 0 15180 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1696364841
transform 1 0 368 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1696364841
transform 1 0 1104 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1696364841
transform 1 0 1748 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_25
timestamp 1696364841
transform 1 0 2392 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1696364841
transform 1 0 2852 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1696364841
transform 1 0 3220 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1696364841
transform 1 0 3772 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1696364841
transform 1 0 4416 0 1 3264
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1696364841
transform 1 0 5612 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1696364841
transform 1 0 6348 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1696364841
transform 1 0 6716 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1696364841
transform 1 0 7268 0 1 3264
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1696364841
transform 1 0 8096 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1696364841
transform 1 0 8832 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1696364841
transform 1 0 9936 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1696364841
transform 1 0 10672 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_5_122
timestamp 1696364841
transform 1 0 11316 0 1 3264
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1696364841
transform 1 0 12144 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1696364841
transform 1 0 12880 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1696364841
transform 1 0 13340 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_5_148
timestamp 1696364841
transform 1 0 13708 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1696364841
transform 1 0 14260 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1696364841
transform 1 0 14996 0 1 3264
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1696364841
transform 1 0 368 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1696364841
transform 1 0 736 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_6_28
timestamp 1696364841
transform 1 0 2668 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1696364841
transform 1 0 3036 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1696364841
transform 1 0 3680 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_6_51
timestamp 1696364841
transform 1 0 4784 0 -1 4272
box -38 -88 590 552
use sky130_fd_sc_hd__decap_6  FILLER_6_58
timestamp 1696364841
transform 1 0 5428 0 -1 4272
box -38 -88 590 552
use sky130_fd_sc_hd__decap_8  FILLER_6_70
timestamp 1696364841
transform 1 0 6532 0 -1 4272
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1696364841
transform 1 0 7268 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1696364841
transform 1 0 7820 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1696364841
transform 1 0 9016 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1696364841
transform 1 0 10120 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1696364841
transform 1 0 10488 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1696364841
transform 1 0 10672 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_6_122
timestamp 1696364841
transform 1 0 11316 0 -1 4272
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1696364841
transform 1 0 12144 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 1696364841
transform 1 0 14352 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1696364841
transform 1 0 14720 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1696364841
transform 1 0 15180 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1696364841
transform 1 0 368 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1696364841
transform 1 0 1104 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_7_23
timestamp 1696364841
transform 1 0 2208 0 1 4352
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1696364841
transform 1 0 2852 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_7_43
timestamp 1696364841
transform 1 0 4048 0 1 4352
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1696364841
transform 1 0 4784 0 1 4352
box -38 -88 222 552
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1696364841
transform 1 0 5796 0 1 4352
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1696364841
transform 1 0 6532 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1696364841
transform 1 0 7268 0 1 4352
box -38 -88 774 552
use sky130_fd_sc_hd__decap_6  FILLER_7_87
timestamp 1696364841
transform 1 0 8096 0 1 4352
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1696364841
transform 1 0 8648 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_7_114
timestamp 1696364841
transform 1 0 10580 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1696364841
transform 1 0 11408 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_7_130
timestamp 1696364841
transform 1 0 12052 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_7_134
timestamp 1696364841
transform 1 0 12420 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1696364841
transform 1 0 12880 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_7_144
timestamp 1696364841
transform 1 0 13340 0 1 4352
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1696364841
transform 1 0 14352 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1696364841
transform 1 0 15088 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1696364841
transform 1 0 15456 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1696364841
transform 1 0 368 0 -1 5360
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_8_28
timestamp 1696364841
transform 1 0 2668 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1696364841
transform 1 0 3588 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_8_51
timestamp 1696364841
transform 1 0 4784 0 -1 5360
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1696364841
transform 1 0 5428 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1696364841
transform 1 0 6624 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_8_82
timestamp 1696364841
transform 1 0 7636 0 -1 5360
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_8_88
timestamp 1696364841
transform 1 0 8188 0 -1 5360
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1696364841
transform 1 0 9016 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1696364841
transform 1 0 10212 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1696364841
transform 1 0 10672 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_8_128
timestamp 1696364841
transform 1 0 11868 0 -1 5360
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_8_134
timestamp 1696364841
transform 1 0 12420 0 -1 5360
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 1696364841
transform 1 0 14352 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1696364841
transform 1 0 15180 0 -1 5360
box -38 -88 406 552
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1696364841
transform 1 0 368 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1696364841
transform 1 0 920 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1696364841
transform 1 0 1656 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1696364841
transform 1 0 2392 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1696364841
transform 1 0 2852 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1696364841
transform 1 0 3220 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1696364841
transform 1 0 3864 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_54
timestamp 1696364841
transform 1 0 5060 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_67
timestamp 1696364841
transform 1 0 6256 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1696364841
transform 1 0 7268 0 1 5440
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1696364841
transform 1 0 8096 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_94
timestamp 1696364841
transform 1 0 8740 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 1696364841
transform 1 0 9108 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_9_119
timestamp 1696364841
transform 1 0 11040 0 1 5440
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1696364841
transform 1 0 11776 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1696364841
transform 1 0 12144 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1696364841
transform 1 0 12788 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1696364841
transform 1 0 13156 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_9_144
timestamp 1696364841
transform 1 0 13340 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_9_151
timestamp 1696364841
transform 1 0 13984 0 1 5440
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1696364841
transform 1 0 14720 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1696364841
transform 1 0 15180 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1696364841
transform 1 0 368 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1696364841
transform 1 0 2760 0 -1 6448
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_10_44
timestamp 1696364841
transform 1 0 4140 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1696364841
transform 1 0 4968 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_10_58
timestamp 1696364841
transform 1 0 5428 0 -1 6448
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1696364841
transform 1 0 6256 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1696364841
transform 1 0 8464 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1696364841
transform 1 0 9292 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_10_108
timestamp 1696364841
transform 1 0 10028 0 -1 6448
box -38 -88 590 552
use sky130_fd_sc_hd__decap_8  FILLER_10_115
timestamp 1696364841
transform 1 0 10672 0 -1 6448
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1696364841
transform 1 0 11684 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_10_133
timestamp 1696364841
transform 1 0 12328 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1696364841
transform 1 0 13340 0 -1 6448
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1696364841
transform 1 0 14076 0 -1 6448
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1696364841
transform 1 0 14536 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1696364841
transform 1 0 15180 0 -1 6448
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1696364841
transform 1 0 368 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1696364841
transform 1 0 1104 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1696364841
transform 1 0 1748 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_25
timestamp 1696364841
transform 1 0 2392 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1696364841
transform 1 0 2852 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1696364841
transform 1 0 3680 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1696364841
transform 1 0 5980 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 1696364841
transform 1 0 7084 0 1 6528
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1696364841
transform 1 0 7820 0 1 6528
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_11_87
timestamp 1696364841
transform 1 0 8096 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_11_96
timestamp 1696364841
transform 1 0 8924 0 1 6528
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_11_102
timestamp 1696364841
transform 1 0 9476 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_11_115
timestamp 1696364841
transform 1 0 10672 0 1 6528
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_11_123
timestamp 1696364841
transform 1 0 11408 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1696364841
transform 1 0 12144 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1696364841
transform 1 0 12512 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1696364841
transform 1 0 12880 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1696364841
transform 1 0 13340 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1696364841
transform 1 0 14352 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1696364841
transform 1 0 15088 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1696364841
transform 1 0 15456 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1696364841
transform 1 0 368 0 -1 7536
box -38 -88 130 552
use sky130_fd_sc_hd__decap_6  FILLER_12_24
timestamp 1696364841
transform 1 0 2300 0 -1 7536
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1696364841
transform 1 0 2852 0 -1 7536
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1696364841
transform 1 0 3220 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_12_47
timestamp 1696364841
transform 1 0 4416 0 -1 7536
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1696364841
transform 1 0 5152 0 -1 7536
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1696364841
transform 1 0 5428 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1696364841
transform 1 0 6440 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_12_77
timestamp 1696364841
transform 1 0 7176 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1696364841
transform 1 0 9384 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1696364841
transform 1 0 10212 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1696364841
transform 1 0 10672 0 -1 7536
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_12_128
timestamp 1696364841
transform 1 0 11868 0 -1 7536
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_12_136
timestamp 1696364841
transform 1 0 12604 0 -1 7536
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1696364841
transform 1 0 14628 0 -1 7536
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1696364841
transform 1 0 15364 0 -1 7536
box -38 -88 222 552
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1696364841
transform 1 0 368 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_13_8
timestamp 1696364841
transform 1 0 828 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1696364841
transform 1 0 1656 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1696364841
transform 1 0 2392 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_13_30
timestamp 1696364841
transform 1 0 2852 0 1 7616
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1696364841
transform 1 0 3680 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1696364841
transform 1 0 4324 0 1 7616
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1696364841
transform 1 0 5060 0 1 7616
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1696364841
transform 1 0 6072 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_73
timestamp 1696364841
transform 1 0 6808 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp 1696364841
transform 1 0 7176 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1696364841
transform 1 0 7636 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_87
timestamp 1696364841
transform 1 0 8096 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1696364841
transform 1 0 10304 0 1 7616
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1696364841
transform 1 0 11776 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1696364841
transform 1 0 12880 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1696364841
transform 1 0 13340 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1696364841
transform 1 0 14352 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1696364841
transform 1 0 15088 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1696364841
transform 1 0 15456 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1696364841
transform 1 0 368 0 -1 8624
box -38 -88 314 552
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1696364841
transform 1 0 2484 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_14_35
timestamp 1696364841
transform 1 0 3312 0 -1 8624
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1696364841
transform 1 0 4048 0 -1 8624
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1696364841
transform 1 0 4968 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1696364841
transform 1 0 5428 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_14_83
timestamp 1696364841
transform 1 0 7728 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_14_90
timestamp 1696364841
transform 1 0 8372 0 -1 8624
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1696364841
transform 1 0 9108 0 -1 8624
box -38 -88 222 552
use sky130_fd_sc_hd__decap_6  FILLER_14_108
timestamp 1696364841
transform 1 0 10028 0 -1 8624
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1696364841
transform 1 0 10672 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1696364841
transform 1 0 11316 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_14_133
timestamp 1696364841
transform 1 0 12328 0 -1 8624
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1696364841
transform 1 0 14628 0 -1 8624
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1696364841
transform 1 0 15364 0 -1 8624
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1696364841
transform 1 0 368 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_15_11
timestamp 1696364841
transform 1 0 1104 0 1 8704
box -38 -88 774 552
use sky130_fd_sc_hd__decap_6  FILLER_15_23
timestamp 1696364841
transform 1 0 2208 0 1 8704
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1696364841
transform 1 0 2852 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_15_38
timestamp 1696364841
transform 1 0 3588 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_15_42
timestamp 1696364841
transform 1 0 3956 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1696364841
transform 1 0 4784 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1696364841
transform 1 0 6992 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_15_82
timestamp 1696364841
transform 1 0 7636 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1696364841
transform 1 0 8096 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1696364841
transform 1 0 8464 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_15_95
timestamp 1696364841
transform 1 0 8832 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1696364841
transform 1 0 9476 0 1 8704
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1696364841
transform 1 0 10212 0 1 8704
box -38 -88 222 552
use sky130_fd_sc_hd__decap_8  FILLER_15_133
timestamp 1696364841
transform 1 0 12328 0 1 8704
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1696364841
transform 1 0 13064 0 1 8704
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1696364841
transform 1 0 13340 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_15_155
timestamp 1696364841
transform 1 0 14352 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_15_159
timestamp 1696364841
transform 1 0 14720 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1696364841
transform 1 0 15180 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1696364841
transform 1 0 368 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1696364841
transform 1 0 1104 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_16_35
timestamp 1696364841
transform 1 0 3312 0 -1 9712
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1696364841
transform 1 0 4048 0 -1 9712
box -38 -88 222 552
use sky130_fd_sc_hd__decap_6  FILLER_16_50
timestamp 1696364841
transform 1 0 4692 0 -1 9712
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_16_56
timestamp 1696364841
transform 1 0 5244 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1696364841
transform 1 0 5428 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_16_70
timestamp 1696364841
transform 1 0 6532 0 -1 9712
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_16_76
timestamp 1696364841
transform 1 0 7084 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1696364841
transform 1 0 7912 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1696364841
transform 1 0 8556 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_16_99
timestamp 1696364841
transform 1 0 9200 0 -1 9712
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1696364841
transform 1 0 10212 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_16_115
timestamp 1696364841
transform 1 0 10672 0 -1 9712
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1696364841
transform 1 0 11868 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1696364841
transform 1 0 12512 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_16_142
timestamp 1696364841
transform 1 0 13156 0 -1 9712
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_16_150
timestamp 1696364841
transform 1 0 13892 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1696364841
transform 1 0 14260 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_16_161
timestamp 1696364841
transform 1 0 14904 0 -1 9712
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1696364841
transform 1 0 15456 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1696364841
transform 1 0 368 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1696364841
transform 1 0 736 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_17_14
timestamp 1696364841
transform 1 0 1380 0 1 9792
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_17_20
timestamp 1696364841
transform 1 0 1932 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1696364841
transform 1 0 2392 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1696364841
transform 1 0 2852 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_17_38
timestamp 1696364841
transform 1 0 3588 0 1 9792
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_17_44
timestamp 1696364841
transform 1 0 4140 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_65
timestamp 1696364841
transform 1 0 6072 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1696364841
transform 1 0 7544 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp 1696364841
transform 1 0 7912 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_87
timestamp 1696364841
transform 1 0 8096 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_17_96
timestamp 1696364841
transform 1 0 8924 0 1 9792
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_17_106
timestamp 1696364841
transform 1 0 9844 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1696364841
transform 1 0 10488 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 1696364841
transform 1 0 11132 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_17_127
timestamp 1696364841
transform 1 0 11776 0 1 9792
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1696364841
transform 1 0 12512 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1696364841
transform 1 0 12880 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_17_144
timestamp 1696364841
transform 1 0 13340 0 1 9792
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1696364841
transform 1 0 14076 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1696364841
transform 1 0 14444 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1696364841
transform 1 0 15180 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1696364841
transform 1 0 368 0 -1 10800
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1696364841
transform 1 0 2760 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_37
timestamp 1696364841
transform 1 0 3496 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1696364841
transform 1 0 3864 0 -1 10800
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1696364841
transform 1 0 4232 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1696364841
transform 1 0 4968 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1696364841
transform 1 0 5428 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1696364841
transform 1 0 6440 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1696364841
transform 1 0 8648 0 -1 10800
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1696364841
transform 1 0 9200 0 -1 10800
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1696364841
transform 1 0 9660 0 -1 10800
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_18_112
timestamp 1696364841
transform 1 0 10396 0 -1 10800
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1696364841
transform 1 0 10672 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1696364841
transform 1 0 11500 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1696364841
transform 1 0 12144 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_12  FILLER_18_138
timestamp 1696364841
transform 1 0 12788 0 -1 10800
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_8  FILLER_18_150
timestamp 1696364841
transform 1 0 13892 0 -1 10800
box -38 -88 774 552
use sky130_fd_sc_hd__decap_3  FILLER_18_158
timestamp 1696364841
transform 1 0 14628 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1696364841
transform 1 0 15180 0 -1 10800
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1696364841
transform 1 0 368 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_19_11
timestamp 1696364841
transform 1 0 1104 0 1 10880
box -38 -88 774 552
use sky130_fd_sc_hd__decap_6  FILLER_19_22
timestamp 1696364841
transform 1 0 2116 0 1 10880
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1696364841
transform 1 0 2668 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1696364841
transform 1 0 2852 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1696364841
transform 1 0 3588 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_46
timestamp 1696364841
transform 1 0 4324 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1696364841
transform 1 0 6532 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1696364841
transform 1 0 7636 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_87
timestamp 1696364841
transform 1 0 8096 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_19_99
timestamp 1696364841
transform 1 0 9200 0 1 10880
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1696364841
transform 1 0 9752 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__decap_12  FILLER_19_126
timestamp 1696364841
transform 1 0 11684 0 1 10880
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1696364841
transform 1 0 12788 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_19_142
timestamp 1696364841
transform 1 0 13156 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_19_144
timestamp 1696364841
transform 1 0 13340 0 1 10880
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 1696364841
transform 1 0 14076 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1696364841
transform 1 0 14444 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1696364841
transform 1 0 15180 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1696364841
transform 1 0 368 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_20_11
timestamp 1696364841
transform 1 0 1104 0 -1 11888
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_20_17
timestamp 1696364841
transform 1 0 1656 0 -1 11888
box -38 -88 130 552
use sky130_fd_sc_hd__decap_8  FILLER_20_38
timestamp 1696364841
transform 1 0 3588 0 -1 11888
box -38 -88 774 552
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1696364841
transform 1 0 4324 0 -1 11888
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1696364841
transform 1 0 4968 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1696364841
transform 1 0 5428 0 -1 11888
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_20_86
timestamp 1696364841
transform 1 0 8004 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1696364841
transform 1 0 10212 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1696364841
transform 1 0 10672 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__decap_12  FILLER_20_122
timestamp 1696364841
transform 1 0 11316 0 -1 11888
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_12  FILLER_20_134
timestamp 1696364841
transform 1 0 12420 0 -1 11888
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_8  FILLER_20_146
timestamp 1696364841
transform 1 0 13524 0 -1 11888
box -38 -88 774 552
use sky130_fd_sc_hd__decap_8  FILLER_20_157
timestamp 1696364841
transform 1 0 14536 0 -1 11888
box -38 -88 774 552
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1696364841
transform 1 0 15272 0 -1 11888
box -38 -88 314 552
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1696364841
transform 1 0 368 0 1 11968
box -38 -88 222 552
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1696364841
transform 1 0 2392 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1696364841
transform 1 0 2852 0 1 11968
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1696364841
transform 1 0 3404 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1696364841
transform 1 0 3956 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_21_49
timestamp 1696364841
transform 1 0 4600 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1696364841
transform 1 0 6808 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_21_80
timestamp 1696364841
transform 1 0 7452 0 1 11968
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1696364841
transform 1 0 8096 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1696364841
transform 1 0 9200 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1696364841
transform 1 0 9568 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__decap_12  FILLER_21_124
timestamp 1696364841
transform 1 0 11500 0 1 11968
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_6  FILLER_21_136
timestamp 1696364841
transform 1 0 12604 0 1 11968
box -38 -88 590 552
use sky130_fd_sc_hd__fill_1  FILLER_21_142
timestamp 1696364841
transform 1 0 13156 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__decap_12  FILLER_21_144
timestamp 1696364841
transform 1 0 13340 0 1 11968
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1696364841
transform 1 0 14444 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1696364841
transform 1 0 15180 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1696364841
transform 1 0 368 0 -1 12976
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1696364841
transform 1 0 1288 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_22_21
timestamp 1696364841
transform 1 0 2024 0 -1 12976
box -38 -88 774 552
use sky130_fd_sc_hd__decap_4  FILLER_22_30
timestamp 1696364841
transform 1 0 2852 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1696364841
transform 1 0 3588 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1696364841
transform 1 0 4324 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1696364841
transform 1 0 5060 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 1696364841
transform 1 0 5520 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_22_66
timestamp 1696364841
transform 1 0 6164 0 -1 12976
box -38 -88 774 552
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1696364841
transform 1 0 7268 0 -1 12976
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_22_86
timestamp 1696364841
transform 1 0 8004 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__decap_6  FILLER_22_88
timestamp 1696364841
transform 1 0 8188 0 -1 12976
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1696364841
transform 1 0 9200 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_8  FILLER_22_107
timestamp 1696364841
transform 1 0 9936 0 -1 12976
box -38 -88 774 552
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1696364841
transform 1 0 10672 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1696364841
transform 1 0 10856 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1696364841
transform 1 0 11592 0 -1 12976
box -38 -88 1142 552
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1696364841
transform 1 0 13064 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_6  FILLER_22_146
timestamp 1696364841
transform 1 0 13524 0 -1 12976
box -38 -88 590 552
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1696364841
transform 1 0 14444 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1696364841
transform 1 0 15180 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1696364841
transform 1 0 11684 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__buf_1  input2
timestamp 1696364841
transform -1 0 15180 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1696364841
transform 1 0 736 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__buf_1  input4
timestamp 1696364841
transform -1 0 10396 0 -1 1008
box -38 -88 314 552
use sky130_fd_sc_hd__buf_1  output5
timestamp 1696364841
transform 1 0 14904 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1696364841
transform -1 0 1288 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1696364841
transform -1 0 3588 0 1 1088
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1696364841
transform 1 0 14812 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1696364841
transform 1 0 12696 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1696364841
transform -1 0 11592 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1696364841
transform 1 0 7360 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1696364841
transform -1 0 7544 0 1 2176
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1696364841
transform 1 0 2024 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1696364841
transform -1 0 1288 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output15
timestamp 1696364841
transform -1 0 3588 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output16
timestamp 1696364841
transform 1 0 14812 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output17
timestamp 1696364841
transform 1 0 12696 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output18
timestamp 1696364841
transform -1 0 11592 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output19
timestamp 1696364841
transform -1 0 9936 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output20
timestamp 1696364841
transform -1 0 7268 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output21
timestamp 1696364841
transform 1 0 4692 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output22
timestamp 1696364841
transform -1 0 1104 0 1 6528
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output23
timestamp 1696364841
transform -1 0 828 0 1 7616
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output24
timestamp 1696364841
transform -1 0 1104 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output25
timestamp 1696364841
transform -1 0 1104 0 -1 9712
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output26
timestamp 1696364841
transform -1 0 1104 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output27
timestamp 1696364841
transform -1 0 1104 0 -1 11888
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output28
timestamp 1696364841
transform -1 0 2024 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output29
timestamp 1696364841
transform -1 0 4324 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output30
timestamp 1696364841
transform -1 0 1104 0 1 4352
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output31
timestamp 1696364841
transform 1 0 14812 0 -1 3184
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output32
timestamp 1696364841
transform 1 0 14812 0 -1 4272
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output33
timestamp 1696364841
transform 1 0 14812 0 -1 2096
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output34
timestamp 1696364841
transform 1 0 14076 0 -1 1008
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output35
timestamp 1696364841
transform 1 0 14812 0 1 5440
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output36
timestamp 1696364841
transform 1 0 14812 0 1 10880
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output37
timestamp 1696364841
transform 1 0 14812 0 1 9792
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output38
timestamp 1696364841
transform 1 0 14812 0 1 11968
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1696364841
transform 1 0 14076 0 -1 12976
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1696364841
transform 1 0 14812 0 1 8704
box -38 -88 406 552
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1696364841
transform -1 0 1104 0 1 3264
box -38 -88 406 552
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1696364841
transform 1 0 92 0 -1 1008
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1696364841
transform -1 0 15824 0 -1 1008
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1696364841
transform 1 0 92 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1696364841
transform -1 0 15824 0 1 1088
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1696364841
transform 1 0 92 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1696364841
transform -1 0 15824 0 -1 2096
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1696364841
transform 1 0 92 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1696364841
transform -1 0 15824 0 1 2176
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1696364841
transform 1 0 92 0 -1 3184
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1696364841
transform -1 0 15824 0 -1 3184
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1696364841
transform 1 0 92 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1696364841
transform -1 0 15824 0 1 3264
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1696364841
transform 1 0 92 0 -1 4272
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1696364841
transform -1 0 15824 0 -1 4272
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1696364841
transform 1 0 92 0 1 4352
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1696364841
transform -1 0 15824 0 1 4352
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1696364841
transform 1 0 92 0 -1 5360
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1696364841
transform -1 0 15824 0 -1 5360
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1696364841
transform 1 0 92 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1696364841
transform -1 0 15824 0 1 5440
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1696364841
transform 1 0 92 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1696364841
transform -1 0 15824 0 -1 6448
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1696364841
transform 1 0 92 0 1 6528
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1696364841
transform -1 0 15824 0 1 6528
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1696364841
transform 1 0 92 0 -1 7536
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1696364841
transform -1 0 15824 0 -1 7536
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1696364841
transform 1 0 92 0 1 7616
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1696364841
transform -1 0 15824 0 1 7616
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1696364841
transform 1 0 92 0 -1 8624
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1696364841
transform -1 0 15824 0 -1 8624
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1696364841
transform 1 0 92 0 1 8704
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1696364841
transform -1 0 15824 0 1 8704
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1696364841
transform 1 0 92 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1696364841
transform -1 0 15824 0 -1 9712
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1696364841
transform 1 0 92 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1696364841
transform -1 0 15824 0 1 9792
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1696364841
transform 1 0 92 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1696364841
transform -1 0 15824 0 -1 10800
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1696364841
transform 1 0 92 0 1 10880
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1696364841
transform -1 0 15824 0 1 10880
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1696364841
transform 1 0 92 0 -1 11888
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1696364841
transform -1 0 15824 0 -1 11888
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1696364841
transform 1 0 92 0 1 11968
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1696364841
transform -1 0 15824 0 1 11968
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1696364841
transform 1 0 92 0 -1 12976
box -38 -88 314 552
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1696364841
transform -1 0 15824 0 -1 12976
box -38 -88 314 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1696364841
transform 1 0 2760 0 -1 1008
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1696364841
transform 1 0 5428 0 -1 1008
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1696364841
transform 1 0 8096 0 -1 1008
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1696364841
transform 1 0 10764 0 -1 1008
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1696364841
transform 1 0 13432 0 -1 1008
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1696364841
transform 1 0 2760 0 1 1088
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1696364841
transform 1 0 8004 0 1 1088
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1696364841
transform 1 0 13248 0 1 1088
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1696364841
transform 1 0 5336 0 -1 2096
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1696364841
transform 1 0 10580 0 -1 2096
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1696364841
transform 1 0 2760 0 1 2176
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1696364841
transform 1 0 8004 0 1 2176
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1696364841
transform 1 0 13248 0 1 2176
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1696364841
transform 1 0 5336 0 -1 3184
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1696364841
transform 1 0 10580 0 -1 3184
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1696364841
transform 1 0 2760 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1696364841
transform 1 0 8004 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1696364841
transform 1 0 13248 0 1 3264
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1696364841
transform 1 0 5336 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1696364841
transform 1 0 10580 0 -1 4272
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1696364841
transform 1 0 2760 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1696364841
transform 1 0 8004 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1696364841
transform 1 0 13248 0 1 4352
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1696364841
transform 1 0 5336 0 -1 5360
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1696364841
transform 1 0 10580 0 -1 5360
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1696364841
transform 1 0 2760 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1696364841
transform 1 0 8004 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1696364841
transform 1 0 13248 0 1 5440
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1696364841
transform 1 0 5336 0 -1 6448
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1696364841
transform 1 0 10580 0 -1 6448
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1696364841
transform 1 0 2760 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1696364841
transform 1 0 8004 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1696364841
transform 1 0 13248 0 1 6528
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1696364841
transform 1 0 5336 0 -1 7536
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1696364841
transform 1 0 10580 0 -1 7536
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1696364841
transform 1 0 2760 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1696364841
transform 1 0 8004 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1696364841
transform 1 0 13248 0 1 7616
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1696364841
transform 1 0 5336 0 -1 8624
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1696364841
transform 1 0 10580 0 -1 8624
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1696364841
transform 1 0 2760 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1696364841
transform 1 0 8004 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1696364841
transform 1 0 13248 0 1 8704
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1696364841
transform 1 0 5336 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1696364841
transform 1 0 10580 0 -1 9712
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1696364841
transform 1 0 2760 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1696364841
transform 1 0 8004 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1696364841
transform 1 0 13248 0 1 9792
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1696364841
transform 1 0 5336 0 -1 10800
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1696364841
transform 1 0 10580 0 -1 10800
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1696364841
transform 1 0 2760 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1696364841
transform 1 0 8004 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1696364841
transform 1 0 13248 0 1 10880
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1696364841
transform 1 0 5336 0 -1 11888
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1696364841
transform 1 0 10580 0 -1 11888
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1696364841
transform 1 0 2760 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1696364841
transform 1 0 8004 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1696364841
transform 1 0 13248 0 1 11968
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1696364841
transform 1 0 2760 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1696364841
transform 1 0 5428 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1696364841
transform 1 0 8096 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1696364841
transform 1 0 10764 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1696364841
transform 1 0 13432 0 -1 12976
box -38 -88 130 552
use sky130_fd_sc_hd__buf_8  repeater42
timestamp 1696364841
transform 1 0 6440 0 1 9792
box -38 -88 1142 552
use sky130_fd_sc_hd__buf_8  repeater43
timestamp 1696364841
transform -1 0 2392 0 1 1088
box -38 -88 1142 552
<< labels >>
rlabel metal2 s 938 -40 994 160 4 ctln[0]
port 3 nsew
rlabel metal2 s 2870 -40 2926 160 4 ctln[1]
port 5 nsew
rlabel metal2 s 14922 -40 14978 160 4 ctln[2]
port 7 nsew
rlabel metal2 s 12898 -40 12954 160 4 ctln[3]
port 9 nsew
rlabel metal2 s 10874 -40 10930 160 4 ctln[4]
port 11 nsew
rlabel metal2 s 8942 -40 8998 160 4 ctln[5]
port 13 nsew
rlabel metal2 s 6918 -40 6974 160 4 ctln[6]
port 15 nsew
rlabel metal2 s 4894 -40 4950 160 4 ctln[7]
port 17 nsew
rlabel metal2 s 938 13760 994 13960 4 ctlp[0]
port 19 nsew
rlabel metal2 s 2870 13760 2926 13960 4 ctlp[1]
port 21 nsew
rlabel metal2 s 14922 13760 14978 13960 4 ctlp[2]
port 23 nsew
rlabel metal2 s 12898 13760 12954 13960 4 ctlp[3]
port 25 nsew
rlabel metal2 s 10874 13760 10930 13960 4 ctlp[4]
port 27 nsew
rlabel metal2 s 8942 13760 8998 13960 4 ctlp[5]
port 29 nsew
rlabel metal2 s 6918 13760 6974 13960 4 ctlp[6]
port 31 nsew
rlabel metal2 s 4894 13760 4950 13960 4 ctlp[7]
port 33 nsew
rlabel metal3 s 0 3398 200 3458 4 cal
port 36 nsew
rlabel metal3 s 0 1358 200 1418 4 clk
port 38 nsew
rlabel metal3 s 15800 6254 16000 6314 4 clkc
port 40 nsew
rlabel metal3 s 15800 7478 16000 7538 4 comp
port 42 nsew
rlabel metal3 s 0 2310 200 2370 4 en
port 44 nsew
rlabel metal3 s 0 6390 200 6450 4 result[0]
port 46 nsew
rlabel metal3 s 0 7342 200 7402 4 result[1]
port 48 nsew
rlabel metal3 s 0 8294 200 8354 4 result[2]
port 50 nsew
rlabel metal3 s 0 9382 200 9442 4 result[3]
port 52 nsew
rlabel metal3 s 0 10334 200 10394 4 result[4]
port 54 nsew
rlabel metal3 s 0 11286 200 11346 4 result[5]
port 56 nsew
rlabel metal3 s 0 12374 200 12434 4 result[6]
port 58 nsew
rlabel metal3 s 0 13326 200 13386 4 result[7]
port 60 nsew
rlabel metal3 s 0 406 200 466 4 rstn
port 62 nsew
rlabel metal3 s 0 5302 200 5362 4 sample
port 64 nsew
rlabel metal3 s 15800 2854 16000 2914 4 trim[0]
port 66 nsew
rlabel metal3 s 15800 3942 16000 4002 4 trim[1]
port 68 nsew
rlabel metal3 s 15800 1630 16000 1690 4 trim[2]
port 70 nsew
rlabel metal3 s 15800 542 16000 602 4 trim[3]
port 72 nsew
rlabel metal3 s 15800 5166 16000 5226 4 trim[4]
port 74 nsew
rlabel metal3 s 15800 11014 16000 11074 4 trimb[0]
port 76 nsew
rlabel metal3 s 15800 9790 16000 9850 4 trimb[1]
port 78 nsew
rlabel metal3 s 15800 12102 16000 12162 4 trimb[2]
port 80 nsew
rlabel metal3 s 15800 13326 16000 13386 4 trimb[3]
port 82 nsew
rlabel metal3 s 15800 8702 16000 8762 4 trimb[4]
port 84 nsew
rlabel metal3 s 0 4350 200 4410 4 valid
port 86 nsew
rlabel metal4 s 13112 456 13432 13064 4 VPWR
port 89 nsew
rlabel metal4 s 7840 456 8160 13064 4 VPWR
port 89 nsew
rlabel metal4 s 2568 456 2888 13064 4 VPWR
port 89 nsew
rlabel metal4 s 10476 456 10796 13064 4 VGND
port 91 nsew
rlabel metal4 s 5204 456 5524 13064 4 VGND
port 91 nsew
rlabel metal5 s 92 11056 15824 11376 4 VPWR
port 89 nsew
rlabel metal5 s 92 6752 15824 7072 4 VPWR
port 89 nsew
rlabel metal5 s 92 2448 15824 2768 4 VPWR
port 89 nsew
rlabel metal5 s 92 8904 15824 9224 4 VGND
port 91 nsew
rlabel metal5 s 92 4600 15824 4920 4 VGND
port 91 nsew
<< properties >>
string FIXED_BBOX 0 -40 16000 13960
<< end >>
