magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 866 542
<< pwell >>
rect 1 -19 808 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
rect 247 7 277 137
rect 437 7 467 137
rect 521 7 551 137
rect 605 7 635 137
rect 689 7 719 137
<< scpmoshvt >>
rect 79 257 109 457
rect 163 257 193 457
rect 247 257 277 457
rect 437 257 467 457
rect 521 257 551 457
rect 605 257 635 457
rect 689 257 719 457
<< ndiff >>
rect 27 125 79 137
rect 27 91 35 125
rect 69 91 79 125
rect 27 57 79 91
rect 27 23 35 57
rect 69 23 79 57
rect 27 7 79 23
rect 109 55 163 137
rect 109 21 119 55
rect 153 21 163 55
rect 109 7 163 21
rect 193 125 247 137
rect 193 91 203 125
rect 237 91 247 125
rect 193 57 247 91
rect 193 23 203 57
rect 237 23 247 57
rect 193 7 247 23
rect 277 55 437 137
rect 277 21 287 55
rect 321 21 393 55
rect 427 21 437 55
rect 277 7 437 21
rect 467 123 521 137
rect 467 89 477 123
rect 511 89 521 123
rect 467 55 521 89
rect 467 21 477 55
rect 511 21 521 55
rect 467 7 521 21
rect 551 55 605 137
rect 551 21 561 55
rect 595 21 605 55
rect 551 7 605 21
rect 635 123 689 137
rect 635 89 645 123
rect 679 89 689 123
rect 635 55 689 89
rect 635 21 645 55
rect 679 21 689 55
rect 635 7 689 21
rect 719 55 782 137
rect 719 21 729 55
rect 763 21 782 55
rect 719 7 782 21
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 257 163 457
rect 193 257 247 457
rect 277 445 437 457
rect 277 411 300 445
rect 334 411 393 445
rect 427 411 437 445
rect 277 377 437 411
rect 277 343 300 377
rect 334 343 393 377
rect 427 343 437 377
rect 277 257 437 343
rect 467 437 521 457
rect 467 403 477 437
rect 511 403 521 437
rect 467 369 521 403
rect 467 335 477 369
rect 511 335 521 369
rect 467 301 521 335
rect 467 267 477 301
rect 511 267 521 301
rect 467 257 521 267
rect 551 437 605 457
rect 551 403 561 437
rect 595 403 605 437
rect 551 369 605 403
rect 551 335 561 369
rect 595 335 605 369
rect 551 257 605 335
rect 635 437 689 457
rect 635 403 645 437
rect 679 403 689 437
rect 635 369 689 403
rect 635 335 645 369
rect 679 335 689 369
rect 635 301 689 335
rect 635 267 645 301
rect 679 267 689 301
rect 635 257 689 267
rect 719 437 791 457
rect 719 403 729 437
rect 763 403 791 437
rect 719 369 791 403
rect 719 335 729 369
rect 763 335 791 369
rect 719 257 791 335
<< ndiffc >>
rect 35 91 69 125
rect 35 23 69 57
rect 119 21 153 55
rect 203 91 237 125
rect 203 23 237 57
rect 287 21 321 55
rect 393 21 427 55
rect 477 89 511 123
rect 477 21 511 55
rect 561 21 595 55
rect 645 89 679 123
rect 645 21 679 55
rect 729 21 763 55
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 300 411 334 445
rect 393 411 427 445
rect 300 343 334 377
rect 393 343 427 377
rect 477 403 511 437
rect 477 335 511 369
rect 477 267 511 301
rect 561 403 595 437
rect 561 335 595 369
rect 645 403 679 437
rect 645 335 679 369
rect 645 267 679 301
rect 729 403 763 437
rect 729 335 763 369
<< poly >>
rect 79 457 109 483
rect 163 457 193 483
rect 247 457 277 483
rect 437 457 467 483
rect 521 457 551 483
rect 605 457 635 483
rect 689 457 719 483
rect 79 225 109 257
rect 163 225 193 257
rect 247 225 277 257
rect 437 225 467 257
rect 521 225 551 257
rect 605 225 635 257
rect 689 225 719 257
rect 25 209 109 225
rect 25 175 35 209
rect 69 175 109 209
rect 25 159 109 175
rect 151 209 205 225
rect 151 175 161 209
rect 195 175 205 209
rect 151 159 205 175
rect 247 209 305 225
rect 247 175 261 209
rect 295 175 305 209
rect 247 159 305 175
rect 380 209 719 225
rect 380 175 396 209
rect 430 175 464 209
rect 498 175 532 209
rect 566 175 600 209
rect 634 175 668 209
rect 702 175 719 209
rect 380 159 719 175
rect 79 137 109 159
rect 163 137 193 159
rect 247 137 277 159
rect 437 137 467 159
rect 521 137 551 159
rect 605 137 635 159
rect 689 137 719 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 247 -19 277 7
rect 437 -19 467 7
rect 521 -19 551 7
rect 605 -19 635 7
rect 689 -19 719 7
<< polycont >>
rect 35 175 69 209
rect 161 175 195 209
rect 261 175 295 209
rect 396 175 430 209
rect 464 175 498 209
rect 532 175 566 209
rect 600 175 634 209
rect 668 175 702 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 17 445 253 453
rect 17 411 35 445
rect 69 419 253 445
rect 69 411 85 419
rect 17 377 85 411
rect 17 343 35 377
rect 69 343 85 377
rect 17 309 85 343
rect 17 275 35 309
rect 69 275 85 309
rect 17 259 85 275
rect 119 225 166 370
rect 200 293 253 419
rect 287 445 427 487
rect 287 411 300 445
rect 334 411 393 445
rect 287 377 427 411
rect 287 343 300 377
rect 334 343 393 377
rect 287 327 427 343
rect 469 437 519 453
rect 469 403 477 437
rect 511 403 519 437
rect 469 369 519 403
rect 469 335 477 369
rect 511 335 519 369
rect 469 301 519 335
rect 553 437 603 487
rect 553 403 561 437
rect 595 403 603 437
rect 553 369 603 403
rect 553 335 561 369
rect 595 335 603 369
rect 553 319 603 335
rect 637 437 687 453
rect 637 403 645 437
rect 679 403 687 437
rect 637 369 687 403
rect 637 335 645 369
rect 679 335 687 369
rect 200 259 418 293
rect 17 209 85 225
rect 17 175 35 209
rect 69 175 85 209
rect 119 209 211 225
rect 119 175 161 209
rect 195 175 211 209
rect 245 209 340 225
rect 245 175 261 209
rect 295 175 340 209
rect 374 209 418 259
rect 469 267 477 301
rect 511 285 519 301
rect 637 301 687 335
rect 721 437 771 487
rect 721 403 729 437
rect 763 403 771 437
rect 721 369 771 403
rect 721 335 729 369
rect 763 335 771 369
rect 721 319 771 335
rect 637 285 645 301
rect 511 267 645 285
rect 679 285 687 301
rect 679 267 811 285
rect 469 251 811 267
rect 374 175 396 209
rect 430 175 464 209
rect 498 175 532 209
rect 566 175 600 209
rect 634 175 668 209
rect 702 175 719 209
rect 374 141 418 175
rect 753 141 811 251
rect 17 125 418 141
rect 17 91 35 125
rect 69 105 203 125
rect 69 91 85 105
rect 17 57 85 91
rect 187 91 203 105
rect 237 105 418 125
rect 461 123 811 141
rect 237 91 253 105
rect 17 23 35 57
rect 69 23 85 57
rect 17 11 85 23
rect 119 55 153 71
rect 119 -23 153 21
rect 187 57 253 91
rect 461 89 477 123
rect 511 107 645 123
rect 511 89 527 107
rect 187 23 203 57
rect 237 23 253 57
rect 187 11 253 23
rect 287 55 427 71
rect 321 21 393 55
rect 287 -23 427 21
rect 461 55 527 89
rect 629 89 645 107
rect 679 107 811 123
rect 679 89 695 107
rect 461 21 477 55
rect 511 21 527 55
rect 461 13 527 21
rect 561 55 595 71
rect 561 -23 595 21
rect 629 55 695 89
rect 629 21 645 55
rect 679 21 695 55
rect 629 13 695 21
rect 729 55 763 71
rect 729 -23 763 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
<< metal1 >>
rect 0 521 828 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 0 456 828 487
rect 0 -23 828 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
rect 0 -88 828 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or3_4
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 306 181 340 215 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 766 113 800 147 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 122 317 156 351 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 C
port 8 nsew
flabel locali s 122 249 156 283 0 FreeSans 400 0 0 0 B
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 828 504
string path 0.000 -1.000 20.700 -1.000 
<< end >>
