magic
tech sky130B
magscale 1 2
timestamp 1698189341
<< locali >>
rect 34394 15115 34440 15131
rect 30074 15069 34440 15115
rect 34394 13427 34440 15069
rect 35061 13427 35107 13438
rect 33700 13381 35107 13427
rect 33700 12057 33746 13381
rect 35061 13246 35107 13381
rect 33413 12006 33746 12057
rect 33413 12005 33685 12006
rect 29404 10483 29536 10517
rect 34402 10508 34436 11065
rect 29404 8879 29438 10483
rect 33758 10474 34436 10508
rect 29404 8845 29556 8879
<< metal1 >>
rect 29492 18054 32575 18149
rect 32670 18054 32676 18149
rect 29492 17891 29587 18054
rect 30038 17946 33465 17988
rect 30038 17894 30243 17946
rect 30295 17894 33465 17946
rect 30038 17893 33465 17894
rect 33560 17893 33566 17988
rect 952 17829 1046 17835
rect 396 17763 490 17769
rect 396 15856 490 17669
rect 952 16394 1046 17735
rect 952 16300 1351 16394
rect 396 15762 1430 15856
rect 30701 15019 30747 15218
rect 31943 15024 31987 15218
rect 33031 15037 33077 15218
rect 33550 15004 33594 15218
rect 34284 14855 34334 15218
rect 151 14508 1417 14544
rect 34019 13528 34071 13534
rect 34071 13486 35033 13518
rect 34019 13470 34071 13476
rect 35001 13216 35033 13486
rect 32447 12492 32499 12498
rect 32447 12434 32499 12440
rect 32457 12277 32489 12434
rect 35656 12121 35759 12181
rect 31249 12061 31255 12113
rect 31307 12061 31313 12113
rect 31241 11940 31247 12000
rect 31307 11940 31313 12000
rect 32439 11570 32471 11777
rect 32429 11564 32481 11570
rect 32429 11506 32481 11512
rect 34989 11046 34995 11098
rect 35047 11046 35053 11098
rect 185 9426 1477 9462
rect 30724 8709 30770 8918
rect 31966 8694 32010 8919
rect 33054 8703 33100 8945
rect 33573 8700 33617 8958
rect 34307 8683 34357 9013
rect 388 8114 1434 8208
rect 388 6737 482 8114
rect 388 6637 482 6643
rect 950 7576 1351 7670
rect 950 6737 1044 7576
rect 950 6637 1044 6643
rect 29492 5938 29587 6079
rect 33213 6077 33308 6083
rect 30038 5982 33213 6077
rect 33213 5976 33308 5982
rect 32655 5938 32750 5944
rect 29492 5912 32655 5938
rect 29492 5860 30195 5912
rect 30247 5860 32655 5912
rect 29492 5843 32655 5860
rect 32655 5837 32750 5843
<< via1 >>
rect 32575 18054 32670 18149
rect 30243 17894 30295 17946
rect 33465 17893 33560 17988
rect 396 17669 490 17763
rect 952 17735 1046 17829
rect 34019 13476 34071 13528
rect 32447 12440 32499 12492
rect 31255 12061 31307 12113
rect 31247 11940 31307 12000
rect 32429 11512 32481 11564
rect 34995 11046 35047 11098
rect 388 6643 482 6737
rect 950 6643 1044 6737
rect 33213 5982 33308 6077
rect 30195 5860 30247 5912
rect 32655 5843 32750 5938
<< metal2 >>
rect 32575 18149 32670 18155
rect 32566 18054 32575 18149
rect 32670 18054 32679 18149
rect 32575 18048 32670 18054
rect 33465 17988 33560 17994
rect 30243 17946 30295 17952
rect 30243 17888 30295 17894
rect 33456 17893 33465 17988
rect 33560 17893 33569 17988
rect 952 17829 1046 17838
rect 387 17669 396 17763
rect 490 17669 499 17763
rect 946 17735 952 17829
rect 1046 17735 1052 17829
rect 952 17726 1046 17735
rect 30252 17689 30285 17888
rect 33465 17887 33560 17893
rect 30208 17656 30285 17689
rect 30180 17377 30304 17411
rect 30186 17106 30302 17140
rect 30194 16829 30302 16863
rect 30188 16555 30302 16589
rect 1305 7510 1346 16462
rect 30184 16280 30302 16314
rect 30186 16004 30304 16038
rect 30192 15729 30296 15763
rect 30198 15455 30290 15489
rect 34013 13518 34019 13528
rect 32457 13486 34019 13518
rect 32457 12492 32489 13486
rect 34013 13476 34019 13486
rect 34071 13476 34077 13528
rect 34239 13442 35733 13470
rect 30409 12442 30465 12451
rect 32441 12440 32447 12492
rect 32499 12440 32505 12492
rect 30465 12397 31298 12432
rect 30409 12377 30465 12386
rect 31263 12119 31298 12397
rect 31255 12113 31307 12119
rect 31255 12055 31307 12061
rect 31247 12000 31307 12006
rect 31247 11936 31307 11940
rect 31240 11880 31249 11936
rect 31305 11880 31314 11936
rect 31247 11878 31307 11880
rect 34239 11628 34267 13442
rect 33485 11598 34268 11628
rect 32423 11512 32429 11564
rect 32481 11512 32487 11564
rect 32439 10914 32471 11512
rect 34995 11098 35047 11104
rect 34995 11040 35047 11046
rect 35005 10914 35037 11040
rect 32439 10882 35037 10914
rect 30190 8481 30300 8515
rect 30182 8207 30300 8241
rect 30184 7932 30300 7966
rect 30188 7656 30298 7690
rect 30196 7381 30294 7415
rect 30182 7107 30288 7141
rect 30192 6830 30286 6864
rect 388 6737 482 6746
rect 950 6737 1044 6746
rect 382 6643 388 6737
rect 482 6643 488 6737
rect 944 6643 950 6737
rect 1044 6643 1050 6737
rect 388 6634 482 6643
rect 950 6634 1044 6643
rect 30184 6559 30290 6593
rect 30204 5918 30238 6315
rect 33213 6077 33308 6086
rect 33207 5982 33213 6077
rect 33308 5982 33314 6077
rect 33213 5973 33308 5982
rect 32655 5938 32750 5947
rect 30195 5912 30247 5918
rect 30195 5854 30247 5860
rect 32649 5843 32655 5938
rect 32750 5843 32756 5938
rect 32655 5834 32750 5843
<< via2 >>
rect 32575 18054 32670 18149
rect 33465 17893 33560 17988
rect 396 17669 490 17763
rect 952 17735 1046 17829
rect 30409 12386 30465 12442
rect 31249 11880 31305 11936
rect 388 6643 482 6737
rect 950 6643 1044 6737
rect 33213 5982 33308 6077
rect 32655 5843 32750 5938
<< metal3 >>
rect 32570 18149 32580 18154
rect 32570 18054 32575 18149
rect 32570 18049 32580 18054
rect 32675 18049 32681 18154
rect 33460 17988 33470 17993
rect 33460 17893 33465 17988
rect 33460 17888 33470 17893
rect 33565 17888 33571 17993
rect 947 17834 1051 17840
rect 391 17768 495 17774
rect 947 17735 952 17740
rect 1046 17735 1051 17740
rect 947 17730 1051 17735
rect 391 17669 396 17674
rect 490 17669 495 17674
rect 391 17664 495 17669
rect 30383 12446 30481 12460
rect 30383 12382 30405 12446
rect 30469 12382 30481 12446
rect 30383 12362 30481 12382
rect 31237 11940 31313 12000
rect 31237 11876 31245 11940
rect 31309 11876 31313 11940
rect 31237 11870 31313 11876
rect 383 6737 487 6742
rect 383 6732 388 6737
rect 482 6732 487 6737
rect 383 6632 487 6638
rect 945 6737 1049 6742
rect 945 6732 950 6737
rect 1044 6732 1049 6737
rect 945 6632 1049 6638
rect 33208 6082 33313 6088
rect 33208 5982 33213 5987
rect 33308 5982 33313 5987
rect 33208 5977 33313 5982
rect 32650 5943 32755 5949
rect 32650 5843 32655 5848
rect 32750 5843 32755 5848
rect 32650 5838 32755 5843
<< via3 >>
rect 32580 18149 32675 18154
rect 32580 18054 32670 18149
rect 32670 18054 32675 18149
rect 32580 18049 32675 18054
rect 33470 17988 33565 17993
rect 33470 17893 33560 17988
rect 33560 17893 33565 17988
rect 33470 17888 33565 17893
rect 947 17829 1051 17834
rect 391 17763 495 17768
rect 391 17674 396 17763
rect 396 17674 490 17763
rect 490 17674 495 17763
rect 947 17740 952 17829
rect 952 17740 1046 17829
rect 1046 17740 1051 17829
rect 30405 12442 30469 12446
rect 30405 12386 30409 12442
rect 30409 12386 30465 12442
rect 30465 12386 30469 12442
rect 30405 12382 30469 12386
rect 31245 11936 31309 11940
rect 31245 11880 31249 11936
rect 31249 11880 31305 11936
rect 31305 11880 31309 11936
rect 31245 11876 31309 11880
rect 383 6643 388 6732
rect 388 6643 482 6732
rect 482 6643 487 6732
rect 383 6638 487 6643
rect 945 6643 950 6732
rect 950 6643 1044 6732
rect 1044 6643 1049 6732
rect 945 6638 1049 6643
rect 33208 6077 33313 6082
rect 33208 5987 33213 6077
rect 33213 5987 33308 6077
rect 33308 5987 33313 6077
rect 32650 5938 32755 5943
rect 32650 5848 32655 5938
rect 32655 5848 32750 5938
rect 32750 5848 32755 5938
<< metal4 >>
rect 323 18688 563 23652
rect 323 17768 563 18368
rect 323 17674 391 17768
rect 495 17674 563 17768
rect 323 6732 563 17674
rect 323 6638 383 6732
rect 487 6638 563 6732
rect 323 5662 563 6638
rect 887 17834 1127 21036
rect 32509 18154 32749 21076
rect 33395 18726 33635 23642
rect 32509 18049 32580 18154
rect 32675 18049 32749 18154
rect 32509 18028 32749 18049
rect 887 17740 947 17834
rect 1051 17740 1127 17834
rect 33395 17993 33635 18406
rect 33395 17888 33470 17993
rect 33565 17888 33635 17993
rect 33395 17832 33635 17888
rect 887 6732 1127 17740
rect 30404 12446 30470 12447
rect 30404 12382 30405 12446
rect 30469 12382 30470 12446
rect 30404 12381 30470 12382
rect 27793 12080 27853 12368
rect 30407 12080 30467 12381
rect 27793 12020 30469 12080
rect 31244 11940 31310 11941
rect 31244 11938 31245 11940
rect 27793 11878 31245 11938
rect 27793 11602 27853 11878
rect 31244 11876 31245 11878
rect 31309 11876 31310 11940
rect 31244 11875 31310 11876
rect 887 6638 945 6732
rect 1049 6638 1127 6732
rect 283 520 603 5342
rect 887 3078 1127 6638
rect 33147 6082 33387 6158
rect 33147 5987 33208 6082
rect 33313 5987 33387 6082
rect 32595 5943 32835 5984
rect 32595 5848 32650 5943
rect 32755 5848 32835 5943
rect 32595 3022 32835 5848
rect 33147 5614 33387 5987
rect 33147 450 33387 5294
<< via4 >>
rect 283 23652 603 23972
rect 33355 23642 33675 23962
rect 847 21036 1167 21356
rect 32469 21076 32789 21396
rect 283 18368 603 18688
rect 33355 18406 33675 18726
rect 283 5342 603 5662
rect 847 2758 1167 3078
rect 33107 5294 33427 5614
rect 32555 2702 32875 3022
rect 283 200 603 520
rect 33107 130 33427 450
<< metal5 >>
rect 0 23972 33824 24162
rect 0 23652 283 23972
rect 603 23962 33824 23972
rect 603 23652 33355 23962
rect 0 23642 33355 23652
rect 33675 23642 33824 23962
rect 0 23500 33824 23642
rect 666 21396 32942 21540
rect 666 21356 32469 21396
rect 666 21036 847 21356
rect 1167 21076 32469 21356
rect 32789 21076 32942 21396
rect 1167 21036 32942 21076
rect 666 20878 32942 21036
rect 114 18726 33864 18910
rect 114 18688 33355 18726
rect 114 18368 283 18688
rect 603 18406 33355 18688
rect 33675 18406 33864 18726
rect 603 18368 33864 18406
rect 114 18248 33864 18368
rect 160 5662 33508 5800
rect 160 5342 283 5662
rect 603 5614 33508 5662
rect 603 5342 33107 5614
rect 160 5294 33107 5342
rect 33427 5294 33508 5614
rect 160 5138 33508 5294
rect 731 3078 32908 3224
rect 731 2758 847 3078
rect 1167 3022 32908 3078
rect 1167 2758 32555 3022
rect 731 2702 32555 2758
rect 32875 2702 32908 3022
rect 731 2562 32908 2702
rect 118 520 33570 662
rect 118 200 283 520
rect 603 450 33570 520
rect 603 200 33107 450
rect 118 130 33107 200
rect 33427 130 33570 450
rect 118 0 33570 130
use comparator  comparator_0 comparator
timestamp 1697741630
transform 0 1 31351 1 0 10647
box -1805 -1948 4495 3006
use dac  dac_0 dac
timestamp 1697762684
transform 1 0 1537 0 -1 17966
box -280 -22 28705 5880
use dac  dac_1
timestamp 1697762684
transform 1 0 1537 0 1 6004
box -280 -22 28705 5880
use latch  latch_0 latch
timestamp 1697130564
transform 0 1 34368 -1 0 13304
box 0 -41 2306 1348
use vpp_cap  vpp_cap_0
timestamp 1697748102
transform 1 0 30105 0 1 3040
box 4 4 2286 2342
use vpp_cap  vpp_cap_1
timestamp 1697748102
transform 1 0 30111 0 -1 2728
box 4 4 2286 2342
use vpp_cap  vpp_cap_2
timestamp 1697748102
transform 1 0 27487 0 1 3040
box 4 4 2286 2342
use vpp_cap  vpp_cap_3
timestamp 1697748102
transform 1 0 27493 0 -1 2728
box 4 4 2286 2342
use vpp_cap  vpp_cap_4
timestamp 1697748102
transform 1 0 24875 0 -1 2724
box 4 4 2286 2342
use vpp_cap  vpp_cap_5
timestamp 1697748102
transform 1 0 24869 0 1 3044
box 4 4 2286 2342
use vpp_cap  vpp_cap_6
timestamp 1697748102
transform 1 0 22251 0 1 3044
box 4 4 2286 2342
use vpp_cap  vpp_cap_7
timestamp 1697748102
transform 1 0 22257 0 -1 2724
box 4 4 2286 2342
use vpp_cap  vpp_cap_8
timestamp 1697748102
transform 1 0 6557 0 -1 2720
box 4 4 2286 2342
use vpp_cap  vpp_cap_9
timestamp 1697748102
transform 1 0 9175 0 -1 2720
box 4 4 2286 2342
use vpp_cap  vpp_cap_10
timestamp 1697748102
transform 1 0 1321 0 -1 2716
box 4 4 2286 2342
use vpp_cap  vpp_cap_11
timestamp 1697748102
transform 1 0 3939 0 -1 2716
box 4 4 2286 2342
use vpp_cap  vpp_cap_12
timestamp 1697748102
transform 1 0 6551 0 1 3048
box 4 4 2286 2342
use vpp_cap  vpp_cap_13
timestamp 1697748102
transform 1 0 9169 0 1 3048
box 4 4 2286 2342
use vpp_cap  vpp_cap_14
timestamp 1697748102
transform 1 0 1315 0 1 3052
box 4 4 2286 2342
use vpp_cap  vpp_cap_15
timestamp 1697748102
transform 1 0 3933 0 1 3052
box 4 4 2286 2342
use vpp_cap  vpp_cap_16
timestamp 1697748102
transform 1 0 11785 0 -1 2720
box 4 4 2286 2342
use vpp_cap  vpp_cap_17
timestamp 1697748102
transform 1 0 14403 0 -1 2720
box 4 4 2286 2342
use vpp_cap  vpp_cap_18
timestamp 1697748102
transform 1 0 17021 0 -1 2724
box 4 4 2286 2342
use vpp_cap  vpp_cap_19
timestamp 1697748102
transform 1 0 19639 0 -1 2724
box 4 4 2286 2342
use vpp_cap  vpp_cap_20
timestamp 1697748102
transform 1 0 11779 0 1 3048
box 4 4 2286 2342
use vpp_cap  vpp_cap_21
timestamp 1697748102
transform 1 0 14397 0 1 3048
box 4 4 2286 2342
use vpp_cap  vpp_cap_22
timestamp 1697748102
transform 1 0 17015 0 1 3044
box 4 4 2286 2342
use vpp_cap  vpp_cap_23
timestamp 1697748102
transform 1 0 19633 0 1 3044
box 4 4 2286 2342
use vpp_cap  vpp_cap_24
timestamp 1697748102
transform 1 0 11697 0 -1 21048
box 4 4 2286 2342
use vpp_cap  vpp_cap_25
timestamp 1697748102
transform 1 0 9087 0 -1 21048
box 4 4 2286 2342
use vpp_cap  vpp_cap_26
timestamp 1697748102
transform 1 0 6469 0 -1 21048
box 4 4 2286 2342
use vpp_cap  vpp_cap_27
timestamp 1697748102
transform 1 0 3851 0 -1 21044
box 4 4 2286 2342
use vpp_cap  vpp_cap_28
timestamp 1697748102
transform 1 0 1233 0 -1 21044
box 4 4 2286 2342
use vpp_cap  vpp_cap_29
timestamp 1697748102
transform 1 0 30023 0 -1 21056
box 4 4 2286 2342
use vpp_cap  vpp_cap_30
timestamp 1697748102
transform 1 0 27405 0 -1 21056
box 4 4 2286 2342
use vpp_cap  vpp_cap_31
timestamp 1697748102
transform 1 0 24787 0 -1 21052
box 4 4 2286 2342
use vpp_cap  vpp_cap_32
timestamp 1697748102
transform 1 0 22169 0 -1 21052
box 4 4 2286 2342
use vpp_cap  vpp_cap_33
timestamp 1697748102
transform 1 0 19551 0 -1 21052
box 4 4 2286 2342
use vpp_cap  vpp_cap_34
timestamp 1697748102
transform 1 0 16933 0 -1 21052
box 4 4 2286 2342
use vpp_cap  vpp_cap_35
timestamp 1697748102
transform 1 0 14315 0 -1 21048
box 4 4 2286 2342
use vpp_cap  vpp_cap_36
timestamp 1697748102
transform 1 0 11691 0 1 21376
box 4 4 2286 2342
use vpp_cap  vpp_cap_37
timestamp 1697748102
transform 1 0 9081 0 1 21376
box 4 4 2286 2342
use vpp_cap  vpp_cap_38
timestamp 1697748102
transform 1 0 6463 0 1 21376
box 4 4 2286 2342
use vpp_cap  vpp_cap_39
timestamp 1697748102
transform 1 0 3845 0 1 21380
box 4 4 2286 2342
use vpp_cap  vpp_cap_40
timestamp 1697748102
transform 1 0 1227 0 1 21380
box 4 4 2286 2342
use vpp_cap  vpp_cap_41
timestamp 1697748102
transform 1 0 30017 0 1 21368
box 4 4 2286 2342
use vpp_cap  vpp_cap_42
timestamp 1697748102
transform 1 0 27399 0 1 21368
box 4 4 2286 2342
use vpp_cap  vpp_cap_43
timestamp 1697748102
transform 1 0 24781 0 1 21372
box 4 4 2286 2342
use vpp_cap  vpp_cap_44
timestamp 1697748102
transform 1 0 22163 0 1 21372
box 4 4 2286 2342
use vpp_cap  vpp_cap_45
timestamp 1697748102
transform 1 0 19545 0 1 21372
box 4 4 2286 2342
use vpp_cap  vpp_cap_46
timestamp 1697748102
transform 1 0 16927 0 1 21372
box 4 4 2286 2342
use vpp_cap  vpp_cap_47
timestamp 1697748102
transform 1 0 14309 0 1 21376
box 4 4 2286 2342
<< labels >>
flabel metal1 35699 12121 35759 12181 0 FreeSans 1280 0 0 0 comp
port 30 nsew signal output
flabel metal2 35705 13442 35733 13470 0 FreeSans 1280 0 0 0 clkc
port 31 nsew signal input
flabel metal4 887 6732 1127 17740 0 FreeSans 1280 90 0 0 avss
port 33 nsew ground bidirectional
flabel metal4 323 6732 563 17674 0 FreeSans 1280 90 0 0 avdd
port 32 nsew power bidirectional
flabel metal1 151 14508 187 14544 0 FreeSans 1280 0 0 0 vinp
port 27 nsew signal input
flabel metal1 185 9426 221 9462 0 FreeSans 1280 0 0 0 vinn
port 28 nsew signal input
flabel metal2 30256 15455 30290 15489 0 FreeSans 1280 0 0 0 ctlp7
port 1 nsew signal input
flabel metal2 30262 15729 30296 15763 0 FreeSans 1280 0 0 0 ctlp6
port 2 nsew signal input
flabel metal2 30270 16004 30304 16038 0 FreeSans 1280 0 0 0 ctlp5
port 3 nsew signal input
flabel metal2 30268 16280 30302 16314 0 FreeSans 1280 0 0 0 ctlp4
port 4 nsew signal input
flabel metal2 30268 16555 30302 16589 0 FreeSans 1280 0 0 0 ctlp3
port 5 nsew signal input
flabel metal2 30268 16829 30302 16863 0 FreeSans 1280 0 0 0 ctlp2
port 6 nsew signal input
flabel metal2 30268 17106 30302 17140 0 FreeSans 1280 0 0 0 ctlp1
port 7 nsew signal input
flabel metal2 30270 17377 30304 17411 0 FreeSans 1280 0 0 0 ctlp0
port 8 nsew signal input
flabel metal2 30256 6559 30290 6593 0 FreeSans 1280 0 0 0 ctln0
port 16 nsew signal input
flabel metal2 30252 6830 30286 6864 0 FreeSans 1280 0 0 0 ctln1
port 15 nsew signal input
flabel metal2 30254 7107 30288 7141 0 FreeSans 1280 0 0 0 ctln2
port 14 nsew signal input
flabel metal2 30260 7381 30294 7415 0 FreeSans 1280 0 0 0 ctln3
port 13 nsew signal input
flabel metal2 30264 7656 30298 7690 0 FreeSans 1280 0 0 0 ctln4
port 12 nsew signal input
flabel metal2 30266 7932 30300 7966 0 FreeSans 1280 0 0 0 ctln5
port 11 nsew signal input
flabel metal2 30266 8207 30300 8241 0 FreeSans 1280 0 0 0 ctln6
port 10 nsew signal input
flabel metal2 30266 8481 30300 8515 0 FreeSans 1280 0 0 0 ctln7
port 9 nsew signal input
flabel metal1 30724 8709 30770 8996 0 FreeSans 1280 90 0 0 trim4
port 17 nsew signal input
flabel metal1 31966 8694 32010 8996 0 FreeSans 1280 90 0 0 trim3
port 18 nsew signal input
flabel metal1 33054 8703 33100 9000 0 FreeSans 1280 90 0 0 trim2
port 19 nsew signal input
flabel metal1 33573 8700 33617 9005 0 FreeSans 1280 90 0 0 trim1
port 20 nsew signal input
flabel metal1 34307 8683 34357 8733 0 FreeSans 1280 90 0 0 trim0
port 21 nsew signal input
flabel metal1 34284 15168 34334 15218 0 FreeSans 1280 90 0 0 trimb0
port 26 nsew signal input
flabel metal1 33550 15174 33594 15218 0 FreeSans 1280 90 0 0 trimb1
port 25 nsew signal input
flabel metal1 33031 15172 33077 15218 0 FreeSans 1280 90 0 0 trimb2
port 24 nsew signal input
flabel metal1 31943 15174 31987 15218 0 FreeSans 1280 90 0 0 trimb3
port 23 nsew signal input
flabel metal1 30701 15172 30747 15218 0 FreeSans 1280 90 0 0 trimb4
port 22 nsew signal input
flabel metal2 1305 7510 1346 16462 0 FreeSans 1280 90 0 0 sample
port 29 nsew signal input
<< properties >>
string FIXED_BBOX P��KV
string LEFclass CORE
string LEFsite unithddbl
<< end >>
