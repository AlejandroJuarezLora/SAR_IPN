VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO latch
  CLASS BLOCK ;
  FOREIGN latch ;
  ORIGIN 0.000 0.200 ;
  SIZE 11.530 BY 6.855 ;
  PIN vdd
    ANTENNADIFFAREA 5.865600 ;
    PORT
      LAYER nwell ;
        RECT 0.000 3.285 11.530 6.655 ;
      LAYER li1 ;
        RECT 0.180 6.305 11.350 6.475 ;
        RECT 0.180 3.635 0.350 6.305 ;
        RECT 1.015 4.480 1.185 5.520 ;
        RECT 4.155 4.480 4.325 5.520 ;
        RECT 7.205 4.480 7.375 5.520 ;
        RECT 10.345 4.480 10.515 5.520 ;
        RECT 11.180 3.635 11.350 6.305 ;
        RECT 0.180 3.465 11.350 3.635 ;
      LAYER mcon ;
        RECT 1.835 6.305 2.005 6.475 ;
        RECT 2.195 6.305 2.365 6.475 ;
        RECT 2.835 6.305 3.005 6.475 ;
        RECT 3.195 6.305 3.365 6.475 ;
        RECT 7.835 6.305 8.005 6.475 ;
        RECT 8.195 6.305 8.365 6.475 ;
        RECT 8.835 6.305 9.005 6.475 ;
        RECT 9.195 6.305 9.365 6.475 ;
        RECT 1.015 5.095 1.185 5.265 ;
        RECT 1.015 4.735 1.185 4.905 ;
        RECT 4.155 5.095 4.325 5.265 ;
        RECT 4.155 4.735 4.325 4.905 ;
        RECT 7.205 5.095 7.375 5.265 ;
        RECT 7.205 4.735 7.375 4.905 ;
        RECT 10.345 5.095 10.515 5.265 ;
        RECT 10.345 4.735 10.515 4.905 ;
      LAYER met1 ;
        RECT 0.750 6.240 4.590 6.540 ;
        RECT 6.805 6.240 10.780 6.540 ;
        RECT 0.985 4.500 1.215 6.240 ;
        RECT 4.125 4.500 4.355 6.240 ;
        RECT 7.175 4.500 7.405 6.240 ;
        RECT 10.315 4.500 10.545 6.240 ;
      LAYER via ;
        RECT 0.810 6.260 1.070 6.520 ;
        RECT 1.130 6.260 1.390 6.520 ;
        RECT 3.950 6.260 4.210 6.520 ;
        RECT 4.270 6.260 4.530 6.520 ;
        RECT 7.000 6.260 7.260 6.520 ;
        RECT 7.320 6.260 7.580 6.520 ;
        RECT 10.140 6.260 10.400 6.520 ;
        RECT 10.460 6.260 10.720 6.520 ;
      LAYER met2 ;
        RECT 0.800 6.190 10.730 6.590 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 6.445600 ;
    PORT
      LAYER pwell ;
        RECT 0.050 2.635 11.480 3.065 ;
        RECT 0.050 0.225 0.480 2.635 ;
        RECT 11.050 0.225 11.480 2.635 ;
        RECT 0.050 -0.205 11.480 0.225 ;
      LAYER li1 ;
        RECT 0.180 2.765 11.350 2.935 ;
        RECT 0.180 0.095 0.350 2.765 ;
        RECT 1.015 1.055 1.185 2.095 ;
        RECT 2.585 1.055 2.755 2.095 ;
        RECT 4.155 1.055 4.325 2.095 ;
        RECT 7.205 1.055 7.375 2.095 ;
        RECT 8.775 1.055 8.945 2.095 ;
        RECT 10.345 1.055 10.515 2.095 ;
        RECT 11.180 0.095 11.350 2.765 ;
        RECT 0.180 -0.075 11.350 0.095 ;
      LAYER mcon ;
        RECT 1.015 1.670 1.185 1.840 ;
        RECT 1.015 1.310 1.185 1.480 ;
        RECT 2.585 1.670 2.755 1.840 ;
        RECT 2.585 1.310 2.755 1.480 ;
        RECT 4.155 1.670 4.325 1.840 ;
        RECT 4.155 1.310 4.325 1.480 ;
        RECT 7.205 1.670 7.375 1.840 ;
        RECT 7.205 1.310 7.375 1.480 ;
        RECT 8.775 1.670 8.945 1.840 ;
        RECT 8.775 1.310 8.945 1.480 ;
        RECT 10.345 1.670 10.515 1.840 ;
        RECT 10.345 1.310 10.515 1.480 ;
        RECT 2.270 -0.075 2.440 0.095 ;
        RECT 2.630 -0.075 2.800 0.095 ;
        RECT 3.270 -0.075 3.440 0.095 ;
        RECT 3.630 -0.075 3.800 0.095 ;
        RECT 4.270 -0.075 4.440 0.095 ;
        RECT 4.630 -0.075 4.800 0.095 ;
        RECT 5.270 -0.075 5.440 0.095 ;
        RECT 5.630 -0.075 5.800 0.095 ;
        RECT 6.270 -0.075 6.440 0.095 ;
        RECT 6.630 -0.075 6.800 0.095 ;
        RECT 7.270 -0.075 7.440 0.095 ;
        RECT 7.630 -0.075 7.800 0.095 ;
        RECT 8.270 -0.075 8.440 0.095 ;
        RECT 8.630 -0.075 8.800 0.095 ;
      LAYER met1 ;
        RECT 0.985 0.160 1.215 2.075 ;
        RECT 2.555 0.160 2.785 2.075 ;
        RECT 4.125 0.160 4.355 2.075 ;
        RECT 7.175 0.160 7.405 2.075 ;
        RECT 8.745 0.160 8.975 2.075 ;
        RECT 10.315 0.160 10.545 2.075 ;
        RECT 0.750 -0.140 10.780 0.160 ;
      LAYER via ;
        RECT 0.810 -0.120 1.070 0.140 ;
        RECT 1.130 -0.120 1.390 0.140 ;
        RECT 2.380 -0.120 2.640 0.140 ;
        RECT 2.700 -0.120 2.960 0.140 ;
        RECT 3.950 -0.120 4.210 0.140 ;
        RECT 4.270 -0.120 4.530 0.140 ;
        RECT 7.000 -0.120 7.260 0.140 ;
        RECT 7.320 -0.120 7.580 0.140 ;
        RECT 8.570 -0.120 8.830 0.140 ;
        RECT 8.890 -0.120 9.150 0.140 ;
        RECT 10.140 -0.120 10.400 0.140 ;
        RECT 10.460 -0.120 10.720 0.140 ;
      LAYER met2 ;
        RECT 0.800 -0.190 10.730 0.210 ;
    END
  END vss
  PIN Qn
    ANTENNAGATEAREA 0.800000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 6.515 4.480 6.685 5.520 ;
        RECT 4.385 4.095 4.785 4.265 ;
        RECT 4.385 2.265 4.785 2.435 ;
        RECT 3.275 1.055 3.445 2.095 ;
        RECT 6.515 1.055 6.685 2.095 ;
      LAYER mcon ;
        RECT 6.515 5.095 6.685 5.265 ;
        RECT 6.515 4.735 6.685 4.905 ;
        RECT 4.500 4.095 4.670 4.265 ;
        RECT 4.500 2.265 4.670 2.435 ;
        RECT 3.275 1.670 3.445 1.840 ;
        RECT 3.275 1.310 3.445 1.480 ;
        RECT 6.515 1.670 6.685 1.840 ;
        RECT 6.515 1.310 6.685 1.480 ;
      LAYER met1 ;
        RECT 6.485 5.350 6.715 5.500 ;
        RECT 6.415 4.650 6.715 5.350 ;
        RECT 6.485 4.500 6.715 4.650 ;
        RECT 4.405 3.415 4.765 4.295 ;
        RECT 3.625 3.115 4.765 3.415 ;
        RECT 3.625 2.075 3.925 3.115 ;
        RECT 4.405 2.465 4.765 3.115 ;
        RECT 6.100 2.915 6.400 3.615 ;
        RECT 6.130 2.465 6.360 2.915 ;
        RECT 4.405 2.235 6.360 2.465 ;
        RECT 3.245 1.775 3.925 2.075 ;
        RECT 6.485 1.925 6.715 2.075 ;
        RECT 3.245 1.075 3.475 1.775 ;
        RECT 6.415 1.225 6.715 1.925 ;
        RECT 6.485 1.075 6.715 1.225 ;
      LAYER via ;
        RECT 6.435 5.030 6.695 5.290 ;
        RECT 6.435 4.710 6.695 4.970 ;
        RECT 6.120 3.295 6.380 3.555 ;
        RECT 6.120 2.975 6.380 3.235 ;
        RECT 6.435 1.605 6.695 1.865 ;
        RECT 6.435 1.285 6.695 1.545 ;
      LAYER met2 ;
        RECT 6.365 4.700 6.765 5.300 ;
        RECT 6.450 3.565 6.680 4.700 ;
        RECT 6.050 2.965 6.680 3.565 ;
        RECT 6.450 1.875 6.680 2.965 ;
        RECT 6.365 1.275 6.765 1.875 ;
    END
  END Qn
  PIN S
    ANTENNAGATEAREA 0.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.245 4.095 1.645 4.265 ;
        RECT 1.245 2.265 1.645 2.435 ;
      LAYER mcon ;
        RECT 1.360 4.095 1.530 4.265 ;
        RECT 1.360 2.265 1.530 2.435 ;
      LAYER met1 ;
        RECT 1.265 3.415 1.625 4.295 ;
        RECT 0.265 3.115 1.625 3.415 ;
        RECT 1.265 2.235 1.625 3.115 ;
    END
  END S
  PIN R
    ANTENNAGATEAREA 0.800000 ;
    PORT
      LAYER li1 ;
        RECT 9.885 4.095 10.285 4.265 ;
        RECT 9.885 2.265 10.285 2.435 ;
      LAYER mcon ;
        RECT 10.000 4.095 10.170 4.265 ;
        RECT 10.000 2.265 10.170 2.435 ;
      LAYER met1 ;
        RECT 9.905 3.415 10.265 4.295 ;
        RECT 9.905 3.115 11.265 3.415 ;
        RECT 9.905 2.235 10.265 3.115 ;
    END
  END R
  PIN Q
    ANTENNAGATEAREA 0.800000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 4.845 4.480 5.015 5.520 ;
        RECT 6.745 4.095 7.145 4.265 ;
        RECT 6.745 2.265 7.145 2.435 ;
        RECT 4.845 1.055 5.015 2.095 ;
        RECT 8.085 1.055 8.255 2.095 ;
      LAYER mcon ;
        RECT 4.845 5.095 5.015 5.265 ;
        RECT 4.845 4.735 5.015 4.905 ;
        RECT 6.860 4.095 7.030 4.265 ;
        RECT 6.860 2.265 7.030 2.435 ;
        RECT 4.845 1.670 5.015 1.840 ;
        RECT 4.845 1.310 5.015 1.480 ;
        RECT 8.085 1.670 8.255 1.840 ;
        RECT 8.085 1.310 8.255 1.480 ;
      LAYER met1 ;
        RECT 4.815 5.350 5.045 5.500 ;
        RECT 4.815 4.650 5.115 5.350 ;
        RECT 4.815 4.500 5.045 4.650 ;
        RECT 5.615 4.295 5.915 6.740 ;
        RECT 5.165 4.065 7.125 4.295 ;
        RECT 5.165 3.615 5.395 4.065 ;
        RECT 5.130 2.915 5.430 3.615 ;
        RECT 6.765 3.415 7.125 4.065 ;
        RECT 6.765 3.115 7.905 3.415 ;
        RECT 6.765 2.235 7.125 3.115 ;
        RECT 7.605 2.075 7.905 3.115 ;
        RECT 4.815 1.925 5.045 2.075 ;
        RECT 4.815 1.225 5.115 1.925 ;
        RECT 7.605 1.775 8.285 2.075 ;
        RECT 4.815 1.075 5.045 1.225 ;
        RECT 8.055 1.075 8.285 1.775 ;
      LAYER via ;
        RECT 4.835 5.030 5.095 5.290 ;
        RECT 4.835 4.710 5.095 4.970 ;
        RECT 5.150 3.295 5.410 3.555 ;
        RECT 5.150 2.975 5.410 3.235 ;
        RECT 4.835 1.605 5.095 1.865 ;
        RECT 4.835 1.285 5.095 1.545 ;
      LAYER met2 ;
        RECT 4.765 4.700 5.165 5.300 ;
        RECT 4.850 3.565 5.080 4.700 ;
        RECT 4.850 2.965 5.480 3.565 ;
        RECT 4.850 1.875 5.080 2.965 ;
        RECT 4.765 1.275 5.165 1.875 ;
    END
  END Q
  OBS
      LAYER pwell ;
        RECT 0.825 0.945 2.065 2.205 ;
        RECT 2.395 0.945 3.635 2.205 ;
        RECT 3.965 0.945 5.205 2.205 ;
        RECT 6.325 0.945 7.565 2.205 ;
        RECT 7.895 0.945 9.135 2.205 ;
        RECT 9.465 0.945 10.705 2.205 ;
      LAYER li1 ;
        RECT 1.705 4.480 1.875 5.520 ;
        RECT 9.655 4.480 9.825 5.520 ;
        RECT 2.815 2.265 3.215 2.435 ;
        RECT 8.315 2.265 8.715 2.435 ;
        RECT 1.705 1.055 1.875 2.095 ;
        RECT 9.655 1.055 9.825 2.095 ;
      LAYER mcon ;
        RECT 1.705 5.095 1.875 5.265 ;
        RECT 1.705 4.735 1.875 4.905 ;
        RECT 9.655 5.095 9.825 5.265 ;
        RECT 9.655 4.735 9.825 4.905 ;
        RECT 2.930 2.265 3.100 2.435 ;
        RECT 8.430 2.265 8.600 2.435 ;
        RECT 1.705 1.670 1.875 1.840 ;
        RECT 1.705 1.310 1.875 1.480 ;
        RECT 9.655 1.670 9.825 1.840 ;
        RECT 9.655 1.310 9.825 1.480 ;
      LAYER met1 ;
        RECT 1.675 5.350 1.905 5.500 ;
        RECT 9.625 5.350 9.855 5.500 ;
        RECT 1.675 4.650 1.975 5.350 ;
        RECT 9.555 4.650 9.855 5.350 ;
        RECT 1.675 4.500 1.905 4.650 ;
        RECT 9.625 4.500 9.855 4.650 ;
        RECT 1.990 3.415 2.290 3.615 ;
        RECT 9.240 3.415 9.540 3.615 ;
        RECT 1.990 3.115 3.165 3.415 ;
        RECT 1.990 2.915 2.290 3.115 ;
        RECT 2.865 2.465 3.165 3.115 ;
        RECT 8.365 3.115 9.540 3.415 ;
        RECT 8.365 2.465 8.665 3.115 ;
        RECT 9.240 2.915 9.540 3.115 ;
        RECT 2.835 2.235 3.195 2.465 ;
        RECT 8.335 2.235 8.695 2.465 ;
        RECT 1.675 1.925 1.905 2.075 ;
        RECT 9.625 1.925 9.855 2.075 ;
        RECT 1.675 1.225 1.975 1.925 ;
        RECT 9.555 1.225 9.855 1.925 ;
        RECT 1.675 1.075 1.905 1.225 ;
        RECT 9.625 1.075 9.855 1.225 ;
      LAYER via ;
        RECT 1.695 5.030 1.955 5.290 ;
        RECT 1.695 4.710 1.955 4.970 ;
        RECT 9.575 5.030 9.835 5.290 ;
        RECT 9.575 4.710 9.835 4.970 ;
        RECT 2.010 3.295 2.270 3.555 ;
        RECT 2.010 2.975 2.270 3.235 ;
        RECT 9.260 3.295 9.520 3.555 ;
        RECT 9.260 2.975 9.520 3.235 ;
        RECT 1.695 1.605 1.955 1.865 ;
        RECT 1.695 1.285 1.955 1.545 ;
        RECT 9.575 1.605 9.835 1.865 ;
        RECT 9.575 1.285 9.835 1.545 ;
      LAYER met2 ;
        RECT 1.625 4.700 2.025 5.300 ;
        RECT 9.505 4.700 9.905 5.300 ;
        RECT 1.710 3.565 1.940 4.700 ;
        RECT 9.590 3.565 9.820 4.700 ;
        RECT 1.710 2.965 2.340 3.565 ;
        RECT 9.190 2.965 9.820 3.565 ;
        RECT 1.710 1.875 1.940 2.965 ;
        RECT 9.590 1.875 9.820 2.965 ;
        RECT 1.625 1.275 2.025 1.875 ;
        RECT 9.505 1.275 9.905 1.875 ;
  END
END latch
END LIBRARY

