magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 682 542
<< pwell >>
rect 1 -19 643 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 267 7 297 137
rect 351 7 381 137
rect 451 7 481 137
rect 535 7 565 137
<< scpmoshvt >>
rect 83 257 113 457
rect 262 257 292 457
rect 339 257 369 457
rect 463 257 493 457
rect 535 257 565 457
<< ndiff >>
rect 27 96 79 137
rect 27 62 35 96
rect 69 62 79 96
rect 27 7 79 62
rect 109 53 161 137
rect 109 19 119 53
rect 153 19 161 53
rect 109 7 161 19
rect 215 55 267 137
rect 215 21 223 55
rect 257 21 267 55
rect 215 7 267 21
rect 297 123 351 137
rect 297 89 307 123
rect 341 89 351 123
rect 297 7 351 89
rect 381 123 451 137
rect 381 89 407 123
rect 441 89 451 123
rect 381 55 451 89
rect 381 21 407 55
rect 441 21 451 55
rect 381 7 451 21
rect 481 49 535 137
rect 481 15 491 49
rect 525 15 535 49
rect 481 7 535 15
rect 565 123 617 137
rect 565 89 575 123
rect 609 89 617 123
rect 565 55 617 89
rect 565 21 575 55
rect 609 21 617 55
rect 565 7 617 21
<< pdiff >>
rect 27 437 83 457
rect 27 403 39 437
rect 73 403 83 437
rect 27 369 83 403
rect 27 335 39 369
rect 73 335 83 369
rect 27 301 83 335
rect 27 267 39 301
rect 73 267 83 301
rect 27 257 83 267
rect 113 437 262 457
rect 113 403 127 437
rect 161 403 218 437
rect 252 403 262 437
rect 113 369 262 403
rect 113 335 127 369
rect 161 335 218 369
rect 252 335 262 369
rect 113 257 262 335
rect 292 257 339 457
rect 369 437 463 457
rect 369 403 379 437
rect 413 403 463 437
rect 369 369 463 403
rect 369 335 379 369
rect 413 335 463 369
rect 369 301 463 335
rect 369 267 379 301
rect 413 267 463 301
rect 369 257 463 267
rect 493 257 535 457
rect 565 445 617 457
rect 565 411 575 445
rect 609 411 617 445
rect 565 377 617 411
rect 565 343 575 377
rect 609 343 617 377
rect 565 309 617 343
rect 565 275 575 309
rect 609 275 617 309
rect 565 257 617 275
<< ndiffc >>
rect 35 62 69 96
rect 119 19 153 53
rect 223 21 257 55
rect 307 89 341 123
rect 407 89 441 123
rect 407 21 441 55
rect 491 15 525 49
rect 575 89 609 123
rect 575 21 609 55
<< pdiffc >>
rect 39 403 73 437
rect 39 335 73 369
rect 39 267 73 301
rect 127 403 161 437
rect 218 403 252 437
rect 127 335 161 369
rect 218 335 252 369
rect 379 403 413 437
rect 379 335 413 369
rect 379 267 413 301
rect 575 411 609 445
rect 575 343 609 377
rect 575 275 609 309
<< poly >>
rect 83 457 113 483
rect 262 457 292 483
rect 339 457 369 483
rect 463 457 493 483
rect 535 457 565 483
rect 83 225 113 257
rect 262 225 292 257
rect 78 209 165 225
rect 78 175 121 209
rect 155 175 165 209
rect 78 159 165 175
rect 207 224 292 225
rect 339 225 369 257
rect 463 225 493 257
rect 207 209 297 224
rect 207 175 217 209
rect 251 175 297 209
rect 207 159 297 175
rect 339 209 393 225
rect 339 175 349 209
rect 383 175 393 209
rect 339 159 393 175
rect 435 209 493 225
rect 435 175 449 209
rect 483 175 493 209
rect 435 159 493 175
rect 535 225 565 257
rect 535 209 603 225
rect 535 175 550 209
rect 584 175 603 209
rect 535 159 603 175
rect 79 137 109 159
rect 267 137 297 159
rect 351 137 381 159
rect 451 137 481 159
rect 535 137 565 159
rect 79 -19 109 7
rect 267 -19 297 7
rect 351 -19 381 7
rect 451 -19 481 7
rect 535 -19 565 7
<< polycont >>
rect 121 175 155 209
rect 217 175 251 209
rect 349 175 383 209
rect 449 175 483 209
rect 550 175 584 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 17 437 73 453
rect 17 403 39 437
rect 17 369 73 403
rect 17 335 39 369
rect 111 437 268 487
rect 111 403 127 437
rect 161 403 218 437
rect 252 403 268 437
rect 111 369 268 403
rect 111 335 127 369
rect 161 335 218 369
rect 252 335 268 369
rect 347 437 424 453
rect 563 445 627 487
rect 347 403 379 437
rect 413 403 424 437
rect 347 369 424 403
rect 347 335 379 369
rect 413 335 424 369
rect 17 301 73 335
rect 347 321 424 335
rect 347 301 429 321
rect 17 267 39 301
rect 17 96 73 267
rect 107 267 379 301
rect 413 267 429 301
rect 489 283 529 441
rect 107 259 429 267
rect 107 209 162 259
rect 463 249 529 283
rect 563 411 575 445
rect 609 411 627 445
rect 563 377 627 411
rect 563 343 575 377
rect 609 343 627 377
rect 563 309 627 343
rect 563 275 575 309
rect 609 275 627 309
rect 563 251 627 275
rect 463 225 499 249
rect 107 175 121 209
rect 155 175 162 209
rect 196 209 267 225
rect 196 175 217 209
rect 251 175 267 209
rect 306 209 399 225
rect 306 175 349 209
rect 383 175 399 209
rect 433 209 499 225
rect 433 175 449 209
rect 483 175 499 209
rect 534 209 627 215
rect 534 175 550 209
rect 584 175 627 209
rect 107 139 162 175
rect 107 123 357 139
rect 107 103 307 123
rect 17 62 35 96
rect 69 62 73 96
rect 284 89 307 103
rect 341 89 357 123
rect 391 123 627 133
rect 391 89 407 123
rect 441 99 575 123
rect 441 89 457 99
rect 17 33 73 62
rect 119 53 153 69
rect 391 55 457 89
rect 559 89 575 99
rect 609 89 627 123
rect 207 21 223 55
rect 257 21 407 55
rect 441 21 457 55
rect 207 19 457 21
rect 491 49 525 65
rect 119 -23 153 19
rect 559 55 627 89
rect 559 21 575 55
rect 609 21 627 55
rect 559 16 627 21
rect 491 -23 525 15
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
<< metal1 >>
rect 0 521 644 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 0 456 644 487
rect 0 -23 644 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
rect 0 -88 644 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o22a_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 489 317 523 351 0 FreeSans 400 0 0 0 A2
port 8 nsew
flabel locali s 29 385 63 419 0 FreeSans 400 0 0 0 X
port 11 nsew
flabel locali s 213 181 247 215 0 FreeSans 400 0 0 0 B1
port 10 nsew
flabel locali s 581 181 615 215 0 FreeSans 400 0 0 0 A1
port 9 nsew
flabel locali s 310 181 344 215 0 FreeSans 400 0 0 0 B2
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 644 504
string path 0.000 -1.000 16.100 -1.000 
<< end >>
