VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sar_analog
  CLASS CORE ;
  FOREIGN sar_analog ;
  ORIGIN 0.000 0.000 ;
  SIZE 178.795 BY 120.810 ;
  SITE unithddbl ;
  PIN ctlp7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 77.155 149.035 77.485 ;
      LAYER mcon ;
        RECT 148.790 77.260 148.990 77.460 ;
      LAYER met1 ;
        RECT 148.760 77.200 149.020 77.520 ;
      LAYER via ;
        RECT 148.760 77.230 149.020 77.490 ;
      LAYER met2 ;
        RECT 148.730 77.445 149.050 77.490 ;
        RECT 148.730 77.275 151.450 77.445 ;
        RECT 148.730 77.230 149.050 77.275 ;
    END
  END ctlp7
  PIN ctlp6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 78.530 149.035 78.860 ;
      LAYER mcon ;
        RECT 148.805 78.630 149.005 78.830 ;
      LAYER met1 ;
        RECT 148.775 78.570 149.035 78.890 ;
      LAYER via ;
        RECT 148.775 78.600 149.035 78.860 ;
      LAYER met2 ;
        RECT 148.745 78.815 149.065 78.860 ;
        RECT 148.745 78.645 151.480 78.815 ;
        RECT 148.745 78.600 149.065 78.645 ;
    END
  END ctlp6
  PIN ctlp5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 79.900 149.035 80.230 ;
      LAYER mcon ;
        RECT 148.795 80.005 148.995 80.205 ;
      LAYER met1 ;
        RECT 148.765 79.945 149.025 80.265 ;
      LAYER via ;
        RECT 148.765 79.975 149.025 80.235 ;
      LAYER met2 ;
        RECT 148.735 80.190 149.055 80.235 ;
        RECT 148.735 80.020 151.520 80.190 ;
        RECT 148.735 79.975 149.055 80.020 ;
    END
  END ctlp5
  PIN ctlp4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 81.275 149.035 81.605 ;
      LAYER mcon ;
        RECT 148.790 81.385 148.990 81.585 ;
      LAYER met1 ;
        RECT 148.760 81.325 149.020 81.645 ;
      LAYER via ;
        RECT 148.760 81.355 149.020 81.615 ;
      LAYER met2 ;
        RECT 148.730 81.570 149.050 81.615 ;
        RECT 148.730 81.400 151.510 81.570 ;
        RECT 148.730 81.355 149.050 81.400 ;
    END
  END ctlp4
  PIN ctlp3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 82.650 149.035 82.980 ;
      LAYER mcon ;
        RECT 148.795 82.760 148.995 82.960 ;
      LAYER met1 ;
        RECT 148.765 82.700 149.025 83.020 ;
      LAYER via ;
        RECT 148.765 82.730 149.025 82.990 ;
      LAYER met2 ;
        RECT 148.735 82.945 149.055 82.990 ;
        RECT 148.735 82.775 151.510 82.945 ;
        RECT 148.735 82.730 149.055 82.775 ;
    END
  END ctlp3
  PIN ctlp2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 84.030 149.035 84.360 ;
      LAYER mcon ;
        RECT 148.795 84.130 148.995 84.330 ;
      LAYER met1 ;
        RECT 148.765 84.070 149.025 84.390 ;
      LAYER via ;
        RECT 148.765 84.100 149.025 84.360 ;
      LAYER met2 ;
        RECT 148.735 84.315 149.055 84.360 ;
        RECT 148.735 84.145 151.510 84.315 ;
        RECT 148.735 84.100 149.055 84.145 ;
    END
  END ctlp2
  PIN ctlp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 85.405 149.035 85.735 ;
      LAYER mcon ;
        RECT 148.795 85.515 148.995 85.715 ;
      LAYER met1 ;
        RECT 148.765 85.455 149.025 85.775 ;
      LAYER via ;
        RECT 148.765 85.485 149.025 85.745 ;
      LAYER met2 ;
        RECT 148.735 85.700 149.055 85.745 ;
        RECT 148.735 85.530 151.510 85.700 ;
        RECT 148.735 85.485 149.055 85.530 ;
    END
  END ctlp1
  PIN ctlp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 86.775 149.035 87.105 ;
      LAYER mcon ;
        RECT 148.810 86.870 149.010 87.070 ;
      LAYER met1 ;
        RECT 148.780 86.810 149.040 87.130 ;
      LAYER via ;
        RECT 148.780 86.840 149.040 87.100 ;
      LAYER met2 ;
        RECT 148.750 87.055 149.070 87.100 ;
        RECT 148.750 86.885 151.520 87.055 ;
        RECT 148.750 86.840 149.070 86.885 ;
    END
  END ctlp0
  PIN ctln7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 42.365 149.035 42.695 ;
      LAYER mcon ;
        RECT 148.790 42.390 148.990 42.590 ;
      LAYER met1 ;
        RECT 148.760 42.330 149.020 42.650 ;
      LAYER via ;
        RECT 148.760 42.360 149.020 42.620 ;
      LAYER met2 ;
        RECT 148.730 42.575 149.050 42.620 ;
        RECT 148.730 42.405 151.500 42.575 ;
        RECT 148.730 42.360 149.050 42.405 ;
    END
  END ctln7
  PIN ctln6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 40.990 149.035 41.320 ;
      LAYER mcon ;
        RECT 148.805 41.020 149.005 41.220 ;
      LAYER met1 ;
        RECT 148.775 40.960 149.035 41.280 ;
      LAYER via ;
        RECT 148.775 40.990 149.035 41.250 ;
      LAYER met2 ;
        RECT 148.745 41.205 149.065 41.250 ;
        RECT 148.745 41.035 151.500 41.205 ;
        RECT 148.745 40.990 149.065 41.035 ;
    END
  END ctln6
  PIN ctln5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 39.620 149.035 39.950 ;
      LAYER mcon ;
        RECT 148.795 39.645 148.995 39.845 ;
      LAYER met1 ;
        RECT 148.765 39.585 149.025 39.905 ;
      LAYER via ;
        RECT 148.765 39.615 149.025 39.875 ;
      LAYER met2 ;
        RECT 148.735 39.830 149.055 39.875 ;
        RECT 148.735 39.660 151.500 39.830 ;
        RECT 148.735 39.615 149.055 39.660 ;
    END
  END ctln5
  PIN ctln4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 38.245 149.035 38.575 ;
      LAYER mcon ;
        RECT 148.790 38.265 148.990 38.465 ;
      LAYER met1 ;
        RECT 148.760 38.205 149.020 38.525 ;
      LAYER via ;
        RECT 148.760 38.235 149.020 38.495 ;
      LAYER met2 ;
        RECT 148.730 38.450 149.050 38.495 ;
        RECT 148.730 38.280 151.490 38.450 ;
        RECT 148.730 38.235 149.050 38.280 ;
    END
  END ctln4
  PIN ctln3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 36.870 149.035 37.200 ;
      LAYER mcon ;
        RECT 148.795 36.890 148.995 37.090 ;
      LAYER met1 ;
        RECT 148.765 36.830 149.025 37.150 ;
      LAYER via ;
        RECT 148.765 36.860 149.025 37.120 ;
      LAYER met2 ;
        RECT 148.735 37.075 149.055 37.120 ;
        RECT 148.735 36.905 151.470 37.075 ;
        RECT 148.735 36.860 149.055 36.905 ;
    END
  END ctln3
  PIN ctln2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 35.490 149.035 35.820 ;
      LAYER mcon ;
        RECT 148.795 35.520 148.995 35.720 ;
      LAYER met1 ;
        RECT 148.765 35.460 149.025 35.780 ;
      LAYER via ;
        RECT 148.765 35.490 149.025 35.750 ;
      LAYER met2 ;
        RECT 148.735 35.705 149.055 35.750 ;
        RECT 148.735 35.535 151.440 35.705 ;
        RECT 148.735 35.490 149.055 35.535 ;
    END
  END ctln2
  PIN ctln1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 34.115 149.035 34.445 ;
      LAYER mcon ;
        RECT 148.795 34.135 148.995 34.335 ;
      LAYER met1 ;
        RECT 148.765 34.075 149.025 34.395 ;
      LAYER via ;
        RECT 148.765 34.105 149.025 34.365 ;
      LAYER met2 ;
        RECT 148.735 34.320 149.055 34.365 ;
        RECT 148.735 34.150 151.430 34.320 ;
        RECT 148.735 34.105 149.055 34.150 ;
    END
  END ctln1
  PIN ctln0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 148.785 32.745 149.035 33.075 ;
      LAYER mcon ;
        RECT 148.810 32.780 149.010 32.980 ;
      LAYER met1 ;
        RECT 148.780 32.720 149.040 33.040 ;
      LAYER via ;
        RECT 148.780 32.750 149.040 33.010 ;
      LAYER met2 ;
        RECT 148.750 32.965 149.070 33.010 ;
        RECT 148.750 32.795 151.450 32.965 ;
        RECT 148.750 32.750 149.070 32.795 ;
    END
  END ctln0
  PIN trim4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER li1 ;
        RECT 150.920 50.665 151.250 50.835 ;
        RECT 151.510 50.665 151.840 50.835 ;
        RECT 152.100 50.665 152.430 50.835 ;
        RECT 152.690 50.665 153.020 50.835 ;
        RECT 153.280 50.665 153.610 50.835 ;
        RECT 153.870 50.665 154.200 50.835 ;
        RECT 154.460 50.665 154.790 50.835 ;
        RECT 155.050 50.665 155.380 50.835 ;
        RECT 153.620 44.950 153.850 50.165 ;
      LAYER mcon ;
        RECT 151.000 50.665 151.170 50.835 ;
        RECT 151.590 50.665 151.760 50.835 ;
        RECT 152.180 50.665 152.350 50.835 ;
        RECT 152.770 50.665 152.940 50.835 ;
        RECT 153.360 50.665 153.530 50.835 ;
        RECT 153.950 50.665 154.120 50.835 ;
        RECT 154.540 50.665 154.710 50.835 ;
        RECT 155.130 50.665 155.300 50.835 ;
        RECT 153.650 49.965 153.820 50.135 ;
        RECT 153.620 44.980 153.850 45.210 ;
      LAYER met1 ;
        RECT 150.940 50.635 155.375 50.865 ;
        RECT 153.620 49.905 153.850 50.635 ;
        RECT 153.590 44.920 153.880 45.270 ;
        RECT 153.620 43.545 153.850 44.920 ;
    END
  END trim4
  PIN trim3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 158.910 50.665 159.240 50.835 ;
        RECT 159.500 50.665 159.830 50.835 ;
        RECT 160.090 50.665 160.420 50.835 ;
        RECT 160.680 50.665 161.010 50.835 ;
        RECT 159.830 44.980 160.060 46.320 ;
      LAYER mcon ;
        RECT 158.990 50.665 159.160 50.835 ;
        RECT 159.580 50.665 159.750 50.835 ;
        RECT 160.170 50.665 160.340 50.835 ;
        RECT 160.760 50.665 160.930 50.835 ;
        RECT 159.860 46.120 160.030 46.290 ;
      LAYER met1 ;
        RECT 158.930 50.635 160.990 50.865 ;
        RECT 159.830 46.060 160.060 50.635 ;
        RECT 159.800 44.920 160.080 45.270 ;
        RECT 159.830 43.470 160.050 44.920 ;
    END
  END trim3
  PIN trim2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 163.815 50.665 164.145 50.835 ;
        RECT 164.405 50.665 164.735 50.835 ;
        RECT 165.270 45.000 165.500 47.735 ;
      LAYER mcon ;
        RECT 163.895 50.665 164.065 50.835 ;
        RECT 164.485 50.665 164.655 50.835 ;
        RECT 165.300 47.535 165.470 47.705 ;
      LAYER met1 ;
        RECT 163.825 50.860 164.130 50.900 ;
        RECT 164.415 50.860 164.720 50.895 ;
        RECT 163.825 50.630 165.500 50.860 ;
        RECT 163.825 50.600 164.130 50.630 ;
        RECT 164.415 50.595 164.720 50.630 ;
        RECT 165.270 47.475 165.500 50.630 ;
        RECT 165.240 44.940 165.530 45.290 ;
        RECT 165.270 43.515 165.500 44.940 ;
    END
  END trim2
  PIN trim1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 167.900 51.140 168.070 51.470 ;
        RECT 167.865 45.025 168.085 47.810 ;
      LAYER mcon ;
        RECT 167.900 51.220 168.070 51.390 ;
        RECT 167.890 47.615 168.060 47.785 ;
      LAYER met1 ;
        RECT 167.845 51.155 168.135 51.455 ;
        RECT 167.865 47.845 168.085 51.155 ;
        RECT 167.860 47.555 168.090 47.845 ;
        RECT 167.805 44.995 168.145 45.275 ;
        RECT 167.865 43.500 168.085 44.995 ;
    END
  END trim1
  PIN trim0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 170.695 51.075 170.865 51.405 ;
      LAYER mcon ;
        RECT 170.695 51.155 170.865 51.325 ;
      LAYER met1 ;
        RECT 170.640 51.370 170.930 51.390 ;
        RECT 170.640 51.120 171.785 51.370 ;
        RECT 170.640 51.090 170.930 51.120 ;
        RECT 171.535 43.415 171.785 51.120 ;
    END
  END trim0
  PIN trimb4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER li1 ;
        RECT 153.505 69.815 153.735 75.030 ;
        RECT 150.805 69.145 151.135 69.315 ;
        RECT 151.395 69.145 151.725 69.315 ;
        RECT 151.985 69.145 152.315 69.315 ;
        RECT 152.575 69.145 152.905 69.315 ;
        RECT 153.165 69.145 153.495 69.315 ;
        RECT 153.755 69.145 154.085 69.315 ;
        RECT 154.345 69.145 154.675 69.315 ;
        RECT 154.935 69.145 155.265 69.315 ;
      LAYER mcon ;
        RECT 153.505 74.770 153.735 75.000 ;
        RECT 153.535 69.845 153.705 70.015 ;
        RECT 150.885 69.145 151.055 69.315 ;
        RECT 151.475 69.145 151.645 69.315 ;
        RECT 152.065 69.145 152.235 69.315 ;
        RECT 152.655 69.145 152.825 69.315 ;
        RECT 153.245 69.145 153.415 69.315 ;
        RECT 153.835 69.145 154.005 69.315 ;
        RECT 154.425 69.145 154.595 69.315 ;
        RECT 155.015 69.145 155.185 69.315 ;
      LAYER met1 ;
        RECT 153.505 75.060 153.735 76.090 ;
        RECT 153.475 74.710 153.765 75.060 ;
        RECT 153.505 69.345 153.735 70.075 ;
        RECT 150.825 69.115 155.260 69.345 ;
    END
  END trimb4
  PIN trimb3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 159.715 73.660 159.945 75.000 ;
        RECT 158.795 69.145 159.125 69.315 ;
        RECT 159.385 69.145 159.715 69.315 ;
        RECT 159.975 69.145 160.305 69.315 ;
        RECT 160.565 69.145 160.895 69.315 ;
      LAYER mcon ;
        RECT 159.715 74.770 159.935 75.000 ;
        RECT 159.745 73.690 159.915 73.860 ;
        RECT 158.875 69.145 159.045 69.315 ;
        RECT 159.465 69.145 159.635 69.315 ;
        RECT 160.055 69.145 160.225 69.315 ;
        RECT 160.645 69.145 160.815 69.315 ;
      LAYER met1 ;
        RECT 159.715 75.060 159.935 76.090 ;
        RECT 159.685 74.710 159.965 75.060 ;
        RECT 159.715 69.345 159.945 73.920 ;
        RECT 158.815 69.115 160.875 69.345 ;
    END
  END trimb3
  PIN trimb2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 165.155 72.245 165.385 74.980 ;
        RECT 163.700 69.145 164.030 69.315 ;
        RECT 164.290 69.145 164.620 69.315 ;
      LAYER mcon ;
        RECT 165.155 74.750 165.385 74.980 ;
        RECT 165.185 72.275 165.355 72.445 ;
        RECT 163.780 69.145 163.950 69.315 ;
        RECT 164.370 69.145 164.540 69.315 ;
      LAYER met1 ;
        RECT 165.155 75.040 165.385 76.090 ;
        RECT 165.125 74.690 165.415 75.040 ;
        RECT 163.710 69.350 164.015 69.380 ;
        RECT 164.300 69.350 164.605 69.385 ;
        RECT 165.155 69.350 165.385 72.505 ;
        RECT 163.710 69.120 165.385 69.350 ;
        RECT 163.710 69.080 164.015 69.120 ;
        RECT 164.300 69.085 164.605 69.120 ;
    END
  END trimb2
  PIN trimb1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 167.750 72.170 167.970 74.955 ;
        RECT 167.785 68.510 167.955 68.840 ;
      LAYER mcon ;
        RECT 167.750 74.735 167.970 74.955 ;
        RECT 167.775 72.195 167.945 72.365 ;
        RECT 167.785 68.590 167.955 68.760 ;
      LAYER met1 ;
        RECT 167.750 74.985 167.970 76.090 ;
        RECT 167.690 74.705 168.030 74.985 ;
        RECT 167.745 72.135 167.975 72.425 ;
        RECT 167.750 68.825 167.970 72.135 ;
        RECT 167.730 68.525 168.020 68.825 ;
    END
  END trimb1
  PIN trimb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 170.580 68.575 170.750 68.905 ;
      LAYER mcon ;
        RECT 170.580 68.655 170.750 68.825 ;
      LAYER met1 ;
        RECT 170.525 68.860 170.815 68.890 ;
        RECT 171.420 68.860 171.670 76.090 ;
        RECT 170.525 68.610 171.670 68.860 ;
        RECT 170.525 68.590 170.815 68.610 ;
    END
  END trimb0
  PIN vinp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.920000 ;
    PORT
      LAYER li1 ;
        RECT 12.185 76.370 12.355 77.230 ;
        RECT 13.365 76.370 13.535 77.230 ;
        RECT 14.545 76.370 14.715 77.230 ;
        RECT 15.725 76.370 15.895 77.230 ;
        RECT 16.905 76.370 17.075 77.230 ;
        RECT 18.085 76.370 18.255 77.230 ;
        RECT 21.800 76.370 21.970 77.230 ;
        RECT 22.980 76.370 23.150 77.230 ;
        RECT 24.160 76.370 24.330 77.230 ;
        RECT 25.340 76.370 25.510 77.230 ;
        RECT 26.520 76.370 26.690 77.230 ;
        RECT 27.700 76.370 27.870 77.230 ;
        RECT 31.415 76.370 31.585 77.230 ;
        RECT 32.595 76.370 32.765 77.230 ;
        RECT 33.775 76.370 33.945 77.230 ;
        RECT 34.955 76.370 35.125 77.230 ;
        RECT 36.135 76.370 36.305 77.230 ;
        RECT 37.315 76.370 37.485 77.230 ;
        RECT 41.030 76.370 41.200 77.230 ;
        RECT 42.210 76.370 42.380 77.230 ;
        RECT 43.390 76.370 43.560 77.230 ;
        RECT 44.570 76.370 44.740 77.230 ;
        RECT 45.750 76.370 45.920 77.230 ;
        RECT 46.930 76.370 47.100 77.230 ;
        RECT 12.195 73.885 12.365 74.745 ;
        RECT 13.375 73.885 13.545 74.745 ;
        RECT 14.555 73.885 14.725 74.745 ;
        RECT 15.735 73.885 15.905 74.745 ;
        RECT 16.915 73.885 17.085 74.745 ;
        RECT 18.095 73.885 18.265 74.745 ;
        RECT 21.810 73.885 21.980 74.745 ;
        RECT 22.990 73.885 23.160 74.745 ;
        RECT 24.170 73.885 24.340 74.745 ;
        RECT 25.350 73.885 25.520 74.745 ;
        RECT 26.530 73.885 26.700 74.745 ;
        RECT 27.710 73.885 27.880 74.745 ;
        RECT 31.425 73.885 31.595 74.745 ;
        RECT 32.605 73.885 32.775 74.745 ;
        RECT 33.785 73.885 33.955 74.745 ;
        RECT 34.965 73.885 35.135 74.745 ;
        RECT 36.145 73.885 36.315 74.745 ;
        RECT 37.325 73.885 37.495 74.745 ;
        RECT 41.040 73.885 41.210 74.745 ;
        RECT 42.220 73.885 42.390 74.745 ;
        RECT 43.400 73.885 43.570 74.745 ;
        RECT 44.580 73.885 44.750 74.745 ;
        RECT 45.760 73.885 45.930 74.745 ;
        RECT 46.940 73.885 47.110 74.745 ;
      LAYER mcon ;
        RECT 12.185 76.450 12.355 77.150 ;
        RECT 13.365 76.450 13.535 77.150 ;
        RECT 14.545 76.450 14.715 77.150 ;
        RECT 15.725 76.450 15.895 77.150 ;
        RECT 16.905 76.450 17.075 77.150 ;
        RECT 18.085 76.450 18.255 77.150 ;
        RECT 21.800 76.450 21.970 77.150 ;
        RECT 22.980 76.450 23.150 77.150 ;
        RECT 24.160 76.450 24.330 77.150 ;
        RECT 25.340 76.450 25.510 77.150 ;
        RECT 26.520 76.450 26.690 77.150 ;
        RECT 27.700 76.450 27.870 77.150 ;
        RECT 31.415 76.450 31.585 77.150 ;
        RECT 32.595 76.450 32.765 77.150 ;
        RECT 33.775 76.450 33.945 77.150 ;
        RECT 34.955 76.450 35.125 77.150 ;
        RECT 36.135 76.450 36.305 77.150 ;
        RECT 37.315 76.450 37.485 77.150 ;
        RECT 41.030 76.450 41.200 77.150 ;
        RECT 42.210 76.450 42.380 77.150 ;
        RECT 43.390 76.450 43.560 77.150 ;
        RECT 44.570 76.450 44.740 77.150 ;
        RECT 45.750 76.450 45.920 77.150 ;
        RECT 46.930 76.450 47.100 77.150 ;
        RECT 12.195 73.965 12.365 74.665 ;
        RECT 13.375 73.965 13.545 74.665 ;
        RECT 14.555 73.965 14.725 74.665 ;
        RECT 15.735 73.965 15.905 74.665 ;
        RECT 16.915 73.965 17.085 74.665 ;
        RECT 18.095 73.965 18.265 74.665 ;
        RECT 21.810 73.965 21.980 74.665 ;
        RECT 22.990 73.965 23.160 74.665 ;
        RECT 24.170 73.965 24.340 74.665 ;
        RECT 25.350 73.965 25.520 74.665 ;
        RECT 26.530 73.965 26.700 74.665 ;
        RECT 27.710 73.965 27.880 74.665 ;
        RECT 31.425 73.965 31.595 74.665 ;
        RECT 32.605 73.965 32.775 74.665 ;
        RECT 33.785 73.965 33.955 74.665 ;
        RECT 34.965 73.965 35.135 74.665 ;
        RECT 36.145 73.965 36.315 74.665 ;
        RECT 37.325 73.965 37.495 74.665 ;
        RECT 41.040 73.965 41.210 74.665 ;
        RECT 42.220 73.965 42.390 74.665 ;
        RECT 43.400 73.965 43.570 74.665 ;
        RECT 44.580 73.965 44.750 74.665 ;
        RECT 45.760 73.965 45.930 74.665 ;
        RECT 46.940 73.965 47.110 74.665 ;
      LAYER met1 ;
        RECT 12.155 76.390 12.385 77.210 ;
        RECT 13.335 76.390 13.565 77.210 ;
        RECT 14.515 76.390 14.745 77.210 ;
        RECT 15.695 76.390 15.925 77.210 ;
        RECT 16.875 76.390 17.105 77.210 ;
        RECT 18.055 76.390 18.285 77.210 ;
        RECT 21.770 76.390 22.000 77.210 ;
        RECT 22.950 76.390 23.180 77.210 ;
        RECT 24.130 76.390 24.360 77.210 ;
        RECT 25.310 76.390 25.540 77.210 ;
        RECT 26.490 76.390 26.720 77.210 ;
        RECT 27.670 76.390 27.900 77.210 ;
        RECT 31.385 76.390 31.615 77.210 ;
        RECT 32.565 76.390 32.795 77.210 ;
        RECT 33.745 76.390 33.975 77.210 ;
        RECT 34.925 76.390 35.155 77.210 ;
        RECT 36.105 76.390 36.335 77.210 ;
        RECT 37.285 76.390 37.515 77.210 ;
        RECT 41.000 76.390 41.230 77.210 ;
        RECT 42.180 76.390 42.410 77.210 ;
        RECT 43.360 76.390 43.590 77.210 ;
        RECT 44.540 76.390 44.770 77.210 ;
        RECT 45.720 76.390 45.950 77.210 ;
        RECT 46.900 76.390 47.130 77.210 ;
        RECT 10.865 75.655 11.575 75.665 ;
        RECT 12.180 75.655 12.360 76.390 ;
        RECT 13.355 75.655 13.535 76.390 ;
        RECT 14.540 75.655 14.720 76.390 ;
        RECT 15.715 75.655 15.895 76.390 ;
        RECT 16.915 75.655 17.095 76.390 ;
        RECT 18.080 75.655 18.260 76.390 ;
        RECT 21.795 75.655 21.975 76.390 ;
        RECT 22.970 75.655 23.150 76.390 ;
        RECT 24.155 75.655 24.335 76.390 ;
        RECT 25.330 75.655 25.510 76.390 ;
        RECT 26.530 75.655 26.710 76.390 ;
        RECT 27.695 75.655 27.875 76.390 ;
        RECT 31.410 75.655 31.590 76.390 ;
        RECT 32.585 75.655 32.765 76.390 ;
        RECT 33.770 75.655 33.950 76.390 ;
        RECT 34.945 75.655 35.125 76.390 ;
        RECT 36.145 75.655 36.325 76.390 ;
        RECT 37.310 75.655 37.490 76.390 ;
        RECT 41.025 75.655 41.205 76.390 ;
        RECT 42.200 75.655 42.380 76.390 ;
        RECT 43.385 75.655 43.565 76.390 ;
        RECT 44.560 75.655 44.740 76.390 ;
        RECT 45.760 75.655 45.940 76.390 ;
        RECT 46.925 75.655 47.105 76.390 ;
        RECT 10.865 75.485 18.260 75.655 ;
        RECT 20.965 75.650 27.875 75.655 ;
        RECT 30.580 75.650 37.490 75.655 ;
        RECT 10.865 72.720 11.045 75.485 ;
        RECT 11.350 75.475 18.260 75.485 ;
        RECT 12.180 75.470 18.260 75.475 ;
        RECT 12.180 75.465 13.535 75.470 ;
        RECT 12.180 74.725 12.360 75.465 ;
        RECT 13.355 74.725 13.535 75.465 ;
        RECT 14.540 74.725 14.720 75.470 ;
        RECT 15.715 74.725 15.895 75.470 ;
        RECT 16.915 74.725 17.095 75.470 ;
        RECT 18.080 74.725 18.260 75.470 ;
        RECT 20.955 75.475 27.875 75.650 ;
        RECT 12.165 73.905 12.395 74.725 ;
        RECT 13.345 73.905 13.575 74.725 ;
        RECT 14.525 73.905 14.755 74.725 ;
        RECT 15.705 73.905 15.935 74.725 ;
        RECT 16.885 73.905 17.115 74.725 ;
        RECT 18.065 73.905 18.295 74.725 ;
        RECT 20.955 72.720 21.135 75.475 ;
        RECT 21.795 75.470 27.875 75.475 ;
        RECT 21.795 75.465 23.150 75.470 ;
        RECT 21.795 74.725 21.975 75.465 ;
        RECT 22.970 74.725 23.150 75.465 ;
        RECT 24.155 74.725 24.335 75.470 ;
        RECT 25.330 74.725 25.510 75.470 ;
        RECT 26.530 74.725 26.710 75.470 ;
        RECT 27.695 74.725 27.875 75.470 ;
        RECT 30.575 75.475 37.490 75.650 ;
        RECT 21.780 73.905 22.010 74.725 ;
        RECT 22.960 73.905 23.190 74.725 ;
        RECT 24.140 73.905 24.370 74.725 ;
        RECT 25.320 73.905 25.550 74.725 ;
        RECT 26.500 73.905 26.730 74.725 ;
        RECT 27.680 73.905 27.910 74.725 ;
        RECT 30.575 72.720 30.755 75.475 ;
        RECT 31.410 75.470 37.490 75.475 ;
        RECT 31.410 75.465 32.765 75.470 ;
        RECT 31.410 74.725 31.590 75.465 ;
        RECT 32.585 74.725 32.765 75.465 ;
        RECT 33.770 74.725 33.950 75.470 ;
        RECT 34.945 74.725 35.125 75.470 ;
        RECT 36.145 74.725 36.325 75.470 ;
        RECT 37.310 74.725 37.490 75.470 ;
        RECT 40.195 75.475 47.105 75.655 ;
        RECT 31.395 73.905 31.625 74.725 ;
        RECT 32.575 73.905 32.805 74.725 ;
        RECT 33.755 73.905 33.985 74.725 ;
        RECT 34.935 73.905 35.165 74.725 ;
        RECT 36.115 73.905 36.345 74.725 ;
        RECT 37.295 73.905 37.525 74.725 ;
        RECT 40.195 72.720 40.375 75.475 ;
        RECT 41.025 75.470 47.105 75.475 ;
        RECT 41.025 75.465 42.380 75.470 ;
        RECT 41.025 74.725 41.205 75.465 ;
        RECT 42.200 74.725 42.380 75.465 ;
        RECT 43.385 74.725 43.565 75.470 ;
        RECT 44.560 74.725 44.740 75.470 ;
        RECT 45.760 74.725 45.940 75.470 ;
        RECT 46.925 74.725 47.105 75.470 ;
        RECT 41.010 73.905 41.240 74.725 ;
        RECT 42.190 73.905 42.420 74.725 ;
        RECT 43.370 73.905 43.600 74.725 ;
        RECT 44.550 73.905 44.780 74.725 ;
        RECT 45.730 73.905 45.960 74.725 ;
        RECT 46.910 73.905 47.140 74.725 ;
        RECT 0.755 72.540 40.375 72.720 ;
    END
  END vinp
  PIN vinn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.920000 ;
    PORT
      LAYER li1 ;
        RECT 12.195 45.105 12.365 45.965 ;
        RECT 13.375 45.105 13.545 45.965 ;
        RECT 14.555 45.105 14.725 45.965 ;
        RECT 15.735 45.105 15.905 45.965 ;
        RECT 16.915 45.105 17.085 45.965 ;
        RECT 18.095 45.105 18.265 45.965 ;
        RECT 21.810 45.105 21.980 45.965 ;
        RECT 22.990 45.105 23.160 45.965 ;
        RECT 24.170 45.105 24.340 45.965 ;
        RECT 25.350 45.105 25.520 45.965 ;
        RECT 26.530 45.105 26.700 45.965 ;
        RECT 27.710 45.105 27.880 45.965 ;
        RECT 31.425 45.105 31.595 45.965 ;
        RECT 32.605 45.105 32.775 45.965 ;
        RECT 33.785 45.105 33.955 45.965 ;
        RECT 34.965 45.105 35.135 45.965 ;
        RECT 36.145 45.105 36.315 45.965 ;
        RECT 37.325 45.105 37.495 45.965 ;
        RECT 41.040 45.105 41.210 45.965 ;
        RECT 42.220 45.105 42.390 45.965 ;
        RECT 43.400 45.105 43.570 45.965 ;
        RECT 44.580 45.105 44.750 45.965 ;
        RECT 45.760 45.105 45.930 45.965 ;
        RECT 46.940 45.105 47.110 45.965 ;
        RECT 12.185 42.620 12.355 43.480 ;
        RECT 13.365 42.620 13.535 43.480 ;
        RECT 14.545 42.620 14.715 43.480 ;
        RECT 15.725 42.620 15.895 43.480 ;
        RECT 16.905 42.620 17.075 43.480 ;
        RECT 18.085 42.620 18.255 43.480 ;
        RECT 21.800 42.620 21.970 43.480 ;
        RECT 22.980 42.620 23.150 43.480 ;
        RECT 24.160 42.620 24.330 43.480 ;
        RECT 25.340 42.620 25.510 43.480 ;
        RECT 26.520 42.620 26.690 43.480 ;
        RECT 27.700 42.620 27.870 43.480 ;
        RECT 31.415 42.620 31.585 43.480 ;
        RECT 32.595 42.620 32.765 43.480 ;
        RECT 33.775 42.620 33.945 43.480 ;
        RECT 34.955 42.620 35.125 43.480 ;
        RECT 36.135 42.620 36.305 43.480 ;
        RECT 37.315 42.620 37.485 43.480 ;
        RECT 41.030 42.620 41.200 43.480 ;
        RECT 42.210 42.620 42.380 43.480 ;
        RECT 43.390 42.620 43.560 43.480 ;
        RECT 44.570 42.620 44.740 43.480 ;
        RECT 45.750 42.620 45.920 43.480 ;
        RECT 46.930 42.620 47.100 43.480 ;
      LAYER mcon ;
        RECT 12.195 45.185 12.365 45.885 ;
        RECT 13.375 45.185 13.545 45.885 ;
        RECT 14.555 45.185 14.725 45.885 ;
        RECT 15.735 45.185 15.905 45.885 ;
        RECT 16.915 45.185 17.085 45.885 ;
        RECT 18.095 45.185 18.265 45.885 ;
        RECT 21.810 45.185 21.980 45.885 ;
        RECT 22.990 45.185 23.160 45.885 ;
        RECT 24.170 45.185 24.340 45.885 ;
        RECT 25.350 45.185 25.520 45.885 ;
        RECT 26.530 45.185 26.700 45.885 ;
        RECT 27.710 45.185 27.880 45.885 ;
        RECT 31.425 45.185 31.595 45.885 ;
        RECT 32.605 45.185 32.775 45.885 ;
        RECT 33.785 45.185 33.955 45.885 ;
        RECT 34.965 45.185 35.135 45.885 ;
        RECT 36.145 45.185 36.315 45.885 ;
        RECT 37.325 45.185 37.495 45.885 ;
        RECT 41.040 45.185 41.210 45.885 ;
        RECT 42.220 45.185 42.390 45.885 ;
        RECT 43.400 45.185 43.570 45.885 ;
        RECT 44.580 45.185 44.750 45.885 ;
        RECT 45.760 45.185 45.930 45.885 ;
        RECT 46.940 45.185 47.110 45.885 ;
        RECT 12.185 42.700 12.355 43.400 ;
        RECT 13.365 42.700 13.535 43.400 ;
        RECT 14.545 42.700 14.715 43.400 ;
        RECT 15.725 42.700 15.895 43.400 ;
        RECT 16.905 42.700 17.075 43.400 ;
        RECT 18.085 42.700 18.255 43.400 ;
        RECT 21.800 42.700 21.970 43.400 ;
        RECT 22.980 42.700 23.150 43.400 ;
        RECT 24.160 42.700 24.330 43.400 ;
        RECT 25.340 42.700 25.510 43.400 ;
        RECT 26.520 42.700 26.690 43.400 ;
        RECT 27.700 42.700 27.870 43.400 ;
        RECT 31.415 42.700 31.585 43.400 ;
        RECT 32.595 42.700 32.765 43.400 ;
        RECT 33.775 42.700 33.945 43.400 ;
        RECT 34.955 42.700 35.125 43.400 ;
        RECT 36.135 42.700 36.305 43.400 ;
        RECT 37.315 42.700 37.485 43.400 ;
        RECT 41.030 42.700 41.200 43.400 ;
        RECT 42.210 42.700 42.380 43.400 ;
        RECT 43.390 42.700 43.560 43.400 ;
        RECT 44.570 42.700 44.740 43.400 ;
        RECT 45.750 42.700 45.920 43.400 ;
        RECT 46.930 42.700 47.100 43.400 ;
      LAYER met1 ;
        RECT 0.925 47.130 40.375 47.310 ;
        RECT 10.865 44.365 11.045 47.130 ;
        RECT 12.165 45.125 12.395 45.945 ;
        RECT 13.345 45.125 13.575 45.945 ;
        RECT 14.525 45.125 14.755 45.945 ;
        RECT 15.705 45.125 15.935 45.945 ;
        RECT 16.885 45.125 17.115 45.945 ;
        RECT 18.065 45.125 18.295 45.945 ;
        RECT 12.180 44.385 12.360 45.125 ;
        RECT 13.355 44.385 13.535 45.125 ;
        RECT 12.180 44.380 13.535 44.385 ;
        RECT 14.540 44.380 14.720 45.125 ;
        RECT 15.715 44.380 15.895 45.125 ;
        RECT 16.915 44.380 17.095 45.125 ;
        RECT 18.080 44.380 18.260 45.125 ;
        RECT 12.180 44.375 18.260 44.380 ;
        RECT 11.350 44.365 18.260 44.375 ;
        RECT 10.865 44.195 18.260 44.365 ;
        RECT 20.955 44.375 21.135 47.130 ;
        RECT 21.780 45.125 22.010 45.945 ;
        RECT 22.960 45.125 23.190 45.945 ;
        RECT 24.140 45.125 24.370 45.945 ;
        RECT 25.320 45.125 25.550 45.945 ;
        RECT 26.500 45.125 26.730 45.945 ;
        RECT 27.680 45.125 27.910 45.945 ;
        RECT 21.795 44.385 21.975 45.125 ;
        RECT 22.970 44.385 23.150 45.125 ;
        RECT 21.795 44.380 23.150 44.385 ;
        RECT 24.155 44.380 24.335 45.125 ;
        RECT 25.330 44.380 25.510 45.125 ;
        RECT 26.530 44.380 26.710 45.125 ;
        RECT 27.695 44.380 27.875 45.125 ;
        RECT 21.795 44.375 27.875 44.380 ;
        RECT 20.955 44.200 27.875 44.375 ;
        RECT 30.575 44.375 30.755 47.130 ;
        RECT 31.395 45.125 31.625 45.945 ;
        RECT 32.575 45.125 32.805 45.945 ;
        RECT 33.755 45.125 33.985 45.945 ;
        RECT 34.935 45.125 35.165 45.945 ;
        RECT 36.115 45.125 36.345 45.945 ;
        RECT 37.295 45.125 37.525 45.945 ;
        RECT 31.410 44.385 31.590 45.125 ;
        RECT 32.585 44.385 32.765 45.125 ;
        RECT 31.410 44.380 32.765 44.385 ;
        RECT 33.770 44.380 33.950 45.125 ;
        RECT 34.945 44.380 35.125 45.125 ;
        RECT 36.145 44.380 36.325 45.125 ;
        RECT 37.310 44.380 37.490 45.125 ;
        RECT 31.410 44.375 37.490 44.380 ;
        RECT 30.575 44.200 37.490 44.375 ;
        RECT 20.965 44.195 27.875 44.200 ;
        RECT 30.580 44.195 37.490 44.200 ;
        RECT 40.195 44.375 40.375 47.130 ;
        RECT 41.010 45.125 41.240 45.945 ;
        RECT 42.190 45.125 42.420 45.945 ;
        RECT 43.370 45.125 43.600 45.945 ;
        RECT 44.550 45.125 44.780 45.945 ;
        RECT 45.730 45.125 45.960 45.945 ;
        RECT 46.910 45.125 47.140 45.945 ;
        RECT 41.025 44.385 41.205 45.125 ;
        RECT 42.200 44.385 42.380 45.125 ;
        RECT 41.025 44.380 42.380 44.385 ;
        RECT 43.385 44.380 43.565 45.125 ;
        RECT 44.560 44.380 44.740 45.125 ;
        RECT 45.760 44.380 45.940 45.125 ;
        RECT 46.925 44.380 47.105 45.125 ;
        RECT 41.025 44.375 47.105 44.380 ;
        RECT 40.195 44.195 47.105 44.375 ;
        RECT 10.865 44.185 11.575 44.195 ;
        RECT 12.180 43.460 12.360 44.195 ;
        RECT 13.355 43.460 13.535 44.195 ;
        RECT 14.540 43.460 14.720 44.195 ;
        RECT 15.715 43.460 15.895 44.195 ;
        RECT 16.915 43.460 17.095 44.195 ;
        RECT 18.080 43.460 18.260 44.195 ;
        RECT 21.795 43.460 21.975 44.195 ;
        RECT 22.970 43.460 23.150 44.195 ;
        RECT 24.155 43.460 24.335 44.195 ;
        RECT 25.330 43.460 25.510 44.195 ;
        RECT 26.530 43.460 26.710 44.195 ;
        RECT 27.695 43.460 27.875 44.195 ;
        RECT 31.410 43.460 31.590 44.195 ;
        RECT 32.585 43.460 32.765 44.195 ;
        RECT 33.770 43.460 33.950 44.195 ;
        RECT 34.945 43.460 35.125 44.195 ;
        RECT 36.145 43.460 36.325 44.195 ;
        RECT 37.310 43.460 37.490 44.195 ;
        RECT 41.025 43.460 41.205 44.195 ;
        RECT 42.200 43.460 42.380 44.195 ;
        RECT 43.385 43.460 43.565 44.195 ;
        RECT 44.560 43.460 44.740 44.195 ;
        RECT 45.760 43.460 45.940 44.195 ;
        RECT 46.925 43.460 47.105 44.195 ;
        RECT 12.155 42.640 12.385 43.460 ;
        RECT 13.335 42.640 13.565 43.460 ;
        RECT 14.515 42.640 14.745 43.460 ;
        RECT 15.695 42.640 15.925 43.460 ;
        RECT 16.875 42.640 17.105 43.460 ;
        RECT 18.055 42.640 18.285 43.460 ;
        RECT 21.770 42.640 22.000 43.460 ;
        RECT 22.950 42.640 23.180 43.460 ;
        RECT 24.130 42.640 24.360 43.460 ;
        RECT 25.310 42.640 25.540 43.460 ;
        RECT 26.490 42.640 26.720 43.460 ;
        RECT 27.670 42.640 27.900 43.460 ;
        RECT 31.385 42.640 31.615 43.460 ;
        RECT 32.565 42.640 32.795 43.460 ;
        RECT 33.745 42.640 33.975 43.460 ;
        RECT 34.925 42.640 35.155 43.460 ;
        RECT 36.105 42.640 36.335 43.460 ;
        RECT 37.285 42.640 37.515 43.460 ;
        RECT 41.000 42.640 41.230 43.460 ;
        RECT 42.180 42.640 42.410 43.460 ;
        RECT 43.360 42.640 43.590 43.460 ;
        RECT 44.540 42.640 44.770 43.460 ;
        RECT 45.720 42.640 45.950 43.460 ;
        RECT 46.900 42.640 47.130 43.460 ;
    END
  END vinn
  PIN sample
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.920000 ;
    PORT
      LAYER li1 ;
        RECT 14.520 80.425 16.150 80.675 ;
        RECT 24.135 80.425 25.765 80.675 ;
        RECT 33.750 80.425 35.380 80.675 ;
        RECT 43.365 80.425 44.995 80.675 ;
        RECT 14.520 39.175 16.150 39.425 ;
        RECT 24.135 39.175 25.765 39.425 ;
        RECT 33.750 39.175 35.380 39.425 ;
        RECT 43.365 39.175 44.995 39.425 ;
      LAYER mcon ;
        RECT 14.590 80.455 14.790 80.655 ;
        RECT 24.205 80.455 24.405 80.655 ;
        RECT 33.820 80.455 34.020 80.655 ;
        RECT 43.435 80.455 43.635 80.655 ;
        RECT 14.590 39.195 14.790 39.395 ;
        RECT 24.205 39.195 24.405 39.395 ;
        RECT 33.820 39.195 34.020 39.395 ;
        RECT 43.435 39.195 43.635 39.395 ;
      LAYER met1 ;
        RECT 14.530 80.425 14.850 80.685 ;
        RECT 24.145 80.425 24.465 80.685 ;
        RECT 33.760 80.425 34.080 80.685 ;
        RECT 43.375 80.425 43.695 80.685 ;
        RECT 14.530 39.165 14.850 39.425 ;
        RECT 24.145 39.165 24.465 39.425 ;
        RECT 33.760 39.165 34.080 39.425 ;
        RECT 43.375 39.165 43.695 39.425 ;
      LAYER via ;
        RECT 14.560 80.425 14.820 80.685 ;
        RECT 24.175 80.425 24.435 80.685 ;
        RECT 33.790 80.425 34.050 80.685 ;
        RECT 43.405 80.425 43.665 80.685 ;
        RECT 14.560 39.165 14.820 39.425 ;
        RECT 24.175 39.165 24.435 39.425 ;
        RECT 33.790 39.165 34.050 39.425 ;
        RECT 43.405 39.165 43.665 39.425 ;
      LAYER met2 ;
        RECT 6.525 82.105 43.655 82.310 ;
        RECT 6.525 37.745 6.730 82.105 ;
        RECT 14.585 80.715 14.790 82.105 ;
        RECT 24.200 80.715 24.405 82.105 ;
        RECT 33.815 80.715 34.020 82.105 ;
        RECT 43.430 80.715 43.635 82.105 ;
        RECT 14.560 80.395 14.820 80.715 ;
        RECT 24.175 80.395 24.435 80.715 ;
        RECT 33.790 80.395 34.050 80.715 ;
        RECT 43.405 80.395 43.665 80.715 ;
        RECT 14.560 39.135 14.820 39.455 ;
        RECT 24.175 39.135 24.435 39.455 ;
        RECT 33.790 39.135 34.050 39.455 ;
        RECT 43.405 39.135 43.665 39.455 ;
        RECT 14.585 37.745 14.790 39.135 ;
        RECT 24.200 37.745 24.405 39.135 ;
        RECT 33.815 37.745 34.020 39.135 ;
        RECT 43.430 37.745 43.635 39.135 ;
        RECT 6.525 37.540 43.655 37.745 ;
    END
  END sample
  PIN comp
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.800000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 172.895 61.505 173.935 61.675 ;
        RECT 176.320 61.505 177.360 61.675 ;
        RECT 174.105 59.375 174.275 59.775 ;
        RECT 175.935 59.375 176.105 59.775 ;
        RECT 172.895 58.265 173.935 58.435 ;
      LAYER mcon ;
        RECT 173.150 61.505 173.320 61.675 ;
        RECT 173.510 61.505 173.680 61.675 ;
        RECT 176.575 61.505 176.745 61.675 ;
        RECT 176.935 61.505 177.105 61.675 ;
        RECT 174.105 59.490 174.275 59.660 ;
        RECT 175.935 59.490 176.105 59.660 ;
        RECT 173.150 58.265 173.320 58.435 ;
        RECT 173.510 58.265 173.680 58.435 ;
      LAYER met1 ;
        RECT 172.915 61.475 173.915 61.705 ;
        RECT 176.340 61.475 177.340 61.705 ;
        RECT 173.065 61.405 173.765 61.475 ;
        RECT 176.490 61.405 177.190 61.475 ;
        RECT 174.755 61.355 175.455 61.390 ;
        RECT 174.755 61.125 176.135 61.355 ;
        RECT 174.755 61.090 175.455 61.125 ;
        RECT 175.905 60.905 176.135 61.125 ;
        RECT 175.905 60.605 178.795 60.905 ;
        RECT 175.905 59.755 176.135 60.605 ;
        RECT 174.075 59.395 176.135 59.755 ;
        RECT 174.955 58.915 175.255 59.395 ;
        RECT 173.615 58.615 175.255 58.915 ;
        RECT 173.615 58.465 173.915 58.615 ;
        RECT 172.915 58.235 173.915 58.465 ;
      LAYER via ;
        RECT 173.125 61.425 173.385 61.685 ;
        RECT 173.445 61.425 173.705 61.685 ;
        RECT 176.550 61.425 176.810 61.685 ;
        RECT 176.870 61.425 177.130 61.685 ;
        RECT 174.815 61.110 175.075 61.370 ;
        RECT 175.135 61.110 175.395 61.370 ;
      LAYER met2 ;
        RECT 173.115 61.670 173.715 61.755 ;
        RECT 176.540 61.670 177.140 61.755 ;
        RECT 173.115 61.440 177.140 61.670 ;
        RECT 173.115 61.355 173.715 61.440 ;
        RECT 174.805 61.040 175.405 61.440 ;
        RECT 176.540 61.355 177.140 61.440 ;
    END
  END comp
  PIN clkc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 163.655 60.890 163.825 61.220 ;
        RECT 165.480 60.890 165.650 61.220 ;
        RECT 153.920 60.325 154.250 60.495 ;
        RECT 153.920 59.745 154.250 59.915 ;
        RECT 163.655 59.095 163.825 59.425 ;
        RECT 165.480 59.095 165.650 59.425 ;
      LAYER mcon ;
        RECT 163.655 60.970 163.825 61.140 ;
        RECT 165.480 60.970 165.650 61.140 ;
        RECT 154.000 60.325 154.170 60.495 ;
        RECT 154.000 59.745 154.170 59.915 ;
        RECT 163.655 59.175 163.825 59.345 ;
        RECT 165.480 59.175 165.650 59.345 ;
      LAYER met1 ;
        RECT 163.660 61.205 163.810 61.240 ;
        RECT 163.590 60.905 163.870 61.205 ;
        RECT 165.430 60.905 165.710 61.205 ;
        RECT 153.935 60.260 154.235 60.560 ;
        RECT 153.990 59.980 154.140 60.260 ;
        RECT 153.935 59.960 154.235 59.980 ;
        RECT 153.905 59.700 154.235 59.960 ;
        RECT 153.935 59.680 154.235 59.700 ;
        RECT 163.660 59.410 163.810 60.905 ;
        RECT 165.470 59.410 165.620 60.905 ;
        RECT 163.590 59.385 163.870 59.410 ;
        RECT 165.430 59.400 165.710 59.410 ;
        RECT 163.575 59.125 163.895 59.385 ;
        RECT 165.385 59.140 165.710 59.400 ;
        RECT 163.590 59.110 163.870 59.125 ;
        RECT 165.430 59.110 165.710 59.140 ;
      LAYER via ;
        RECT 153.935 59.700 154.195 59.960 ;
        RECT 163.605 59.125 163.865 59.385 ;
        RECT 165.415 59.140 165.675 59.400 ;
      LAYER met2 ;
        RECT 171.195 67.210 178.665 67.350 ;
        RECT 153.935 59.670 154.195 59.990 ;
        RECT 153.990 58.140 154.140 59.670 ;
        RECT 163.605 59.095 163.865 59.415 ;
        RECT 165.415 59.110 165.675 59.430 ;
        RECT 163.660 58.140 163.810 59.095 ;
        RECT 165.470 58.140 165.620 59.110 ;
        RECT 171.195 58.140 171.335 67.210 ;
        RECT 153.990 57.990 171.340 58.140 ;
    END
  END clkc
  PIN avdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 9.635 78.840 50.315 80.445 ;
        RECT 10.555 78.350 49.400 78.840 ;
        RECT 11.445 72.715 19.015 75.555 ;
        RECT 21.060 72.715 28.630 75.555 ;
        RECT 30.675 72.715 38.245 75.555 ;
        RECT 40.290 72.715 47.860 75.555 ;
        RECT 159.855 58.080 166.345 62.235 ;
        RECT 175.125 54.990 178.495 66.520 ;
        RECT 11.445 44.295 19.015 47.135 ;
        RECT 21.060 44.295 28.630 47.135 ;
        RECT 30.675 44.295 38.245 47.135 ;
        RECT 40.290 44.295 47.860 47.135 ;
        RECT 10.555 41.010 49.400 41.500 ;
        RECT 9.635 39.405 50.315 41.010 ;
      LAYER li1 ;
        RECT 148.785 88.150 149.035 88.480 ;
        RECT 150.345 88.460 150.515 89.490 ;
        RECT 149.205 88.230 150.515 88.460 ;
        RECT 150.345 87.560 150.515 88.230 ;
        RECT 149.205 87.350 150.515 87.560 ;
        RECT 150.345 87.085 150.515 87.350 ;
        RECT 149.205 86.855 150.515 87.085 ;
        RECT 150.345 86.185 150.515 86.855 ;
        RECT 149.205 85.975 150.515 86.185 ;
        RECT 150.345 85.715 150.515 85.975 ;
        RECT 149.205 85.485 150.515 85.715 ;
        RECT 150.345 84.815 150.515 85.485 ;
        RECT 149.205 84.605 150.515 84.815 ;
        RECT 150.345 84.340 150.515 84.605 ;
        RECT 149.205 84.110 150.515 84.340 ;
        RECT 150.345 83.440 150.515 84.110 ;
        RECT 149.205 83.230 150.515 83.440 ;
        RECT 150.345 82.960 150.515 83.230 ;
        RECT 149.205 82.730 150.515 82.960 ;
        RECT 150.345 82.060 150.515 82.730 ;
        RECT 149.205 81.850 150.515 82.060 ;
        RECT 150.345 81.585 150.515 81.850 ;
        RECT 149.205 81.355 150.515 81.585 ;
        RECT 9.910 79.295 10.660 80.280 ;
        RECT 12.650 80.205 14.340 80.725 ;
        RECT 10.830 79.115 14.340 80.205 ;
        RECT 14.545 79.115 14.810 80.255 ;
        RECT 15.480 79.115 15.650 79.915 ;
        RECT 16.320 79.115 16.530 79.575 ;
        RECT 16.810 79.115 17.075 80.255 ;
        RECT 19.755 80.205 20.275 80.745 ;
        RECT 22.265 80.205 23.955 80.725 ;
        RECT 17.745 79.115 17.915 79.915 ;
        RECT 18.585 79.115 18.795 79.575 ;
        RECT 19.065 79.115 20.275 80.205 ;
        RECT 20.445 79.115 23.955 80.205 ;
        RECT 24.160 79.115 24.425 80.255 ;
        RECT 25.095 79.115 25.265 79.915 ;
        RECT 25.935 79.115 26.145 79.575 ;
        RECT 26.425 79.115 26.690 80.255 ;
        RECT 29.370 80.205 29.890 80.745 ;
        RECT 31.880 80.205 33.570 80.725 ;
        RECT 27.360 79.115 27.530 79.915 ;
        RECT 28.200 79.115 28.410 79.575 ;
        RECT 28.680 79.115 29.890 80.205 ;
        RECT 30.060 79.115 33.570 80.205 ;
        RECT 33.775 79.115 34.040 80.255 ;
        RECT 34.710 79.115 34.880 79.915 ;
        RECT 35.550 79.115 35.760 79.575 ;
        RECT 36.040 79.115 36.305 80.255 ;
        RECT 38.985 80.205 39.505 80.745 ;
        RECT 41.495 80.205 43.185 80.725 ;
        RECT 36.975 79.115 37.145 79.915 ;
        RECT 37.815 79.115 38.025 79.575 ;
        RECT 38.295 79.115 39.505 80.205 ;
        RECT 39.675 79.115 43.185 80.205 ;
        RECT 43.390 79.115 43.655 80.255 ;
        RECT 44.325 79.115 44.495 79.915 ;
        RECT 45.165 79.115 45.375 79.575 ;
        RECT 45.655 79.115 45.920 80.255 ;
        RECT 48.600 80.205 49.120 80.745 ;
        RECT 150.345 80.685 150.515 81.355 ;
        RECT 149.205 80.475 150.515 80.685 ;
        RECT 46.590 79.115 46.760 79.915 ;
        RECT 47.430 79.115 47.640 79.575 ;
        RECT 47.910 79.115 49.120 80.205 ;
        RECT 49.290 79.295 50.040 80.280 ;
        RECT 150.345 80.210 150.515 80.475 ;
        RECT 149.205 79.980 150.515 80.210 ;
        RECT 150.345 79.310 150.515 79.980 ;
        RECT 9.825 78.945 50.125 79.115 ;
        RECT 149.205 79.100 150.515 79.310 ;
        RECT 11.605 78.560 13.015 78.945 ;
        RECT 21.220 78.560 22.630 78.945 ;
        RECT 30.835 78.560 32.245 78.945 ;
        RECT 40.450 78.560 41.860 78.945 ;
        RECT 150.345 78.840 150.515 79.100 ;
        RECT 149.205 78.610 150.515 78.840 ;
        RECT 150.345 77.940 150.515 78.610 ;
        RECT 149.205 77.730 150.515 77.940 ;
        RECT 150.345 77.465 150.515 77.730 ;
        RECT 149.205 77.235 150.515 77.465 ;
        RECT 150.345 76.565 150.515 77.235 ;
        RECT 149.205 76.355 150.515 76.565 ;
        RECT 150.345 75.575 150.515 76.355 ;
        RECT 171.970 75.575 172.200 75.655 ;
        RECT 150.345 75.345 172.200 75.575 ;
        RECT 150.345 75.305 150.515 75.345 ;
        RECT 11.625 73.450 11.795 74.820 ;
        RECT 18.665 74.390 18.835 74.820 ;
        RECT 18.660 73.735 18.835 74.390 ;
        RECT 18.665 73.450 18.835 73.735 ;
        RECT 21.240 73.450 21.410 74.820 ;
        RECT 28.280 74.390 28.450 74.820 ;
        RECT 28.275 73.735 28.450 74.390 ;
        RECT 28.280 73.450 28.450 73.735 ;
        RECT 30.855 73.450 31.025 74.820 ;
        RECT 37.895 74.390 38.065 74.820 ;
        RECT 37.890 73.735 38.065 74.390 ;
        RECT 37.895 73.450 38.065 73.735 ;
        RECT 40.470 73.450 40.640 74.820 ;
        RECT 47.510 74.390 47.680 74.820 ;
        RECT 47.505 73.735 47.680 74.390 ;
        RECT 47.510 73.450 47.680 73.735 ;
        RECT 12.650 72.895 17.810 73.065 ;
        RECT 22.265 72.895 27.425 73.065 ;
        RECT 31.880 72.895 37.040 73.065 ;
        RECT 41.495 72.895 46.655 73.065 ;
        RECT 171.970 67.135 172.200 75.345 ;
        RECT 175.305 67.135 175.535 67.190 ;
        RECT 168.500 66.905 175.535 67.135 ;
        RECT 160.985 60.675 161.845 60.845 ;
        RECT 162.490 60.675 163.350 60.845 ;
        RECT 164.315 60.675 165.175 60.845 ;
        RECT 161.360 60.285 161.620 60.675 ;
        RECT 162.805 60.285 163.065 60.675 ;
        RECT 164.645 60.285 164.905 60.675 ;
        RECT 168.500 60.285 168.730 66.905 ;
        RECT 161.090 60.030 168.730 60.285 ;
        RECT 175.305 66.340 175.535 66.905 ;
        RECT 175.305 66.170 178.315 66.340 ;
        RECT 161.090 60.025 168.425 60.030 ;
        RECT 161.360 60.015 164.905 60.025 ;
        RECT 161.360 59.640 161.620 60.015 ;
        RECT 162.805 59.995 164.905 60.015 ;
        RECT 162.805 59.640 163.065 59.995 ;
        RECT 164.645 59.640 164.905 59.995 ;
        RECT 160.985 59.470 161.845 59.640 ;
        RECT 162.490 59.470 163.350 59.640 ;
        RECT 164.315 59.470 165.175 59.640 ;
        RECT 175.305 55.340 175.475 66.170 ;
        RECT 176.320 65.335 177.360 65.505 ;
        RECT 176.320 62.195 177.360 62.365 ;
        RECT 176.320 59.145 177.360 59.315 ;
        RECT 176.320 56.005 177.360 56.175 ;
        RECT 178.145 55.340 178.315 66.170 ;
        RECT 175.305 55.170 178.315 55.340 ;
        RECT 12.650 46.785 17.810 46.955 ;
        RECT 22.265 46.785 27.425 46.955 ;
        RECT 31.880 46.785 37.040 46.955 ;
        RECT 41.495 46.785 46.655 46.955 ;
        RECT 11.625 45.030 11.795 46.400 ;
        RECT 18.665 46.115 18.835 46.400 ;
        RECT 18.660 45.460 18.835 46.115 ;
        RECT 18.665 45.030 18.835 45.460 ;
        RECT 21.240 45.030 21.410 46.400 ;
        RECT 28.280 46.115 28.450 46.400 ;
        RECT 28.275 45.460 28.450 46.115 ;
        RECT 28.280 45.030 28.450 45.460 ;
        RECT 30.855 45.030 31.025 46.400 ;
        RECT 37.895 46.115 38.065 46.400 ;
        RECT 37.890 45.460 38.065 46.115 ;
        RECT 37.895 45.030 38.065 45.460 ;
        RECT 40.470 45.030 40.640 46.400 ;
        RECT 47.510 46.115 47.680 46.400 ;
        RECT 47.505 45.460 47.680 46.115 ;
        RECT 47.510 45.030 47.680 45.460 ;
        RECT 150.345 43.495 150.515 44.545 ;
        RECT 149.205 43.285 150.515 43.495 ;
        RECT 150.345 42.615 150.515 43.285 ;
        RECT 149.205 42.385 150.515 42.615 ;
        RECT 150.345 42.120 150.515 42.385 ;
        RECT 149.205 41.910 150.515 42.120 ;
        RECT 11.605 40.905 13.015 41.290 ;
        RECT 21.220 40.905 22.630 41.290 ;
        RECT 30.835 40.905 32.245 41.290 ;
        RECT 40.450 40.905 41.860 41.290 ;
        RECT 150.345 41.240 150.515 41.910 ;
        RECT 149.205 41.010 150.515 41.240 ;
        RECT 9.825 40.735 50.125 40.905 ;
        RECT 150.345 40.750 150.515 41.010 ;
        RECT 9.910 39.570 10.660 40.555 ;
        RECT 10.830 39.645 14.340 40.735 ;
        RECT 12.650 39.125 14.340 39.645 ;
        RECT 14.545 39.595 14.810 40.735 ;
        RECT 15.480 39.935 15.650 40.735 ;
        RECT 16.320 40.275 16.530 40.735 ;
        RECT 16.810 39.595 17.075 40.735 ;
        RECT 17.745 39.935 17.915 40.735 ;
        RECT 18.585 40.275 18.795 40.735 ;
        RECT 19.065 39.645 20.275 40.735 ;
        RECT 20.445 39.645 23.955 40.735 ;
        RECT 19.755 39.105 20.275 39.645 ;
        RECT 22.265 39.125 23.955 39.645 ;
        RECT 24.160 39.595 24.425 40.735 ;
        RECT 25.095 39.935 25.265 40.735 ;
        RECT 25.935 40.275 26.145 40.735 ;
        RECT 26.425 39.595 26.690 40.735 ;
        RECT 27.360 39.935 27.530 40.735 ;
        RECT 28.200 40.275 28.410 40.735 ;
        RECT 28.680 39.645 29.890 40.735 ;
        RECT 30.060 39.645 33.570 40.735 ;
        RECT 29.370 39.105 29.890 39.645 ;
        RECT 31.880 39.125 33.570 39.645 ;
        RECT 33.775 39.595 34.040 40.735 ;
        RECT 34.710 39.935 34.880 40.735 ;
        RECT 35.550 40.275 35.760 40.735 ;
        RECT 36.040 39.595 36.305 40.735 ;
        RECT 36.975 39.935 37.145 40.735 ;
        RECT 37.815 40.275 38.025 40.735 ;
        RECT 38.295 39.645 39.505 40.735 ;
        RECT 39.675 39.645 43.185 40.735 ;
        RECT 38.985 39.105 39.505 39.645 ;
        RECT 41.495 39.125 43.185 39.645 ;
        RECT 43.390 39.595 43.655 40.735 ;
        RECT 44.325 39.935 44.495 40.735 ;
        RECT 45.165 40.275 45.375 40.735 ;
        RECT 45.655 39.595 45.920 40.735 ;
        RECT 46.590 39.935 46.760 40.735 ;
        RECT 47.430 40.275 47.640 40.735 ;
        RECT 47.910 39.645 49.120 40.735 ;
        RECT 48.600 39.105 49.120 39.645 ;
        RECT 49.290 39.570 50.040 40.555 ;
        RECT 149.205 40.540 150.515 40.750 ;
        RECT 150.345 39.870 150.515 40.540 ;
        RECT 149.205 39.640 150.515 39.870 ;
        RECT 150.345 39.375 150.515 39.640 ;
        RECT 149.205 39.165 150.515 39.375 ;
        RECT 150.345 38.495 150.515 39.165 ;
        RECT 149.205 38.265 150.515 38.495 ;
        RECT 150.345 38.000 150.515 38.265 ;
        RECT 149.205 37.790 150.515 38.000 ;
        RECT 150.345 37.120 150.515 37.790 ;
        RECT 149.205 36.890 150.515 37.120 ;
        RECT 150.345 36.620 150.515 36.890 ;
        RECT 149.205 36.410 150.515 36.620 ;
        RECT 150.345 35.740 150.515 36.410 ;
        RECT 149.205 35.510 150.515 35.740 ;
        RECT 150.345 35.245 150.515 35.510 ;
        RECT 149.205 35.035 150.515 35.245 ;
        RECT 150.345 34.365 150.515 35.035 ;
        RECT 149.205 34.135 150.515 34.365 ;
        RECT 150.345 33.875 150.515 34.135 ;
        RECT 149.205 33.665 150.515 33.875 ;
        RECT 150.345 32.995 150.515 33.665 ;
        RECT 149.205 32.765 150.515 32.995 ;
        RECT 150.345 32.500 150.515 32.765 ;
        RECT 149.205 32.290 150.515 32.500 ;
        RECT 150.345 31.620 150.515 32.290 ;
        RECT 149.205 31.390 150.515 31.620 ;
        RECT 150.345 30.360 150.515 31.390 ;
      LAYER mcon ;
        RECT 150.345 89.175 150.515 89.345 ;
        RECT 150.345 88.715 150.515 88.885 ;
        RECT 148.810 88.260 149.010 88.460 ;
        RECT 150.345 88.270 150.515 88.440 ;
        RECT 150.345 87.810 150.515 87.980 ;
        RECT 150.345 87.350 150.515 87.520 ;
        RECT 150.345 86.895 150.515 87.065 ;
        RECT 150.345 86.435 150.515 86.605 ;
        RECT 150.345 85.975 150.515 86.145 ;
        RECT 150.345 85.525 150.515 85.695 ;
        RECT 150.345 85.065 150.515 85.235 ;
        RECT 150.345 84.605 150.515 84.775 ;
        RECT 150.345 84.150 150.515 84.320 ;
        RECT 150.345 83.690 150.515 83.860 ;
        RECT 150.345 83.230 150.515 83.400 ;
        RECT 150.345 82.770 150.515 82.940 ;
        RECT 150.345 82.310 150.515 82.480 ;
        RECT 150.345 81.850 150.515 82.020 ;
        RECT 150.345 81.395 150.515 81.565 ;
        RECT 150.345 80.935 150.515 81.105 ;
        RECT 150.345 80.475 150.515 80.645 ;
        RECT 150.345 80.020 150.515 80.190 ;
        RECT 150.345 79.560 150.515 79.730 ;
        RECT 9.970 78.945 10.140 79.115 ;
        RECT 10.430 78.945 10.600 79.115 ;
        RECT 10.890 78.945 11.060 79.115 ;
        RECT 11.350 78.945 11.520 79.115 ;
        RECT 11.810 78.945 11.980 79.115 ;
        RECT 12.270 78.945 12.440 79.115 ;
        RECT 12.730 78.945 12.900 79.115 ;
        RECT 13.190 78.945 13.360 79.115 ;
        RECT 13.650 78.945 13.820 79.115 ;
        RECT 14.110 78.945 14.280 79.115 ;
        RECT 14.560 78.945 14.730 79.115 ;
        RECT 15.020 78.945 15.190 79.115 ;
        RECT 15.480 78.945 15.650 79.115 ;
        RECT 15.940 78.945 16.110 79.115 ;
        RECT 16.400 78.945 16.570 79.115 ;
        RECT 16.825 78.945 16.995 79.115 ;
        RECT 17.285 78.945 17.455 79.115 ;
        RECT 17.745 78.945 17.915 79.115 ;
        RECT 18.205 78.945 18.375 79.115 ;
        RECT 18.665 78.945 18.835 79.115 ;
        RECT 19.125 78.945 19.295 79.115 ;
        RECT 19.585 78.945 19.755 79.115 ;
        RECT 20.045 78.945 20.215 79.115 ;
        RECT 20.505 78.945 20.675 79.115 ;
        RECT 20.965 78.945 21.135 79.115 ;
        RECT 21.425 78.945 21.595 79.115 ;
        RECT 21.885 78.945 22.055 79.115 ;
        RECT 22.345 78.945 22.515 79.115 ;
        RECT 22.805 78.945 22.975 79.115 ;
        RECT 23.265 78.945 23.435 79.115 ;
        RECT 23.725 78.945 23.895 79.115 ;
        RECT 24.175 78.945 24.345 79.115 ;
        RECT 24.635 78.945 24.805 79.115 ;
        RECT 25.095 78.945 25.265 79.115 ;
        RECT 25.555 78.945 25.725 79.115 ;
        RECT 26.015 78.945 26.185 79.115 ;
        RECT 26.440 78.945 26.610 79.115 ;
        RECT 26.900 78.945 27.070 79.115 ;
        RECT 27.360 78.945 27.530 79.115 ;
        RECT 27.820 78.945 27.990 79.115 ;
        RECT 28.280 78.945 28.450 79.115 ;
        RECT 28.740 78.945 28.910 79.115 ;
        RECT 29.200 78.945 29.370 79.115 ;
        RECT 29.660 78.945 29.830 79.115 ;
        RECT 30.120 78.945 30.290 79.115 ;
        RECT 30.580 78.945 30.750 79.115 ;
        RECT 31.040 78.945 31.210 79.115 ;
        RECT 31.500 78.945 31.670 79.115 ;
        RECT 31.960 78.945 32.130 79.115 ;
        RECT 32.420 78.945 32.590 79.115 ;
        RECT 32.880 78.945 33.050 79.115 ;
        RECT 33.340 78.945 33.510 79.115 ;
        RECT 33.790 78.945 33.960 79.115 ;
        RECT 34.250 78.945 34.420 79.115 ;
        RECT 34.710 78.945 34.880 79.115 ;
        RECT 35.170 78.945 35.340 79.115 ;
        RECT 35.630 78.945 35.800 79.115 ;
        RECT 36.055 78.945 36.225 79.115 ;
        RECT 36.515 78.945 36.685 79.115 ;
        RECT 36.975 78.945 37.145 79.115 ;
        RECT 37.435 78.945 37.605 79.115 ;
        RECT 37.895 78.945 38.065 79.115 ;
        RECT 38.355 78.945 38.525 79.115 ;
        RECT 38.815 78.945 38.985 79.115 ;
        RECT 39.275 78.945 39.445 79.115 ;
        RECT 39.735 78.945 39.905 79.115 ;
        RECT 40.195 78.945 40.365 79.115 ;
        RECT 40.655 78.945 40.825 79.115 ;
        RECT 41.115 78.945 41.285 79.115 ;
        RECT 41.575 78.945 41.745 79.115 ;
        RECT 42.035 78.945 42.205 79.115 ;
        RECT 42.495 78.945 42.665 79.115 ;
        RECT 42.955 78.945 43.125 79.115 ;
        RECT 43.405 78.945 43.575 79.115 ;
        RECT 43.865 78.945 44.035 79.115 ;
        RECT 44.325 78.945 44.495 79.115 ;
        RECT 44.785 78.945 44.955 79.115 ;
        RECT 45.245 78.945 45.415 79.115 ;
        RECT 45.670 78.945 45.840 79.115 ;
        RECT 46.130 78.945 46.300 79.115 ;
        RECT 46.590 78.945 46.760 79.115 ;
        RECT 47.050 78.945 47.220 79.115 ;
        RECT 47.510 78.945 47.680 79.115 ;
        RECT 47.970 78.945 48.140 79.115 ;
        RECT 48.430 78.945 48.600 79.115 ;
        RECT 48.890 78.945 49.060 79.115 ;
        RECT 49.350 78.945 49.520 79.115 ;
        RECT 49.810 78.945 49.980 79.115 ;
        RECT 150.345 79.100 150.515 79.270 ;
        RECT 150.345 78.650 150.515 78.820 ;
        RECT 150.345 78.190 150.515 78.360 ;
        RECT 150.345 77.730 150.515 77.900 ;
        RECT 150.345 77.275 150.515 77.445 ;
        RECT 150.345 76.815 150.515 76.985 ;
        RECT 150.345 76.355 150.515 76.525 ;
        RECT 150.345 75.910 150.515 76.080 ;
        RECT 150.345 75.450 150.515 75.620 ;
        RECT 18.660 74.220 18.830 74.390 ;
        RECT 28.275 74.220 28.445 74.390 ;
        RECT 37.890 74.220 38.060 74.390 ;
        RECT 47.505 74.220 47.675 74.390 ;
        RECT 161.150 60.675 161.680 60.845 ;
        RECT 162.655 60.675 163.185 60.845 ;
        RECT 164.480 60.675 165.010 60.845 ;
        RECT 161.150 59.470 161.680 59.640 ;
        RECT 162.655 59.470 163.185 59.640 ;
        RECT 164.480 59.470 165.010 59.640 ;
        RECT 176.575 65.335 176.745 65.505 ;
        RECT 176.935 65.335 177.105 65.505 ;
        RECT 178.145 64.515 178.315 64.685 ;
        RECT 178.145 64.155 178.315 64.325 ;
        RECT 178.145 63.515 178.315 63.685 ;
        RECT 178.145 63.155 178.315 63.325 ;
        RECT 176.575 62.195 176.745 62.365 ;
        RECT 176.935 62.195 177.105 62.365 ;
        RECT 176.575 59.145 176.745 59.315 ;
        RECT 176.935 59.145 177.105 59.315 ;
        RECT 178.145 58.515 178.315 58.685 ;
        RECT 178.145 58.155 178.315 58.325 ;
        RECT 178.145 57.515 178.315 57.685 ;
        RECT 178.145 57.155 178.315 57.325 ;
        RECT 176.575 56.005 176.745 56.175 ;
        RECT 176.935 56.005 177.105 56.175 ;
        RECT 18.660 45.460 18.830 45.630 ;
        RECT 28.275 45.460 28.445 45.630 ;
        RECT 37.890 45.460 38.060 45.630 ;
        RECT 47.505 45.460 47.675 45.630 ;
        RECT 150.345 44.230 150.515 44.400 ;
        RECT 150.345 43.770 150.515 43.940 ;
        RECT 150.345 43.325 150.515 43.495 ;
        RECT 150.345 42.865 150.515 43.035 ;
        RECT 150.345 42.405 150.515 42.575 ;
        RECT 150.345 41.950 150.515 42.120 ;
        RECT 150.345 41.490 150.515 41.660 ;
        RECT 150.345 41.030 150.515 41.200 ;
        RECT 9.970 40.735 10.140 40.905 ;
        RECT 10.430 40.735 10.600 40.905 ;
        RECT 10.890 40.735 11.060 40.905 ;
        RECT 11.350 40.735 11.520 40.905 ;
        RECT 11.810 40.735 11.980 40.905 ;
        RECT 12.270 40.735 12.440 40.905 ;
        RECT 12.730 40.735 12.900 40.905 ;
        RECT 13.190 40.735 13.360 40.905 ;
        RECT 13.650 40.735 13.820 40.905 ;
        RECT 14.110 40.735 14.280 40.905 ;
        RECT 14.560 40.735 14.730 40.905 ;
        RECT 15.020 40.735 15.190 40.905 ;
        RECT 15.480 40.735 15.650 40.905 ;
        RECT 15.940 40.735 16.110 40.905 ;
        RECT 16.400 40.735 16.570 40.905 ;
        RECT 16.825 40.735 16.995 40.905 ;
        RECT 17.285 40.735 17.455 40.905 ;
        RECT 17.745 40.735 17.915 40.905 ;
        RECT 18.205 40.735 18.375 40.905 ;
        RECT 18.665 40.735 18.835 40.905 ;
        RECT 19.125 40.735 19.295 40.905 ;
        RECT 19.585 40.735 19.755 40.905 ;
        RECT 20.045 40.735 20.215 40.905 ;
        RECT 20.505 40.735 20.675 40.905 ;
        RECT 20.965 40.735 21.135 40.905 ;
        RECT 21.425 40.735 21.595 40.905 ;
        RECT 21.885 40.735 22.055 40.905 ;
        RECT 22.345 40.735 22.515 40.905 ;
        RECT 22.805 40.735 22.975 40.905 ;
        RECT 23.265 40.735 23.435 40.905 ;
        RECT 23.725 40.735 23.895 40.905 ;
        RECT 24.175 40.735 24.345 40.905 ;
        RECT 24.635 40.735 24.805 40.905 ;
        RECT 25.095 40.735 25.265 40.905 ;
        RECT 25.555 40.735 25.725 40.905 ;
        RECT 26.015 40.735 26.185 40.905 ;
        RECT 26.440 40.735 26.610 40.905 ;
        RECT 26.900 40.735 27.070 40.905 ;
        RECT 27.360 40.735 27.530 40.905 ;
        RECT 27.820 40.735 27.990 40.905 ;
        RECT 28.280 40.735 28.450 40.905 ;
        RECT 28.740 40.735 28.910 40.905 ;
        RECT 29.200 40.735 29.370 40.905 ;
        RECT 29.660 40.735 29.830 40.905 ;
        RECT 30.120 40.735 30.290 40.905 ;
        RECT 30.580 40.735 30.750 40.905 ;
        RECT 31.040 40.735 31.210 40.905 ;
        RECT 31.500 40.735 31.670 40.905 ;
        RECT 31.960 40.735 32.130 40.905 ;
        RECT 32.420 40.735 32.590 40.905 ;
        RECT 32.880 40.735 33.050 40.905 ;
        RECT 33.340 40.735 33.510 40.905 ;
        RECT 33.790 40.735 33.960 40.905 ;
        RECT 34.250 40.735 34.420 40.905 ;
        RECT 34.710 40.735 34.880 40.905 ;
        RECT 35.170 40.735 35.340 40.905 ;
        RECT 35.630 40.735 35.800 40.905 ;
        RECT 36.055 40.735 36.225 40.905 ;
        RECT 36.515 40.735 36.685 40.905 ;
        RECT 36.975 40.735 37.145 40.905 ;
        RECT 37.435 40.735 37.605 40.905 ;
        RECT 37.895 40.735 38.065 40.905 ;
        RECT 38.355 40.735 38.525 40.905 ;
        RECT 38.815 40.735 38.985 40.905 ;
        RECT 39.275 40.735 39.445 40.905 ;
        RECT 39.735 40.735 39.905 40.905 ;
        RECT 40.195 40.735 40.365 40.905 ;
        RECT 40.655 40.735 40.825 40.905 ;
        RECT 41.115 40.735 41.285 40.905 ;
        RECT 41.575 40.735 41.745 40.905 ;
        RECT 42.035 40.735 42.205 40.905 ;
        RECT 42.495 40.735 42.665 40.905 ;
        RECT 42.955 40.735 43.125 40.905 ;
        RECT 43.405 40.735 43.575 40.905 ;
        RECT 43.865 40.735 44.035 40.905 ;
        RECT 44.325 40.735 44.495 40.905 ;
        RECT 44.785 40.735 44.955 40.905 ;
        RECT 45.245 40.735 45.415 40.905 ;
        RECT 45.670 40.735 45.840 40.905 ;
        RECT 46.130 40.735 46.300 40.905 ;
        RECT 46.590 40.735 46.760 40.905 ;
        RECT 47.050 40.735 47.220 40.905 ;
        RECT 47.510 40.735 47.680 40.905 ;
        RECT 47.970 40.735 48.140 40.905 ;
        RECT 48.430 40.735 48.600 40.905 ;
        RECT 48.890 40.735 49.060 40.905 ;
        RECT 49.350 40.735 49.520 40.905 ;
        RECT 49.810 40.735 49.980 40.905 ;
        RECT 150.345 40.580 150.515 40.750 ;
        RECT 150.345 40.120 150.515 40.290 ;
        RECT 150.345 39.660 150.515 39.830 ;
        RECT 150.345 39.205 150.515 39.375 ;
        RECT 150.345 38.745 150.515 38.915 ;
        RECT 150.345 38.285 150.515 38.455 ;
        RECT 150.345 37.830 150.515 38.000 ;
        RECT 150.345 37.370 150.515 37.540 ;
        RECT 150.345 36.910 150.515 37.080 ;
        RECT 150.345 36.450 150.515 36.620 ;
        RECT 150.345 35.990 150.515 36.160 ;
        RECT 150.345 35.530 150.515 35.700 ;
        RECT 150.345 35.075 150.515 35.245 ;
        RECT 150.345 34.615 150.515 34.785 ;
        RECT 150.345 34.155 150.515 34.325 ;
        RECT 150.345 33.705 150.515 33.875 ;
        RECT 150.345 33.245 150.515 33.415 ;
        RECT 150.345 32.785 150.515 32.955 ;
        RECT 150.345 32.330 150.515 32.500 ;
        RECT 150.345 31.870 150.515 32.040 ;
        RECT 150.345 31.410 150.515 31.580 ;
        RECT 150.345 30.965 150.515 31.135 ;
        RECT 150.345 30.505 150.515 30.675 ;
      LAYER met1 ;
        RECT 6.155 118.280 17.565 118.610 ;
        RECT 6.155 107.390 6.295 118.280 ;
        RECT 6.715 107.390 6.855 118.280 ;
        RECT 7.275 107.390 7.415 118.280 ;
        RECT 7.835 107.390 7.975 118.280 ;
        RECT 8.395 107.390 8.535 118.280 ;
        RECT 8.955 107.390 9.095 118.280 ;
        RECT 9.515 107.390 9.655 118.280 ;
        RECT 10.075 107.390 10.215 118.280 ;
        RECT 10.635 107.390 10.775 118.280 ;
        RECT 11.195 107.390 11.335 118.280 ;
        RECT 11.755 107.390 11.895 118.280 ;
        RECT 12.315 107.390 12.455 118.280 ;
        RECT 12.875 107.390 13.015 118.280 ;
        RECT 13.435 107.390 13.575 118.280 ;
        RECT 13.995 107.390 14.135 118.280 ;
        RECT 14.555 107.390 14.695 118.280 ;
        RECT 15.115 107.390 15.255 118.280 ;
        RECT 15.675 107.390 15.815 118.280 ;
        RECT 16.235 107.390 16.375 118.280 ;
        RECT 16.795 107.390 16.935 118.280 ;
        RECT 17.355 107.390 17.565 118.280 ;
        RECT 19.245 118.280 30.655 118.610 ;
        RECT 19.245 107.390 19.385 118.280 ;
        RECT 19.805 107.390 19.945 118.280 ;
        RECT 20.365 107.390 20.505 118.280 ;
        RECT 20.925 107.390 21.065 118.280 ;
        RECT 21.485 107.390 21.625 118.280 ;
        RECT 22.045 107.390 22.185 118.280 ;
        RECT 22.605 107.390 22.745 118.280 ;
        RECT 23.165 107.390 23.305 118.280 ;
        RECT 23.725 107.390 23.865 118.280 ;
        RECT 24.285 107.390 24.425 118.280 ;
        RECT 24.845 107.390 24.985 118.280 ;
        RECT 25.405 107.390 25.545 118.280 ;
        RECT 25.965 107.390 26.105 118.280 ;
        RECT 26.525 107.390 26.665 118.280 ;
        RECT 27.085 107.390 27.225 118.280 ;
        RECT 27.645 107.390 27.785 118.280 ;
        RECT 28.205 107.390 28.345 118.280 ;
        RECT 28.765 107.390 28.905 118.280 ;
        RECT 29.325 107.390 29.465 118.280 ;
        RECT 29.885 107.390 30.025 118.280 ;
        RECT 30.445 107.390 30.655 118.280 ;
        RECT 32.335 118.260 43.745 118.590 ;
        RECT 32.335 107.370 32.475 118.260 ;
        RECT 32.895 107.370 33.035 118.260 ;
        RECT 33.455 107.370 33.595 118.260 ;
        RECT 34.015 107.370 34.155 118.260 ;
        RECT 34.575 107.370 34.715 118.260 ;
        RECT 35.135 107.370 35.275 118.260 ;
        RECT 35.695 107.370 35.835 118.260 ;
        RECT 36.255 107.370 36.395 118.260 ;
        RECT 36.815 107.370 36.955 118.260 ;
        RECT 37.375 107.370 37.515 118.260 ;
        RECT 37.935 107.370 38.075 118.260 ;
        RECT 38.495 107.370 38.635 118.260 ;
        RECT 39.055 107.370 39.195 118.260 ;
        RECT 39.615 107.370 39.755 118.260 ;
        RECT 40.175 107.370 40.315 118.260 ;
        RECT 40.735 107.370 40.875 118.260 ;
        RECT 41.295 107.370 41.435 118.260 ;
        RECT 41.855 107.370 41.995 118.260 ;
        RECT 42.415 107.370 42.555 118.260 ;
        RECT 42.975 107.370 43.115 118.260 ;
        RECT 43.535 107.370 43.745 118.260 ;
        RECT 45.425 118.260 56.835 118.590 ;
        RECT 45.425 107.370 45.565 118.260 ;
        RECT 45.985 107.370 46.125 118.260 ;
        RECT 46.545 107.370 46.685 118.260 ;
        RECT 47.105 107.370 47.245 118.260 ;
        RECT 47.665 107.370 47.805 118.260 ;
        RECT 48.225 107.370 48.365 118.260 ;
        RECT 48.785 107.370 48.925 118.260 ;
        RECT 49.345 107.370 49.485 118.260 ;
        RECT 49.905 107.370 50.045 118.260 ;
        RECT 50.465 107.370 50.605 118.260 ;
        RECT 51.025 107.370 51.165 118.260 ;
        RECT 51.585 107.370 51.725 118.260 ;
        RECT 52.145 107.370 52.285 118.260 ;
        RECT 52.705 107.370 52.845 118.260 ;
        RECT 53.265 107.370 53.405 118.260 ;
        RECT 53.825 107.370 53.965 118.260 ;
        RECT 54.385 107.370 54.525 118.260 ;
        RECT 54.945 107.370 55.085 118.260 ;
        RECT 55.505 107.370 55.645 118.260 ;
        RECT 56.065 107.370 56.205 118.260 ;
        RECT 56.625 107.370 56.835 118.260 ;
        RECT 58.475 118.260 69.885 118.590 ;
        RECT 58.475 107.370 58.615 118.260 ;
        RECT 59.035 107.370 59.175 118.260 ;
        RECT 59.595 107.370 59.735 118.260 ;
        RECT 60.155 107.370 60.295 118.260 ;
        RECT 60.715 107.370 60.855 118.260 ;
        RECT 61.275 107.370 61.415 118.260 ;
        RECT 61.835 107.370 61.975 118.260 ;
        RECT 62.395 107.370 62.535 118.260 ;
        RECT 62.955 107.370 63.095 118.260 ;
        RECT 63.515 107.370 63.655 118.260 ;
        RECT 64.075 107.370 64.215 118.260 ;
        RECT 64.635 107.370 64.775 118.260 ;
        RECT 65.195 107.370 65.335 118.260 ;
        RECT 65.755 107.370 65.895 118.260 ;
        RECT 66.315 107.370 66.455 118.260 ;
        RECT 66.875 107.370 67.015 118.260 ;
        RECT 67.435 107.370 67.575 118.260 ;
        RECT 67.995 107.370 68.135 118.260 ;
        RECT 68.555 107.370 68.695 118.260 ;
        RECT 69.115 107.370 69.255 118.260 ;
        RECT 69.675 107.370 69.885 118.260 ;
        RECT 71.565 118.260 82.975 118.590 ;
        RECT 71.565 107.370 71.705 118.260 ;
        RECT 72.125 107.370 72.265 118.260 ;
        RECT 72.685 107.370 72.825 118.260 ;
        RECT 73.245 107.370 73.385 118.260 ;
        RECT 73.805 107.370 73.945 118.260 ;
        RECT 74.365 107.370 74.505 118.260 ;
        RECT 74.925 107.370 75.065 118.260 ;
        RECT 75.485 107.370 75.625 118.260 ;
        RECT 76.045 107.370 76.185 118.260 ;
        RECT 76.605 107.370 76.745 118.260 ;
        RECT 77.165 107.370 77.305 118.260 ;
        RECT 77.725 107.370 77.865 118.260 ;
        RECT 78.285 107.370 78.425 118.260 ;
        RECT 78.845 107.370 78.985 118.260 ;
        RECT 79.405 107.370 79.545 118.260 ;
        RECT 79.965 107.370 80.105 118.260 ;
        RECT 80.525 107.370 80.665 118.260 ;
        RECT 81.085 107.370 81.225 118.260 ;
        RECT 81.645 107.370 81.785 118.260 ;
        RECT 82.205 107.370 82.345 118.260 ;
        RECT 82.765 107.370 82.975 118.260 ;
        RECT 84.655 118.240 96.065 118.570 ;
        RECT 84.655 107.350 84.795 118.240 ;
        RECT 85.215 107.350 85.355 118.240 ;
        RECT 85.775 107.350 85.915 118.240 ;
        RECT 86.335 107.350 86.475 118.240 ;
        RECT 86.895 107.350 87.035 118.240 ;
        RECT 87.455 107.350 87.595 118.240 ;
        RECT 88.015 107.350 88.155 118.240 ;
        RECT 88.575 107.350 88.715 118.240 ;
        RECT 89.135 107.350 89.275 118.240 ;
        RECT 89.695 107.350 89.835 118.240 ;
        RECT 90.255 107.350 90.395 118.240 ;
        RECT 90.815 107.350 90.955 118.240 ;
        RECT 91.375 107.350 91.515 118.240 ;
        RECT 91.935 107.350 92.075 118.240 ;
        RECT 92.495 107.350 92.635 118.240 ;
        RECT 93.055 107.350 93.195 118.240 ;
        RECT 93.615 107.350 93.755 118.240 ;
        RECT 94.175 107.350 94.315 118.240 ;
        RECT 94.735 107.350 94.875 118.240 ;
        RECT 95.295 107.350 95.435 118.240 ;
        RECT 95.855 107.350 96.065 118.240 ;
        RECT 97.745 118.240 109.155 118.570 ;
        RECT 97.745 107.350 97.885 118.240 ;
        RECT 98.305 107.350 98.445 118.240 ;
        RECT 98.865 107.350 99.005 118.240 ;
        RECT 99.425 107.350 99.565 118.240 ;
        RECT 99.985 107.350 100.125 118.240 ;
        RECT 100.545 107.350 100.685 118.240 ;
        RECT 101.105 107.350 101.245 118.240 ;
        RECT 101.665 107.350 101.805 118.240 ;
        RECT 102.225 107.350 102.365 118.240 ;
        RECT 102.785 107.350 102.925 118.240 ;
        RECT 103.345 107.350 103.485 118.240 ;
        RECT 103.905 107.350 104.045 118.240 ;
        RECT 104.465 107.350 104.605 118.240 ;
        RECT 105.025 107.350 105.165 118.240 ;
        RECT 105.585 107.350 105.725 118.240 ;
        RECT 106.145 107.350 106.285 118.240 ;
        RECT 106.705 107.350 106.845 118.240 ;
        RECT 107.265 107.350 107.405 118.240 ;
        RECT 107.825 107.350 107.965 118.240 ;
        RECT 108.385 107.350 108.525 118.240 ;
        RECT 108.945 107.350 109.155 118.240 ;
        RECT 110.835 118.240 122.245 118.570 ;
        RECT 110.835 107.350 110.975 118.240 ;
        RECT 111.395 107.350 111.535 118.240 ;
        RECT 111.955 107.350 112.095 118.240 ;
        RECT 112.515 107.350 112.655 118.240 ;
        RECT 113.075 107.350 113.215 118.240 ;
        RECT 113.635 107.350 113.775 118.240 ;
        RECT 114.195 107.350 114.335 118.240 ;
        RECT 114.755 107.350 114.895 118.240 ;
        RECT 115.315 107.350 115.455 118.240 ;
        RECT 115.875 107.350 116.015 118.240 ;
        RECT 116.435 107.350 116.575 118.240 ;
        RECT 116.995 107.350 117.135 118.240 ;
        RECT 117.555 107.350 117.695 118.240 ;
        RECT 118.115 107.350 118.255 118.240 ;
        RECT 118.675 107.350 118.815 118.240 ;
        RECT 119.235 107.350 119.375 118.240 ;
        RECT 119.795 107.350 119.935 118.240 ;
        RECT 120.355 107.350 120.495 118.240 ;
        RECT 120.915 107.350 121.055 118.240 ;
        RECT 121.475 107.350 121.615 118.240 ;
        RECT 122.035 107.350 122.245 118.240 ;
        RECT 123.925 118.240 135.335 118.570 ;
        RECT 123.925 107.350 124.065 118.240 ;
        RECT 124.485 107.350 124.625 118.240 ;
        RECT 125.045 107.350 125.185 118.240 ;
        RECT 125.605 107.350 125.745 118.240 ;
        RECT 126.165 107.350 126.305 118.240 ;
        RECT 126.725 107.350 126.865 118.240 ;
        RECT 127.285 107.350 127.425 118.240 ;
        RECT 127.845 107.350 127.985 118.240 ;
        RECT 128.405 107.350 128.545 118.240 ;
        RECT 128.965 107.350 129.105 118.240 ;
        RECT 129.525 107.350 129.665 118.240 ;
        RECT 130.085 107.350 130.225 118.240 ;
        RECT 130.645 107.350 130.785 118.240 ;
        RECT 131.205 107.350 131.345 118.240 ;
        RECT 131.765 107.350 131.905 118.240 ;
        RECT 132.325 107.350 132.465 118.240 ;
        RECT 132.885 107.350 133.025 118.240 ;
        RECT 133.445 107.350 133.585 118.240 ;
        RECT 134.005 107.350 134.145 118.240 ;
        RECT 134.565 107.350 134.705 118.240 ;
        RECT 135.125 107.350 135.335 118.240 ;
        RECT 137.015 118.220 148.425 118.550 ;
        RECT 137.015 107.330 137.155 118.220 ;
        RECT 137.575 107.330 137.715 118.220 ;
        RECT 138.135 107.330 138.275 118.220 ;
        RECT 138.695 107.330 138.835 118.220 ;
        RECT 139.255 107.330 139.395 118.220 ;
        RECT 139.815 107.330 139.955 118.220 ;
        RECT 140.375 107.330 140.515 118.220 ;
        RECT 140.935 107.330 141.075 118.220 ;
        RECT 141.495 107.330 141.635 118.220 ;
        RECT 142.055 107.330 142.195 118.220 ;
        RECT 142.615 107.330 142.755 118.220 ;
        RECT 143.175 107.330 143.315 118.220 ;
        RECT 143.735 107.330 143.875 118.220 ;
        RECT 144.295 107.330 144.435 118.220 ;
        RECT 144.855 107.330 144.995 118.220 ;
        RECT 145.415 107.330 145.555 118.220 ;
        RECT 145.975 107.330 146.115 118.220 ;
        RECT 146.535 107.330 146.675 118.220 ;
        RECT 147.095 107.330 147.235 118.220 ;
        RECT 147.655 107.330 147.795 118.220 ;
        RECT 148.215 107.330 148.425 118.220 ;
        RECT 150.105 118.220 161.515 118.550 ;
        RECT 150.105 107.330 150.245 118.220 ;
        RECT 150.665 107.330 150.805 118.220 ;
        RECT 151.225 107.330 151.365 118.220 ;
        RECT 151.785 107.330 151.925 118.220 ;
        RECT 152.345 107.330 152.485 118.220 ;
        RECT 152.905 107.330 153.045 118.220 ;
        RECT 153.465 107.330 153.605 118.220 ;
        RECT 154.025 107.330 154.165 118.220 ;
        RECT 154.585 107.330 154.725 118.220 ;
        RECT 155.145 107.330 155.285 118.220 ;
        RECT 155.705 107.330 155.845 118.220 ;
        RECT 156.265 107.330 156.405 118.220 ;
        RECT 156.825 107.330 156.965 118.220 ;
        RECT 157.385 107.330 157.525 118.220 ;
        RECT 157.945 107.330 158.085 118.220 ;
        RECT 158.505 107.330 158.645 118.220 ;
        RECT 159.065 107.330 159.205 118.220 ;
        RECT 159.625 107.330 159.765 118.220 ;
        RECT 160.185 107.330 160.325 118.220 ;
        RECT 160.745 107.330 160.885 118.220 ;
        RECT 161.305 107.330 161.515 118.220 ;
        RECT 6.185 93.840 6.325 104.730 ;
        RECT 6.745 93.840 6.885 104.730 ;
        RECT 7.305 93.840 7.445 104.730 ;
        RECT 7.865 93.840 8.005 104.730 ;
        RECT 8.425 93.840 8.565 104.730 ;
        RECT 8.985 93.840 9.125 104.730 ;
        RECT 9.545 93.840 9.685 104.730 ;
        RECT 10.105 93.840 10.245 104.730 ;
        RECT 10.665 93.840 10.805 104.730 ;
        RECT 11.225 93.840 11.365 104.730 ;
        RECT 11.785 93.840 11.925 104.730 ;
        RECT 12.345 93.840 12.485 104.730 ;
        RECT 12.905 93.840 13.045 104.730 ;
        RECT 13.465 93.840 13.605 104.730 ;
        RECT 14.025 93.840 14.165 104.730 ;
        RECT 14.585 93.840 14.725 104.730 ;
        RECT 15.145 93.840 15.285 104.730 ;
        RECT 15.705 93.840 15.845 104.730 ;
        RECT 16.265 93.840 16.405 104.730 ;
        RECT 16.825 93.840 16.965 104.730 ;
        RECT 17.385 93.840 17.595 104.730 ;
        RECT 6.185 93.510 17.595 93.840 ;
        RECT 19.275 93.840 19.415 104.730 ;
        RECT 19.835 93.840 19.975 104.730 ;
        RECT 20.395 93.840 20.535 104.730 ;
        RECT 20.955 93.840 21.095 104.730 ;
        RECT 21.515 93.840 21.655 104.730 ;
        RECT 22.075 93.840 22.215 104.730 ;
        RECT 22.635 93.840 22.775 104.730 ;
        RECT 23.195 93.840 23.335 104.730 ;
        RECT 23.755 93.840 23.895 104.730 ;
        RECT 24.315 93.840 24.455 104.730 ;
        RECT 24.875 93.840 25.015 104.730 ;
        RECT 25.435 93.840 25.575 104.730 ;
        RECT 25.995 93.840 26.135 104.730 ;
        RECT 26.555 93.840 26.695 104.730 ;
        RECT 27.115 93.840 27.255 104.730 ;
        RECT 27.675 93.840 27.815 104.730 ;
        RECT 28.235 93.840 28.375 104.730 ;
        RECT 28.795 93.840 28.935 104.730 ;
        RECT 29.355 93.840 29.495 104.730 ;
        RECT 29.915 93.840 30.055 104.730 ;
        RECT 30.475 93.840 30.685 104.730 ;
        RECT 19.275 93.510 30.685 93.840 ;
        RECT 32.365 93.860 32.505 104.750 ;
        RECT 32.925 93.860 33.065 104.750 ;
        RECT 33.485 93.860 33.625 104.750 ;
        RECT 34.045 93.860 34.185 104.750 ;
        RECT 34.605 93.860 34.745 104.750 ;
        RECT 35.165 93.860 35.305 104.750 ;
        RECT 35.725 93.860 35.865 104.750 ;
        RECT 36.285 93.860 36.425 104.750 ;
        RECT 36.845 93.860 36.985 104.750 ;
        RECT 37.405 93.860 37.545 104.750 ;
        RECT 37.965 93.860 38.105 104.750 ;
        RECT 38.525 93.860 38.665 104.750 ;
        RECT 39.085 93.860 39.225 104.750 ;
        RECT 39.645 93.860 39.785 104.750 ;
        RECT 40.205 93.860 40.345 104.750 ;
        RECT 40.765 93.860 40.905 104.750 ;
        RECT 41.325 93.860 41.465 104.750 ;
        RECT 41.885 93.860 42.025 104.750 ;
        RECT 42.445 93.860 42.585 104.750 ;
        RECT 43.005 93.860 43.145 104.750 ;
        RECT 43.565 93.860 43.775 104.750 ;
        RECT 32.365 93.530 43.775 93.860 ;
        RECT 45.455 93.860 45.595 104.750 ;
        RECT 46.015 93.860 46.155 104.750 ;
        RECT 46.575 93.860 46.715 104.750 ;
        RECT 47.135 93.860 47.275 104.750 ;
        RECT 47.695 93.860 47.835 104.750 ;
        RECT 48.255 93.860 48.395 104.750 ;
        RECT 48.815 93.860 48.955 104.750 ;
        RECT 49.375 93.860 49.515 104.750 ;
        RECT 49.935 93.860 50.075 104.750 ;
        RECT 50.495 93.860 50.635 104.750 ;
        RECT 51.055 93.860 51.195 104.750 ;
        RECT 51.615 93.860 51.755 104.750 ;
        RECT 52.175 93.860 52.315 104.750 ;
        RECT 52.735 93.860 52.875 104.750 ;
        RECT 53.295 93.860 53.435 104.750 ;
        RECT 53.855 93.860 53.995 104.750 ;
        RECT 54.415 93.860 54.555 104.750 ;
        RECT 54.975 93.860 55.115 104.750 ;
        RECT 55.535 93.860 55.675 104.750 ;
        RECT 56.095 93.860 56.235 104.750 ;
        RECT 56.655 93.860 56.865 104.750 ;
        RECT 45.455 93.530 56.865 93.860 ;
        RECT 58.505 93.860 58.645 104.750 ;
        RECT 59.065 93.860 59.205 104.750 ;
        RECT 59.625 93.860 59.765 104.750 ;
        RECT 60.185 93.860 60.325 104.750 ;
        RECT 60.745 93.860 60.885 104.750 ;
        RECT 61.305 93.860 61.445 104.750 ;
        RECT 61.865 93.860 62.005 104.750 ;
        RECT 62.425 93.860 62.565 104.750 ;
        RECT 62.985 93.860 63.125 104.750 ;
        RECT 63.545 93.860 63.685 104.750 ;
        RECT 64.105 93.860 64.245 104.750 ;
        RECT 64.665 93.860 64.805 104.750 ;
        RECT 65.225 93.860 65.365 104.750 ;
        RECT 65.785 93.860 65.925 104.750 ;
        RECT 66.345 93.860 66.485 104.750 ;
        RECT 66.905 93.860 67.045 104.750 ;
        RECT 67.465 93.860 67.605 104.750 ;
        RECT 68.025 93.860 68.165 104.750 ;
        RECT 68.585 93.860 68.725 104.750 ;
        RECT 69.145 93.860 69.285 104.750 ;
        RECT 69.705 93.860 69.915 104.750 ;
        RECT 58.505 93.530 69.915 93.860 ;
        RECT 71.595 93.860 71.735 104.750 ;
        RECT 72.155 93.860 72.295 104.750 ;
        RECT 72.715 93.860 72.855 104.750 ;
        RECT 73.275 93.860 73.415 104.750 ;
        RECT 73.835 93.860 73.975 104.750 ;
        RECT 74.395 93.860 74.535 104.750 ;
        RECT 74.955 93.860 75.095 104.750 ;
        RECT 75.515 93.860 75.655 104.750 ;
        RECT 76.075 93.860 76.215 104.750 ;
        RECT 76.635 93.860 76.775 104.750 ;
        RECT 77.195 93.860 77.335 104.750 ;
        RECT 77.755 93.860 77.895 104.750 ;
        RECT 78.315 93.860 78.455 104.750 ;
        RECT 78.875 93.860 79.015 104.750 ;
        RECT 79.435 93.860 79.575 104.750 ;
        RECT 79.995 93.860 80.135 104.750 ;
        RECT 80.555 93.860 80.695 104.750 ;
        RECT 81.115 93.860 81.255 104.750 ;
        RECT 81.675 93.860 81.815 104.750 ;
        RECT 82.235 93.860 82.375 104.750 ;
        RECT 82.795 93.860 83.005 104.750 ;
        RECT 71.595 93.530 83.005 93.860 ;
        RECT 84.685 93.880 84.825 104.770 ;
        RECT 85.245 93.880 85.385 104.770 ;
        RECT 85.805 93.880 85.945 104.770 ;
        RECT 86.365 93.880 86.505 104.770 ;
        RECT 86.925 93.880 87.065 104.770 ;
        RECT 87.485 93.880 87.625 104.770 ;
        RECT 88.045 93.880 88.185 104.770 ;
        RECT 88.605 93.880 88.745 104.770 ;
        RECT 89.165 93.880 89.305 104.770 ;
        RECT 89.725 93.880 89.865 104.770 ;
        RECT 90.285 93.880 90.425 104.770 ;
        RECT 90.845 93.880 90.985 104.770 ;
        RECT 91.405 93.880 91.545 104.770 ;
        RECT 91.965 93.880 92.105 104.770 ;
        RECT 92.525 93.880 92.665 104.770 ;
        RECT 93.085 93.880 93.225 104.770 ;
        RECT 93.645 93.880 93.785 104.770 ;
        RECT 94.205 93.880 94.345 104.770 ;
        RECT 94.765 93.880 94.905 104.770 ;
        RECT 95.325 93.880 95.465 104.770 ;
        RECT 95.885 93.880 96.095 104.770 ;
        RECT 84.685 93.550 96.095 93.880 ;
        RECT 97.775 93.880 97.915 104.770 ;
        RECT 98.335 93.880 98.475 104.770 ;
        RECT 98.895 93.880 99.035 104.770 ;
        RECT 99.455 93.880 99.595 104.770 ;
        RECT 100.015 93.880 100.155 104.770 ;
        RECT 100.575 93.880 100.715 104.770 ;
        RECT 101.135 93.880 101.275 104.770 ;
        RECT 101.695 93.880 101.835 104.770 ;
        RECT 102.255 93.880 102.395 104.770 ;
        RECT 102.815 93.880 102.955 104.770 ;
        RECT 103.375 93.880 103.515 104.770 ;
        RECT 103.935 93.880 104.075 104.770 ;
        RECT 104.495 93.880 104.635 104.770 ;
        RECT 105.055 93.880 105.195 104.770 ;
        RECT 105.615 93.880 105.755 104.770 ;
        RECT 106.175 93.880 106.315 104.770 ;
        RECT 106.735 93.880 106.875 104.770 ;
        RECT 107.295 93.880 107.435 104.770 ;
        RECT 107.855 93.880 107.995 104.770 ;
        RECT 108.415 93.880 108.555 104.770 ;
        RECT 108.975 93.880 109.185 104.770 ;
        RECT 97.775 93.550 109.185 93.880 ;
        RECT 110.865 93.880 111.005 104.770 ;
        RECT 111.425 93.880 111.565 104.770 ;
        RECT 111.985 93.880 112.125 104.770 ;
        RECT 112.545 93.880 112.685 104.770 ;
        RECT 113.105 93.880 113.245 104.770 ;
        RECT 113.665 93.880 113.805 104.770 ;
        RECT 114.225 93.880 114.365 104.770 ;
        RECT 114.785 93.880 114.925 104.770 ;
        RECT 115.345 93.880 115.485 104.770 ;
        RECT 115.905 93.880 116.045 104.770 ;
        RECT 116.465 93.880 116.605 104.770 ;
        RECT 117.025 93.880 117.165 104.770 ;
        RECT 117.585 93.880 117.725 104.770 ;
        RECT 118.145 93.880 118.285 104.770 ;
        RECT 118.705 93.880 118.845 104.770 ;
        RECT 119.265 93.880 119.405 104.770 ;
        RECT 119.825 93.880 119.965 104.770 ;
        RECT 120.385 93.880 120.525 104.770 ;
        RECT 120.945 93.880 121.085 104.770 ;
        RECT 121.505 93.880 121.645 104.770 ;
        RECT 122.065 93.880 122.275 104.770 ;
        RECT 110.865 93.550 122.275 93.880 ;
        RECT 123.955 93.880 124.095 104.770 ;
        RECT 124.515 93.880 124.655 104.770 ;
        RECT 125.075 93.880 125.215 104.770 ;
        RECT 125.635 93.880 125.775 104.770 ;
        RECT 126.195 93.880 126.335 104.770 ;
        RECT 126.755 93.880 126.895 104.770 ;
        RECT 127.315 93.880 127.455 104.770 ;
        RECT 127.875 93.880 128.015 104.770 ;
        RECT 128.435 93.880 128.575 104.770 ;
        RECT 128.995 93.880 129.135 104.770 ;
        RECT 129.555 93.880 129.695 104.770 ;
        RECT 130.115 93.880 130.255 104.770 ;
        RECT 130.675 93.880 130.815 104.770 ;
        RECT 131.235 93.880 131.375 104.770 ;
        RECT 131.795 93.880 131.935 104.770 ;
        RECT 132.355 93.880 132.495 104.770 ;
        RECT 132.915 93.880 133.055 104.770 ;
        RECT 133.475 93.880 133.615 104.770 ;
        RECT 134.035 93.880 134.175 104.770 ;
        RECT 134.595 93.880 134.735 104.770 ;
        RECT 135.155 93.880 135.365 104.770 ;
        RECT 123.955 93.550 135.365 93.880 ;
        RECT 137.045 93.900 137.185 104.790 ;
        RECT 137.605 93.900 137.745 104.790 ;
        RECT 138.165 93.900 138.305 104.790 ;
        RECT 138.725 93.900 138.865 104.790 ;
        RECT 139.285 93.900 139.425 104.790 ;
        RECT 139.845 93.900 139.985 104.790 ;
        RECT 140.405 93.900 140.545 104.790 ;
        RECT 140.965 93.900 141.105 104.790 ;
        RECT 141.525 93.900 141.665 104.790 ;
        RECT 142.085 93.900 142.225 104.790 ;
        RECT 142.645 93.900 142.785 104.790 ;
        RECT 143.205 93.900 143.345 104.790 ;
        RECT 143.765 93.900 143.905 104.790 ;
        RECT 144.325 93.900 144.465 104.790 ;
        RECT 144.885 93.900 145.025 104.790 ;
        RECT 145.445 93.900 145.585 104.790 ;
        RECT 146.005 93.900 146.145 104.790 ;
        RECT 146.565 93.900 146.705 104.790 ;
        RECT 147.125 93.900 147.265 104.790 ;
        RECT 147.685 93.900 147.825 104.790 ;
        RECT 148.245 93.900 148.455 104.790 ;
        RECT 137.045 93.570 148.455 93.900 ;
        RECT 150.135 93.900 150.275 104.790 ;
        RECT 150.695 93.900 150.835 104.790 ;
        RECT 151.255 93.900 151.395 104.790 ;
        RECT 151.815 93.900 151.955 104.790 ;
        RECT 152.375 93.900 152.515 104.790 ;
        RECT 152.935 93.900 153.075 104.790 ;
        RECT 153.495 93.900 153.635 104.790 ;
        RECT 154.055 93.900 154.195 104.790 ;
        RECT 154.615 93.900 154.755 104.790 ;
        RECT 155.175 93.900 155.315 104.790 ;
        RECT 155.735 93.900 155.875 104.790 ;
        RECT 156.295 93.900 156.435 104.790 ;
        RECT 156.855 93.900 156.995 104.790 ;
        RECT 157.415 93.900 157.555 104.790 ;
        RECT 157.975 93.900 158.115 104.790 ;
        RECT 158.535 93.900 158.675 104.790 ;
        RECT 159.095 93.900 159.235 104.790 ;
        RECT 159.655 93.900 159.795 104.790 ;
        RECT 160.215 93.900 160.355 104.790 ;
        RECT 160.775 93.900 160.915 104.790 ;
        RECT 161.335 93.900 161.545 104.790 ;
        RECT 150.135 93.570 161.545 93.900 ;
        RECT 150.190 89.465 167.830 89.940 ;
        RECT 1.980 79.280 2.450 88.845 ;
        RECT 148.780 88.200 149.040 88.520 ;
        RECT 1.980 79.270 10.815 79.280 ;
        RECT 1.980 78.810 50.125 79.270 ;
        RECT 9.825 78.790 50.125 78.810 ;
        RECT 18.600 74.390 18.890 74.420 ;
        RECT 19.115 74.390 19.285 78.790 ;
        RECT 18.600 74.220 19.285 74.390 ;
        RECT 28.215 74.390 28.505 74.420 ;
        RECT 28.730 74.390 28.900 78.790 ;
        RECT 28.215 74.220 28.900 74.390 ;
        RECT 37.830 74.390 38.120 74.420 ;
        RECT 38.345 74.390 38.515 78.790 ;
        RECT 37.830 74.220 38.515 74.390 ;
        RECT 47.445 74.390 47.735 74.420 ;
        RECT 47.960 74.390 48.130 78.790 ;
        RECT 150.190 75.305 150.670 89.465 ;
        RECT 47.445 74.220 48.130 74.390 ;
        RECT 18.600 74.190 18.890 74.220 ;
        RECT 28.215 74.190 28.505 74.220 ;
        RECT 37.830 74.190 38.120 74.220 ;
        RECT 47.445 74.190 47.735 74.220 ;
        RECT 178.080 65.535 178.380 65.770 ;
        RECT 176.340 65.305 178.380 65.535 ;
        RECT 178.080 62.395 178.380 65.305 ;
        RECT 176.340 62.165 178.380 62.395 ;
        RECT 178.080 61.930 178.380 62.165 ;
        RECT 161.090 60.645 161.740 60.875 ;
        RECT 162.595 60.645 163.245 60.875 ;
        RECT 164.420 60.645 165.070 60.875 ;
        RECT 161.090 59.440 161.740 59.670 ;
        RECT 162.595 59.440 163.245 59.670 ;
        RECT 164.420 59.440 165.070 59.670 ;
        RECT 178.080 59.345 178.380 59.715 ;
        RECT 176.340 59.115 178.380 59.345 ;
        RECT 178.080 56.205 178.380 59.115 ;
        RECT 176.340 55.975 178.380 56.205 ;
        RECT 178.080 55.740 178.380 55.975 ;
        RECT 18.600 45.630 18.890 45.660 ;
        RECT 28.215 45.630 28.505 45.660 ;
        RECT 37.830 45.630 38.120 45.660 ;
        RECT 47.445 45.630 47.735 45.660 ;
        RECT 18.600 45.460 19.285 45.630 ;
        RECT 18.600 45.430 18.890 45.460 ;
        RECT 19.115 41.060 19.285 45.460 ;
        RECT 28.215 45.460 28.900 45.630 ;
        RECT 28.215 45.430 28.505 45.460 ;
        RECT 28.730 41.060 28.900 45.460 ;
        RECT 37.830 45.460 38.515 45.630 ;
        RECT 37.830 45.430 38.120 45.460 ;
        RECT 38.345 41.060 38.515 45.460 ;
        RECT 47.445 45.460 48.130 45.630 ;
        RECT 47.445 45.430 47.735 45.460 ;
        RECT 47.960 41.060 48.130 45.460 ;
        RECT 9.825 41.040 50.125 41.060 ;
        RECT 1.940 40.580 50.125 41.040 ;
        RECT 1.940 40.570 10.815 40.580 ;
        RECT 1.940 33.185 2.410 40.570 ;
        RECT 150.190 30.385 150.670 44.545 ;
        RECT 166.065 30.385 166.540 30.415 ;
        RECT 150.190 29.910 166.540 30.385 ;
        RECT 166.065 29.880 166.540 29.910 ;
        RECT 6.595 26.640 18.005 26.970 ;
        RECT 6.595 15.750 6.735 26.640 ;
        RECT 7.155 15.750 7.295 26.640 ;
        RECT 7.715 15.750 7.855 26.640 ;
        RECT 8.275 15.750 8.415 26.640 ;
        RECT 8.835 15.750 8.975 26.640 ;
        RECT 9.395 15.750 9.535 26.640 ;
        RECT 9.955 15.750 10.095 26.640 ;
        RECT 10.515 15.750 10.655 26.640 ;
        RECT 11.075 15.750 11.215 26.640 ;
        RECT 11.635 15.750 11.775 26.640 ;
        RECT 12.195 15.750 12.335 26.640 ;
        RECT 12.755 15.750 12.895 26.640 ;
        RECT 13.315 15.750 13.455 26.640 ;
        RECT 13.875 15.750 14.015 26.640 ;
        RECT 14.435 15.750 14.575 26.640 ;
        RECT 14.995 15.750 15.135 26.640 ;
        RECT 15.555 15.750 15.695 26.640 ;
        RECT 16.115 15.750 16.255 26.640 ;
        RECT 16.675 15.750 16.815 26.640 ;
        RECT 17.235 15.750 17.375 26.640 ;
        RECT 17.795 15.750 18.005 26.640 ;
        RECT 19.685 26.640 31.095 26.970 ;
        RECT 19.685 15.750 19.825 26.640 ;
        RECT 20.245 15.750 20.385 26.640 ;
        RECT 20.805 15.750 20.945 26.640 ;
        RECT 21.365 15.750 21.505 26.640 ;
        RECT 21.925 15.750 22.065 26.640 ;
        RECT 22.485 15.750 22.625 26.640 ;
        RECT 23.045 15.750 23.185 26.640 ;
        RECT 23.605 15.750 23.745 26.640 ;
        RECT 24.165 15.750 24.305 26.640 ;
        RECT 24.725 15.750 24.865 26.640 ;
        RECT 25.285 15.750 25.425 26.640 ;
        RECT 25.845 15.750 25.985 26.640 ;
        RECT 26.405 15.750 26.545 26.640 ;
        RECT 26.965 15.750 27.105 26.640 ;
        RECT 27.525 15.750 27.665 26.640 ;
        RECT 28.085 15.750 28.225 26.640 ;
        RECT 28.645 15.750 28.785 26.640 ;
        RECT 29.205 15.750 29.345 26.640 ;
        RECT 29.765 15.750 29.905 26.640 ;
        RECT 30.325 15.750 30.465 26.640 ;
        RECT 30.885 15.750 31.095 26.640 ;
        RECT 32.775 26.620 44.185 26.950 ;
        RECT 32.775 15.730 32.915 26.620 ;
        RECT 33.335 15.730 33.475 26.620 ;
        RECT 33.895 15.730 34.035 26.620 ;
        RECT 34.455 15.730 34.595 26.620 ;
        RECT 35.015 15.730 35.155 26.620 ;
        RECT 35.575 15.730 35.715 26.620 ;
        RECT 36.135 15.730 36.275 26.620 ;
        RECT 36.695 15.730 36.835 26.620 ;
        RECT 37.255 15.730 37.395 26.620 ;
        RECT 37.815 15.730 37.955 26.620 ;
        RECT 38.375 15.730 38.515 26.620 ;
        RECT 38.935 15.730 39.075 26.620 ;
        RECT 39.495 15.730 39.635 26.620 ;
        RECT 40.055 15.730 40.195 26.620 ;
        RECT 40.615 15.730 40.755 26.620 ;
        RECT 41.175 15.730 41.315 26.620 ;
        RECT 41.735 15.730 41.875 26.620 ;
        RECT 42.295 15.730 42.435 26.620 ;
        RECT 42.855 15.730 42.995 26.620 ;
        RECT 43.415 15.730 43.555 26.620 ;
        RECT 43.975 15.730 44.185 26.620 ;
        RECT 45.865 26.620 57.275 26.950 ;
        RECT 45.865 15.730 46.005 26.620 ;
        RECT 46.425 15.730 46.565 26.620 ;
        RECT 46.985 15.730 47.125 26.620 ;
        RECT 47.545 15.730 47.685 26.620 ;
        RECT 48.105 15.730 48.245 26.620 ;
        RECT 48.665 15.730 48.805 26.620 ;
        RECT 49.225 15.730 49.365 26.620 ;
        RECT 49.785 15.730 49.925 26.620 ;
        RECT 50.345 15.730 50.485 26.620 ;
        RECT 50.905 15.730 51.045 26.620 ;
        RECT 51.465 15.730 51.605 26.620 ;
        RECT 52.025 15.730 52.165 26.620 ;
        RECT 52.585 15.730 52.725 26.620 ;
        RECT 53.145 15.730 53.285 26.620 ;
        RECT 53.705 15.730 53.845 26.620 ;
        RECT 54.265 15.730 54.405 26.620 ;
        RECT 54.825 15.730 54.965 26.620 ;
        RECT 55.385 15.730 55.525 26.620 ;
        RECT 55.945 15.730 56.085 26.620 ;
        RECT 56.505 15.730 56.645 26.620 ;
        RECT 57.065 15.730 57.275 26.620 ;
        RECT 58.915 26.620 70.325 26.950 ;
        RECT 58.915 15.730 59.055 26.620 ;
        RECT 59.475 15.730 59.615 26.620 ;
        RECT 60.035 15.730 60.175 26.620 ;
        RECT 60.595 15.730 60.735 26.620 ;
        RECT 61.155 15.730 61.295 26.620 ;
        RECT 61.715 15.730 61.855 26.620 ;
        RECT 62.275 15.730 62.415 26.620 ;
        RECT 62.835 15.730 62.975 26.620 ;
        RECT 63.395 15.730 63.535 26.620 ;
        RECT 63.955 15.730 64.095 26.620 ;
        RECT 64.515 15.730 64.655 26.620 ;
        RECT 65.075 15.730 65.215 26.620 ;
        RECT 65.635 15.730 65.775 26.620 ;
        RECT 66.195 15.730 66.335 26.620 ;
        RECT 66.755 15.730 66.895 26.620 ;
        RECT 67.315 15.730 67.455 26.620 ;
        RECT 67.875 15.730 68.015 26.620 ;
        RECT 68.435 15.730 68.575 26.620 ;
        RECT 68.995 15.730 69.135 26.620 ;
        RECT 69.555 15.730 69.695 26.620 ;
        RECT 70.115 15.730 70.325 26.620 ;
        RECT 72.005 26.620 83.415 26.950 ;
        RECT 72.005 15.730 72.145 26.620 ;
        RECT 72.565 15.730 72.705 26.620 ;
        RECT 73.125 15.730 73.265 26.620 ;
        RECT 73.685 15.730 73.825 26.620 ;
        RECT 74.245 15.730 74.385 26.620 ;
        RECT 74.805 15.730 74.945 26.620 ;
        RECT 75.365 15.730 75.505 26.620 ;
        RECT 75.925 15.730 76.065 26.620 ;
        RECT 76.485 15.730 76.625 26.620 ;
        RECT 77.045 15.730 77.185 26.620 ;
        RECT 77.605 15.730 77.745 26.620 ;
        RECT 78.165 15.730 78.305 26.620 ;
        RECT 78.725 15.730 78.865 26.620 ;
        RECT 79.285 15.730 79.425 26.620 ;
        RECT 79.845 15.730 79.985 26.620 ;
        RECT 80.405 15.730 80.545 26.620 ;
        RECT 80.965 15.730 81.105 26.620 ;
        RECT 81.525 15.730 81.665 26.620 ;
        RECT 82.085 15.730 82.225 26.620 ;
        RECT 82.645 15.730 82.785 26.620 ;
        RECT 83.205 15.730 83.415 26.620 ;
        RECT 85.095 26.600 96.505 26.930 ;
        RECT 85.095 15.710 85.235 26.600 ;
        RECT 85.655 15.710 85.795 26.600 ;
        RECT 86.215 15.710 86.355 26.600 ;
        RECT 86.775 15.710 86.915 26.600 ;
        RECT 87.335 15.710 87.475 26.600 ;
        RECT 87.895 15.710 88.035 26.600 ;
        RECT 88.455 15.710 88.595 26.600 ;
        RECT 89.015 15.710 89.155 26.600 ;
        RECT 89.575 15.710 89.715 26.600 ;
        RECT 90.135 15.710 90.275 26.600 ;
        RECT 90.695 15.710 90.835 26.600 ;
        RECT 91.255 15.710 91.395 26.600 ;
        RECT 91.815 15.710 91.955 26.600 ;
        RECT 92.375 15.710 92.515 26.600 ;
        RECT 92.935 15.710 93.075 26.600 ;
        RECT 93.495 15.710 93.635 26.600 ;
        RECT 94.055 15.710 94.195 26.600 ;
        RECT 94.615 15.710 94.755 26.600 ;
        RECT 95.175 15.710 95.315 26.600 ;
        RECT 95.735 15.710 95.875 26.600 ;
        RECT 96.295 15.710 96.505 26.600 ;
        RECT 98.185 26.600 109.595 26.930 ;
        RECT 98.185 15.710 98.325 26.600 ;
        RECT 98.745 15.710 98.885 26.600 ;
        RECT 99.305 15.710 99.445 26.600 ;
        RECT 99.865 15.710 100.005 26.600 ;
        RECT 100.425 15.710 100.565 26.600 ;
        RECT 100.985 15.710 101.125 26.600 ;
        RECT 101.545 15.710 101.685 26.600 ;
        RECT 102.105 15.710 102.245 26.600 ;
        RECT 102.665 15.710 102.805 26.600 ;
        RECT 103.225 15.710 103.365 26.600 ;
        RECT 103.785 15.710 103.925 26.600 ;
        RECT 104.345 15.710 104.485 26.600 ;
        RECT 104.905 15.710 105.045 26.600 ;
        RECT 105.465 15.710 105.605 26.600 ;
        RECT 106.025 15.710 106.165 26.600 ;
        RECT 106.585 15.710 106.725 26.600 ;
        RECT 107.145 15.710 107.285 26.600 ;
        RECT 107.705 15.710 107.845 26.600 ;
        RECT 108.265 15.710 108.405 26.600 ;
        RECT 108.825 15.710 108.965 26.600 ;
        RECT 109.385 15.710 109.595 26.600 ;
        RECT 111.275 26.600 122.685 26.930 ;
        RECT 111.275 15.710 111.415 26.600 ;
        RECT 111.835 15.710 111.975 26.600 ;
        RECT 112.395 15.710 112.535 26.600 ;
        RECT 112.955 15.710 113.095 26.600 ;
        RECT 113.515 15.710 113.655 26.600 ;
        RECT 114.075 15.710 114.215 26.600 ;
        RECT 114.635 15.710 114.775 26.600 ;
        RECT 115.195 15.710 115.335 26.600 ;
        RECT 115.755 15.710 115.895 26.600 ;
        RECT 116.315 15.710 116.455 26.600 ;
        RECT 116.875 15.710 117.015 26.600 ;
        RECT 117.435 15.710 117.575 26.600 ;
        RECT 117.995 15.710 118.135 26.600 ;
        RECT 118.555 15.710 118.695 26.600 ;
        RECT 119.115 15.710 119.255 26.600 ;
        RECT 119.675 15.710 119.815 26.600 ;
        RECT 120.235 15.710 120.375 26.600 ;
        RECT 120.795 15.710 120.935 26.600 ;
        RECT 121.355 15.710 121.495 26.600 ;
        RECT 121.915 15.710 122.055 26.600 ;
        RECT 122.475 15.710 122.685 26.600 ;
        RECT 124.365 26.600 135.775 26.930 ;
        RECT 124.365 15.710 124.505 26.600 ;
        RECT 124.925 15.710 125.065 26.600 ;
        RECT 125.485 15.710 125.625 26.600 ;
        RECT 126.045 15.710 126.185 26.600 ;
        RECT 126.605 15.710 126.745 26.600 ;
        RECT 127.165 15.710 127.305 26.600 ;
        RECT 127.725 15.710 127.865 26.600 ;
        RECT 128.285 15.710 128.425 26.600 ;
        RECT 128.845 15.710 128.985 26.600 ;
        RECT 129.405 15.710 129.545 26.600 ;
        RECT 129.965 15.710 130.105 26.600 ;
        RECT 130.525 15.710 130.665 26.600 ;
        RECT 131.085 15.710 131.225 26.600 ;
        RECT 131.645 15.710 131.785 26.600 ;
        RECT 132.205 15.710 132.345 26.600 ;
        RECT 132.765 15.710 132.905 26.600 ;
        RECT 133.325 15.710 133.465 26.600 ;
        RECT 133.885 15.710 134.025 26.600 ;
        RECT 134.445 15.710 134.585 26.600 ;
        RECT 135.005 15.710 135.145 26.600 ;
        RECT 135.565 15.710 135.775 26.600 ;
        RECT 137.455 26.580 148.865 26.910 ;
        RECT 137.455 15.690 137.595 26.580 ;
        RECT 138.015 15.690 138.155 26.580 ;
        RECT 138.575 15.690 138.715 26.580 ;
        RECT 139.135 15.690 139.275 26.580 ;
        RECT 139.695 15.690 139.835 26.580 ;
        RECT 140.255 15.690 140.395 26.580 ;
        RECT 140.815 15.690 140.955 26.580 ;
        RECT 141.375 15.690 141.515 26.580 ;
        RECT 141.935 15.690 142.075 26.580 ;
        RECT 142.495 15.690 142.635 26.580 ;
        RECT 143.055 15.690 143.195 26.580 ;
        RECT 143.615 15.690 143.755 26.580 ;
        RECT 144.175 15.690 144.315 26.580 ;
        RECT 144.735 15.690 144.875 26.580 ;
        RECT 145.295 15.690 145.435 26.580 ;
        RECT 145.855 15.690 145.995 26.580 ;
        RECT 146.415 15.690 146.555 26.580 ;
        RECT 146.975 15.690 147.115 26.580 ;
        RECT 147.535 15.690 147.675 26.580 ;
        RECT 148.095 15.690 148.235 26.580 ;
        RECT 148.655 15.690 148.865 26.580 ;
        RECT 150.545 26.580 161.955 26.910 ;
        RECT 150.545 15.690 150.685 26.580 ;
        RECT 151.105 15.690 151.245 26.580 ;
        RECT 151.665 15.690 151.805 26.580 ;
        RECT 152.225 15.690 152.365 26.580 ;
        RECT 152.785 15.690 152.925 26.580 ;
        RECT 153.345 15.690 153.485 26.580 ;
        RECT 153.905 15.690 154.045 26.580 ;
        RECT 154.465 15.690 154.605 26.580 ;
        RECT 155.025 15.690 155.165 26.580 ;
        RECT 155.585 15.690 155.725 26.580 ;
        RECT 156.145 15.690 156.285 26.580 ;
        RECT 156.705 15.690 156.845 26.580 ;
        RECT 157.265 15.690 157.405 26.580 ;
        RECT 157.825 15.690 157.965 26.580 ;
        RECT 158.385 15.690 158.525 26.580 ;
        RECT 158.945 15.690 159.085 26.580 ;
        RECT 159.505 15.690 159.645 26.580 ;
        RECT 160.065 15.690 160.205 26.580 ;
        RECT 160.625 15.690 160.765 26.580 ;
        RECT 161.185 15.690 161.325 26.580 ;
        RECT 161.745 15.690 161.955 26.580 ;
        RECT 6.625 2.200 6.765 13.090 ;
        RECT 7.185 2.200 7.325 13.090 ;
        RECT 7.745 2.200 7.885 13.090 ;
        RECT 8.305 2.200 8.445 13.090 ;
        RECT 8.865 2.200 9.005 13.090 ;
        RECT 9.425 2.200 9.565 13.090 ;
        RECT 9.985 2.200 10.125 13.090 ;
        RECT 10.545 2.200 10.685 13.090 ;
        RECT 11.105 2.200 11.245 13.090 ;
        RECT 11.665 2.200 11.805 13.090 ;
        RECT 12.225 2.200 12.365 13.090 ;
        RECT 12.785 2.200 12.925 13.090 ;
        RECT 13.345 2.200 13.485 13.090 ;
        RECT 13.905 2.200 14.045 13.090 ;
        RECT 14.465 2.200 14.605 13.090 ;
        RECT 15.025 2.200 15.165 13.090 ;
        RECT 15.585 2.200 15.725 13.090 ;
        RECT 16.145 2.200 16.285 13.090 ;
        RECT 16.705 2.200 16.845 13.090 ;
        RECT 17.265 2.200 17.405 13.090 ;
        RECT 17.825 2.200 18.035 13.090 ;
        RECT 6.625 1.870 18.035 2.200 ;
        RECT 19.715 2.200 19.855 13.090 ;
        RECT 20.275 2.200 20.415 13.090 ;
        RECT 20.835 2.200 20.975 13.090 ;
        RECT 21.395 2.200 21.535 13.090 ;
        RECT 21.955 2.200 22.095 13.090 ;
        RECT 22.515 2.200 22.655 13.090 ;
        RECT 23.075 2.200 23.215 13.090 ;
        RECT 23.635 2.200 23.775 13.090 ;
        RECT 24.195 2.200 24.335 13.090 ;
        RECT 24.755 2.200 24.895 13.090 ;
        RECT 25.315 2.200 25.455 13.090 ;
        RECT 25.875 2.200 26.015 13.090 ;
        RECT 26.435 2.200 26.575 13.090 ;
        RECT 26.995 2.200 27.135 13.090 ;
        RECT 27.555 2.200 27.695 13.090 ;
        RECT 28.115 2.200 28.255 13.090 ;
        RECT 28.675 2.200 28.815 13.090 ;
        RECT 29.235 2.200 29.375 13.090 ;
        RECT 29.795 2.200 29.935 13.090 ;
        RECT 30.355 2.200 30.495 13.090 ;
        RECT 30.915 2.200 31.125 13.090 ;
        RECT 19.715 1.870 31.125 2.200 ;
        RECT 32.805 2.220 32.945 13.110 ;
        RECT 33.365 2.220 33.505 13.110 ;
        RECT 33.925 2.220 34.065 13.110 ;
        RECT 34.485 2.220 34.625 13.110 ;
        RECT 35.045 2.220 35.185 13.110 ;
        RECT 35.605 2.220 35.745 13.110 ;
        RECT 36.165 2.220 36.305 13.110 ;
        RECT 36.725 2.220 36.865 13.110 ;
        RECT 37.285 2.220 37.425 13.110 ;
        RECT 37.845 2.220 37.985 13.110 ;
        RECT 38.405 2.220 38.545 13.110 ;
        RECT 38.965 2.220 39.105 13.110 ;
        RECT 39.525 2.220 39.665 13.110 ;
        RECT 40.085 2.220 40.225 13.110 ;
        RECT 40.645 2.220 40.785 13.110 ;
        RECT 41.205 2.220 41.345 13.110 ;
        RECT 41.765 2.220 41.905 13.110 ;
        RECT 42.325 2.220 42.465 13.110 ;
        RECT 42.885 2.220 43.025 13.110 ;
        RECT 43.445 2.220 43.585 13.110 ;
        RECT 44.005 2.220 44.215 13.110 ;
        RECT 32.805 1.890 44.215 2.220 ;
        RECT 45.895 2.220 46.035 13.110 ;
        RECT 46.455 2.220 46.595 13.110 ;
        RECT 47.015 2.220 47.155 13.110 ;
        RECT 47.575 2.220 47.715 13.110 ;
        RECT 48.135 2.220 48.275 13.110 ;
        RECT 48.695 2.220 48.835 13.110 ;
        RECT 49.255 2.220 49.395 13.110 ;
        RECT 49.815 2.220 49.955 13.110 ;
        RECT 50.375 2.220 50.515 13.110 ;
        RECT 50.935 2.220 51.075 13.110 ;
        RECT 51.495 2.220 51.635 13.110 ;
        RECT 52.055 2.220 52.195 13.110 ;
        RECT 52.615 2.220 52.755 13.110 ;
        RECT 53.175 2.220 53.315 13.110 ;
        RECT 53.735 2.220 53.875 13.110 ;
        RECT 54.295 2.220 54.435 13.110 ;
        RECT 54.855 2.220 54.995 13.110 ;
        RECT 55.415 2.220 55.555 13.110 ;
        RECT 55.975 2.220 56.115 13.110 ;
        RECT 56.535 2.220 56.675 13.110 ;
        RECT 57.095 2.220 57.305 13.110 ;
        RECT 45.895 1.890 57.305 2.220 ;
        RECT 58.945 2.220 59.085 13.110 ;
        RECT 59.505 2.220 59.645 13.110 ;
        RECT 60.065 2.220 60.205 13.110 ;
        RECT 60.625 2.220 60.765 13.110 ;
        RECT 61.185 2.220 61.325 13.110 ;
        RECT 61.745 2.220 61.885 13.110 ;
        RECT 62.305 2.220 62.445 13.110 ;
        RECT 62.865 2.220 63.005 13.110 ;
        RECT 63.425 2.220 63.565 13.110 ;
        RECT 63.985 2.220 64.125 13.110 ;
        RECT 64.545 2.220 64.685 13.110 ;
        RECT 65.105 2.220 65.245 13.110 ;
        RECT 65.665 2.220 65.805 13.110 ;
        RECT 66.225 2.220 66.365 13.110 ;
        RECT 66.785 2.220 66.925 13.110 ;
        RECT 67.345 2.220 67.485 13.110 ;
        RECT 67.905 2.220 68.045 13.110 ;
        RECT 68.465 2.220 68.605 13.110 ;
        RECT 69.025 2.220 69.165 13.110 ;
        RECT 69.585 2.220 69.725 13.110 ;
        RECT 70.145 2.220 70.355 13.110 ;
        RECT 58.945 1.890 70.355 2.220 ;
        RECT 72.035 2.220 72.175 13.110 ;
        RECT 72.595 2.220 72.735 13.110 ;
        RECT 73.155 2.220 73.295 13.110 ;
        RECT 73.715 2.220 73.855 13.110 ;
        RECT 74.275 2.220 74.415 13.110 ;
        RECT 74.835 2.220 74.975 13.110 ;
        RECT 75.395 2.220 75.535 13.110 ;
        RECT 75.955 2.220 76.095 13.110 ;
        RECT 76.515 2.220 76.655 13.110 ;
        RECT 77.075 2.220 77.215 13.110 ;
        RECT 77.635 2.220 77.775 13.110 ;
        RECT 78.195 2.220 78.335 13.110 ;
        RECT 78.755 2.220 78.895 13.110 ;
        RECT 79.315 2.220 79.455 13.110 ;
        RECT 79.875 2.220 80.015 13.110 ;
        RECT 80.435 2.220 80.575 13.110 ;
        RECT 80.995 2.220 81.135 13.110 ;
        RECT 81.555 2.220 81.695 13.110 ;
        RECT 82.115 2.220 82.255 13.110 ;
        RECT 82.675 2.220 82.815 13.110 ;
        RECT 83.235 2.220 83.445 13.110 ;
        RECT 72.035 1.890 83.445 2.220 ;
        RECT 85.125 2.240 85.265 13.130 ;
        RECT 85.685 2.240 85.825 13.130 ;
        RECT 86.245 2.240 86.385 13.130 ;
        RECT 86.805 2.240 86.945 13.130 ;
        RECT 87.365 2.240 87.505 13.130 ;
        RECT 87.925 2.240 88.065 13.130 ;
        RECT 88.485 2.240 88.625 13.130 ;
        RECT 89.045 2.240 89.185 13.130 ;
        RECT 89.605 2.240 89.745 13.130 ;
        RECT 90.165 2.240 90.305 13.130 ;
        RECT 90.725 2.240 90.865 13.130 ;
        RECT 91.285 2.240 91.425 13.130 ;
        RECT 91.845 2.240 91.985 13.130 ;
        RECT 92.405 2.240 92.545 13.130 ;
        RECT 92.965 2.240 93.105 13.130 ;
        RECT 93.525 2.240 93.665 13.130 ;
        RECT 94.085 2.240 94.225 13.130 ;
        RECT 94.645 2.240 94.785 13.130 ;
        RECT 95.205 2.240 95.345 13.130 ;
        RECT 95.765 2.240 95.905 13.130 ;
        RECT 96.325 2.240 96.535 13.130 ;
        RECT 85.125 1.910 96.535 2.240 ;
        RECT 98.215 2.240 98.355 13.130 ;
        RECT 98.775 2.240 98.915 13.130 ;
        RECT 99.335 2.240 99.475 13.130 ;
        RECT 99.895 2.240 100.035 13.130 ;
        RECT 100.455 2.240 100.595 13.130 ;
        RECT 101.015 2.240 101.155 13.130 ;
        RECT 101.575 2.240 101.715 13.130 ;
        RECT 102.135 2.240 102.275 13.130 ;
        RECT 102.695 2.240 102.835 13.130 ;
        RECT 103.255 2.240 103.395 13.130 ;
        RECT 103.815 2.240 103.955 13.130 ;
        RECT 104.375 2.240 104.515 13.130 ;
        RECT 104.935 2.240 105.075 13.130 ;
        RECT 105.495 2.240 105.635 13.130 ;
        RECT 106.055 2.240 106.195 13.130 ;
        RECT 106.615 2.240 106.755 13.130 ;
        RECT 107.175 2.240 107.315 13.130 ;
        RECT 107.735 2.240 107.875 13.130 ;
        RECT 108.295 2.240 108.435 13.130 ;
        RECT 108.855 2.240 108.995 13.130 ;
        RECT 109.415 2.240 109.625 13.130 ;
        RECT 98.215 1.910 109.625 2.240 ;
        RECT 111.305 2.240 111.445 13.130 ;
        RECT 111.865 2.240 112.005 13.130 ;
        RECT 112.425 2.240 112.565 13.130 ;
        RECT 112.985 2.240 113.125 13.130 ;
        RECT 113.545 2.240 113.685 13.130 ;
        RECT 114.105 2.240 114.245 13.130 ;
        RECT 114.665 2.240 114.805 13.130 ;
        RECT 115.225 2.240 115.365 13.130 ;
        RECT 115.785 2.240 115.925 13.130 ;
        RECT 116.345 2.240 116.485 13.130 ;
        RECT 116.905 2.240 117.045 13.130 ;
        RECT 117.465 2.240 117.605 13.130 ;
        RECT 118.025 2.240 118.165 13.130 ;
        RECT 118.585 2.240 118.725 13.130 ;
        RECT 119.145 2.240 119.285 13.130 ;
        RECT 119.705 2.240 119.845 13.130 ;
        RECT 120.265 2.240 120.405 13.130 ;
        RECT 120.825 2.240 120.965 13.130 ;
        RECT 121.385 2.240 121.525 13.130 ;
        RECT 121.945 2.240 122.085 13.130 ;
        RECT 122.505 2.240 122.715 13.130 ;
        RECT 111.305 1.910 122.715 2.240 ;
        RECT 124.395 2.240 124.535 13.130 ;
        RECT 124.955 2.240 125.095 13.130 ;
        RECT 125.515 2.240 125.655 13.130 ;
        RECT 126.075 2.240 126.215 13.130 ;
        RECT 126.635 2.240 126.775 13.130 ;
        RECT 127.195 2.240 127.335 13.130 ;
        RECT 127.755 2.240 127.895 13.130 ;
        RECT 128.315 2.240 128.455 13.130 ;
        RECT 128.875 2.240 129.015 13.130 ;
        RECT 129.435 2.240 129.575 13.130 ;
        RECT 129.995 2.240 130.135 13.130 ;
        RECT 130.555 2.240 130.695 13.130 ;
        RECT 131.115 2.240 131.255 13.130 ;
        RECT 131.675 2.240 131.815 13.130 ;
        RECT 132.235 2.240 132.375 13.130 ;
        RECT 132.795 2.240 132.935 13.130 ;
        RECT 133.355 2.240 133.495 13.130 ;
        RECT 133.915 2.240 134.055 13.130 ;
        RECT 134.475 2.240 134.615 13.130 ;
        RECT 135.035 2.240 135.175 13.130 ;
        RECT 135.595 2.240 135.805 13.130 ;
        RECT 124.395 1.910 135.805 2.240 ;
        RECT 137.485 2.260 137.625 13.150 ;
        RECT 138.045 2.260 138.185 13.150 ;
        RECT 138.605 2.260 138.745 13.150 ;
        RECT 139.165 2.260 139.305 13.150 ;
        RECT 139.725 2.260 139.865 13.150 ;
        RECT 140.285 2.260 140.425 13.150 ;
        RECT 140.845 2.260 140.985 13.150 ;
        RECT 141.405 2.260 141.545 13.150 ;
        RECT 141.965 2.260 142.105 13.150 ;
        RECT 142.525 2.260 142.665 13.150 ;
        RECT 143.085 2.260 143.225 13.150 ;
        RECT 143.645 2.260 143.785 13.150 ;
        RECT 144.205 2.260 144.345 13.150 ;
        RECT 144.765 2.260 144.905 13.150 ;
        RECT 145.325 2.260 145.465 13.150 ;
        RECT 145.885 2.260 146.025 13.150 ;
        RECT 146.445 2.260 146.585 13.150 ;
        RECT 147.005 2.260 147.145 13.150 ;
        RECT 147.565 2.260 147.705 13.150 ;
        RECT 148.125 2.260 148.265 13.150 ;
        RECT 148.685 2.260 148.895 13.150 ;
        RECT 137.485 1.930 148.895 2.260 ;
        RECT 150.575 2.260 150.715 13.150 ;
        RECT 151.135 2.260 151.275 13.150 ;
        RECT 151.695 2.260 151.835 13.150 ;
        RECT 152.255 2.260 152.395 13.150 ;
        RECT 152.815 2.260 152.955 13.150 ;
        RECT 153.375 2.260 153.515 13.150 ;
        RECT 153.935 2.260 154.075 13.150 ;
        RECT 154.495 2.260 154.635 13.150 ;
        RECT 155.055 2.260 155.195 13.150 ;
        RECT 155.615 2.260 155.755 13.150 ;
        RECT 156.175 2.260 156.315 13.150 ;
        RECT 156.735 2.260 156.875 13.150 ;
        RECT 157.295 2.260 157.435 13.150 ;
        RECT 157.855 2.260 157.995 13.150 ;
        RECT 158.415 2.260 158.555 13.150 ;
        RECT 158.975 2.260 159.115 13.150 ;
        RECT 159.535 2.260 159.675 13.150 ;
        RECT 160.095 2.260 160.235 13.150 ;
        RECT 160.655 2.260 160.795 13.150 ;
        RECT 161.215 2.260 161.355 13.150 ;
        RECT 161.775 2.260 161.985 13.150 ;
        RECT 150.575 1.930 161.985 2.260 ;
      LAYER via ;
        RECT 6.495 118.315 6.755 118.575 ;
        RECT 6.815 118.315 7.075 118.575 ;
        RECT 7.615 118.315 7.875 118.575 ;
        RECT 7.935 118.315 8.195 118.575 ;
        RECT 8.735 118.315 8.995 118.575 ;
        RECT 9.055 118.315 9.315 118.575 ;
        RECT 9.855 118.315 10.115 118.575 ;
        RECT 10.175 118.315 10.435 118.575 ;
        RECT 10.975 118.315 11.235 118.575 ;
        RECT 11.295 118.315 11.555 118.575 ;
        RECT 12.095 118.315 12.355 118.575 ;
        RECT 12.415 118.315 12.675 118.575 ;
        RECT 13.215 118.315 13.475 118.575 ;
        RECT 13.535 118.315 13.795 118.575 ;
        RECT 14.335 118.315 14.595 118.575 ;
        RECT 14.655 118.315 14.915 118.575 ;
        RECT 15.455 118.315 15.715 118.575 ;
        RECT 15.775 118.315 16.035 118.575 ;
        RECT 16.575 118.315 16.835 118.575 ;
        RECT 16.895 118.315 17.155 118.575 ;
        RECT 19.585 118.315 19.845 118.575 ;
        RECT 19.905 118.315 20.165 118.575 ;
        RECT 20.705 118.315 20.965 118.575 ;
        RECT 21.025 118.315 21.285 118.575 ;
        RECT 21.825 118.315 22.085 118.575 ;
        RECT 22.145 118.315 22.405 118.575 ;
        RECT 22.945 118.315 23.205 118.575 ;
        RECT 23.265 118.315 23.525 118.575 ;
        RECT 24.065 118.315 24.325 118.575 ;
        RECT 24.385 118.315 24.645 118.575 ;
        RECT 25.185 118.315 25.445 118.575 ;
        RECT 25.505 118.315 25.765 118.575 ;
        RECT 26.305 118.315 26.565 118.575 ;
        RECT 26.625 118.315 26.885 118.575 ;
        RECT 27.425 118.315 27.685 118.575 ;
        RECT 27.745 118.315 28.005 118.575 ;
        RECT 28.545 118.315 28.805 118.575 ;
        RECT 28.865 118.315 29.125 118.575 ;
        RECT 29.665 118.315 29.925 118.575 ;
        RECT 29.985 118.315 30.245 118.575 ;
        RECT 32.675 118.295 32.935 118.555 ;
        RECT 32.995 118.295 33.255 118.555 ;
        RECT 33.795 118.295 34.055 118.555 ;
        RECT 34.115 118.295 34.375 118.555 ;
        RECT 34.915 118.295 35.175 118.555 ;
        RECT 35.235 118.295 35.495 118.555 ;
        RECT 36.035 118.295 36.295 118.555 ;
        RECT 36.355 118.295 36.615 118.555 ;
        RECT 37.155 118.295 37.415 118.555 ;
        RECT 37.475 118.295 37.735 118.555 ;
        RECT 38.275 118.295 38.535 118.555 ;
        RECT 38.595 118.295 38.855 118.555 ;
        RECT 39.395 118.295 39.655 118.555 ;
        RECT 39.715 118.295 39.975 118.555 ;
        RECT 40.515 118.295 40.775 118.555 ;
        RECT 40.835 118.295 41.095 118.555 ;
        RECT 41.635 118.295 41.895 118.555 ;
        RECT 41.955 118.295 42.215 118.555 ;
        RECT 42.755 118.295 43.015 118.555 ;
        RECT 43.075 118.295 43.335 118.555 ;
        RECT 45.765 118.295 46.025 118.555 ;
        RECT 46.085 118.295 46.345 118.555 ;
        RECT 46.885 118.295 47.145 118.555 ;
        RECT 47.205 118.295 47.465 118.555 ;
        RECT 48.005 118.295 48.265 118.555 ;
        RECT 48.325 118.295 48.585 118.555 ;
        RECT 49.125 118.295 49.385 118.555 ;
        RECT 49.445 118.295 49.705 118.555 ;
        RECT 50.245 118.295 50.505 118.555 ;
        RECT 50.565 118.295 50.825 118.555 ;
        RECT 51.365 118.295 51.625 118.555 ;
        RECT 51.685 118.295 51.945 118.555 ;
        RECT 52.485 118.295 52.745 118.555 ;
        RECT 52.805 118.295 53.065 118.555 ;
        RECT 53.605 118.295 53.865 118.555 ;
        RECT 53.925 118.295 54.185 118.555 ;
        RECT 54.725 118.295 54.985 118.555 ;
        RECT 55.045 118.295 55.305 118.555 ;
        RECT 55.845 118.295 56.105 118.555 ;
        RECT 56.165 118.295 56.425 118.555 ;
        RECT 58.815 118.295 59.075 118.555 ;
        RECT 59.135 118.295 59.395 118.555 ;
        RECT 59.935 118.295 60.195 118.555 ;
        RECT 60.255 118.295 60.515 118.555 ;
        RECT 61.055 118.295 61.315 118.555 ;
        RECT 61.375 118.295 61.635 118.555 ;
        RECT 62.175 118.295 62.435 118.555 ;
        RECT 62.495 118.295 62.755 118.555 ;
        RECT 63.295 118.295 63.555 118.555 ;
        RECT 63.615 118.295 63.875 118.555 ;
        RECT 64.415 118.295 64.675 118.555 ;
        RECT 64.735 118.295 64.995 118.555 ;
        RECT 65.535 118.295 65.795 118.555 ;
        RECT 65.855 118.295 66.115 118.555 ;
        RECT 66.655 118.295 66.915 118.555 ;
        RECT 66.975 118.295 67.235 118.555 ;
        RECT 67.775 118.295 68.035 118.555 ;
        RECT 68.095 118.295 68.355 118.555 ;
        RECT 68.895 118.295 69.155 118.555 ;
        RECT 69.215 118.295 69.475 118.555 ;
        RECT 71.905 118.295 72.165 118.555 ;
        RECT 72.225 118.295 72.485 118.555 ;
        RECT 73.025 118.295 73.285 118.555 ;
        RECT 73.345 118.295 73.605 118.555 ;
        RECT 74.145 118.295 74.405 118.555 ;
        RECT 74.465 118.295 74.725 118.555 ;
        RECT 75.265 118.295 75.525 118.555 ;
        RECT 75.585 118.295 75.845 118.555 ;
        RECT 76.385 118.295 76.645 118.555 ;
        RECT 76.705 118.295 76.965 118.555 ;
        RECT 77.505 118.295 77.765 118.555 ;
        RECT 77.825 118.295 78.085 118.555 ;
        RECT 78.625 118.295 78.885 118.555 ;
        RECT 78.945 118.295 79.205 118.555 ;
        RECT 79.745 118.295 80.005 118.555 ;
        RECT 80.065 118.295 80.325 118.555 ;
        RECT 80.865 118.295 81.125 118.555 ;
        RECT 81.185 118.295 81.445 118.555 ;
        RECT 81.985 118.295 82.245 118.555 ;
        RECT 82.305 118.295 82.565 118.555 ;
        RECT 84.995 118.275 85.255 118.535 ;
        RECT 85.315 118.275 85.575 118.535 ;
        RECT 86.115 118.275 86.375 118.535 ;
        RECT 86.435 118.275 86.695 118.535 ;
        RECT 87.235 118.275 87.495 118.535 ;
        RECT 87.555 118.275 87.815 118.535 ;
        RECT 88.355 118.275 88.615 118.535 ;
        RECT 88.675 118.275 88.935 118.535 ;
        RECT 89.475 118.275 89.735 118.535 ;
        RECT 89.795 118.275 90.055 118.535 ;
        RECT 90.595 118.275 90.855 118.535 ;
        RECT 90.915 118.275 91.175 118.535 ;
        RECT 91.715 118.275 91.975 118.535 ;
        RECT 92.035 118.275 92.295 118.535 ;
        RECT 92.835 118.275 93.095 118.535 ;
        RECT 93.155 118.275 93.415 118.535 ;
        RECT 93.955 118.275 94.215 118.535 ;
        RECT 94.275 118.275 94.535 118.535 ;
        RECT 95.075 118.275 95.335 118.535 ;
        RECT 95.395 118.275 95.655 118.535 ;
        RECT 98.085 118.275 98.345 118.535 ;
        RECT 98.405 118.275 98.665 118.535 ;
        RECT 99.205 118.275 99.465 118.535 ;
        RECT 99.525 118.275 99.785 118.535 ;
        RECT 100.325 118.275 100.585 118.535 ;
        RECT 100.645 118.275 100.905 118.535 ;
        RECT 101.445 118.275 101.705 118.535 ;
        RECT 101.765 118.275 102.025 118.535 ;
        RECT 102.565 118.275 102.825 118.535 ;
        RECT 102.885 118.275 103.145 118.535 ;
        RECT 103.685 118.275 103.945 118.535 ;
        RECT 104.005 118.275 104.265 118.535 ;
        RECT 104.805 118.275 105.065 118.535 ;
        RECT 105.125 118.275 105.385 118.535 ;
        RECT 105.925 118.275 106.185 118.535 ;
        RECT 106.245 118.275 106.505 118.535 ;
        RECT 107.045 118.275 107.305 118.535 ;
        RECT 107.365 118.275 107.625 118.535 ;
        RECT 108.165 118.275 108.425 118.535 ;
        RECT 108.485 118.275 108.745 118.535 ;
        RECT 111.175 118.275 111.435 118.535 ;
        RECT 111.495 118.275 111.755 118.535 ;
        RECT 112.295 118.275 112.555 118.535 ;
        RECT 112.615 118.275 112.875 118.535 ;
        RECT 113.415 118.275 113.675 118.535 ;
        RECT 113.735 118.275 113.995 118.535 ;
        RECT 114.535 118.275 114.795 118.535 ;
        RECT 114.855 118.275 115.115 118.535 ;
        RECT 115.655 118.275 115.915 118.535 ;
        RECT 115.975 118.275 116.235 118.535 ;
        RECT 116.775 118.275 117.035 118.535 ;
        RECT 117.095 118.275 117.355 118.535 ;
        RECT 117.895 118.275 118.155 118.535 ;
        RECT 118.215 118.275 118.475 118.535 ;
        RECT 119.015 118.275 119.275 118.535 ;
        RECT 119.335 118.275 119.595 118.535 ;
        RECT 120.135 118.275 120.395 118.535 ;
        RECT 120.455 118.275 120.715 118.535 ;
        RECT 121.255 118.275 121.515 118.535 ;
        RECT 121.575 118.275 121.835 118.535 ;
        RECT 124.265 118.275 124.525 118.535 ;
        RECT 124.585 118.275 124.845 118.535 ;
        RECT 125.385 118.275 125.645 118.535 ;
        RECT 125.705 118.275 125.965 118.535 ;
        RECT 126.505 118.275 126.765 118.535 ;
        RECT 126.825 118.275 127.085 118.535 ;
        RECT 127.625 118.275 127.885 118.535 ;
        RECT 127.945 118.275 128.205 118.535 ;
        RECT 128.745 118.275 129.005 118.535 ;
        RECT 129.065 118.275 129.325 118.535 ;
        RECT 129.865 118.275 130.125 118.535 ;
        RECT 130.185 118.275 130.445 118.535 ;
        RECT 130.985 118.275 131.245 118.535 ;
        RECT 131.305 118.275 131.565 118.535 ;
        RECT 132.105 118.275 132.365 118.535 ;
        RECT 132.425 118.275 132.685 118.535 ;
        RECT 133.225 118.275 133.485 118.535 ;
        RECT 133.545 118.275 133.805 118.535 ;
        RECT 134.345 118.275 134.605 118.535 ;
        RECT 134.665 118.275 134.925 118.535 ;
        RECT 137.355 118.255 137.615 118.515 ;
        RECT 137.675 118.255 137.935 118.515 ;
        RECT 138.475 118.255 138.735 118.515 ;
        RECT 138.795 118.255 139.055 118.515 ;
        RECT 139.595 118.255 139.855 118.515 ;
        RECT 139.915 118.255 140.175 118.515 ;
        RECT 140.715 118.255 140.975 118.515 ;
        RECT 141.035 118.255 141.295 118.515 ;
        RECT 141.835 118.255 142.095 118.515 ;
        RECT 142.155 118.255 142.415 118.515 ;
        RECT 142.955 118.255 143.215 118.515 ;
        RECT 143.275 118.255 143.535 118.515 ;
        RECT 144.075 118.255 144.335 118.515 ;
        RECT 144.395 118.255 144.655 118.515 ;
        RECT 145.195 118.255 145.455 118.515 ;
        RECT 145.515 118.255 145.775 118.515 ;
        RECT 146.315 118.255 146.575 118.515 ;
        RECT 146.635 118.255 146.895 118.515 ;
        RECT 147.435 118.255 147.695 118.515 ;
        RECT 147.755 118.255 148.015 118.515 ;
        RECT 150.445 118.255 150.705 118.515 ;
        RECT 150.765 118.255 151.025 118.515 ;
        RECT 151.565 118.255 151.825 118.515 ;
        RECT 151.885 118.255 152.145 118.515 ;
        RECT 152.685 118.255 152.945 118.515 ;
        RECT 153.005 118.255 153.265 118.515 ;
        RECT 153.805 118.255 154.065 118.515 ;
        RECT 154.125 118.255 154.385 118.515 ;
        RECT 154.925 118.255 155.185 118.515 ;
        RECT 155.245 118.255 155.505 118.515 ;
        RECT 156.045 118.255 156.305 118.515 ;
        RECT 156.365 118.255 156.625 118.515 ;
        RECT 157.165 118.255 157.425 118.515 ;
        RECT 157.485 118.255 157.745 118.515 ;
        RECT 158.285 118.255 158.545 118.515 ;
        RECT 158.605 118.255 158.865 118.515 ;
        RECT 159.405 118.255 159.665 118.515 ;
        RECT 159.725 118.255 159.985 118.515 ;
        RECT 160.525 118.255 160.785 118.515 ;
        RECT 160.845 118.255 161.105 118.515 ;
        RECT 6.525 93.545 6.785 93.805 ;
        RECT 6.845 93.545 7.105 93.805 ;
        RECT 7.645 93.545 7.905 93.805 ;
        RECT 7.965 93.545 8.225 93.805 ;
        RECT 8.765 93.545 9.025 93.805 ;
        RECT 9.085 93.545 9.345 93.805 ;
        RECT 9.885 93.545 10.145 93.805 ;
        RECT 10.205 93.545 10.465 93.805 ;
        RECT 11.005 93.545 11.265 93.805 ;
        RECT 11.325 93.545 11.585 93.805 ;
        RECT 12.125 93.545 12.385 93.805 ;
        RECT 12.445 93.545 12.705 93.805 ;
        RECT 13.245 93.545 13.505 93.805 ;
        RECT 13.565 93.545 13.825 93.805 ;
        RECT 14.365 93.545 14.625 93.805 ;
        RECT 14.685 93.545 14.945 93.805 ;
        RECT 15.485 93.545 15.745 93.805 ;
        RECT 15.805 93.545 16.065 93.805 ;
        RECT 16.605 93.545 16.865 93.805 ;
        RECT 16.925 93.545 17.185 93.805 ;
        RECT 19.615 93.545 19.875 93.805 ;
        RECT 19.935 93.545 20.195 93.805 ;
        RECT 20.735 93.545 20.995 93.805 ;
        RECT 21.055 93.545 21.315 93.805 ;
        RECT 21.855 93.545 22.115 93.805 ;
        RECT 22.175 93.545 22.435 93.805 ;
        RECT 22.975 93.545 23.235 93.805 ;
        RECT 23.295 93.545 23.555 93.805 ;
        RECT 24.095 93.545 24.355 93.805 ;
        RECT 24.415 93.545 24.675 93.805 ;
        RECT 25.215 93.545 25.475 93.805 ;
        RECT 25.535 93.545 25.795 93.805 ;
        RECT 26.335 93.545 26.595 93.805 ;
        RECT 26.655 93.545 26.915 93.805 ;
        RECT 27.455 93.545 27.715 93.805 ;
        RECT 27.775 93.545 28.035 93.805 ;
        RECT 28.575 93.545 28.835 93.805 ;
        RECT 28.895 93.545 29.155 93.805 ;
        RECT 29.695 93.545 29.955 93.805 ;
        RECT 30.015 93.545 30.275 93.805 ;
        RECT 32.705 93.565 32.965 93.825 ;
        RECT 33.025 93.565 33.285 93.825 ;
        RECT 33.825 93.565 34.085 93.825 ;
        RECT 34.145 93.565 34.405 93.825 ;
        RECT 34.945 93.565 35.205 93.825 ;
        RECT 35.265 93.565 35.525 93.825 ;
        RECT 36.065 93.565 36.325 93.825 ;
        RECT 36.385 93.565 36.645 93.825 ;
        RECT 37.185 93.565 37.445 93.825 ;
        RECT 37.505 93.565 37.765 93.825 ;
        RECT 38.305 93.565 38.565 93.825 ;
        RECT 38.625 93.565 38.885 93.825 ;
        RECT 39.425 93.565 39.685 93.825 ;
        RECT 39.745 93.565 40.005 93.825 ;
        RECT 40.545 93.565 40.805 93.825 ;
        RECT 40.865 93.565 41.125 93.825 ;
        RECT 41.665 93.565 41.925 93.825 ;
        RECT 41.985 93.565 42.245 93.825 ;
        RECT 42.785 93.565 43.045 93.825 ;
        RECT 43.105 93.565 43.365 93.825 ;
        RECT 45.795 93.565 46.055 93.825 ;
        RECT 46.115 93.565 46.375 93.825 ;
        RECT 46.915 93.565 47.175 93.825 ;
        RECT 47.235 93.565 47.495 93.825 ;
        RECT 48.035 93.565 48.295 93.825 ;
        RECT 48.355 93.565 48.615 93.825 ;
        RECT 49.155 93.565 49.415 93.825 ;
        RECT 49.475 93.565 49.735 93.825 ;
        RECT 50.275 93.565 50.535 93.825 ;
        RECT 50.595 93.565 50.855 93.825 ;
        RECT 51.395 93.565 51.655 93.825 ;
        RECT 51.715 93.565 51.975 93.825 ;
        RECT 52.515 93.565 52.775 93.825 ;
        RECT 52.835 93.565 53.095 93.825 ;
        RECT 53.635 93.565 53.895 93.825 ;
        RECT 53.955 93.565 54.215 93.825 ;
        RECT 54.755 93.565 55.015 93.825 ;
        RECT 55.075 93.565 55.335 93.825 ;
        RECT 55.875 93.565 56.135 93.825 ;
        RECT 56.195 93.565 56.455 93.825 ;
        RECT 58.845 93.565 59.105 93.825 ;
        RECT 59.165 93.565 59.425 93.825 ;
        RECT 59.965 93.565 60.225 93.825 ;
        RECT 60.285 93.565 60.545 93.825 ;
        RECT 61.085 93.565 61.345 93.825 ;
        RECT 61.405 93.565 61.665 93.825 ;
        RECT 62.205 93.565 62.465 93.825 ;
        RECT 62.525 93.565 62.785 93.825 ;
        RECT 63.325 93.565 63.585 93.825 ;
        RECT 63.645 93.565 63.905 93.825 ;
        RECT 64.445 93.565 64.705 93.825 ;
        RECT 64.765 93.565 65.025 93.825 ;
        RECT 65.565 93.565 65.825 93.825 ;
        RECT 65.885 93.565 66.145 93.825 ;
        RECT 66.685 93.565 66.945 93.825 ;
        RECT 67.005 93.565 67.265 93.825 ;
        RECT 67.805 93.565 68.065 93.825 ;
        RECT 68.125 93.565 68.385 93.825 ;
        RECT 68.925 93.565 69.185 93.825 ;
        RECT 69.245 93.565 69.505 93.825 ;
        RECT 71.935 93.565 72.195 93.825 ;
        RECT 72.255 93.565 72.515 93.825 ;
        RECT 73.055 93.565 73.315 93.825 ;
        RECT 73.375 93.565 73.635 93.825 ;
        RECT 74.175 93.565 74.435 93.825 ;
        RECT 74.495 93.565 74.755 93.825 ;
        RECT 75.295 93.565 75.555 93.825 ;
        RECT 75.615 93.565 75.875 93.825 ;
        RECT 76.415 93.565 76.675 93.825 ;
        RECT 76.735 93.565 76.995 93.825 ;
        RECT 77.535 93.565 77.795 93.825 ;
        RECT 77.855 93.565 78.115 93.825 ;
        RECT 78.655 93.565 78.915 93.825 ;
        RECT 78.975 93.565 79.235 93.825 ;
        RECT 79.775 93.565 80.035 93.825 ;
        RECT 80.095 93.565 80.355 93.825 ;
        RECT 80.895 93.565 81.155 93.825 ;
        RECT 81.215 93.565 81.475 93.825 ;
        RECT 82.015 93.565 82.275 93.825 ;
        RECT 82.335 93.565 82.595 93.825 ;
        RECT 85.025 93.585 85.285 93.845 ;
        RECT 85.345 93.585 85.605 93.845 ;
        RECT 86.145 93.585 86.405 93.845 ;
        RECT 86.465 93.585 86.725 93.845 ;
        RECT 87.265 93.585 87.525 93.845 ;
        RECT 87.585 93.585 87.845 93.845 ;
        RECT 88.385 93.585 88.645 93.845 ;
        RECT 88.705 93.585 88.965 93.845 ;
        RECT 89.505 93.585 89.765 93.845 ;
        RECT 89.825 93.585 90.085 93.845 ;
        RECT 90.625 93.585 90.885 93.845 ;
        RECT 90.945 93.585 91.205 93.845 ;
        RECT 91.745 93.585 92.005 93.845 ;
        RECT 92.065 93.585 92.325 93.845 ;
        RECT 92.865 93.585 93.125 93.845 ;
        RECT 93.185 93.585 93.445 93.845 ;
        RECT 93.985 93.585 94.245 93.845 ;
        RECT 94.305 93.585 94.565 93.845 ;
        RECT 95.105 93.585 95.365 93.845 ;
        RECT 95.425 93.585 95.685 93.845 ;
        RECT 98.115 93.585 98.375 93.845 ;
        RECT 98.435 93.585 98.695 93.845 ;
        RECT 99.235 93.585 99.495 93.845 ;
        RECT 99.555 93.585 99.815 93.845 ;
        RECT 100.355 93.585 100.615 93.845 ;
        RECT 100.675 93.585 100.935 93.845 ;
        RECT 101.475 93.585 101.735 93.845 ;
        RECT 101.795 93.585 102.055 93.845 ;
        RECT 102.595 93.585 102.855 93.845 ;
        RECT 102.915 93.585 103.175 93.845 ;
        RECT 103.715 93.585 103.975 93.845 ;
        RECT 104.035 93.585 104.295 93.845 ;
        RECT 104.835 93.585 105.095 93.845 ;
        RECT 105.155 93.585 105.415 93.845 ;
        RECT 105.955 93.585 106.215 93.845 ;
        RECT 106.275 93.585 106.535 93.845 ;
        RECT 107.075 93.585 107.335 93.845 ;
        RECT 107.395 93.585 107.655 93.845 ;
        RECT 108.195 93.585 108.455 93.845 ;
        RECT 108.515 93.585 108.775 93.845 ;
        RECT 111.205 93.585 111.465 93.845 ;
        RECT 111.525 93.585 111.785 93.845 ;
        RECT 112.325 93.585 112.585 93.845 ;
        RECT 112.645 93.585 112.905 93.845 ;
        RECT 113.445 93.585 113.705 93.845 ;
        RECT 113.765 93.585 114.025 93.845 ;
        RECT 114.565 93.585 114.825 93.845 ;
        RECT 114.885 93.585 115.145 93.845 ;
        RECT 115.685 93.585 115.945 93.845 ;
        RECT 116.005 93.585 116.265 93.845 ;
        RECT 116.805 93.585 117.065 93.845 ;
        RECT 117.125 93.585 117.385 93.845 ;
        RECT 117.925 93.585 118.185 93.845 ;
        RECT 118.245 93.585 118.505 93.845 ;
        RECT 119.045 93.585 119.305 93.845 ;
        RECT 119.365 93.585 119.625 93.845 ;
        RECT 120.165 93.585 120.425 93.845 ;
        RECT 120.485 93.585 120.745 93.845 ;
        RECT 121.285 93.585 121.545 93.845 ;
        RECT 121.605 93.585 121.865 93.845 ;
        RECT 124.295 93.585 124.555 93.845 ;
        RECT 124.615 93.585 124.875 93.845 ;
        RECT 125.415 93.585 125.675 93.845 ;
        RECT 125.735 93.585 125.995 93.845 ;
        RECT 126.535 93.585 126.795 93.845 ;
        RECT 126.855 93.585 127.115 93.845 ;
        RECT 127.655 93.585 127.915 93.845 ;
        RECT 127.975 93.585 128.235 93.845 ;
        RECT 128.775 93.585 129.035 93.845 ;
        RECT 129.095 93.585 129.355 93.845 ;
        RECT 129.895 93.585 130.155 93.845 ;
        RECT 130.215 93.585 130.475 93.845 ;
        RECT 131.015 93.585 131.275 93.845 ;
        RECT 131.335 93.585 131.595 93.845 ;
        RECT 132.135 93.585 132.395 93.845 ;
        RECT 132.455 93.585 132.715 93.845 ;
        RECT 133.255 93.585 133.515 93.845 ;
        RECT 133.575 93.585 133.835 93.845 ;
        RECT 134.375 93.585 134.635 93.845 ;
        RECT 134.695 93.585 134.955 93.845 ;
        RECT 137.385 93.605 137.645 93.865 ;
        RECT 137.705 93.605 137.965 93.865 ;
        RECT 138.505 93.605 138.765 93.865 ;
        RECT 138.825 93.605 139.085 93.865 ;
        RECT 139.625 93.605 139.885 93.865 ;
        RECT 139.945 93.605 140.205 93.865 ;
        RECT 140.745 93.605 141.005 93.865 ;
        RECT 141.065 93.605 141.325 93.865 ;
        RECT 141.865 93.605 142.125 93.865 ;
        RECT 142.185 93.605 142.445 93.865 ;
        RECT 142.985 93.605 143.245 93.865 ;
        RECT 143.305 93.605 143.565 93.865 ;
        RECT 144.105 93.605 144.365 93.865 ;
        RECT 144.425 93.605 144.685 93.865 ;
        RECT 145.225 93.605 145.485 93.865 ;
        RECT 145.545 93.605 145.805 93.865 ;
        RECT 146.345 93.605 146.605 93.865 ;
        RECT 146.665 93.605 146.925 93.865 ;
        RECT 147.465 93.605 147.725 93.865 ;
        RECT 147.785 93.605 148.045 93.865 ;
        RECT 150.475 93.605 150.735 93.865 ;
        RECT 150.795 93.605 151.055 93.865 ;
        RECT 151.595 93.605 151.855 93.865 ;
        RECT 151.915 93.605 152.175 93.865 ;
        RECT 152.715 93.605 152.975 93.865 ;
        RECT 153.035 93.605 153.295 93.865 ;
        RECT 153.835 93.605 154.095 93.865 ;
        RECT 154.155 93.605 154.415 93.865 ;
        RECT 154.955 93.605 155.215 93.865 ;
        RECT 155.275 93.605 155.535 93.865 ;
        RECT 156.075 93.605 156.335 93.865 ;
        RECT 156.395 93.605 156.655 93.865 ;
        RECT 157.195 93.605 157.455 93.865 ;
        RECT 157.515 93.605 157.775 93.865 ;
        RECT 158.315 93.605 158.575 93.865 ;
        RECT 158.635 93.605 158.895 93.865 ;
        RECT 159.435 93.605 159.695 93.865 ;
        RECT 159.755 93.605 160.015 93.865 ;
        RECT 160.555 93.605 160.815 93.865 ;
        RECT 160.875 93.605 161.135 93.865 ;
        RECT 151.215 89.470 151.475 89.730 ;
        RECT 167.325 89.465 167.800 89.940 ;
        RECT 1.980 88.345 2.450 88.815 ;
        RECT 148.780 88.230 149.040 88.490 ;
        RECT 178.100 65.450 178.360 65.710 ;
        RECT 178.100 65.130 178.360 65.390 ;
        RECT 178.100 62.310 178.360 62.570 ;
        RECT 178.100 61.990 178.360 62.250 ;
        RECT 178.100 59.260 178.360 59.520 ;
        RECT 178.100 58.940 178.360 59.200 ;
        RECT 178.100 56.120 178.360 56.380 ;
        RECT 178.100 55.800 178.360 56.060 ;
        RECT 1.940 33.215 2.410 33.685 ;
        RECT 166.065 29.910 166.540 30.385 ;
        RECT 6.935 26.675 7.195 26.935 ;
        RECT 7.255 26.675 7.515 26.935 ;
        RECT 8.055 26.675 8.315 26.935 ;
        RECT 8.375 26.675 8.635 26.935 ;
        RECT 9.175 26.675 9.435 26.935 ;
        RECT 9.495 26.675 9.755 26.935 ;
        RECT 10.295 26.675 10.555 26.935 ;
        RECT 10.615 26.675 10.875 26.935 ;
        RECT 11.415 26.675 11.675 26.935 ;
        RECT 11.735 26.675 11.995 26.935 ;
        RECT 12.535 26.675 12.795 26.935 ;
        RECT 12.855 26.675 13.115 26.935 ;
        RECT 13.655 26.675 13.915 26.935 ;
        RECT 13.975 26.675 14.235 26.935 ;
        RECT 14.775 26.675 15.035 26.935 ;
        RECT 15.095 26.675 15.355 26.935 ;
        RECT 15.895 26.675 16.155 26.935 ;
        RECT 16.215 26.675 16.475 26.935 ;
        RECT 17.015 26.675 17.275 26.935 ;
        RECT 17.335 26.675 17.595 26.935 ;
        RECT 20.025 26.675 20.285 26.935 ;
        RECT 20.345 26.675 20.605 26.935 ;
        RECT 21.145 26.675 21.405 26.935 ;
        RECT 21.465 26.675 21.725 26.935 ;
        RECT 22.265 26.675 22.525 26.935 ;
        RECT 22.585 26.675 22.845 26.935 ;
        RECT 23.385 26.675 23.645 26.935 ;
        RECT 23.705 26.675 23.965 26.935 ;
        RECT 24.505 26.675 24.765 26.935 ;
        RECT 24.825 26.675 25.085 26.935 ;
        RECT 25.625 26.675 25.885 26.935 ;
        RECT 25.945 26.675 26.205 26.935 ;
        RECT 26.745 26.675 27.005 26.935 ;
        RECT 27.065 26.675 27.325 26.935 ;
        RECT 27.865 26.675 28.125 26.935 ;
        RECT 28.185 26.675 28.445 26.935 ;
        RECT 28.985 26.675 29.245 26.935 ;
        RECT 29.305 26.675 29.565 26.935 ;
        RECT 30.105 26.675 30.365 26.935 ;
        RECT 30.425 26.675 30.685 26.935 ;
        RECT 33.115 26.655 33.375 26.915 ;
        RECT 33.435 26.655 33.695 26.915 ;
        RECT 34.235 26.655 34.495 26.915 ;
        RECT 34.555 26.655 34.815 26.915 ;
        RECT 35.355 26.655 35.615 26.915 ;
        RECT 35.675 26.655 35.935 26.915 ;
        RECT 36.475 26.655 36.735 26.915 ;
        RECT 36.795 26.655 37.055 26.915 ;
        RECT 37.595 26.655 37.855 26.915 ;
        RECT 37.915 26.655 38.175 26.915 ;
        RECT 38.715 26.655 38.975 26.915 ;
        RECT 39.035 26.655 39.295 26.915 ;
        RECT 39.835 26.655 40.095 26.915 ;
        RECT 40.155 26.655 40.415 26.915 ;
        RECT 40.955 26.655 41.215 26.915 ;
        RECT 41.275 26.655 41.535 26.915 ;
        RECT 42.075 26.655 42.335 26.915 ;
        RECT 42.395 26.655 42.655 26.915 ;
        RECT 43.195 26.655 43.455 26.915 ;
        RECT 43.515 26.655 43.775 26.915 ;
        RECT 46.205 26.655 46.465 26.915 ;
        RECT 46.525 26.655 46.785 26.915 ;
        RECT 47.325 26.655 47.585 26.915 ;
        RECT 47.645 26.655 47.905 26.915 ;
        RECT 48.445 26.655 48.705 26.915 ;
        RECT 48.765 26.655 49.025 26.915 ;
        RECT 49.565 26.655 49.825 26.915 ;
        RECT 49.885 26.655 50.145 26.915 ;
        RECT 50.685 26.655 50.945 26.915 ;
        RECT 51.005 26.655 51.265 26.915 ;
        RECT 51.805 26.655 52.065 26.915 ;
        RECT 52.125 26.655 52.385 26.915 ;
        RECT 52.925 26.655 53.185 26.915 ;
        RECT 53.245 26.655 53.505 26.915 ;
        RECT 54.045 26.655 54.305 26.915 ;
        RECT 54.365 26.655 54.625 26.915 ;
        RECT 55.165 26.655 55.425 26.915 ;
        RECT 55.485 26.655 55.745 26.915 ;
        RECT 56.285 26.655 56.545 26.915 ;
        RECT 56.605 26.655 56.865 26.915 ;
        RECT 59.255 26.655 59.515 26.915 ;
        RECT 59.575 26.655 59.835 26.915 ;
        RECT 60.375 26.655 60.635 26.915 ;
        RECT 60.695 26.655 60.955 26.915 ;
        RECT 61.495 26.655 61.755 26.915 ;
        RECT 61.815 26.655 62.075 26.915 ;
        RECT 62.615 26.655 62.875 26.915 ;
        RECT 62.935 26.655 63.195 26.915 ;
        RECT 63.735 26.655 63.995 26.915 ;
        RECT 64.055 26.655 64.315 26.915 ;
        RECT 64.855 26.655 65.115 26.915 ;
        RECT 65.175 26.655 65.435 26.915 ;
        RECT 65.975 26.655 66.235 26.915 ;
        RECT 66.295 26.655 66.555 26.915 ;
        RECT 67.095 26.655 67.355 26.915 ;
        RECT 67.415 26.655 67.675 26.915 ;
        RECT 68.215 26.655 68.475 26.915 ;
        RECT 68.535 26.655 68.795 26.915 ;
        RECT 69.335 26.655 69.595 26.915 ;
        RECT 69.655 26.655 69.915 26.915 ;
        RECT 72.345 26.655 72.605 26.915 ;
        RECT 72.665 26.655 72.925 26.915 ;
        RECT 73.465 26.655 73.725 26.915 ;
        RECT 73.785 26.655 74.045 26.915 ;
        RECT 74.585 26.655 74.845 26.915 ;
        RECT 74.905 26.655 75.165 26.915 ;
        RECT 75.705 26.655 75.965 26.915 ;
        RECT 76.025 26.655 76.285 26.915 ;
        RECT 76.825 26.655 77.085 26.915 ;
        RECT 77.145 26.655 77.405 26.915 ;
        RECT 77.945 26.655 78.205 26.915 ;
        RECT 78.265 26.655 78.525 26.915 ;
        RECT 79.065 26.655 79.325 26.915 ;
        RECT 79.385 26.655 79.645 26.915 ;
        RECT 80.185 26.655 80.445 26.915 ;
        RECT 80.505 26.655 80.765 26.915 ;
        RECT 81.305 26.655 81.565 26.915 ;
        RECT 81.625 26.655 81.885 26.915 ;
        RECT 82.425 26.655 82.685 26.915 ;
        RECT 82.745 26.655 83.005 26.915 ;
        RECT 85.435 26.635 85.695 26.895 ;
        RECT 85.755 26.635 86.015 26.895 ;
        RECT 86.555 26.635 86.815 26.895 ;
        RECT 86.875 26.635 87.135 26.895 ;
        RECT 87.675 26.635 87.935 26.895 ;
        RECT 87.995 26.635 88.255 26.895 ;
        RECT 88.795 26.635 89.055 26.895 ;
        RECT 89.115 26.635 89.375 26.895 ;
        RECT 89.915 26.635 90.175 26.895 ;
        RECT 90.235 26.635 90.495 26.895 ;
        RECT 91.035 26.635 91.295 26.895 ;
        RECT 91.355 26.635 91.615 26.895 ;
        RECT 92.155 26.635 92.415 26.895 ;
        RECT 92.475 26.635 92.735 26.895 ;
        RECT 93.275 26.635 93.535 26.895 ;
        RECT 93.595 26.635 93.855 26.895 ;
        RECT 94.395 26.635 94.655 26.895 ;
        RECT 94.715 26.635 94.975 26.895 ;
        RECT 95.515 26.635 95.775 26.895 ;
        RECT 95.835 26.635 96.095 26.895 ;
        RECT 98.525 26.635 98.785 26.895 ;
        RECT 98.845 26.635 99.105 26.895 ;
        RECT 99.645 26.635 99.905 26.895 ;
        RECT 99.965 26.635 100.225 26.895 ;
        RECT 100.765 26.635 101.025 26.895 ;
        RECT 101.085 26.635 101.345 26.895 ;
        RECT 101.885 26.635 102.145 26.895 ;
        RECT 102.205 26.635 102.465 26.895 ;
        RECT 103.005 26.635 103.265 26.895 ;
        RECT 103.325 26.635 103.585 26.895 ;
        RECT 104.125 26.635 104.385 26.895 ;
        RECT 104.445 26.635 104.705 26.895 ;
        RECT 105.245 26.635 105.505 26.895 ;
        RECT 105.565 26.635 105.825 26.895 ;
        RECT 106.365 26.635 106.625 26.895 ;
        RECT 106.685 26.635 106.945 26.895 ;
        RECT 107.485 26.635 107.745 26.895 ;
        RECT 107.805 26.635 108.065 26.895 ;
        RECT 108.605 26.635 108.865 26.895 ;
        RECT 108.925 26.635 109.185 26.895 ;
        RECT 111.615 26.635 111.875 26.895 ;
        RECT 111.935 26.635 112.195 26.895 ;
        RECT 112.735 26.635 112.995 26.895 ;
        RECT 113.055 26.635 113.315 26.895 ;
        RECT 113.855 26.635 114.115 26.895 ;
        RECT 114.175 26.635 114.435 26.895 ;
        RECT 114.975 26.635 115.235 26.895 ;
        RECT 115.295 26.635 115.555 26.895 ;
        RECT 116.095 26.635 116.355 26.895 ;
        RECT 116.415 26.635 116.675 26.895 ;
        RECT 117.215 26.635 117.475 26.895 ;
        RECT 117.535 26.635 117.795 26.895 ;
        RECT 118.335 26.635 118.595 26.895 ;
        RECT 118.655 26.635 118.915 26.895 ;
        RECT 119.455 26.635 119.715 26.895 ;
        RECT 119.775 26.635 120.035 26.895 ;
        RECT 120.575 26.635 120.835 26.895 ;
        RECT 120.895 26.635 121.155 26.895 ;
        RECT 121.695 26.635 121.955 26.895 ;
        RECT 122.015 26.635 122.275 26.895 ;
        RECT 124.705 26.635 124.965 26.895 ;
        RECT 125.025 26.635 125.285 26.895 ;
        RECT 125.825 26.635 126.085 26.895 ;
        RECT 126.145 26.635 126.405 26.895 ;
        RECT 126.945 26.635 127.205 26.895 ;
        RECT 127.265 26.635 127.525 26.895 ;
        RECT 128.065 26.635 128.325 26.895 ;
        RECT 128.385 26.635 128.645 26.895 ;
        RECT 129.185 26.635 129.445 26.895 ;
        RECT 129.505 26.635 129.765 26.895 ;
        RECT 130.305 26.635 130.565 26.895 ;
        RECT 130.625 26.635 130.885 26.895 ;
        RECT 131.425 26.635 131.685 26.895 ;
        RECT 131.745 26.635 132.005 26.895 ;
        RECT 132.545 26.635 132.805 26.895 ;
        RECT 132.865 26.635 133.125 26.895 ;
        RECT 133.665 26.635 133.925 26.895 ;
        RECT 133.985 26.635 134.245 26.895 ;
        RECT 134.785 26.635 135.045 26.895 ;
        RECT 135.105 26.635 135.365 26.895 ;
        RECT 137.795 26.615 138.055 26.875 ;
        RECT 138.115 26.615 138.375 26.875 ;
        RECT 138.915 26.615 139.175 26.875 ;
        RECT 139.235 26.615 139.495 26.875 ;
        RECT 140.035 26.615 140.295 26.875 ;
        RECT 140.355 26.615 140.615 26.875 ;
        RECT 141.155 26.615 141.415 26.875 ;
        RECT 141.475 26.615 141.735 26.875 ;
        RECT 142.275 26.615 142.535 26.875 ;
        RECT 142.595 26.615 142.855 26.875 ;
        RECT 143.395 26.615 143.655 26.875 ;
        RECT 143.715 26.615 143.975 26.875 ;
        RECT 144.515 26.615 144.775 26.875 ;
        RECT 144.835 26.615 145.095 26.875 ;
        RECT 145.635 26.615 145.895 26.875 ;
        RECT 145.955 26.615 146.215 26.875 ;
        RECT 146.755 26.615 147.015 26.875 ;
        RECT 147.075 26.615 147.335 26.875 ;
        RECT 147.875 26.615 148.135 26.875 ;
        RECT 148.195 26.615 148.455 26.875 ;
        RECT 150.885 26.615 151.145 26.875 ;
        RECT 151.205 26.615 151.465 26.875 ;
        RECT 152.005 26.615 152.265 26.875 ;
        RECT 152.325 26.615 152.585 26.875 ;
        RECT 153.125 26.615 153.385 26.875 ;
        RECT 153.445 26.615 153.705 26.875 ;
        RECT 154.245 26.615 154.505 26.875 ;
        RECT 154.565 26.615 154.825 26.875 ;
        RECT 155.365 26.615 155.625 26.875 ;
        RECT 155.685 26.615 155.945 26.875 ;
        RECT 156.485 26.615 156.745 26.875 ;
        RECT 156.805 26.615 157.065 26.875 ;
        RECT 157.605 26.615 157.865 26.875 ;
        RECT 157.925 26.615 158.185 26.875 ;
        RECT 158.725 26.615 158.985 26.875 ;
        RECT 159.045 26.615 159.305 26.875 ;
        RECT 159.845 26.615 160.105 26.875 ;
        RECT 160.165 26.615 160.425 26.875 ;
        RECT 160.965 26.615 161.225 26.875 ;
        RECT 161.285 26.615 161.545 26.875 ;
        RECT 6.965 1.905 7.225 2.165 ;
        RECT 7.285 1.905 7.545 2.165 ;
        RECT 8.085 1.905 8.345 2.165 ;
        RECT 8.405 1.905 8.665 2.165 ;
        RECT 9.205 1.905 9.465 2.165 ;
        RECT 9.525 1.905 9.785 2.165 ;
        RECT 10.325 1.905 10.585 2.165 ;
        RECT 10.645 1.905 10.905 2.165 ;
        RECT 11.445 1.905 11.705 2.165 ;
        RECT 11.765 1.905 12.025 2.165 ;
        RECT 12.565 1.905 12.825 2.165 ;
        RECT 12.885 1.905 13.145 2.165 ;
        RECT 13.685 1.905 13.945 2.165 ;
        RECT 14.005 1.905 14.265 2.165 ;
        RECT 14.805 1.905 15.065 2.165 ;
        RECT 15.125 1.905 15.385 2.165 ;
        RECT 15.925 1.905 16.185 2.165 ;
        RECT 16.245 1.905 16.505 2.165 ;
        RECT 17.045 1.905 17.305 2.165 ;
        RECT 17.365 1.905 17.625 2.165 ;
        RECT 20.055 1.905 20.315 2.165 ;
        RECT 20.375 1.905 20.635 2.165 ;
        RECT 21.175 1.905 21.435 2.165 ;
        RECT 21.495 1.905 21.755 2.165 ;
        RECT 22.295 1.905 22.555 2.165 ;
        RECT 22.615 1.905 22.875 2.165 ;
        RECT 23.415 1.905 23.675 2.165 ;
        RECT 23.735 1.905 23.995 2.165 ;
        RECT 24.535 1.905 24.795 2.165 ;
        RECT 24.855 1.905 25.115 2.165 ;
        RECT 25.655 1.905 25.915 2.165 ;
        RECT 25.975 1.905 26.235 2.165 ;
        RECT 26.775 1.905 27.035 2.165 ;
        RECT 27.095 1.905 27.355 2.165 ;
        RECT 27.895 1.905 28.155 2.165 ;
        RECT 28.215 1.905 28.475 2.165 ;
        RECT 29.015 1.905 29.275 2.165 ;
        RECT 29.335 1.905 29.595 2.165 ;
        RECT 30.135 1.905 30.395 2.165 ;
        RECT 30.455 1.905 30.715 2.165 ;
        RECT 33.145 1.925 33.405 2.185 ;
        RECT 33.465 1.925 33.725 2.185 ;
        RECT 34.265 1.925 34.525 2.185 ;
        RECT 34.585 1.925 34.845 2.185 ;
        RECT 35.385 1.925 35.645 2.185 ;
        RECT 35.705 1.925 35.965 2.185 ;
        RECT 36.505 1.925 36.765 2.185 ;
        RECT 36.825 1.925 37.085 2.185 ;
        RECT 37.625 1.925 37.885 2.185 ;
        RECT 37.945 1.925 38.205 2.185 ;
        RECT 38.745 1.925 39.005 2.185 ;
        RECT 39.065 1.925 39.325 2.185 ;
        RECT 39.865 1.925 40.125 2.185 ;
        RECT 40.185 1.925 40.445 2.185 ;
        RECT 40.985 1.925 41.245 2.185 ;
        RECT 41.305 1.925 41.565 2.185 ;
        RECT 42.105 1.925 42.365 2.185 ;
        RECT 42.425 1.925 42.685 2.185 ;
        RECT 43.225 1.925 43.485 2.185 ;
        RECT 43.545 1.925 43.805 2.185 ;
        RECT 46.235 1.925 46.495 2.185 ;
        RECT 46.555 1.925 46.815 2.185 ;
        RECT 47.355 1.925 47.615 2.185 ;
        RECT 47.675 1.925 47.935 2.185 ;
        RECT 48.475 1.925 48.735 2.185 ;
        RECT 48.795 1.925 49.055 2.185 ;
        RECT 49.595 1.925 49.855 2.185 ;
        RECT 49.915 1.925 50.175 2.185 ;
        RECT 50.715 1.925 50.975 2.185 ;
        RECT 51.035 1.925 51.295 2.185 ;
        RECT 51.835 1.925 52.095 2.185 ;
        RECT 52.155 1.925 52.415 2.185 ;
        RECT 52.955 1.925 53.215 2.185 ;
        RECT 53.275 1.925 53.535 2.185 ;
        RECT 54.075 1.925 54.335 2.185 ;
        RECT 54.395 1.925 54.655 2.185 ;
        RECT 55.195 1.925 55.455 2.185 ;
        RECT 55.515 1.925 55.775 2.185 ;
        RECT 56.315 1.925 56.575 2.185 ;
        RECT 56.635 1.925 56.895 2.185 ;
        RECT 59.285 1.925 59.545 2.185 ;
        RECT 59.605 1.925 59.865 2.185 ;
        RECT 60.405 1.925 60.665 2.185 ;
        RECT 60.725 1.925 60.985 2.185 ;
        RECT 61.525 1.925 61.785 2.185 ;
        RECT 61.845 1.925 62.105 2.185 ;
        RECT 62.645 1.925 62.905 2.185 ;
        RECT 62.965 1.925 63.225 2.185 ;
        RECT 63.765 1.925 64.025 2.185 ;
        RECT 64.085 1.925 64.345 2.185 ;
        RECT 64.885 1.925 65.145 2.185 ;
        RECT 65.205 1.925 65.465 2.185 ;
        RECT 66.005 1.925 66.265 2.185 ;
        RECT 66.325 1.925 66.585 2.185 ;
        RECT 67.125 1.925 67.385 2.185 ;
        RECT 67.445 1.925 67.705 2.185 ;
        RECT 68.245 1.925 68.505 2.185 ;
        RECT 68.565 1.925 68.825 2.185 ;
        RECT 69.365 1.925 69.625 2.185 ;
        RECT 69.685 1.925 69.945 2.185 ;
        RECT 72.375 1.925 72.635 2.185 ;
        RECT 72.695 1.925 72.955 2.185 ;
        RECT 73.495 1.925 73.755 2.185 ;
        RECT 73.815 1.925 74.075 2.185 ;
        RECT 74.615 1.925 74.875 2.185 ;
        RECT 74.935 1.925 75.195 2.185 ;
        RECT 75.735 1.925 75.995 2.185 ;
        RECT 76.055 1.925 76.315 2.185 ;
        RECT 76.855 1.925 77.115 2.185 ;
        RECT 77.175 1.925 77.435 2.185 ;
        RECT 77.975 1.925 78.235 2.185 ;
        RECT 78.295 1.925 78.555 2.185 ;
        RECT 79.095 1.925 79.355 2.185 ;
        RECT 79.415 1.925 79.675 2.185 ;
        RECT 80.215 1.925 80.475 2.185 ;
        RECT 80.535 1.925 80.795 2.185 ;
        RECT 81.335 1.925 81.595 2.185 ;
        RECT 81.655 1.925 81.915 2.185 ;
        RECT 82.455 1.925 82.715 2.185 ;
        RECT 82.775 1.925 83.035 2.185 ;
        RECT 85.465 1.945 85.725 2.205 ;
        RECT 85.785 1.945 86.045 2.205 ;
        RECT 86.585 1.945 86.845 2.205 ;
        RECT 86.905 1.945 87.165 2.205 ;
        RECT 87.705 1.945 87.965 2.205 ;
        RECT 88.025 1.945 88.285 2.205 ;
        RECT 88.825 1.945 89.085 2.205 ;
        RECT 89.145 1.945 89.405 2.205 ;
        RECT 89.945 1.945 90.205 2.205 ;
        RECT 90.265 1.945 90.525 2.205 ;
        RECT 91.065 1.945 91.325 2.205 ;
        RECT 91.385 1.945 91.645 2.205 ;
        RECT 92.185 1.945 92.445 2.205 ;
        RECT 92.505 1.945 92.765 2.205 ;
        RECT 93.305 1.945 93.565 2.205 ;
        RECT 93.625 1.945 93.885 2.205 ;
        RECT 94.425 1.945 94.685 2.205 ;
        RECT 94.745 1.945 95.005 2.205 ;
        RECT 95.545 1.945 95.805 2.205 ;
        RECT 95.865 1.945 96.125 2.205 ;
        RECT 98.555 1.945 98.815 2.205 ;
        RECT 98.875 1.945 99.135 2.205 ;
        RECT 99.675 1.945 99.935 2.205 ;
        RECT 99.995 1.945 100.255 2.205 ;
        RECT 100.795 1.945 101.055 2.205 ;
        RECT 101.115 1.945 101.375 2.205 ;
        RECT 101.915 1.945 102.175 2.205 ;
        RECT 102.235 1.945 102.495 2.205 ;
        RECT 103.035 1.945 103.295 2.205 ;
        RECT 103.355 1.945 103.615 2.205 ;
        RECT 104.155 1.945 104.415 2.205 ;
        RECT 104.475 1.945 104.735 2.205 ;
        RECT 105.275 1.945 105.535 2.205 ;
        RECT 105.595 1.945 105.855 2.205 ;
        RECT 106.395 1.945 106.655 2.205 ;
        RECT 106.715 1.945 106.975 2.205 ;
        RECT 107.515 1.945 107.775 2.205 ;
        RECT 107.835 1.945 108.095 2.205 ;
        RECT 108.635 1.945 108.895 2.205 ;
        RECT 108.955 1.945 109.215 2.205 ;
        RECT 111.645 1.945 111.905 2.205 ;
        RECT 111.965 1.945 112.225 2.205 ;
        RECT 112.765 1.945 113.025 2.205 ;
        RECT 113.085 1.945 113.345 2.205 ;
        RECT 113.885 1.945 114.145 2.205 ;
        RECT 114.205 1.945 114.465 2.205 ;
        RECT 115.005 1.945 115.265 2.205 ;
        RECT 115.325 1.945 115.585 2.205 ;
        RECT 116.125 1.945 116.385 2.205 ;
        RECT 116.445 1.945 116.705 2.205 ;
        RECT 117.245 1.945 117.505 2.205 ;
        RECT 117.565 1.945 117.825 2.205 ;
        RECT 118.365 1.945 118.625 2.205 ;
        RECT 118.685 1.945 118.945 2.205 ;
        RECT 119.485 1.945 119.745 2.205 ;
        RECT 119.805 1.945 120.065 2.205 ;
        RECT 120.605 1.945 120.865 2.205 ;
        RECT 120.925 1.945 121.185 2.205 ;
        RECT 121.725 1.945 121.985 2.205 ;
        RECT 122.045 1.945 122.305 2.205 ;
        RECT 124.735 1.945 124.995 2.205 ;
        RECT 125.055 1.945 125.315 2.205 ;
        RECT 125.855 1.945 126.115 2.205 ;
        RECT 126.175 1.945 126.435 2.205 ;
        RECT 126.975 1.945 127.235 2.205 ;
        RECT 127.295 1.945 127.555 2.205 ;
        RECT 128.095 1.945 128.355 2.205 ;
        RECT 128.415 1.945 128.675 2.205 ;
        RECT 129.215 1.945 129.475 2.205 ;
        RECT 129.535 1.945 129.795 2.205 ;
        RECT 130.335 1.945 130.595 2.205 ;
        RECT 130.655 1.945 130.915 2.205 ;
        RECT 131.455 1.945 131.715 2.205 ;
        RECT 131.775 1.945 132.035 2.205 ;
        RECT 132.575 1.945 132.835 2.205 ;
        RECT 132.895 1.945 133.155 2.205 ;
        RECT 133.695 1.945 133.955 2.205 ;
        RECT 134.015 1.945 134.275 2.205 ;
        RECT 134.815 1.945 135.075 2.205 ;
        RECT 135.135 1.945 135.395 2.205 ;
        RECT 137.825 1.965 138.085 2.225 ;
        RECT 138.145 1.965 138.405 2.225 ;
        RECT 138.945 1.965 139.205 2.225 ;
        RECT 139.265 1.965 139.525 2.225 ;
        RECT 140.065 1.965 140.325 2.225 ;
        RECT 140.385 1.965 140.645 2.225 ;
        RECT 141.185 1.965 141.445 2.225 ;
        RECT 141.505 1.965 141.765 2.225 ;
        RECT 142.305 1.965 142.565 2.225 ;
        RECT 142.625 1.965 142.885 2.225 ;
        RECT 143.425 1.965 143.685 2.225 ;
        RECT 143.745 1.965 144.005 2.225 ;
        RECT 144.545 1.965 144.805 2.225 ;
        RECT 144.865 1.965 145.125 2.225 ;
        RECT 145.665 1.965 145.925 2.225 ;
        RECT 145.985 1.965 146.245 2.225 ;
        RECT 146.785 1.965 147.045 2.225 ;
        RECT 147.105 1.965 147.365 2.225 ;
        RECT 147.905 1.965 148.165 2.225 ;
        RECT 148.225 1.965 148.485 2.225 ;
        RECT 150.915 1.965 151.175 2.225 ;
        RECT 151.235 1.965 151.495 2.225 ;
        RECT 152.035 1.965 152.295 2.225 ;
        RECT 152.355 1.965 152.615 2.225 ;
        RECT 153.155 1.965 153.415 2.225 ;
        RECT 153.475 1.965 153.735 2.225 ;
        RECT 154.275 1.965 154.535 2.225 ;
        RECT 154.595 1.965 154.855 2.225 ;
        RECT 155.395 1.965 155.655 2.225 ;
        RECT 155.715 1.965 155.975 2.225 ;
        RECT 156.515 1.965 156.775 2.225 ;
        RECT 156.835 1.965 157.095 2.225 ;
        RECT 157.635 1.965 157.895 2.225 ;
        RECT 157.955 1.965 158.215 2.225 ;
        RECT 158.755 1.965 159.015 2.225 ;
        RECT 159.075 1.965 159.335 2.225 ;
        RECT 159.875 1.965 160.135 2.225 ;
        RECT 160.195 1.965 160.455 2.225 ;
        RECT 160.995 1.965 161.255 2.225 ;
        RECT 161.315 1.965 161.575 2.225 ;
      LAYER met2 ;
        RECT 6.435 118.280 7.135 118.610 ;
        RECT 6.435 107.390 6.575 118.280 ;
        RECT 6.995 106.920 7.135 118.280 ;
        RECT 7.555 118.280 8.255 118.610 ;
        RECT 7.555 107.390 7.695 118.280 ;
        RECT 8.115 106.920 8.255 118.280 ;
        RECT 8.675 118.280 9.375 118.610 ;
        RECT 8.675 107.390 8.815 118.280 ;
        RECT 9.235 106.920 9.375 118.280 ;
        RECT 9.795 118.280 10.495 118.610 ;
        RECT 9.795 107.390 9.935 118.280 ;
        RECT 10.355 106.920 10.495 118.280 ;
        RECT 10.915 118.280 11.615 118.610 ;
        RECT 10.915 107.390 11.055 118.280 ;
        RECT 11.475 106.920 11.615 118.280 ;
        RECT 12.035 118.280 12.735 118.610 ;
        RECT 12.035 107.390 12.175 118.280 ;
        RECT 12.595 106.920 12.735 118.280 ;
        RECT 13.155 118.280 13.855 118.610 ;
        RECT 13.155 107.390 13.295 118.280 ;
        RECT 13.715 106.920 13.855 118.280 ;
        RECT 14.275 118.280 14.975 118.610 ;
        RECT 14.275 107.390 14.415 118.280 ;
        RECT 14.835 106.920 14.975 118.280 ;
        RECT 15.395 118.280 17.565 118.610 ;
        RECT 19.525 118.280 20.225 118.610 ;
        RECT 15.395 107.390 15.535 118.280 ;
        RECT 15.955 106.920 16.095 118.280 ;
        RECT 16.515 107.390 16.655 118.280 ;
        RECT 17.075 107.390 17.215 118.280 ;
        RECT 19.525 107.390 19.665 118.280 ;
        RECT 20.085 106.920 20.225 118.280 ;
        RECT 20.645 118.280 21.345 118.610 ;
        RECT 20.645 107.390 20.785 118.280 ;
        RECT 21.205 106.920 21.345 118.280 ;
        RECT 21.765 118.280 22.465 118.610 ;
        RECT 21.765 107.390 21.905 118.280 ;
        RECT 22.325 106.920 22.465 118.280 ;
        RECT 22.885 118.280 23.585 118.610 ;
        RECT 22.885 107.390 23.025 118.280 ;
        RECT 23.445 106.920 23.585 118.280 ;
        RECT 24.005 118.280 24.705 118.610 ;
        RECT 24.005 107.390 24.145 118.280 ;
        RECT 24.565 106.920 24.705 118.280 ;
        RECT 25.125 118.280 25.825 118.610 ;
        RECT 25.125 107.390 25.265 118.280 ;
        RECT 25.685 106.920 25.825 118.280 ;
        RECT 26.245 118.280 26.945 118.610 ;
        RECT 26.245 107.390 26.385 118.280 ;
        RECT 26.805 106.920 26.945 118.280 ;
        RECT 27.365 118.280 28.065 118.610 ;
        RECT 27.365 107.390 27.505 118.280 ;
        RECT 27.925 106.920 28.065 118.280 ;
        RECT 28.485 118.280 30.655 118.610 ;
        RECT 28.485 107.390 28.625 118.280 ;
        RECT 29.045 106.920 29.185 118.280 ;
        RECT 29.605 107.390 29.745 118.280 ;
        RECT 30.165 107.390 30.305 118.280 ;
        RECT 32.615 118.260 33.315 118.590 ;
        RECT 32.615 107.370 32.755 118.260 ;
        RECT 33.175 106.900 33.315 118.260 ;
        RECT 33.735 118.260 34.435 118.590 ;
        RECT 33.735 107.370 33.875 118.260 ;
        RECT 34.295 106.900 34.435 118.260 ;
        RECT 34.855 118.260 35.555 118.590 ;
        RECT 34.855 107.370 34.995 118.260 ;
        RECT 35.415 106.900 35.555 118.260 ;
        RECT 35.975 118.260 36.675 118.590 ;
        RECT 35.975 107.370 36.115 118.260 ;
        RECT 36.535 106.900 36.675 118.260 ;
        RECT 37.095 118.260 37.795 118.590 ;
        RECT 37.095 107.370 37.235 118.260 ;
        RECT 37.655 106.900 37.795 118.260 ;
        RECT 38.215 118.260 38.915 118.590 ;
        RECT 38.215 107.370 38.355 118.260 ;
        RECT 38.775 106.900 38.915 118.260 ;
        RECT 39.335 118.260 40.035 118.590 ;
        RECT 39.335 107.370 39.475 118.260 ;
        RECT 39.895 106.900 40.035 118.260 ;
        RECT 40.455 118.260 41.155 118.590 ;
        RECT 40.455 107.370 40.595 118.260 ;
        RECT 41.015 106.900 41.155 118.260 ;
        RECT 41.575 118.260 43.745 118.590 ;
        RECT 45.705 118.260 46.405 118.590 ;
        RECT 41.575 107.370 41.715 118.260 ;
        RECT 42.135 106.900 42.275 118.260 ;
        RECT 42.695 107.370 42.835 118.260 ;
        RECT 43.255 107.370 43.395 118.260 ;
        RECT 45.705 107.370 45.845 118.260 ;
        RECT 46.265 106.900 46.405 118.260 ;
        RECT 46.825 118.260 47.525 118.590 ;
        RECT 46.825 107.370 46.965 118.260 ;
        RECT 47.385 106.900 47.525 118.260 ;
        RECT 47.945 118.260 48.645 118.590 ;
        RECT 47.945 107.370 48.085 118.260 ;
        RECT 48.505 106.900 48.645 118.260 ;
        RECT 49.065 118.260 49.765 118.590 ;
        RECT 49.065 107.370 49.205 118.260 ;
        RECT 49.625 106.900 49.765 118.260 ;
        RECT 50.185 118.260 50.885 118.590 ;
        RECT 50.185 107.370 50.325 118.260 ;
        RECT 50.745 106.900 50.885 118.260 ;
        RECT 51.305 118.260 52.005 118.590 ;
        RECT 51.305 107.370 51.445 118.260 ;
        RECT 51.865 106.900 52.005 118.260 ;
        RECT 52.425 118.260 53.125 118.590 ;
        RECT 52.425 107.370 52.565 118.260 ;
        RECT 52.985 106.900 53.125 118.260 ;
        RECT 53.545 118.260 54.245 118.590 ;
        RECT 53.545 107.370 53.685 118.260 ;
        RECT 54.105 106.900 54.245 118.260 ;
        RECT 54.665 118.260 56.835 118.590 ;
        RECT 58.755 118.260 59.455 118.590 ;
        RECT 54.665 107.370 54.805 118.260 ;
        RECT 55.225 106.900 55.365 118.260 ;
        RECT 55.785 107.370 55.925 118.260 ;
        RECT 56.345 107.370 56.485 118.260 ;
        RECT 58.755 107.370 58.895 118.260 ;
        RECT 59.315 106.900 59.455 118.260 ;
        RECT 59.875 118.260 60.575 118.590 ;
        RECT 59.875 107.370 60.015 118.260 ;
        RECT 60.435 106.900 60.575 118.260 ;
        RECT 60.995 118.260 61.695 118.590 ;
        RECT 60.995 107.370 61.135 118.260 ;
        RECT 61.555 106.900 61.695 118.260 ;
        RECT 62.115 118.260 62.815 118.590 ;
        RECT 62.115 107.370 62.255 118.260 ;
        RECT 62.675 106.900 62.815 118.260 ;
        RECT 63.235 118.260 63.935 118.590 ;
        RECT 63.235 107.370 63.375 118.260 ;
        RECT 63.795 106.900 63.935 118.260 ;
        RECT 64.355 118.260 65.055 118.590 ;
        RECT 64.355 107.370 64.495 118.260 ;
        RECT 64.915 106.900 65.055 118.260 ;
        RECT 65.475 118.260 66.175 118.590 ;
        RECT 65.475 107.370 65.615 118.260 ;
        RECT 66.035 106.900 66.175 118.260 ;
        RECT 66.595 118.260 67.295 118.590 ;
        RECT 66.595 107.370 66.735 118.260 ;
        RECT 67.155 106.900 67.295 118.260 ;
        RECT 67.715 118.260 69.885 118.590 ;
        RECT 71.845 118.260 72.545 118.590 ;
        RECT 67.715 107.370 67.855 118.260 ;
        RECT 68.275 106.900 68.415 118.260 ;
        RECT 68.835 107.370 68.975 118.260 ;
        RECT 69.395 107.370 69.535 118.260 ;
        RECT 71.845 107.370 71.985 118.260 ;
        RECT 72.405 106.900 72.545 118.260 ;
        RECT 72.965 118.260 73.665 118.590 ;
        RECT 72.965 107.370 73.105 118.260 ;
        RECT 73.525 106.900 73.665 118.260 ;
        RECT 74.085 118.260 74.785 118.590 ;
        RECT 74.085 107.370 74.225 118.260 ;
        RECT 74.645 106.900 74.785 118.260 ;
        RECT 75.205 118.260 75.905 118.590 ;
        RECT 75.205 107.370 75.345 118.260 ;
        RECT 75.765 106.900 75.905 118.260 ;
        RECT 76.325 118.260 77.025 118.590 ;
        RECT 76.325 107.370 76.465 118.260 ;
        RECT 76.885 106.900 77.025 118.260 ;
        RECT 77.445 118.260 78.145 118.590 ;
        RECT 77.445 107.370 77.585 118.260 ;
        RECT 78.005 106.900 78.145 118.260 ;
        RECT 78.565 118.260 79.265 118.590 ;
        RECT 78.565 107.370 78.705 118.260 ;
        RECT 79.125 106.900 79.265 118.260 ;
        RECT 79.685 118.260 80.385 118.590 ;
        RECT 79.685 107.370 79.825 118.260 ;
        RECT 80.245 106.900 80.385 118.260 ;
        RECT 80.805 118.260 82.975 118.590 ;
        RECT 80.805 107.370 80.945 118.260 ;
        RECT 81.365 106.900 81.505 118.260 ;
        RECT 81.925 107.370 82.065 118.260 ;
        RECT 82.485 107.370 82.625 118.260 ;
        RECT 84.935 118.240 85.635 118.570 ;
        RECT 84.935 107.350 85.075 118.240 ;
        RECT 85.495 106.880 85.635 118.240 ;
        RECT 86.055 118.240 86.755 118.570 ;
        RECT 86.055 107.350 86.195 118.240 ;
        RECT 86.615 106.880 86.755 118.240 ;
        RECT 87.175 118.240 87.875 118.570 ;
        RECT 87.175 107.350 87.315 118.240 ;
        RECT 87.735 106.880 87.875 118.240 ;
        RECT 88.295 118.240 88.995 118.570 ;
        RECT 88.295 107.350 88.435 118.240 ;
        RECT 88.855 106.880 88.995 118.240 ;
        RECT 89.415 118.240 90.115 118.570 ;
        RECT 89.415 107.350 89.555 118.240 ;
        RECT 89.975 106.880 90.115 118.240 ;
        RECT 90.535 118.240 91.235 118.570 ;
        RECT 90.535 107.350 90.675 118.240 ;
        RECT 91.095 106.880 91.235 118.240 ;
        RECT 91.655 118.240 92.355 118.570 ;
        RECT 91.655 107.350 91.795 118.240 ;
        RECT 92.215 106.880 92.355 118.240 ;
        RECT 92.775 118.240 93.475 118.570 ;
        RECT 92.775 107.350 92.915 118.240 ;
        RECT 93.335 106.880 93.475 118.240 ;
        RECT 93.895 118.240 96.065 118.570 ;
        RECT 98.025 118.240 98.725 118.570 ;
        RECT 93.895 107.350 94.035 118.240 ;
        RECT 94.455 106.880 94.595 118.240 ;
        RECT 95.015 107.350 95.155 118.240 ;
        RECT 95.575 107.350 95.715 118.240 ;
        RECT 98.025 107.350 98.165 118.240 ;
        RECT 98.585 106.880 98.725 118.240 ;
        RECT 99.145 118.240 99.845 118.570 ;
        RECT 99.145 107.350 99.285 118.240 ;
        RECT 99.705 106.880 99.845 118.240 ;
        RECT 100.265 118.240 100.965 118.570 ;
        RECT 100.265 107.350 100.405 118.240 ;
        RECT 100.825 106.880 100.965 118.240 ;
        RECT 101.385 118.240 102.085 118.570 ;
        RECT 101.385 107.350 101.525 118.240 ;
        RECT 101.945 106.880 102.085 118.240 ;
        RECT 102.505 118.240 103.205 118.570 ;
        RECT 102.505 107.350 102.645 118.240 ;
        RECT 103.065 106.880 103.205 118.240 ;
        RECT 103.625 118.240 104.325 118.570 ;
        RECT 103.625 107.350 103.765 118.240 ;
        RECT 104.185 106.880 104.325 118.240 ;
        RECT 104.745 118.240 105.445 118.570 ;
        RECT 104.745 107.350 104.885 118.240 ;
        RECT 105.305 106.880 105.445 118.240 ;
        RECT 105.865 118.240 106.565 118.570 ;
        RECT 105.865 107.350 106.005 118.240 ;
        RECT 106.425 106.880 106.565 118.240 ;
        RECT 106.985 118.240 109.155 118.570 ;
        RECT 111.115 118.240 111.815 118.570 ;
        RECT 106.985 107.350 107.125 118.240 ;
        RECT 107.545 106.880 107.685 118.240 ;
        RECT 108.105 107.350 108.245 118.240 ;
        RECT 108.665 107.350 108.805 118.240 ;
        RECT 111.115 107.350 111.255 118.240 ;
        RECT 111.675 106.880 111.815 118.240 ;
        RECT 112.235 118.240 112.935 118.570 ;
        RECT 112.235 107.350 112.375 118.240 ;
        RECT 112.795 106.880 112.935 118.240 ;
        RECT 113.355 118.240 114.055 118.570 ;
        RECT 113.355 107.350 113.495 118.240 ;
        RECT 113.915 106.880 114.055 118.240 ;
        RECT 114.475 118.240 115.175 118.570 ;
        RECT 114.475 107.350 114.615 118.240 ;
        RECT 115.035 106.880 115.175 118.240 ;
        RECT 115.595 118.240 116.295 118.570 ;
        RECT 115.595 107.350 115.735 118.240 ;
        RECT 116.155 106.880 116.295 118.240 ;
        RECT 116.715 118.240 117.415 118.570 ;
        RECT 116.715 107.350 116.855 118.240 ;
        RECT 117.275 106.880 117.415 118.240 ;
        RECT 117.835 118.240 118.535 118.570 ;
        RECT 117.835 107.350 117.975 118.240 ;
        RECT 118.395 106.880 118.535 118.240 ;
        RECT 118.955 118.240 119.655 118.570 ;
        RECT 118.955 107.350 119.095 118.240 ;
        RECT 119.515 106.880 119.655 118.240 ;
        RECT 120.075 118.240 122.245 118.570 ;
        RECT 124.205 118.240 124.905 118.570 ;
        RECT 120.075 107.350 120.215 118.240 ;
        RECT 120.635 106.880 120.775 118.240 ;
        RECT 121.195 107.350 121.335 118.240 ;
        RECT 121.755 107.350 121.895 118.240 ;
        RECT 124.205 107.350 124.345 118.240 ;
        RECT 124.765 106.880 124.905 118.240 ;
        RECT 125.325 118.240 126.025 118.570 ;
        RECT 125.325 107.350 125.465 118.240 ;
        RECT 125.885 106.880 126.025 118.240 ;
        RECT 126.445 118.240 127.145 118.570 ;
        RECT 126.445 107.350 126.585 118.240 ;
        RECT 127.005 106.880 127.145 118.240 ;
        RECT 127.565 118.240 128.265 118.570 ;
        RECT 127.565 107.350 127.705 118.240 ;
        RECT 128.125 106.880 128.265 118.240 ;
        RECT 128.685 118.240 129.385 118.570 ;
        RECT 128.685 107.350 128.825 118.240 ;
        RECT 129.245 106.880 129.385 118.240 ;
        RECT 129.805 118.240 130.505 118.570 ;
        RECT 129.805 107.350 129.945 118.240 ;
        RECT 130.365 106.880 130.505 118.240 ;
        RECT 130.925 118.240 131.625 118.570 ;
        RECT 130.925 107.350 131.065 118.240 ;
        RECT 131.485 106.880 131.625 118.240 ;
        RECT 132.045 118.240 132.745 118.570 ;
        RECT 132.045 107.350 132.185 118.240 ;
        RECT 132.605 106.880 132.745 118.240 ;
        RECT 133.165 118.240 135.335 118.570 ;
        RECT 133.165 107.350 133.305 118.240 ;
        RECT 133.725 106.880 133.865 118.240 ;
        RECT 134.285 107.350 134.425 118.240 ;
        RECT 134.845 107.350 134.985 118.240 ;
        RECT 137.295 118.220 137.995 118.550 ;
        RECT 137.295 107.330 137.435 118.220 ;
        RECT 137.855 106.860 137.995 118.220 ;
        RECT 138.415 118.220 139.115 118.550 ;
        RECT 138.415 107.330 138.555 118.220 ;
        RECT 138.975 106.860 139.115 118.220 ;
        RECT 139.535 118.220 140.235 118.550 ;
        RECT 139.535 107.330 139.675 118.220 ;
        RECT 140.095 106.860 140.235 118.220 ;
        RECT 140.655 118.220 141.355 118.550 ;
        RECT 140.655 107.330 140.795 118.220 ;
        RECT 141.215 106.860 141.355 118.220 ;
        RECT 141.775 118.220 142.475 118.550 ;
        RECT 141.775 107.330 141.915 118.220 ;
        RECT 142.335 106.860 142.475 118.220 ;
        RECT 142.895 118.220 143.595 118.550 ;
        RECT 142.895 107.330 143.035 118.220 ;
        RECT 143.455 106.860 143.595 118.220 ;
        RECT 144.015 118.220 144.715 118.550 ;
        RECT 144.015 107.330 144.155 118.220 ;
        RECT 144.575 106.860 144.715 118.220 ;
        RECT 145.135 118.220 145.835 118.550 ;
        RECT 145.135 107.330 145.275 118.220 ;
        RECT 145.695 106.860 145.835 118.220 ;
        RECT 146.255 118.220 148.425 118.550 ;
        RECT 150.385 118.220 151.085 118.550 ;
        RECT 146.255 107.330 146.395 118.220 ;
        RECT 146.815 106.860 146.955 118.220 ;
        RECT 147.375 107.330 147.515 118.220 ;
        RECT 147.935 107.330 148.075 118.220 ;
        RECT 150.385 107.330 150.525 118.220 ;
        RECT 150.945 106.860 151.085 118.220 ;
        RECT 151.505 118.220 152.205 118.550 ;
        RECT 151.505 107.330 151.645 118.220 ;
        RECT 152.065 106.860 152.205 118.220 ;
        RECT 152.625 118.220 153.325 118.550 ;
        RECT 152.625 107.330 152.765 118.220 ;
        RECT 153.185 106.860 153.325 118.220 ;
        RECT 153.745 118.220 154.445 118.550 ;
        RECT 153.745 107.330 153.885 118.220 ;
        RECT 154.305 106.860 154.445 118.220 ;
        RECT 154.865 118.220 155.565 118.550 ;
        RECT 154.865 107.330 155.005 118.220 ;
        RECT 155.425 106.860 155.565 118.220 ;
        RECT 155.985 118.220 156.685 118.550 ;
        RECT 155.985 107.330 156.125 118.220 ;
        RECT 156.545 106.860 156.685 118.220 ;
        RECT 157.105 118.220 157.805 118.550 ;
        RECT 157.105 107.330 157.245 118.220 ;
        RECT 157.665 106.860 157.805 118.220 ;
        RECT 158.225 118.220 158.925 118.550 ;
        RECT 158.225 107.330 158.365 118.220 ;
        RECT 158.785 106.860 158.925 118.220 ;
        RECT 159.345 118.220 161.515 118.550 ;
        RECT 159.345 107.330 159.485 118.220 ;
        RECT 159.905 106.860 160.045 118.220 ;
        RECT 160.465 107.330 160.605 118.220 ;
        RECT 161.025 107.330 161.165 118.220 ;
        RECT 6.465 93.840 6.605 104.730 ;
        RECT 7.025 93.840 7.165 105.200 ;
        RECT 6.465 93.510 7.165 93.840 ;
        RECT 7.585 93.840 7.725 104.730 ;
        RECT 8.145 93.840 8.285 105.200 ;
        RECT 7.585 93.510 8.285 93.840 ;
        RECT 8.705 93.840 8.845 104.730 ;
        RECT 9.265 93.840 9.405 105.200 ;
        RECT 8.705 93.510 9.405 93.840 ;
        RECT 9.825 93.840 9.965 104.730 ;
        RECT 10.385 93.840 10.525 105.200 ;
        RECT 9.825 93.510 10.525 93.840 ;
        RECT 10.945 93.840 11.085 104.730 ;
        RECT 11.505 93.840 11.645 105.200 ;
        RECT 10.945 93.510 11.645 93.840 ;
        RECT 12.065 93.840 12.205 104.730 ;
        RECT 12.625 93.840 12.765 105.200 ;
        RECT 12.065 93.510 12.765 93.840 ;
        RECT 13.185 93.840 13.325 104.730 ;
        RECT 13.745 93.840 13.885 105.200 ;
        RECT 13.185 93.510 13.885 93.840 ;
        RECT 14.305 93.840 14.445 104.730 ;
        RECT 14.865 93.840 15.005 105.200 ;
        RECT 14.305 93.510 15.005 93.840 ;
        RECT 15.425 93.840 15.565 104.730 ;
        RECT 15.985 93.840 16.125 105.200 ;
        RECT 16.545 93.840 16.685 104.730 ;
        RECT 17.105 93.840 17.245 104.730 ;
        RECT 19.555 93.840 19.695 104.730 ;
        RECT 20.115 93.840 20.255 105.200 ;
        RECT 15.425 93.510 17.595 93.840 ;
        RECT 19.555 93.510 20.255 93.840 ;
        RECT 20.675 93.840 20.815 104.730 ;
        RECT 21.235 93.840 21.375 105.200 ;
        RECT 20.675 93.510 21.375 93.840 ;
        RECT 21.795 93.840 21.935 104.730 ;
        RECT 22.355 93.840 22.495 105.200 ;
        RECT 21.795 93.510 22.495 93.840 ;
        RECT 22.915 93.840 23.055 104.730 ;
        RECT 23.475 93.840 23.615 105.200 ;
        RECT 22.915 93.510 23.615 93.840 ;
        RECT 24.035 93.840 24.175 104.730 ;
        RECT 24.595 93.840 24.735 105.200 ;
        RECT 24.035 93.510 24.735 93.840 ;
        RECT 25.155 93.840 25.295 104.730 ;
        RECT 25.715 93.840 25.855 105.200 ;
        RECT 25.155 93.510 25.855 93.840 ;
        RECT 26.275 93.840 26.415 104.730 ;
        RECT 26.835 93.840 26.975 105.200 ;
        RECT 26.275 93.510 26.975 93.840 ;
        RECT 27.395 93.840 27.535 104.730 ;
        RECT 27.955 93.840 28.095 105.200 ;
        RECT 27.395 93.510 28.095 93.840 ;
        RECT 28.515 93.840 28.655 104.730 ;
        RECT 29.075 93.840 29.215 105.200 ;
        RECT 29.635 93.840 29.775 104.730 ;
        RECT 30.195 93.840 30.335 104.730 ;
        RECT 32.645 93.860 32.785 104.750 ;
        RECT 33.205 93.860 33.345 105.220 ;
        RECT 28.515 93.510 30.685 93.840 ;
        RECT 32.645 93.530 33.345 93.860 ;
        RECT 33.765 93.860 33.905 104.750 ;
        RECT 34.325 93.860 34.465 105.220 ;
        RECT 33.765 93.530 34.465 93.860 ;
        RECT 34.885 93.860 35.025 104.750 ;
        RECT 35.445 93.860 35.585 105.220 ;
        RECT 34.885 93.530 35.585 93.860 ;
        RECT 36.005 93.860 36.145 104.750 ;
        RECT 36.565 93.860 36.705 105.220 ;
        RECT 36.005 93.530 36.705 93.860 ;
        RECT 37.125 93.860 37.265 104.750 ;
        RECT 37.685 93.860 37.825 105.220 ;
        RECT 37.125 93.530 37.825 93.860 ;
        RECT 38.245 93.860 38.385 104.750 ;
        RECT 38.805 93.860 38.945 105.220 ;
        RECT 38.245 93.530 38.945 93.860 ;
        RECT 39.365 93.860 39.505 104.750 ;
        RECT 39.925 93.860 40.065 105.220 ;
        RECT 39.365 93.530 40.065 93.860 ;
        RECT 40.485 93.860 40.625 104.750 ;
        RECT 41.045 93.860 41.185 105.220 ;
        RECT 40.485 93.530 41.185 93.860 ;
        RECT 41.605 93.860 41.745 104.750 ;
        RECT 42.165 93.860 42.305 105.220 ;
        RECT 42.725 93.860 42.865 104.750 ;
        RECT 43.285 93.860 43.425 104.750 ;
        RECT 45.735 93.860 45.875 104.750 ;
        RECT 46.295 93.860 46.435 105.220 ;
        RECT 41.605 93.530 43.775 93.860 ;
        RECT 45.735 93.530 46.435 93.860 ;
        RECT 46.855 93.860 46.995 104.750 ;
        RECT 47.415 93.860 47.555 105.220 ;
        RECT 46.855 93.530 47.555 93.860 ;
        RECT 47.975 93.860 48.115 104.750 ;
        RECT 48.535 93.860 48.675 105.220 ;
        RECT 47.975 93.530 48.675 93.860 ;
        RECT 49.095 93.860 49.235 104.750 ;
        RECT 49.655 93.860 49.795 105.220 ;
        RECT 49.095 93.530 49.795 93.860 ;
        RECT 50.215 93.860 50.355 104.750 ;
        RECT 50.775 93.860 50.915 105.220 ;
        RECT 50.215 93.530 50.915 93.860 ;
        RECT 51.335 93.860 51.475 104.750 ;
        RECT 51.895 93.860 52.035 105.220 ;
        RECT 51.335 93.530 52.035 93.860 ;
        RECT 52.455 93.860 52.595 104.750 ;
        RECT 53.015 93.860 53.155 105.220 ;
        RECT 52.455 93.530 53.155 93.860 ;
        RECT 53.575 93.860 53.715 104.750 ;
        RECT 54.135 93.860 54.275 105.220 ;
        RECT 53.575 93.530 54.275 93.860 ;
        RECT 54.695 93.860 54.835 104.750 ;
        RECT 55.255 93.860 55.395 105.220 ;
        RECT 55.815 93.860 55.955 104.750 ;
        RECT 56.375 93.860 56.515 104.750 ;
        RECT 58.785 93.860 58.925 104.750 ;
        RECT 59.345 93.860 59.485 105.220 ;
        RECT 54.695 93.530 56.865 93.860 ;
        RECT 58.785 93.530 59.485 93.860 ;
        RECT 59.905 93.860 60.045 104.750 ;
        RECT 60.465 93.860 60.605 105.220 ;
        RECT 59.905 93.530 60.605 93.860 ;
        RECT 61.025 93.860 61.165 104.750 ;
        RECT 61.585 93.860 61.725 105.220 ;
        RECT 61.025 93.530 61.725 93.860 ;
        RECT 62.145 93.860 62.285 104.750 ;
        RECT 62.705 93.860 62.845 105.220 ;
        RECT 62.145 93.530 62.845 93.860 ;
        RECT 63.265 93.860 63.405 104.750 ;
        RECT 63.825 93.860 63.965 105.220 ;
        RECT 63.265 93.530 63.965 93.860 ;
        RECT 64.385 93.860 64.525 104.750 ;
        RECT 64.945 93.860 65.085 105.220 ;
        RECT 64.385 93.530 65.085 93.860 ;
        RECT 65.505 93.860 65.645 104.750 ;
        RECT 66.065 93.860 66.205 105.220 ;
        RECT 65.505 93.530 66.205 93.860 ;
        RECT 66.625 93.860 66.765 104.750 ;
        RECT 67.185 93.860 67.325 105.220 ;
        RECT 66.625 93.530 67.325 93.860 ;
        RECT 67.745 93.860 67.885 104.750 ;
        RECT 68.305 93.860 68.445 105.220 ;
        RECT 68.865 93.860 69.005 104.750 ;
        RECT 69.425 93.860 69.565 104.750 ;
        RECT 71.875 93.860 72.015 104.750 ;
        RECT 72.435 93.860 72.575 105.220 ;
        RECT 67.745 93.530 69.915 93.860 ;
        RECT 71.875 93.530 72.575 93.860 ;
        RECT 72.995 93.860 73.135 104.750 ;
        RECT 73.555 93.860 73.695 105.220 ;
        RECT 72.995 93.530 73.695 93.860 ;
        RECT 74.115 93.860 74.255 104.750 ;
        RECT 74.675 93.860 74.815 105.220 ;
        RECT 74.115 93.530 74.815 93.860 ;
        RECT 75.235 93.860 75.375 104.750 ;
        RECT 75.795 93.860 75.935 105.220 ;
        RECT 75.235 93.530 75.935 93.860 ;
        RECT 76.355 93.860 76.495 104.750 ;
        RECT 76.915 93.860 77.055 105.220 ;
        RECT 76.355 93.530 77.055 93.860 ;
        RECT 77.475 93.860 77.615 104.750 ;
        RECT 78.035 93.860 78.175 105.220 ;
        RECT 77.475 93.530 78.175 93.860 ;
        RECT 78.595 93.860 78.735 104.750 ;
        RECT 79.155 93.860 79.295 105.220 ;
        RECT 78.595 93.530 79.295 93.860 ;
        RECT 79.715 93.860 79.855 104.750 ;
        RECT 80.275 93.860 80.415 105.220 ;
        RECT 79.715 93.530 80.415 93.860 ;
        RECT 80.835 93.860 80.975 104.750 ;
        RECT 81.395 93.860 81.535 105.220 ;
        RECT 81.955 93.860 82.095 104.750 ;
        RECT 82.515 93.860 82.655 104.750 ;
        RECT 84.965 93.880 85.105 104.770 ;
        RECT 85.525 93.880 85.665 105.240 ;
        RECT 80.835 93.530 83.005 93.860 ;
        RECT 84.965 93.550 85.665 93.880 ;
        RECT 86.085 93.880 86.225 104.770 ;
        RECT 86.645 93.880 86.785 105.240 ;
        RECT 86.085 93.550 86.785 93.880 ;
        RECT 87.205 93.880 87.345 104.770 ;
        RECT 87.765 93.880 87.905 105.240 ;
        RECT 87.205 93.550 87.905 93.880 ;
        RECT 88.325 93.880 88.465 104.770 ;
        RECT 88.885 93.880 89.025 105.240 ;
        RECT 88.325 93.550 89.025 93.880 ;
        RECT 89.445 93.880 89.585 104.770 ;
        RECT 90.005 93.880 90.145 105.240 ;
        RECT 89.445 93.550 90.145 93.880 ;
        RECT 90.565 93.880 90.705 104.770 ;
        RECT 91.125 93.880 91.265 105.240 ;
        RECT 90.565 93.550 91.265 93.880 ;
        RECT 91.685 93.880 91.825 104.770 ;
        RECT 92.245 93.880 92.385 105.240 ;
        RECT 91.685 93.550 92.385 93.880 ;
        RECT 92.805 93.880 92.945 104.770 ;
        RECT 93.365 93.880 93.505 105.240 ;
        RECT 92.805 93.550 93.505 93.880 ;
        RECT 93.925 93.880 94.065 104.770 ;
        RECT 94.485 93.880 94.625 105.240 ;
        RECT 95.045 93.880 95.185 104.770 ;
        RECT 95.605 93.880 95.745 104.770 ;
        RECT 98.055 93.880 98.195 104.770 ;
        RECT 98.615 93.880 98.755 105.240 ;
        RECT 93.925 93.550 96.095 93.880 ;
        RECT 98.055 93.550 98.755 93.880 ;
        RECT 99.175 93.880 99.315 104.770 ;
        RECT 99.735 93.880 99.875 105.240 ;
        RECT 99.175 93.550 99.875 93.880 ;
        RECT 100.295 93.880 100.435 104.770 ;
        RECT 100.855 93.880 100.995 105.240 ;
        RECT 100.295 93.550 100.995 93.880 ;
        RECT 101.415 93.880 101.555 104.770 ;
        RECT 101.975 93.880 102.115 105.240 ;
        RECT 101.415 93.550 102.115 93.880 ;
        RECT 102.535 93.880 102.675 104.770 ;
        RECT 103.095 93.880 103.235 105.240 ;
        RECT 102.535 93.550 103.235 93.880 ;
        RECT 103.655 93.880 103.795 104.770 ;
        RECT 104.215 93.880 104.355 105.240 ;
        RECT 103.655 93.550 104.355 93.880 ;
        RECT 104.775 93.880 104.915 104.770 ;
        RECT 105.335 93.880 105.475 105.240 ;
        RECT 104.775 93.550 105.475 93.880 ;
        RECT 105.895 93.880 106.035 104.770 ;
        RECT 106.455 93.880 106.595 105.240 ;
        RECT 105.895 93.550 106.595 93.880 ;
        RECT 107.015 93.880 107.155 104.770 ;
        RECT 107.575 93.880 107.715 105.240 ;
        RECT 108.135 93.880 108.275 104.770 ;
        RECT 108.695 93.880 108.835 104.770 ;
        RECT 111.145 93.880 111.285 104.770 ;
        RECT 111.705 93.880 111.845 105.240 ;
        RECT 107.015 93.550 109.185 93.880 ;
        RECT 111.145 93.550 111.845 93.880 ;
        RECT 112.265 93.880 112.405 104.770 ;
        RECT 112.825 93.880 112.965 105.240 ;
        RECT 112.265 93.550 112.965 93.880 ;
        RECT 113.385 93.880 113.525 104.770 ;
        RECT 113.945 93.880 114.085 105.240 ;
        RECT 113.385 93.550 114.085 93.880 ;
        RECT 114.505 93.880 114.645 104.770 ;
        RECT 115.065 93.880 115.205 105.240 ;
        RECT 114.505 93.550 115.205 93.880 ;
        RECT 115.625 93.880 115.765 104.770 ;
        RECT 116.185 93.880 116.325 105.240 ;
        RECT 115.625 93.550 116.325 93.880 ;
        RECT 116.745 93.880 116.885 104.770 ;
        RECT 117.305 93.880 117.445 105.240 ;
        RECT 116.745 93.550 117.445 93.880 ;
        RECT 117.865 93.880 118.005 104.770 ;
        RECT 118.425 93.880 118.565 105.240 ;
        RECT 117.865 93.550 118.565 93.880 ;
        RECT 118.985 93.880 119.125 104.770 ;
        RECT 119.545 93.880 119.685 105.240 ;
        RECT 118.985 93.550 119.685 93.880 ;
        RECT 120.105 93.880 120.245 104.770 ;
        RECT 120.665 93.880 120.805 105.240 ;
        RECT 121.225 93.880 121.365 104.770 ;
        RECT 121.785 93.880 121.925 104.770 ;
        RECT 124.235 93.880 124.375 104.770 ;
        RECT 124.795 93.880 124.935 105.240 ;
        RECT 120.105 93.550 122.275 93.880 ;
        RECT 124.235 93.550 124.935 93.880 ;
        RECT 125.355 93.880 125.495 104.770 ;
        RECT 125.915 93.880 126.055 105.240 ;
        RECT 125.355 93.550 126.055 93.880 ;
        RECT 126.475 93.880 126.615 104.770 ;
        RECT 127.035 93.880 127.175 105.240 ;
        RECT 126.475 93.550 127.175 93.880 ;
        RECT 127.595 93.880 127.735 104.770 ;
        RECT 128.155 93.880 128.295 105.240 ;
        RECT 127.595 93.550 128.295 93.880 ;
        RECT 128.715 93.880 128.855 104.770 ;
        RECT 129.275 93.880 129.415 105.240 ;
        RECT 128.715 93.550 129.415 93.880 ;
        RECT 129.835 93.880 129.975 104.770 ;
        RECT 130.395 93.880 130.535 105.240 ;
        RECT 129.835 93.550 130.535 93.880 ;
        RECT 130.955 93.880 131.095 104.770 ;
        RECT 131.515 93.880 131.655 105.240 ;
        RECT 130.955 93.550 131.655 93.880 ;
        RECT 132.075 93.880 132.215 104.770 ;
        RECT 132.635 93.880 132.775 105.240 ;
        RECT 132.075 93.550 132.775 93.880 ;
        RECT 133.195 93.880 133.335 104.770 ;
        RECT 133.755 93.880 133.895 105.240 ;
        RECT 134.315 93.880 134.455 104.770 ;
        RECT 134.875 93.880 135.015 104.770 ;
        RECT 137.325 93.900 137.465 104.790 ;
        RECT 137.885 93.900 138.025 105.260 ;
        RECT 133.195 93.550 135.365 93.880 ;
        RECT 137.325 93.570 138.025 93.900 ;
        RECT 138.445 93.900 138.585 104.790 ;
        RECT 139.005 93.900 139.145 105.260 ;
        RECT 138.445 93.570 139.145 93.900 ;
        RECT 139.565 93.900 139.705 104.790 ;
        RECT 140.125 93.900 140.265 105.260 ;
        RECT 139.565 93.570 140.265 93.900 ;
        RECT 140.685 93.900 140.825 104.790 ;
        RECT 141.245 93.900 141.385 105.260 ;
        RECT 140.685 93.570 141.385 93.900 ;
        RECT 141.805 93.900 141.945 104.790 ;
        RECT 142.365 93.900 142.505 105.260 ;
        RECT 141.805 93.570 142.505 93.900 ;
        RECT 142.925 93.900 143.065 104.790 ;
        RECT 143.485 93.900 143.625 105.260 ;
        RECT 142.925 93.570 143.625 93.900 ;
        RECT 144.045 93.900 144.185 104.790 ;
        RECT 144.605 93.900 144.745 105.260 ;
        RECT 144.045 93.570 144.745 93.900 ;
        RECT 145.165 93.900 145.305 104.790 ;
        RECT 145.725 93.900 145.865 105.260 ;
        RECT 145.165 93.570 145.865 93.900 ;
        RECT 146.285 93.900 146.425 104.790 ;
        RECT 146.845 93.900 146.985 105.260 ;
        RECT 147.405 93.900 147.545 104.790 ;
        RECT 147.965 93.900 148.105 104.790 ;
        RECT 150.415 93.900 150.555 104.790 ;
        RECT 150.975 93.900 151.115 105.260 ;
        RECT 146.285 93.570 148.455 93.900 ;
        RECT 150.415 93.570 151.115 93.900 ;
        RECT 151.535 93.900 151.675 104.790 ;
        RECT 152.095 93.900 152.235 105.260 ;
        RECT 151.535 93.570 152.235 93.900 ;
        RECT 152.655 93.900 152.795 104.790 ;
        RECT 153.215 93.900 153.355 105.260 ;
        RECT 152.655 93.570 153.355 93.900 ;
        RECT 153.775 93.900 153.915 104.790 ;
        RECT 154.335 93.900 154.475 105.260 ;
        RECT 153.775 93.570 154.475 93.900 ;
        RECT 154.895 93.900 155.035 104.790 ;
        RECT 155.455 93.900 155.595 105.260 ;
        RECT 154.895 93.570 155.595 93.900 ;
        RECT 156.015 93.900 156.155 104.790 ;
        RECT 156.575 93.900 156.715 105.260 ;
        RECT 156.015 93.570 156.715 93.900 ;
        RECT 157.135 93.900 157.275 104.790 ;
        RECT 157.695 93.900 157.835 105.260 ;
        RECT 157.135 93.570 157.835 93.900 ;
        RECT 158.255 93.900 158.395 104.790 ;
        RECT 158.815 93.900 158.955 105.260 ;
        RECT 158.255 93.570 158.955 93.900 ;
        RECT 159.375 93.900 159.515 104.790 ;
        RECT 159.935 93.900 160.075 105.260 ;
        RECT 160.495 93.900 160.635 104.790 ;
        RECT 161.055 93.900 161.195 104.790 ;
        RECT 159.375 93.570 161.545 93.900 ;
        RECT 167.325 89.940 167.800 89.970 ;
        RECT 151.215 89.440 151.475 89.760 ;
        RECT 167.280 89.465 167.845 89.940 ;
        RECT 1.935 88.345 2.495 88.815 ;
        RECT 148.750 88.445 149.070 88.490 ;
        RECT 151.260 88.445 151.425 89.440 ;
        RECT 167.325 89.435 167.800 89.465 ;
        RECT 148.750 88.280 151.425 88.445 ;
        RECT 148.750 88.275 151.205 88.280 ;
        RECT 148.750 88.230 149.070 88.275 ;
        RECT 178.030 55.790 178.430 65.720 ;
        RECT 1.940 33.685 2.410 33.730 ;
        RECT 1.910 33.215 2.440 33.685 ;
        RECT 1.940 33.170 2.410 33.215 ;
        RECT 166.065 30.385 166.540 30.430 ;
        RECT 166.035 29.910 166.570 30.385 ;
        RECT 166.065 29.865 166.540 29.910 ;
        RECT 6.875 26.640 7.575 26.970 ;
        RECT 6.875 15.750 7.015 26.640 ;
        RECT 7.435 15.280 7.575 26.640 ;
        RECT 7.995 26.640 8.695 26.970 ;
        RECT 7.995 15.750 8.135 26.640 ;
        RECT 8.555 15.280 8.695 26.640 ;
        RECT 9.115 26.640 9.815 26.970 ;
        RECT 9.115 15.750 9.255 26.640 ;
        RECT 9.675 15.280 9.815 26.640 ;
        RECT 10.235 26.640 10.935 26.970 ;
        RECT 10.235 15.750 10.375 26.640 ;
        RECT 10.795 15.280 10.935 26.640 ;
        RECT 11.355 26.640 12.055 26.970 ;
        RECT 11.355 15.750 11.495 26.640 ;
        RECT 11.915 15.280 12.055 26.640 ;
        RECT 12.475 26.640 13.175 26.970 ;
        RECT 12.475 15.750 12.615 26.640 ;
        RECT 13.035 15.280 13.175 26.640 ;
        RECT 13.595 26.640 14.295 26.970 ;
        RECT 13.595 15.750 13.735 26.640 ;
        RECT 14.155 15.280 14.295 26.640 ;
        RECT 14.715 26.640 15.415 26.970 ;
        RECT 14.715 15.750 14.855 26.640 ;
        RECT 15.275 15.280 15.415 26.640 ;
        RECT 15.835 26.640 18.005 26.970 ;
        RECT 19.965 26.640 20.665 26.970 ;
        RECT 15.835 15.750 15.975 26.640 ;
        RECT 16.395 15.280 16.535 26.640 ;
        RECT 16.955 15.750 17.095 26.640 ;
        RECT 17.515 15.750 17.655 26.640 ;
        RECT 19.965 15.750 20.105 26.640 ;
        RECT 20.525 15.280 20.665 26.640 ;
        RECT 21.085 26.640 21.785 26.970 ;
        RECT 21.085 15.750 21.225 26.640 ;
        RECT 21.645 15.280 21.785 26.640 ;
        RECT 22.205 26.640 22.905 26.970 ;
        RECT 22.205 15.750 22.345 26.640 ;
        RECT 22.765 15.280 22.905 26.640 ;
        RECT 23.325 26.640 24.025 26.970 ;
        RECT 23.325 15.750 23.465 26.640 ;
        RECT 23.885 15.280 24.025 26.640 ;
        RECT 24.445 26.640 25.145 26.970 ;
        RECT 24.445 15.750 24.585 26.640 ;
        RECT 25.005 15.280 25.145 26.640 ;
        RECT 25.565 26.640 26.265 26.970 ;
        RECT 25.565 15.750 25.705 26.640 ;
        RECT 26.125 15.280 26.265 26.640 ;
        RECT 26.685 26.640 27.385 26.970 ;
        RECT 26.685 15.750 26.825 26.640 ;
        RECT 27.245 15.280 27.385 26.640 ;
        RECT 27.805 26.640 28.505 26.970 ;
        RECT 27.805 15.750 27.945 26.640 ;
        RECT 28.365 15.280 28.505 26.640 ;
        RECT 28.925 26.640 31.095 26.970 ;
        RECT 28.925 15.750 29.065 26.640 ;
        RECT 29.485 15.280 29.625 26.640 ;
        RECT 30.045 15.750 30.185 26.640 ;
        RECT 30.605 15.750 30.745 26.640 ;
        RECT 33.055 26.620 33.755 26.950 ;
        RECT 33.055 15.730 33.195 26.620 ;
        RECT 33.615 15.260 33.755 26.620 ;
        RECT 34.175 26.620 34.875 26.950 ;
        RECT 34.175 15.730 34.315 26.620 ;
        RECT 34.735 15.260 34.875 26.620 ;
        RECT 35.295 26.620 35.995 26.950 ;
        RECT 35.295 15.730 35.435 26.620 ;
        RECT 35.855 15.260 35.995 26.620 ;
        RECT 36.415 26.620 37.115 26.950 ;
        RECT 36.415 15.730 36.555 26.620 ;
        RECT 36.975 15.260 37.115 26.620 ;
        RECT 37.535 26.620 38.235 26.950 ;
        RECT 37.535 15.730 37.675 26.620 ;
        RECT 38.095 15.260 38.235 26.620 ;
        RECT 38.655 26.620 39.355 26.950 ;
        RECT 38.655 15.730 38.795 26.620 ;
        RECT 39.215 15.260 39.355 26.620 ;
        RECT 39.775 26.620 40.475 26.950 ;
        RECT 39.775 15.730 39.915 26.620 ;
        RECT 40.335 15.260 40.475 26.620 ;
        RECT 40.895 26.620 41.595 26.950 ;
        RECT 40.895 15.730 41.035 26.620 ;
        RECT 41.455 15.260 41.595 26.620 ;
        RECT 42.015 26.620 44.185 26.950 ;
        RECT 46.145 26.620 46.845 26.950 ;
        RECT 42.015 15.730 42.155 26.620 ;
        RECT 42.575 15.260 42.715 26.620 ;
        RECT 43.135 15.730 43.275 26.620 ;
        RECT 43.695 15.730 43.835 26.620 ;
        RECT 46.145 15.730 46.285 26.620 ;
        RECT 46.705 15.260 46.845 26.620 ;
        RECT 47.265 26.620 47.965 26.950 ;
        RECT 47.265 15.730 47.405 26.620 ;
        RECT 47.825 15.260 47.965 26.620 ;
        RECT 48.385 26.620 49.085 26.950 ;
        RECT 48.385 15.730 48.525 26.620 ;
        RECT 48.945 15.260 49.085 26.620 ;
        RECT 49.505 26.620 50.205 26.950 ;
        RECT 49.505 15.730 49.645 26.620 ;
        RECT 50.065 15.260 50.205 26.620 ;
        RECT 50.625 26.620 51.325 26.950 ;
        RECT 50.625 15.730 50.765 26.620 ;
        RECT 51.185 15.260 51.325 26.620 ;
        RECT 51.745 26.620 52.445 26.950 ;
        RECT 51.745 15.730 51.885 26.620 ;
        RECT 52.305 15.260 52.445 26.620 ;
        RECT 52.865 26.620 53.565 26.950 ;
        RECT 52.865 15.730 53.005 26.620 ;
        RECT 53.425 15.260 53.565 26.620 ;
        RECT 53.985 26.620 54.685 26.950 ;
        RECT 53.985 15.730 54.125 26.620 ;
        RECT 54.545 15.260 54.685 26.620 ;
        RECT 55.105 26.620 57.275 26.950 ;
        RECT 59.195 26.620 59.895 26.950 ;
        RECT 55.105 15.730 55.245 26.620 ;
        RECT 55.665 15.260 55.805 26.620 ;
        RECT 56.225 15.730 56.365 26.620 ;
        RECT 56.785 15.730 56.925 26.620 ;
        RECT 59.195 15.730 59.335 26.620 ;
        RECT 59.755 15.260 59.895 26.620 ;
        RECT 60.315 26.620 61.015 26.950 ;
        RECT 60.315 15.730 60.455 26.620 ;
        RECT 60.875 15.260 61.015 26.620 ;
        RECT 61.435 26.620 62.135 26.950 ;
        RECT 61.435 15.730 61.575 26.620 ;
        RECT 61.995 15.260 62.135 26.620 ;
        RECT 62.555 26.620 63.255 26.950 ;
        RECT 62.555 15.730 62.695 26.620 ;
        RECT 63.115 15.260 63.255 26.620 ;
        RECT 63.675 26.620 64.375 26.950 ;
        RECT 63.675 15.730 63.815 26.620 ;
        RECT 64.235 15.260 64.375 26.620 ;
        RECT 64.795 26.620 65.495 26.950 ;
        RECT 64.795 15.730 64.935 26.620 ;
        RECT 65.355 15.260 65.495 26.620 ;
        RECT 65.915 26.620 66.615 26.950 ;
        RECT 65.915 15.730 66.055 26.620 ;
        RECT 66.475 15.260 66.615 26.620 ;
        RECT 67.035 26.620 67.735 26.950 ;
        RECT 67.035 15.730 67.175 26.620 ;
        RECT 67.595 15.260 67.735 26.620 ;
        RECT 68.155 26.620 70.325 26.950 ;
        RECT 72.285 26.620 72.985 26.950 ;
        RECT 68.155 15.730 68.295 26.620 ;
        RECT 68.715 15.260 68.855 26.620 ;
        RECT 69.275 15.730 69.415 26.620 ;
        RECT 69.835 15.730 69.975 26.620 ;
        RECT 72.285 15.730 72.425 26.620 ;
        RECT 72.845 15.260 72.985 26.620 ;
        RECT 73.405 26.620 74.105 26.950 ;
        RECT 73.405 15.730 73.545 26.620 ;
        RECT 73.965 15.260 74.105 26.620 ;
        RECT 74.525 26.620 75.225 26.950 ;
        RECT 74.525 15.730 74.665 26.620 ;
        RECT 75.085 15.260 75.225 26.620 ;
        RECT 75.645 26.620 76.345 26.950 ;
        RECT 75.645 15.730 75.785 26.620 ;
        RECT 76.205 15.260 76.345 26.620 ;
        RECT 76.765 26.620 77.465 26.950 ;
        RECT 76.765 15.730 76.905 26.620 ;
        RECT 77.325 15.260 77.465 26.620 ;
        RECT 77.885 26.620 78.585 26.950 ;
        RECT 77.885 15.730 78.025 26.620 ;
        RECT 78.445 15.260 78.585 26.620 ;
        RECT 79.005 26.620 79.705 26.950 ;
        RECT 79.005 15.730 79.145 26.620 ;
        RECT 79.565 15.260 79.705 26.620 ;
        RECT 80.125 26.620 80.825 26.950 ;
        RECT 80.125 15.730 80.265 26.620 ;
        RECT 80.685 15.260 80.825 26.620 ;
        RECT 81.245 26.620 83.415 26.950 ;
        RECT 81.245 15.730 81.385 26.620 ;
        RECT 81.805 15.260 81.945 26.620 ;
        RECT 82.365 15.730 82.505 26.620 ;
        RECT 82.925 15.730 83.065 26.620 ;
        RECT 85.375 26.600 86.075 26.930 ;
        RECT 85.375 15.710 85.515 26.600 ;
        RECT 85.935 15.240 86.075 26.600 ;
        RECT 86.495 26.600 87.195 26.930 ;
        RECT 86.495 15.710 86.635 26.600 ;
        RECT 87.055 15.240 87.195 26.600 ;
        RECT 87.615 26.600 88.315 26.930 ;
        RECT 87.615 15.710 87.755 26.600 ;
        RECT 88.175 15.240 88.315 26.600 ;
        RECT 88.735 26.600 89.435 26.930 ;
        RECT 88.735 15.710 88.875 26.600 ;
        RECT 89.295 15.240 89.435 26.600 ;
        RECT 89.855 26.600 90.555 26.930 ;
        RECT 89.855 15.710 89.995 26.600 ;
        RECT 90.415 15.240 90.555 26.600 ;
        RECT 90.975 26.600 91.675 26.930 ;
        RECT 90.975 15.710 91.115 26.600 ;
        RECT 91.535 15.240 91.675 26.600 ;
        RECT 92.095 26.600 92.795 26.930 ;
        RECT 92.095 15.710 92.235 26.600 ;
        RECT 92.655 15.240 92.795 26.600 ;
        RECT 93.215 26.600 93.915 26.930 ;
        RECT 93.215 15.710 93.355 26.600 ;
        RECT 93.775 15.240 93.915 26.600 ;
        RECT 94.335 26.600 96.505 26.930 ;
        RECT 98.465 26.600 99.165 26.930 ;
        RECT 94.335 15.710 94.475 26.600 ;
        RECT 94.895 15.240 95.035 26.600 ;
        RECT 95.455 15.710 95.595 26.600 ;
        RECT 96.015 15.710 96.155 26.600 ;
        RECT 98.465 15.710 98.605 26.600 ;
        RECT 99.025 15.240 99.165 26.600 ;
        RECT 99.585 26.600 100.285 26.930 ;
        RECT 99.585 15.710 99.725 26.600 ;
        RECT 100.145 15.240 100.285 26.600 ;
        RECT 100.705 26.600 101.405 26.930 ;
        RECT 100.705 15.710 100.845 26.600 ;
        RECT 101.265 15.240 101.405 26.600 ;
        RECT 101.825 26.600 102.525 26.930 ;
        RECT 101.825 15.710 101.965 26.600 ;
        RECT 102.385 15.240 102.525 26.600 ;
        RECT 102.945 26.600 103.645 26.930 ;
        RECT 102.945 15.710 103.085 26.600 ;
        RECT 103.505 15.240 103.645 26.600 ;
        RECT 104.065 26.600 104.765 26.930 ;
        RECT 104.065 15.710 104.205 26.600 ;
        RECT 104.625 15.240 104.765 26.600 ;
        RECT 105.185 26.600 105.885 26.930 ;
        RECT 105.185 15.710 105.325 26.600 ;
        RECT 105.745 15.240 105.885 26.600 ;
        RECT 106.305 26.600 107.005 26.930 ;
        RECT 106.305 15.710 106.445 26.600 ;
        RECT 106.865 15.240 107.005 26.600 ;
        RECT 107.425 26.600 109.595 26.930 ;
        RECT 111.555 26.600 112.255 26.930 ;
        RECT 107.425 15.710 107.565 26.600 ;
        RECT 107.985 15.240 108.125 26.600 ;
        RECT 108.545 15.710 108.685 26.600 ;
        RECT 109.105 15.710 109.245 26.600 ;
        RECT 111.555 15.710 111.695 26.600 ;
        RECT 112.115 15.240 112.255 26.600 ;
        RECT 112.675 26.600 113.375 26.930 ;
        RECT 112.675 15.710 112.815 26.600 ;
        RECT 113.235 15.240 113.375 26.600 ;
        RECT 113.795 26.600 114.495 26.930 ;
        RECT 113.795 15.710 113.935 26.600 ;
        RECT 114.355 15.240 114.495 26.600 ;
        RECT 114.915 26.600 115.615 26.930 ;
        RECT 114.915 15.710 115.055 26.600 ;
        RECT 115.475 15.240 115.615 26.600 ;
        RECT 116.035 26.600 116.735 26.930 ;
        RECT 116.035 15.710 116.175 26.600 ;
        RECT 116.595 15.240 116.735 26.600 ;
        RECT 117.155 26.600 117.855 26.930 ;
        RECT 117.155 15.710 117.295 26.600 ;
        RECT 117.715 15.240 117.855 26.600 ;
        RECT 118.275 26.600 118.975 26.930 ;
        RECT 118.275 15.710 118.415 26.600 ;
        RECT 118.835 15.240 118.975 26.600 ;
        RECT 119.395 26.600 120.095 26.930 ;
        RECT 119.395 15.710 119.535 26.600 ;
        RECT 119.955 15.240 120.095 26.600 ;
        RECT 120.515 26.600 122.685 26.930 ;
        RECT 124.645 26.600 125.345 26.930 ;
        RECT 120.515 15.710 120.655 26.600 ;
        RECT 121.075 15.240 121.215 26.600 ;
        RECT 121.635 15.710 121.775 26.600 ;
        RECT 122.195 15.710 122.335 26.600 ;
        RECT 124.645 15.710 124.785 26.600 ;
        RECT 125.205 15.240 125.345 26.600 ;
        RECT 125.765 26.600 126.465 26.930 ;
        RECT 125.765 15.710 125.905 26.600 ;
        RECT 126.325 15.240 126.465 26.600 ;
        RECT 126.885 26.600 127.585 26.930 ;
        RECT 126.885 15.710 127.025 26.600 ;
        RECT 127.445 15.240 127.585 26.600 ;
        RECT 128.005 26.600 128.705 26.930 ;
        RECT 128.005 15.710 128.145 26.600 ;
        RECT 128.565 15.240 128.705 26.600 ;
        RECT 129.125 26.600 129.825 26.930 ;
        RECT 129.125 15.710 129.265 26.600 ;
        RECT 129.685 15.240 129.825 26.600 ;
        RECT 130.245 26.600 130.945 26.930 ;
        RECT 130.245 15.710 130.385 26.600 ;
        RECT 130.805 15.240 130.945 26.600 ;
        RECT 131.365 26.600 132.065 26.930 ;
        RECT 131.365 15.710 131.505 26.600 ;
        RECT 131.925 15.240 132.065 26.600 ;
        RECT 132.485 26.600 133.185 26.930 ;
        RECT 132.485 15.710 132.625 26.600 ;
        RECT 133.045 15.240 133.185 26.600 ;
        RECT 133.605 26.600 135.775 26.930 ;
        RECT 133.605 15.710 133.745 26.600 ;
        RECT 134.165 15.240 134.305 26.600 ;
        RECT 134.725 15.710 134.865 26.600 ;
        RECT 135.285 15.710 135.425 26.600 ;
        RECT 137.735 26.580 138.435 26.910 ;
        RECT 137.735 15.690 137.875 26.580 ;
        RECT 138.295 15.220 138.435 26.580 ;
        RECT 138.855 26.580 139.555 26.910 ;
        RECT 138.855 15.690 138.995 26.580 ;
        RECT 139.415 15.220 139.555 26.580 ;
        RECT 139.975 26.580 140.675 26.910 ;
        RECT 139.975 15.690 140.115 26.580 ;
        RECT 140.535 15.220 140.675 26.580 ;
        RECT 141.095 26.580 141.795 26.910 ;
        RECT 141.095 15.690 141.235 26.580 ;
        RECT 141.655 15.220 141.795 26.580 ;
        RECT 142.215 26.580 142.915 26.910 ;
        RECT 142.215 15.690 142.355 26.580 ;
        RECT 142.775 15.220 142.915 26.580 ;
        RECT 143.335 26.580 144.035 26.910 ;
        RECT 143.335 15.690 143.475 26.580 ;
        RECT 143.895 15.220 144.035 26.580 ;
        RECT 144.455 26.580 145.155 26.910 ;
        RECT 144.455 15.690 144.595 26.580 ;
        RECT 145.015 15.220 145.155 26.580 ;
        RECT 145.575 26.580 146.275 26.910 ;
        RECT 145.575 15.690 145.715 26.580 ;
        RECT 146.135 15.220 146.275 26.580 ;
        RECT 146.695 26.580 148.865 26.910 ;
        RECT 150.825 26.580 151.525 26.910 ;
        RECT 146.695 15.690 146.835 26.580 ;
        RECT 147.255 15.220 147.395 26.580 ;
        RECT 147.815 15.690 147.955 26.580 ;
        RECT 148.375 15.690 148.515 26.580 ;
        RECT 150.825 15.690 150.965 26.580 ;
        RECT 151.385 15.220 151.525 26.580 ;
        RECT 151.945 26.580 152.645 26.910 ;
        RECT 151.945 15.690 152.085 26.580 ;
        RECT 152.505 15.220 152.645 26.580 ;
        RECT 153.065 26.580 153.765 26.910 ;
        RECT 153.065 15.690 153.205 26.580 ;
        RECT 153.625 15.220 153.765 26.580 ;
        RECT 154.185 26.580 154.885 26.910 ;
        RECT 154.185 15.690 154.325 26.580 ;
        RECT 154.745 15.220 154.885 26.580 ;
        RECT 155.305 26.580 156.005 26.910 ;
        RECT 155.305 15.690 155.445 26.580 ;
        RECT 155.865 15.220 156.005 26.580 ;
        RECT 156.425 26.580 157.125 26.910 ;
        RECT 156.425 15.690 156.565 26.580 ;
        RECT 156.985 15.220 157.125 26.580 ;
        RECT 157.545 26.580 158.245 26.910 ;
        RECT 157.545 15.690 157.685 26.580 ;
        RECT 158.105 15.220 158.245 26.580 ;
        RECT 158.665 26.580 159.365 26.910 ;
        RECT 158.665 15.690 158.805 26.580 ;
        RECT 159.225 15.220 159.365 26.580 ;
        RECT 159.785 26.580 161.955 26.910 ;
        RECT 159.785 15.690 159.925 26.580 ;
        RECT 160.345 15.220 160.485 26.580 ;
        RECT 160.905 15.690 161.045 26.580 ;
        RECT 161.465 15.690 161.605 26.580 ;
        RECT 6.905 2.200 7.045 13.090 ;
        RECT 7.465 2.200 7.605 13.560 ;
        RECT 6.905 1.870 7.605 2.200 ;
        RECT 8.025 2.200 8.165 13.090 ;
        RECT 8.585 2.200 8.725 13.560 ;
        RECT 8.025 1.870 8.725 2.200 ;
        RECT 9.145 2.200 9.285 13.090 ;
        RECT 9.705 2.200 9.845 13.560 ;
        RECT 9.145 1.870 9.845 2.200 ;
        RECT 10.265 2.200 10.405 13.090 ;
        RECT 10.825 2.200 10.965 13.560 ;
        RECT 10.265 1.870 10.965 2.200 ;
        RECT 11.385 2.200 11.525 13.090 ;
        RECT 11.945 2.200 12.085 13.560 ;
        RECT 11.385 1.870 12.085 2.200 ;
        RECT 12.505 2.200 12.645 13.090 ;
        RECT 13.065 2.200 13.205 13.560 ;
        RECT 12.505 1.870 13.205 2.200 ;
        RECT 13.625 2.200 13.765 13.090 ;
        RECT 14.185 2.200 14.325 13.560 ;
        RECT 13.625 1.870 14.325 2.200 ;
        RECT 14.745 2.200 14.885 13.090 ;
        RECT 15.305 2.200 15.445 13.560 ;
        RECT 14.745 1.870 15.445 2.200 ;
        RECT 15.865 2.200 16.005 13.090 ;
        RECT 16.425 2.200 16.565 13.560 ;
        RECT 16.985 2.200 17.125 13.090 ;
        RECT 17.545 2.200 17.685 13.090 ;
        RECT 19.995 2.200 20.135 13.090 ;
        RECT 20.555 2.200 20.695 13.560 ;
        RECT 15.865 1.870 18.035 2.200 ;
        RECT 19.995 1.870 20.695 2.200 ;
        RECT 21.115 2.200 21.255 13.090 ;
        RECT 21.675 2.200 21.815 13.560 ;
        RECT 21.115 1.870 21.815 2.200 ;
        RECT 22.235 2.200 22.375 13.090 ;
        RECT 22.795 2.200 22.935 13.560 ;
        RECT 22.235 1.870 22.935 2.200 ;
        RECT 23.355 2.200 23.495 13.090 ;
        RECT 23.915 2.200 24.055 13.560 ;
        RECT 23.355 1.870 24.055 2.200 ;
        RECT 24.475 2.200 24.615 13.090 ;
        RECT 25.035 2.200 25.175 13.560 ;
        RECT 24.475 1.870 25.175 2.200 ;
        RECT 25.595 2.200 25.735 13.090 ;
        RECT 26.155 2.200 26.295 13.560 ;
        RECT 25.595 1.870 26.295 2.200 ;
        RECT 26.715 2.200 26.855 13.090 ;
        RECT 27.275 2.200 27.415 13.560 ;
        RECT 26.715 1.870 27.415 2.200 ;
        RECT 27.835 2.200 27.975 13.090 ;
        RECT 28.395 2.200 28.535 13.560 ;
        RECT 27.835 1.870 28.535 2.200 ;
        RECT 28.955 2.200 29.095 13.090 ;
        RECT 29.515 2.200 29.655 13.560 ;
        RECT 30.075 2.200 30.215 13.090 ;
        RECT 30.635 2.200 30.775 13.090 ;
        RECT 33.085 2.220 33.225 13.110 ;
        RECT 33.645 2.220 33.785 13.580 ;
        RECT 28.955 1.870 31.125 2.200 ;
        RECT 33.085 1.890 33.785 2.220 ;
        RECT 34.205 2.220 34.345 13.110 ;
        RECT 34.765 2.220 34.905 13.580 ;
        RECT 34.205 1.890 34.905 2.220 ;
        RECT 35.325 2.220 35.465 13.110 ;
        RECT 35.885 2.220 36.025 13.580 ;
        RECT 35.325 1.890 36.025 2.220 ;
        RECT 36.445 2.220 36.585 13.110 ;
        RECT 37.005 2.220 37.145 13.580 ;
        RECT 36.445 1.890 37.145 2.220 ;
        RECT 37.565 2.220 37.705 13.110 ;
        RECT 38.125 2.220 38.265 13.580 ;
        RECT 37.565 1.890 38.265 2.220 ;
        RECT 38.685 2.220 38.825 13.110 ;
        RECT 39.245 2.220 39.385 13.580 ;
        RECT 38.685 1.890 39.385 2.220 ;
        RECT 39.805 2.220 39.945 13.110 ;
        RECT 40.365 2.220 40.505 13.580 ;
        RECT 39.805 1.890 40.505 2.220 ;
        RECT 40.925 2.220 41.065 13.110 ;
        RECT 41.485 2.220 41.625 13.580 ;
        RECT 40.925 1.890 41.625 2.220 ;
        RECT 42.045 2.220 42.185 13.110 ;
        RECT 42.605 2.220 42.745 13.580 ;
        RECT 43.165 2.220 43.305 13.110 ;
        RECT 43.725 2.220 43.865 13.110 ;
        RECT 46.175 2.220 46.315 13.110 ;
        RECT 46.735 2.220 46.875 13.580 ;
        RECT 42.045 1.890 44.215 2.220 ;
        RECT 46.175 1.890 46.875 2.220 ;
        RECT 47.295 2.220 47.435 13.110 ;
        RECT 47.855 2.220 47.995 13.580 ;
        RECT 47.295 1.890 47.995 2.220 ;
        RECT 48.415 2.220 48.555 13.110 ;
        RECT 48.975 2.220 49.115 13.580 ;
        RECT 48.415 1.890 49.115 2.220 ;
        RECT 49.535 2.220 49.675 13.110 ;
        RECT 50.095 2.220 50.235 13.580 ;
        RECT 49.535 1.890 50.235 2.220 ;
        RECT 50.655 2.220 50.795 13.110 ;
        RECT 51.215 2.220 51.355 13.580 ;
        RECT 50.655 1.890 51.355 2.220 ;
        RECT 51.775 2.220 51.915 13.110 ;
        RECT 52.335 2.220 52.475 13.580 ;
        RECT 51.775 1.890 52.475 2.220 ;
        RECT 52.895 2.220 53.035 13.110 ;
        RECT 53.455 2.220 53.595 13.580 ;
        RECT 52.895 1.890 53.595 2.220 ;
        RECT 54.015 2.220 54.155 13.110 ;
        RECT 54.575 2.220 54.715 13.580 ;
        RECT 54.015 1.890 54.715 2.220 ;
        RECT 55.135 2.220 55.275 13.110 ;
        RECT 55.695 2.220 55.835 13.580 ;
        RECT 56.255 2.220 56.395 13.110 ;
        RECT 56.815 2.220 56.955 13.110 ;
        RECT 59.225 2.220 59.365 13.110 ;
        RECT 59.785 2.220 59.925 13.580 ;
        RECT 55.135 1.890 57.305 2.220 ;
        RECT 59.225 1.890 59.925 2.220 ;
        RECT 60.345 2.220 60.485 13.110 ;
        RECT 60.905 2.220 61.045 13.580 ;
        RECT 60.345 1.890 61.045 2.220 ;
        RECT 61.465 2.220 61.605 13.110 ;
        RECT 62.025 2.220 62.165 13.580 ;
        RECT 61.465 1.890 62.165 2.220 ;
        RECT 62.585 2.220 62.725 13.110 ;
        RECT 63.145 2.220 63.285 13.580 ;
        RECT 62.585 1.890 63.285 2.220 ;
        RECT 63.705 2.220 63.845 13.110 ;
        RECT 64.265 2.220 64.405 13.580 ;
        RECT 63.705 1.890 64.405 2.220 ;
        RECT 64.825 2.220 64.965 13.110 ;
        RECT 65.385 2.220 65.525 13.580 ;
        RECT 64.825 1.890 65.525 2.220 ;
        RECT 65.945 2.220 66.085 13.110 ;
        RECT 66.505 2.220 66.645 13.580 ;
        RECT 65.945 1.890 66.645 2.220 ;
        RECT 67.065 2.220 67.205 13.110 ;
        RECT 67.625 2.220 67.765 13.580 ;
        RECT 67.065 1.890 67.765 2.220 ;
        RECT 68.185 2.220 68.325 13.110 ;
        RECT 68.745 2.220 68.885 13.580 ;
        RECT 69.305 2.220 69.445 13.110 ;
        RECT 69.865 2.220 70.005 13.110 ;
        RECT 72.315 2.220 72.455 13.110 ;
        RECT 72.875 2.220 73.015 13.580 ;
        RECT 68.185 1.890 70.355 2.220 ;
        RECT 72.315 1.890 73.015 2.220 ;
        RECT 73.435 2.220 73.575 13.110 ;
        RECT 73.995 2.220 74.135 13.580 ;
        RECT 73.435 1.890 74.135 2.220 ;
        RECT 74.555 2.220 74.695 13.110 ;
        RECT 75.115 2.220 75.255 13.580 ;
        RECT 74.555 1.890 75.255 2.220 ;
        RECT 75.675 2.220 75.815 13.110 ;
        RECT 76.235 2.220 76.375 13.580 ;
        RECT 75.675 1.890 76.375 2.220 ;
        RECT 76.795 2.220 76.935 13.110 ;
        RECT 77.355 2.220 77.495 13.580 ;
        RECT 76.795 1.890 77.495 2.220 ;
        RECT 77.915 2.220 78.055 13.110 ;
        RECT 78.475 2.220 78.615 13.580 ;
        RECT 77.915 1.890 78.615 2.220 ;
        RECT 79.035 2.220 79.175 13.110 ;
        RECT 79.595 2.220 79.735 13.580 ;
        RECT 79.035 1.890 79.735 2.220 ;
        RECT 80.155 2.220 80.295 13.110 ;
        RECT 80.715 2.220 80.855 13.580 ;
        RECT 80.155 1.890 80.855 2.220 ;
        RECT 81.275 2.220 81.415 13.110 ;
        RECT 81.835 2.220 81.975 13.580 ;
        RECT 82.395 2.220 82.535 13.110 ;
        RECT 82.955 2.220 83.095 13.110 ;
        RECT 85.405 2.240 85.545 13.130 ;
        RECT 85.965 2.240 86.105 13.600 ;
        RECT 81.275 1.890 83.445 2.220 ;
        RECT 85.405 1.910 86.105 2.240 ;
        RECT 86.525 2.240 86.665 13.130 ;
        RECT 87.085 2.240 87.225 13.600 ;
        RECT 86.525 1.910 87.225 2.240 ;
        RECT 87.645 2.240 87.785 13.130 ;
        RECT 88.205 2.240 88.345 13.600 ;
        RECT 87.645 1.910 88.345 2.240 ;
        RECT 88.765 2.240 88.905 13.130 ;
        RECT 89.325 2.240 89.465 13.600 ;
        RECT 88.765 1.910 89.465 2.240 ;
        RECT 89.885 2.240 90.025 13.130 ;
        RECT 90.445 2.240 90.585 13.600 ;
        RECT 89.885 1.910 90.585 2.240 ;
        RECT 91.005 2.240 91.145 13.130 ;
        RECT 91.565 2.240 91.705 13.600 ;
        RECT 91.005 1.910 91.705 2.240 ;
        RECT 92.125 2.240 92.265 13.130 ;
        RECT 92.685 2.240 92.825 13.600 ;
        RECT 92.125 1.910 92.825 2.240 ;
        RECT 93.245 2.240 93.385 13.130 ;
        RECT 93.805 2.240 93.945 13.600 ;
        RECT 93.245 1.910 93.945 2.240 ;
        RECT 94.365 2.240 94.505 13.130 ;
        RECT 94.925 2.240 95.065 13.600 ;
        RECT 95.485 2.240 95.625 13.130 ;
        RECT 96.045 2.240 96.185 13.130 ;
        RECT 98.495 2.240 98.635 13.130 ;
        RECT 99.055 2.240 99.195 13.600 ;
        RECT 94.365 1.910 96.535 2.240 ;
        RECT 98.495 1.910 99.195 2.240 ;
        RECT 99.615 2.240 99.755 13.130 ;
        RECT 100.175 2.240 100.315 13.600 ;
        RECT 99.615 1.910 100.315 2.240 ;
        RECT 100.735 2.240 100.875 13.130 ;
        RECT 101.295 2.240 101.435 13.600 ;
        RECT 100.735 1.910 101.435 2.240 ;
        RECT 101.855 2.240 101.995 13.130 ;
        RECT 102.415 2.240 102.555 13.600 ;
        RECT 101.855 1.910 102.555 2.240 ;
        RECT 102.975 2.240 103.115 13.130 ;
        RECT 103.535 2.240 103.675 13.600 ;
        RECT 102.975 1.910 103.675 2.240 ;
        RECT 104.095 2.240 104.235 13.130 ;
        RECT 104.655 2.240 104.795 13.600 ;
        RECT 104.095 1.910 104.795 2.240 ;
        RECT 105.215 2.240 105.355 13.130 ;
        RECT 105.775 2.240 105.915 13.600 ;
        RECT 105.215 1.910 105.915 2.240 ;
        RECT 106.335 2.240 106.475 13.130 ;
        RECT 106.895 2.240 107.035 13.600 ;
        RECT 106.335 1.910 107.035 2.240 ;
        RECT 107.455 2.240 107.595 13.130 ;
        RECT 108.015 2.240 108.155 13.600 ;
        RECT 108.575 2.240 108.715 13.130 ;
        RECT 109.135 2.240 109.275 13.130 ;
        RECT 111.585 2.240 111.725 13.130 ;
        RECT 112.145 2.240 112.285 13.600 ;
        RECT 107.455 1.910 109.625 2.240 ;
        RECT 111.585 1.910 112.285 2.240 ;
        RECT 112.705 2.240 112.845 13.130 ;
        RECT 113.265 2.240 113.405 13.600 ;
        RECT 112.705 1.910 113.405 2.240 ;
        RECT 113.825 2.240 113.965 13.130 ;
        RECT 114.385 2.240 114.525 13.600 ;
        RECT 113.825 1.910 114.525 2.240 ;
        RECT 114.945 2.240 115.085 13.130 ;
        RECT 115.505 2.240 115.645 13.600 ;
        RECT 114.945 1.910 115.645 2.240 ;
        RECT 116.065 2.240 116.205 13.130 ;
        RECT 116.625 2.240 116.765 13.600 ;
        RECT 116.065 1.910 116.765 2.240 ;
        RECT 117.185 2.240 117.325 13.130 ;
        RECT 117.745 2.240 117.885 13.600 ;
        RECT 117.185 1.910 117.885 2.240 ;
        RECT 118.305 2.240 118.445 13.130 ;
        RECT 118.865 2.240 119.005 13.600 ;
        RECT 118.305 1.910 119.005 2.240 ;
        RECT 119.425 2.240 119.565 13.130 ;
        RECT 119.985 2.240 120.125 13.600 ;
        RECT 119.425 1.910 120.125 2.240 ;
        RECT 120.545 2.240 120.685 13.130 ;
        RECT 121.105 2.240 121.245 13.600 ;
        RECT 121.665 2.240 121.805 13.130 ;
        RECT 122.225 2.240 122.365 13.130 ;
        RECT 124.675 2.240 124.815 13.130 ;
        RECT 125.235 2.240 125.375 13.600 ;
        RECT 120.545 1.910 122.715 2.240 ;
        RECT 124.675 1.910 125.375 2.240 ;
        RECT 125.795 2.240 125.935 13.130 ;
        RECT 126.355 2.240 126.495 13.600 ;
        RECT 125.795 1.910 126.495 2.240 ;
        RECT 126.915 2.240 127.055 13.130 ;
        RECT 127.475 2.240 127.615 13.600 ;
        RECT 126.915 1.910 127.615 2.240 ;
        RECT 128.035 2.240 128.175 13.130 ;
        RECT 128.595 2.240 128.735 13.600 ;
        RECT 128.035 1.910 128.735 2.240 ;
        RECT 129.155 2.240 129.295 13.130 ;
        RECT 129.715 2.240 129.855 13.600 ;
        RECT 129.155 1.910 129.855 2.240 ;
        RECT 130.275 2.240 130.415 13.130 ;
        RECT 130.835 2.240 130.975 13.600 ;
        RECT 130.275 1.910 130.975 2.240 ;
        RECT 131.395 2.240 131.535 13.130 ;
        RECT 131.955 2.240 132.095 13.600 ;
        RECT 131.395 1.910 132.095 2.240 ;
        RECT 132.515 2.240 132.655 13.130 ;
        RECT 133.075 2.240 133.215 13.600 ;
        RECT 132.515 1.910 133.215 2.240 ;
        RECT 133.635 2.240 133.775 13.130 ;
        RECT 134.195 2.240 134.335 13.600 ;
        RECT 134.755 2.240 134.895 13.130 ;
        RECT 135.315 2.240 135.455 13.130 ;
        RECT 137.765 2.260 137.905 13.150 ;
        RECT 138.325 2.260 138.465 13.620 ;
        RECT 133.635 1.910 135.805 2.240 ;
        RECT 137.765 1.930 138.465 2.260 ;
        RECT 138.885 2.260 139.025 13.150 ;
        RECT 139.445 2.260 139.585 13.620 ;
        RECT 138.885 1.930 139.585 2.260 ;
        RECT 140.005 2.260 140.145 13.150 ;
        RECT 140.565 2.260 140.705 13.620 ;
        RECT 140.005 1.930 140.705 2.260 ;
        RECT 141.125 2.260 141.265 13.150 ;
        RECT 141.685 2.260 141.825 13.620 ;
        RECT 141.125 1.930 141.825 2.260 ;
        RECT 142.245 2.260 142.385 13.150 ;
        RECT 142.805 2.260 142.945 13.620 ;
        RECT 142.245 1.930 142.945 2.260 ;
        RECT 143.365 2.260 143.505 13.150 ;
        RECT 143.925 2.260 144.065 13.620 ;
        RECT 143.365 1.930 144.065 2.260 ;
        RECT 144.485 2.260 144.625 13.150 ;
        RECT 145.045 2.260 145.185 13.620 ;
        RECT 144.485 1.930 145.185 2.260 ;
        RECT 145.605 2.260 145.745 13.150 ;
        RECT 146.165 2.260 146.305 13.620 ;
        RECT 145.605 1.930 146.305 2.260 ;
        RECT 146.725 2.260 146.865 13.150 ;
        RECT 147.285 2.260 147.425 13.620 ;
        RECT 147.845 2.260 147.985 13.150 ;
        RECT 148.405 2.260 148.545 13.150 ;
        RECT 150.855 2.260 150.995 13.150 ;
        RECT 151.415 2.260 151.555 13.620 ;
        RECT 146.725 1.930 148.895 2.260 ;
        RECT 150.855 1.930 151.555 2.260 ;
        RECT 151.975 2.260 152.115 13.150 ;
        RECT 152.535 2.260 152.675 13.620 ;
        RECT 151.975 1.930 152.675 2.260 ;
        RECT 153.095 2.260 153.235 13.150 ;
        RECT 153.655 2.260 153.795 13.620 ;
        RECT 153.095 1.930 153.795 2.260 ;
        RECT 154.215 2.260 154.355 13.150 ;
        RECT 154.775 2.260 154.915 13.620 ;
        RECT 154.215 1.930 154.915 2.260 ;
        RECT 155.335 2.260 155.475 13.150 ;
        RECT 155.895 2.260 156.035 13.620 ;
        RECT 155.335 1.930 156.035 2.260 ;
        RECT 156.455 2.260 156.595 13.150 ;
        RECT 157.015 2.260 157.155 13.620 ;
        RECT 156.455 1.930 157.155 2.260 ;
        RECT 157.575 2.260 157.715 13.150 ;
        RECT 158.135 2.260 158.275 13.620 ;
        RECT 157.575 1.930 158.275 2.260 ;
        RECT 158.695 2.260 158.835 13.150 ;
        RECT 159.255 2.260 159.395 13.620 ;
        RECT 158.695 1.930 159.395 2.260 ;
        RECT 159.815 2.260 159.955 13.150 ;
        RECT 160.375 2.260 160.515 13.620 ;
        RECT 160.935 2.260 161.075 13.150 ;
        RECT 161.495 2.260 161.635 13.150 ;
        RECT 159.815 1.930 161.985 2.260 ;
      LAYER via2 ;
        RECT 6.645 118.305 6.925 118.585 ;
        RECT 7.765 118.305 8.045 118.585 ;
        RECT 8.885 118.305 9.165 118.585 ;
        RECT 10.005 118.305 10.285 118.585 ;
        RECT 11.125 118.305 11.405 118.585 ;
        RECT 12.245 118.305 12.525 118.585 ;
        RECT 13.365 118.305 13.645 118.585 ;
        RECT 14.485 118.305 14.765 118.585 ;
        RECT 15.605 118.305 15.885 118.585 ;
        RECT 16.725 118.305 17.005 118.585 ;
        RECT 19.735 118.305 20.015 118.585 ;
        RECT 20.855 118.305 21.135 118.585 ;
        RECT 21.975 118.305 22.255 118.585 ;
        RECT 23.095 118.305 23.375 118.585 ;
        RECT 24.215 118.305 24.495 118.585 ;
        RECT 25.335 118.305 25.615 118.585 ;
        RECT 26.455 118.305 26.735 118.585 ;
        RECT 27.575 118.305 27.855 118.585 ;
        RECT 28.695 118.305 28.975 118.585 ;
        RECT 29.815 118.305 30.095 118.585 ;
        RECT 32.825 118.285 33.105 118.565 ;
        RECT 33.945 118.285 34.225 118.565 ;
        RECT 35.065 118.285 35.345 118.565 ;
        RECT 36.185 118.285 36.465 118.565 ;
        RECT 37.305 118.285 37.585 118.565 ;
        RECT 38.425 118.285 38.705 118.565 ;
        RECT 39.545 118.285 39.825 118.565 ;
        RECT 40.665 118.285 40.945 118.565 ;
        RECT 41.785 118.285 42.065 118.565 ;
        RECT 42.905 118.285 43.185 118.565 ;
        RECT 45.915 118.285 46.195 118.565 ;
        RECT 47.035 118.285 47.315 118.565 ;
        RECT 48.155 118.285 48.435 118.565 ;
        RECT 49.275 118.285 49.555 118.565 ;
        RECT 50.395 118.285 50.675 118.565 ;
        RECT 51.515 118.285 51.795 118.565 ;
        RECT 52.635 118.285 52.915 118.565 ;
        RECT 53.755 118.285 54.035 118.565 ;
        RECT 54.875 118.285 55.155 118.565 ;
        RECT 55.995 118.285 56.275 118.565 ;
        RECT 58.965 118.285 59.245 118.565 ;
        RECT 60.085 118.285 60.365 118.565 ;
        RECT 61.205 118.285 61.485 118.565 ;
        RECT 62.325 118.285 62.605 118.565 ;
        RECT 63.445 118.285 63.725 118.565 ;
        RECT 64.565 118.285 64.845 118.565 ;
        RECT 65.685 118.285 65.965 118.565 ;
        RECT 66.805 118.285 67.085 118.565 ;
        RECT 67.925 118.285 68.205 118.565 ;
        RECT 69.045 118.285 69.325 118.565 ;
        RECT 72.055 118.285 72.335 118.565 ;
        RECT 73.175 118.285 73.455 118.565 ;
        RECT 74.295 118.285 74.575 118.565 ;
        RECT 75.415 118.285 75.695 118.565 ;
        RECT 76.535 118.285 76.815 118.565 ;
        RECT 77.655 118.285 77.935 118.565 ;
        RECT 78.775 118.285 79.055 118.565 ;
        RECT 79.895 118.285 80.175 118.565 ;
        RECT 81.015 118.285 81.295 118.565 ;
        RECT 82.135 118.285 82.415 118.565 ;
        RECT 85.145 118.265 85.425 118.545 ;
        RECT 86.265 118.265 86.545 118.545 ;
        RECT 87.385 118.265 87.665 118.545 ;
        RECT 88.505 118.265 88.785 118.545 ;
        RECT 89.625 118.265 89.905 118.545 ;
        RECT 90.745 118.265 91.025 118.545 ;
        RECT 91.865 118.265 92.145 118.545 ;
        RECT 92.985 118.265 93.265 118.545 ;
        RECT 94.105 118.265 94.385 118.545 ;
        RECT 95.225 118.265 95.505 118.545 ;
        RECT 98.235 118.265 98.515 118.545 ;
        RECT 99.355 118.265 99.635 118.545 ;
        RECT 100.475 118.265 100.755 118.545 ;
        RECT 101.595 118.265 101.875 118.545 ;
        RECT 102.715 118.265 102.995 118.545 ;
        RECT 103.835 118.265 104.115 118.545 ;
        RECT 104.955 118.265 105.235 118.545 ;
        RECT 106.075 118.265 106.355 118.545 ;
        RECT 107.195 118.265 107.475 118.545 ;
        RECT 108.315 118.265 108.595 118.545 ;
        RECT 111.325 118.265 111.605 118.545 ;
        RECT 112.445 118.265 112.725 118.545 ;
        RECT 113.565 118.265 113.845 118.545 ;
        RECT 114.685 118.265 114.965 118.545 ;
        RECT 115.805 118.265 116.085 118.545 ;
        RECT 116.925 118.265 117.205 118.545 ;
        RECT 118.045 118.265 118.325 118.545 ;
        RECT 119.165 118.265 119.445 118.545 ;
        RECT 120.285 118.265 120.565 118.545 ;
        RECT 121.405 118.265 121.685 118.545 ;
        RECT 124.415 118.265 124.695 118.545 ;
        RECT 125.535 118.265 125.815 118.545 ;
        RECT 126.655 118.265 126.935 118.545 ;
        RECT 127.775 118.265 128.055 118.545 ;
        RECT 128.895 118.265 129.175 118.545 ;
        RECT 130.015 118.265 130.295 118.545 ;
        RECT 131.135 118.265 131.415 118.545 ;
        RECT 132.255 118.265 132.535 118.545 ;
        RECT 133.375 118.265 133.655 118.545 ;
        RECT 134.495 118.265 134.775 118.545 ;
        RECT 137.505 118.245 137.785 118.525 ;
        RECT 138.625 118.245 138.905 118.525 ;
        RECT 139.745 118.245 140.025 118.525 ;
        RECT 140.865 118.245 141.145 118.525 ;
        RECT 141.985 118.245 142.265 118.525 ;
        RECT 143.105 118.245 143.385 118.525 ;
        RECT 144.225 118.245 144.505 118.525 ;
        RECT 145.345 118.245 145.625 118.525 ;
        RECT 146.465 118.245 146.745 118.525 ;
        RECT 147.585 118.245 147.865 118.525 ;
        RECT 150.595 118.245 150.875 118.525 ;
        RECT 151.715 118.245 151.995 118.525 ;
        RECT 152.835 118.245 153.115 118.525 ;
        RECT 153.955 118.245 154.235 118.525 ;
        RECT 155.075 118.245 155.355 118.525 ;
        RECT 156.195 118.245 156.475 118.525 ;
        RECT 157.315 118.245 157.595 118.525 ;
        RECT 158.435 118.245 158.715 118.525 ;
        RECT 159.555 118.245 159.835 118.525 ;
        RECT 160.675 118.245 160.955 118.525 ;
        RECT 6.675 93.535 6.955 93.815 ;
        RECT 7.795 93.535 8.075 93.815 ;
        RECT 8.915 93.535 9.195 93.815 ;
        RECT 10.035 93.535 10.315 93.815 ;
        RECT 11.155 93.535 11.435 93.815 ;
        RECT 12.275 93.535 12.555 93.815 ;
        RECT 13.395 93.535 13.675 93.815 ;
        RECT 14.515 93.535 14.795 93.815 ;
        RECT 15.635 93.535 15.915 93.815 ;
        RECT 16.755 93.535 17.035 93.815 ;
        RECT 19.765 93.535 20.045 93.815 ;
        RECT 20.885 93.535 21.165 93.815 ;
        RECT 22.005 93.535 22.285 93.815 ;
        RECT 23.125 93.535 23.405 93.815 ;
        RECT 24.245 93.535 24.525 93.815 ;
        RECT 25.365 93.535 25.645 93.815 ;
        RECT 26.485 93.535 26.765 93.815 ;
        RECT 27.605 93.535 27.885 93.815 ;
        RECT 28.725 93.535 29.005 93.815 ;
        RECT 29.845 93.535 30.125 93.815 ;
        RECT 32.855 93.555 33.135 93.835 ;
        RECT 33.975 93.555 34.255 93.835 ;
        RECT 35.095 93.555 35.375 93.835 ;
        RECT 36.215 93.555 36.495 93.835 ;
        RECT 37.335 93.555 37.615 93.835 ;
        RECT 38.455 93.555 38.735 93.835 ;
        RECT 39.575 93.555 39.855 93.835 ;
        RECT 40.695 93.555 40.975 93.835 ;
        RECT 41.815 93.555 42.095 93.835 ;
        RECT 42.935 93.555 43.215 93.835 ;
        RECT 45.945 93.555 46.225 93.835 ;
        RECT 47.065 93.555 47.345 93.835 ;
        RECT 48.185 93.555 48.465 93.835 ;
        RECT 49.305 93.555 49.585 93.835 ;
        RECT 50.425 93.555 50.705 93.835 ;
        RECT 51.545 93.555 51.825 93.835 ;
        RECT 52.665 93.555 52.945 93.835 ;
        RECT 53.785 93.555 54.065 93.835 ;
        RECT 54.905 93.555 55.185 93.835 ;
        RECT 56.025 93.555 56.305 93.835 ;
        RECT 58.995 93.555 59.275 93.835 ;
        RECT 60.115 93.555 60.395 93.835 ;
        RECT 61.235 93.555 61.515 93.835 ;
        RECT 62.355 93.555 62.635 93.835 ;
        RECT 63.475 93.555 63.755 93.835 ;
        RECT 64.595 93.555 64.875 93.835 ;
        RECT 65.715 93.555 65.995 93.835 ;
        RECT 66.835 93.555 67.115 93.835 ;
        RECT 67.955 93.555 68.235 93.835 ;
        RECT 69.075 93.555 69.355 93.835 ;
        RECT 72.085 93.555 72.365 93.835 ;
        RECT 73.205 93.555 73.485 93.835 ;
        RECT 74.325 93.555 74.605 93.835 ;
        RECT 75.445 93.555 75.725 93.835 ;
        RECT 76.565 93.555 76.845 93.835 ;
        RECT 77.685 93.555 77.965 93.835 ;
        RECT 78.805 93.555 79.085 93.835 ;
        RECT 79.925 93.555 80.205 93.835 ;
        RECT 81.045 93.555 81.325 93.835 ;
        RECT 82.165 93.555 82.445 93.835 ;
        RECT 85.175 93.575 85.455 93.855 ;
        RECT 86.295 93.575 86.575 93.855 ;
        RECT 87.415 93.575 87.695 93.855 ;
        RECT 88.535 93.575 88.815 93.855 ;
        RECT 89.655 93.575 89.935 93.855 ;
        RECT 90.775 93.575 91.055 93.855 ;
        RECT 91.895 93.575 92.175 93.855 ;
        RECT 93.015 93.575 93.295 93.855 ;
        RECT 94.135 93.575 94.415 93.855 ;
        RECT 95.255 93.575 95.535 93.855 ;
        RECT 98.265 93.575 98.545 93.855 ;
        RECT 99.385 93.575 99.665 93.855 ;
        RECT 100.505 93.575 100.785 93.855 ;
        RECT 101.625 93.575 101.905 93.855 ;
        RECT 102.745 93.575 103.025 93.855 ;
        RECT 103.865 93.575 104.145 93.855 ;
        RECT 104.985 93.575 105.265 93.855 ;
        RECT 106.105 93.575 106.385 93.855 ;
        RECT 107.225 93.575 107.505 93.855 ;
        RECT 108.345 93.575 108.625 93.855 ;
        RECT 111.355 93.575 111.635 93.855 ;
        RECT 112.475 93.575 112.755 93.855 ;
        RECT 113.595 93.575 113.875 93.855 ;
        RECT 114.715 93.575 114.995 93.855 ;
        RECT 115.835 93.575 116.115 93.855 ;
        RECT 116.955 93.575 117.235 93.855 ;
        RECT 118.075 93.575 118.355 93.855 ;
        RECT 119.195 93.575 119.475 93.855 ;
        RECT 120.315 93.575 120.595 93.855 ;
        RECT 121.435 93.575 121.715 93.855 ;
        RECT 124.445 93.575 124.725 93.855 ;
        RECT 125.565 93.575 125.845 93.855 ;
        RECT 126.685 93.575 126.965 93.855 ;
        RECT 127.805 93.575 128.085 93.855 ;
        RECT 128.925 93.575 129.205 93.855 ;
        RECT 130.045 93.575 130.325 93.855 ;
        RECT 131.165 93.575 131.445 93.855 ;
        RECT 132.285 93.575 132.565 93.855 ;
        RECT 133.405 93.575 133.685 93.855 ;
        RECT 134.525 93.575 134.805 93.855 ;
        RECT 137.535 93.595 137.815 93.875 ;
        RECT 138.655 93.595 138.935 93.875 ;
        RECT 139.775 93.595 140.055 93.875 ;
        RECT 140.895 93.595 141.175 93.875 ;
        RECT 142.015 93.595 142.295 93.875 ;
        RECT 143.135 93.595 143.415 93.875 ;
        RECT 144.255 93.595 144.535 93.875 ;
        RECT 145.375 93.595 145.655 93.875 ;
        RECT 146.495 93.595 146.775 93.875 ;
        RECT 147.615 93.595 147.895 93.875 ;
        RECT 150.625 93.595 150.905 93.875 ;
        RECT 151.745 93.595 152.025 93.875 ;
        RECT 152.865 93.595 153.145 93.875 ;
        RECT 153.985 93.595 154.265 93.875 ;
        RECT 155.105 93.595 155.385 93.875 ;
        RECT 156.225 93.595 156.505 93.875 ;
        RECT 157.345 93.595 157.625 93.875 ;
        RECT 158.465 93.595 158.745 93.875 ;
        RECT 159.585 93.595 159.865 93.875 ;
        RECT 160.705 93.595 160.985 93.875 ;
        RECT 167.325 89.465 167.800 89.940 ;
        RECT 1.980 88.345 2.450 88.815 ;
        RECT 1.940 33.215 2.410 33.685 ;
        RECT 166.065 29.910 166.540 30.385 ;
        RECT 7.085 26.665 7.365 26.945 ;
        RECT 8.205 26.665 8.485 26.945 ;
        RECT 9.325 26.665 9.605 26.945 ;
        RECT 10.445 26.665 10.725 26.945 ;
        RECT 11.565 26.665 11.845 26.945 ;
        RECT 12.685 26.665 12.965 26.945 ;
        RECT 13.805 26.665 14.085 26.945 ;
        RECT 14.925 26.665 15.205 26.945 ;
        RECT 16.045 26.665 16.325 26.945 ;
        RECT 17.165 26.665 17.445 26.945 ;
        RECT 20.175 26.665 20.455 26.945 ;
        RECT 21.295 26.665 21.575 26.945 ;
        RECT 22.415 26.665 22.695 26.945 ;
        RECT 23.535 26.665 23.815 26.945 ;
        RECT 24.655 26.665 24.935 26.945 ;
        RECT 25.775 26.665 26.055 26.945 ;
        RECT 26.895 26.665 27.175 26.945 ;
        RECT 28.015 26.665 28.295 26.945 ;
        RECT 29.135 26.665 29.415 26.945 ;
        RECT 30.255 26.665 30.535 26.945 ;
        RECT 33.265 26.645 33.545 26.925 ;
        RECT 34.385 26.645 34.665 26.925 ;
        RECT 35.505 26.645 35.785 26.925 ;
        RECT 36.625 26.645 36.905 26.925 ;
        RECT 37.745 26.645 38.025 26.925 ;
        RECT 38.865 26.645 39.145 26.925 ;
        RECT 39.985 26.645 40.265 26.925 ;
        RECT 41.105 26.645 41.385 26.925 ;
        RECT 42.225 26.645 42.505 26.925 ;
        RECT 43.345 26.645 43.625 26.925 ;
        RECT 46.355 26.645 46.635 26.925 ;
        RECT 47.475 26.645 47.755 26.925 ;
        RECT 48.595 26.645 48.875 26.925 ;
        RECT 49.715 26.645 49.995 26.925 ;
        RECT 50.835 26.645 51.115 26.925 ;
        RECT 51.955 26.645 52.235 26.925 ;
        RECT 53.075 26.645 53.355 26.925 ;
        RECT 54.195 26.645 54.475 26.925 ;
        RECT 55.315 26.645 55.595 26.925 ;
        RECT 56.435 26.645 56.715 26.925 ;
        RECT 59.405 26.645 59.685 26.925 ;
        RECT 60.525 26.645 60.805 26.925 ;
        RECT 61.645 26.645 61.925 26.925 ;
        RECT 62.765 26.645 63.045 26.925 ;
        RECT 63.885 26.645 64.165 26.925 ;
        RECT 65.005 26.645 65.285 26.925 ;
        RECT 66.125 26.645 66.405 26.925 ;
        RECT 67.245 26.645 67.525 26.925 ;
        RECT 68.365 26.645 68.645 26.925 ;
        RECT 69.485 26.645 69.765 26.925 ;
        RECT 72.495 26.645 72.775 26.925 ;
        RECT 73.615 26.645 73.895 26.925 ;
        RECT 74.735 26.645 75.015 26.925 ;
        RECT 75.855 26.645 76.135 26.925 ;
        RECT 76.975 26.645 77.255 26.925 ;
        RECT 78.095 26.645 78.375 26.925 ;
        RECT 79.215 26.645 79.495 26.925 ;
        RECT 80.335 26.645 80.615 26.925 ;
        RECT 81.455 26.645 81.735 26.925 ;
        RECT 82.575 26.645 82.855 26.925 ;
        RECT 85.585 26.625 85.865 26.905 ;
        RECT 86.705 26.625 86.985 26.905 ;
        RECT 87.825 26.625 88.105 26.905 ;
        RECT 88.945 26.625 89.225 26.905 ;
        RECT 90.065 26.625 90.345 26.905 ;
        RECT 91.185 26.625 91.465 26.905 ;
        RECT 92.305 26.625 92.585 26.905 ;
        RECT 93.425 26.625 93.705 26.905 ;
        RECT 94.545 26.625 94.825 26.905 ;
        RECT 95.665 26.625 95.945 26.905 ;
        RECT 98.675 26.625 98.955 26.905 ;
        RECT 99.795 26.625 100.075 26.905 ;
        RECT 100.915 26.625 101.195 26.905 ;
        RECT 102.035 26.625 102.315 26.905 ;
        RECT 103.155 26.625 103.435 26.905 ;
        RECT 104.275 26.625 104.555 26.905 ;
        RECT 105.395 26.625 105.675 26.905 ;
        RECT 106.515 26.625 106.795 26.905 ;
        RECT 107.635 26.625 107.915 26.905 ;
        RECT 108.755 26.625 109.035 26.905 ;
        RECT 111.765 26.625 112.045 26.905 ;
        RECT 112.885 26.625 113.165 26.905 ;
        RECT 114.005 26.625 114.285 26.905 ;
        RECT 115.125 26.625 115.405 26.905 ;
        RECT 116.245 26.625 116.525 26.905 ;
        RECT 117.365 26.625 117.645 26.905 ;
        RECT 118.485 26.625 118.765 26.905 ;
        RECT 119.605 26.625 119.885 26.905 ;
        RECT 120.725 26.625 121.005 26.905 ;
        RECT 121.845 26.625 122.125 26.905 ;
        RECT 124.855 26.625 125.135 26.905 ;
        RECT 125.975 26.625 126.255 26.905 ;
        RECT 127.095 26.625 127.375 26.905 ;
        RECT 128.215 26.625 128.495 26.905 ;
        RECT 129.335 26.625 129.615 26.905 ;
        RECT 130.455 26.625 130.735 26.905 ;
        RECT 131.575 26.625 131.855 26.905 ;
        RECT 132.695 26.625 132.975 26.905 ;
        RECT 133.815 26.625 134.095 26.905 ;
        RECT 134.935 26.625 135.215 26.905 ;
        RECT 137.945 26.605 138.225 26.885 ;
        RECT 139.065 26.605 139.345 26.885 ;
        RECT 140.185 26.605 140.465 26.885 ;
        RECT 141.305 26.605 141.585 26.885 ;
        RECT 142.425 26.605 142.705 26.885 ;
        RECT 143.545 26.605 143.825 26.885 ;
        RECT 144.665 26.605 144.945 26.885 ;
        RECT 145.785 26.605 146.065 26.885 ;
        RECT 146.905 26.605 147.185 26.885 ;
        RECT 148.025 26.605 148.305 26.885 ;
        RECT 151.035 26.605 151.315 26.885 ;
        RECT 152.155 26.605 152.435 26.885 ;
        RECT 153.275 26.605 153.555 26.885 ;
        RECT 154.395 26.605 154.675 26.885 ;
        RECT 155.515 26.605 155.795 26.885 ;
        RECT 156.635 26.605 156.915 26.885 ;
        RECT 157.755 26.605 158.035 26.885 ;
        RECT 158.875 26.605 159.155 26.885 ;
        RECT 159.995 26.605 160.275 26.885 ;
        RECT 161.115 26.605 161.395 26.885 ;
        RECT 7.115 1.895 7.395 2.175 ;
        RECT 8.235 1.895 8.515 2.175 ;
        RECT 9.355 1.895 9.635 2.175 ;
        RECT 10.475 1.895 10.755 2.175 ;
        RECT 11.595 1.895 11.875 2.175 ;
        RECT 12.715 1.895 12.995 2.175 ;
        RECT 13.835 1.895 14.115 2.175 ;
        RECT 14.955 1.895 15.235 2.175 ;
        RECT 16.075 1.895 16.355 2.175 ;
        RECT 17.195 1.895 17.475 2.175 ;
        RECT 20.205 1.895 20.485 2.175 ;
        RECT 21.325 1.895 21.605 2.175 ;
        RECT 22.445 1.895 22.725 2.175 ;
        RECT 23.565 1.895 23.845 2.175 ;
        RECT 24.685 1.895 24.965 2.175 ;
        RECT 25.805 1.895 26.085 2.175 ;
        RECT 26.925 1.895 27.205 2.175 ;
        RECT 28.045 1.895 28.325 2.175 ;
        RECT 29.165 1.895 29.445 2.175 ;
        RECT 30.285 1.895 30.565 2.175 ;
        RECT 33.295 1.915 33.575 2.195 ;
        RECT 34.415 1.915 34.695 2.195 ;
        RECT 35.535 1.915 35.815 2.195 ;
        RECT 36.655 1.915 36.935 2.195 ;
        RECT 37.775 1.915 38.055 2.195 ;
        RECT 38.895 1.915 39.175 2.195 ;
        RECT 40.015 1.915 40.295 2.195 ;
        RECT 41.135 1.915 41.415 2.195 ;
        RECT 42.255 1.915 42.535 2.195 ;
        RECT 43.375 1.915 43.655 2.195 ;
        RECT 46.385 1.915 46.665 2.195 ;
        RECT 47.505 1.915 47.785 2.195 ;
        RECT 48.625 1.915 48.905 2.195 ;
        RECT 49.745 1.915 50.025 2.195 ;
        RECT 50.865 1.915 51.145 2.195 ;
        RECT 51.985 1.915 52.265 2.195 ;
        RECT 53.105 1.915 53.385 2.195 ;
        RECT 54.225 1.915 54.505 2.195 ;
        RECT 55.345 1.915 55.625 2.195 ;
        RECT 56.465 1.915 56.745 2.195 ;
        RECT 59.435 1.915 59.715 2.195 ;
        RECT 60.555 1.915 60.835 2.195 ;
        RECT 61.675 1.915 61.955 2.195 ;
        RECT 62.795 1.915 63.075 2.195 ;
        RECT 63.915 1.915 64.195 2.195 ;
        RECT 65.035 1.915 65.315 2.195 ;
        RECT 66.155 1.915 66.435 2.195 ;
        RECT 67.275 1.915 67.555 2.195 ;
        RECT 68.395 1.915 68.675 2.195 ;
        RECT 69.515 1.915 69.795 2.195 ;
        RECT 72.525 1.915 72.805 2.195 ;
        RECT 73.645 1.915 73.925 2.195 ;
        RECT 74.765 1.915 75.045 2.195 ;
        RECT 75.885 1.915 76.165 2.195 ;
        RECT 77.005 1.915 77.285 2.195 ;
        RECT 78.125 1.915 78.405 2.195 ;
        RECT 79.245 1.915 79.525 2.195 ;
        RECT 80.365 1.915 80.645 2.195 ;
        RECT 81.485 1.915 81.765 2.195 ;
        RECT 82.605 1.915 82.885 2.195 ;
        RECT 85.615 1.935 85.895 2.215 ;
        RECT 86.735 1.935 87.015 2.215 ;
        RECT 87.855 1.935 88.135 2.215 ;
        RECT 88.975 1.935 89.255 2.215 ;
        RECT 90.095 1.935 90.375 2.215 ;
        RECT 91.215 1.935 91.495 2.215 ;
        RECT 92.335 1.935 92.615 2.215 ;
        RECT 93.455 1.935 93.735 2.215 ;
        RECT 94.575 1.935 94.855 2.215 ;
        RECT 95.695 1.935 95.975 2.215 ;
        RECT 98.705 1.935 98.985 2.215 ;
        RECT 99.825 1.935 100.105 2.215 ;
        RECT 100.945 1.935 101.225 2.215 ;
        RECT 102.065 1.935 102.345 2.215 ;
        RECT 103.185 1.935 103.465 2.215 ;
        RECT 104.305 1.935 104.585 2.215 ;
        RECT 105.425 1.935 105.705 2.215 ;
        RECT 106.545 1.935 106.825 2.215 ;
        RECT 107.665 1.935 107.945 2.215 ;
        RECT 108.785 1.935 109.065 2.215 ;
        RECT 111.795 1.935 112.075 2.215 ;
        RECT 112.915 1.935 113.195 2.215 ;
        RECT 114.035 1.935 114.315 2.215 ;
        RECT 115.155 1.935 115.435 2.215 ;
        RECT 116.275 1.935 116.555 2.215 ;
        RECT 117.395 1.935 117.675 2.215 ;
        RECT 118.515 1.935 118.795 2.215 ;
        RECT 119.635 1.935 119.915 2.215 ;
        RECT 120.755 1.935 121.035 2.215 ;
        RECT 121.875 1.935 122.155 2.215 ;
        RECT 124.885 1.935 125.165 2.215 ;
        RECT 126.005 1.935 126.285 2.215 ;
        RECT 127.125 1.935 127.405 2.215 ;
        RECT 128.245 1.935 128.525 2.215 ;
        RECT 129.365 1.935 129.645 2.215 ;
        RECT 130.485 1.935 130.765 2.215 ;
        RECT 131.605 1.935 131.885 2.215 ;
        RECT 132.725 1.935 133.005 2.215 ;
        RECT 133.845 1.935 134.125 2.215 ;
        RECT 134.965 1.935 135.245 2.215 ;
        RECT 137.975 1.955 138.255 2.235 ;
        RECT 139.095 1.955 139.375 2.235 ;
        RECT 140.215 1.955 140.495 2.235 ;
        RECT 141.335 1.955 141.615 2.235 ;
        RECT 142.455 1.955 142.735 2.235 ;
        RECT 143.575 1.955 143.855 2.235 ;
        RECT 144.695 1.955 144.975 2.235 ;
        RECT 145.815 1.955 146.095 2.235 ;
        RECT 146.935 1.955 147.215 2.235 ;
        RECT 148.055 1.955 148.335 2.235 ;
        RECT 151.065 1.955 151.345 2.235 ;
        RECT 152.185 1.955 152.465 2.235 ;
        RECT 153.305 1.955 153.585 2.235 ;
        RECT 154.425 1.955 154.705 2.235 ;
        RECT 155.545 1.955 155.825 2.235 ;
        RECT 156.665 1.955 156.945 2.235 ;
        RECT 157.785 1.955 158.065 2.235 ;
        RECT 158.905 1.955 159.185 2.235 ;
        RECT 160.025 1.955 160.305 2.235 ;
        RECT 161.145 1.955 161.425 2.235 ;
      LAYER met3 ;
        RECT 6.155 118.280 17.565 118.610 ;
        RECT 6.155 107.550 6.455 118.280 ;
        RECT 7.355 107.550 7.655 118.280 ;
        RECT 8.555 107.550 8.855 118.280 ;
        RECT 9.755 107.550 10.055 118.280 ;
        RECT 10.955 107.550 11.255 118.280 ;
        RECT 12.155 107.550 12.455 118.280 ;
        RECT 13.355 107.550 13.655 118.280 ;
        RECT 14.555 107.550 14.855 118.280 ;
        RECT 15.755 107.550 16.055 118.280 ;
        RECT 16.955 107.550 17.565 118.280 ;
        RECT 19.245 118.280 30.655 118.610 ;
        RECT 19.245 107.550 19.545 118.280 ;
        RECT 20.445 107.550 20.745 118.280 ;
        RECT 21.645 107.550 21.945 118.280 ;
        RECT 22.845 107.550 23.145 118.280 ;
        RECT 24.045 107.550 24.345 118.280 ;
        RECT 25.245 107.550 25.545 118.280 ;
        RECT 26.445 107.550 26.745 118.280 ;
        RECT 27.645 107.550 27.945 118.280 ;
        RECT 28.845 107.550 29.145 118.280 ;
        RECT 30.045 107.550 30.655 118.280 ;
        RECT 32.335 118.260 43.745 118.590 ;
        RECT 32.335 107.530 32.635 118.260 ;
        RECT 33.535 107.530 33.835 118.260 ;
        RECT 34.735 107.530 35.035 118.260 ;
        RECT 35.935 107.530 36.235 118.260 ;
        RECT 37.135 107.530 37.435 118.260 ;
        RECT 38.335 107.530 38.635 118.260 ;
        RECT 39.535 107.530 39.835 118.260 ;
        RECT 40.735 107.530 41.035 118.260 ;
        RECT 41.935 107.530 42.235 118.260 ;
        RECT 43.135 107.530 43.745 118.260 ;
        RECT 45.425 118.260 56.835 118.590 ;
        RECT 45.425 107.530 45.725 118.260 ;
        RECT 46.625 107.530 46.925 118.260 ;
        RECT 47.825 107.530 48.125 118.260 ;
        RECT 49.025 107.530 49.325 118.260 ;
        RECT 50.225 107.530 50.525 118.260 ;
        RECT 51.425 107.530 51.725 118.260 ;
        RECT 52.625 107.530 52.925 118.260 ;
        RECT 53.825 107.530 54.125 118.260 ;
        RECT 55.025 107.530 55.325 118.260 ;
        RECT 56.225 107.530 56.835 118.260 ;
        RECT 58.475 118.260 69.885 118.590 ;
        RECT 58.475 107.530 58.775 118.260 ;
        RECT 59.675 107.530 59.975 118.260 ;
        RECT 60.875 107.530 61.175 118.260 ;
        RECT 62.075 107.530 62.375 118.260 ;
        RECT 63.275 107.530 63.575 118.260 ;
        RECT 64.475 107.530 64.775 118.260 ;
        RECT 65.675 107.530 65.975 118.260 ;
        RECT 66.875 107.530 67.175 118.260 ;
        RECT 68.075 107.530 68.375 118.260 ;
        RECT 69.275 107.530 69.885 118.260 ;
        RECT 71.565 118.260 82.975 118.590 ;
        RECT 71.565 107.530 71.865 118.260 ;
        RECT 72.765 107.530 73.065 118.260 ;
        RECT 73.965 107.530 74.265 118.260 ;
        RECT 75.165 107.530 75.465 118.260 ;
        RECT 76.365 107.530 76.665 118.260 ;
        RECT 77.565 107.530 77.865 118.260 ;
        RECT 78.765 107.530 79.065 118.260 ;
        RECT 79.965 107.530 80.265 118.260 ;
        RECT 81.165 107.530 81.465 118.260 ;
        RECT 82.365 107.530 82.975 118.260 ;
        RECT 84.655 118.240 96.065 118.570 ;
        RECT 84.655 107.510 84.955 118.240 ;
        RECT 85.855 107.510 86.155 118.240 ;
        RECT 87.055 107.510 87.355 118.240 ;
        RECT 88.255 107.510 88.555 118.240 ;
        RECT 89.455 107.510 89.755 118.240 ;
        RECT 90.655 107.510 90.955 118.240 ;
        RECT 91.855 107.510 92.155 118.240 ;
        RECT 93.055 107.510 93.355 118.240 ;
        RECT 94.255 107.510 94.555 118.240 ;
        RECT 95.455 107.510 96.065 118.240 ;
        RECT 97.745 118.240 109.155 118.570 ;
        RECT 97.745 107.510 98.045 118.240 ;
        RECT 98.945 107.510 99.245 118.240 ;
        RECT 100.145 107.510 100.445 118.240 ;
        RECT 101.345 107.510 101.645 118.240 ;
        RECT 102.545 107.510 102.845 118.240 ;
        RECT 103.745 107.510 104.045 118.240 ;
        RECT 104.945 107.510 105.245 118.240 ;
        RECT 106.145 107.510 106.445 118.240 ;
        RECT 107.345 107.510 107.645 118.240 ;
        RECT 108.545 107.510 109.155 118.240 ;
        RECT 110.835 118.240 122.245 118.570 ;
        RECT 110.835 107.510 111.135 118.240 ;
        RECT 112.035 107.510 112.335 118.240 ;
        RECT 113.235 107.510 113.535 118.240 ;
        RECT 114.435 107.510 114.735 118.240 ;
        RECT 115.635 107.510 115.935 118.240 ;
        RECT 116.835 107.510 117.135 118.240 ;
        RECT 118.035 107.510 118.335 118.240 ;
        RECT 119.235 107.510 119.535 118.240 ;
        RECT 120.435 107.510 120.735 118.240 ;
        RECT 121.635 107.510 122.245 118.240 ;
        RECT 123.925 118.240 135.335 118.570 ;
        RECT 123.925 107.510 124.225 118.240 ;
        RECT 125.125 107.510 125.425 118.240 ;
        RECT 126.325 107.510 126.625 118.240 ;
        RECT 127.525 107.510 127.825 118.240 ;
        RECT 128.725 107.510 129.025 118.240 ;
        RECT 129.925 107.510 130.225 118.240 ;
        RECT 131.125 107.510 131.425 118.240 ;
        RECT 132.325 107.510 132.625 118.240 ;
        RECT 133.525 107.510 133.825 118.240 ;
        RECT 134.725 107.510 135.335 118.240 ;
        RECT 137.015 118.220 148.425 118.550 ;
        RECT 137.015 107.490 137.315 118.220 ;
        RECT 138.215 107.490 138.515 118.220 ;
        RECT 139.415 107.490 139.715 118.220 ;
        RECT 140.615 107.490 140.915 118.220 ;
        RECT 141.815 107.490 142.115 118.220 ;
        RECT 143.015 107.490 143.315 118.220 ;
        RECT 144.215 107.490 144.515 118.220 ;
        RECT 145.415 107.490 145.715 118.220 ;
        RECT 146.615 107.490 146.915 118.220 ;
        RECT 147.815 107.490 148.425 118.220 ;
        RECT 150.105 118.220 161.515 118.550 ;
        RECT 150.105 107.490 150.405 118.220 ;
        RECT 151.305 107.490 151.605 118.220 ;
        RECT 152.505 107.490 152.805 118.220 ;
        RECT 153.705 107.490 154.005 118.220 ;
        RECT 154.905 107.490 155.205 118.220 ;
        RECT 156.105 107.490 156.405 118.220 ;
        RECT 157.305 107.490 157.605 118.220 ;
        RECT 158.505 107.490 158.805 118.220 ;
        RECT 159.705 107.490 160.005 118.220 ;
        RECT 160.905 107.490 161.515 118.220 ;
        RECT 6.185 93.840 6.485 104.570 ;
        RECT 7.385 93.840 7.685 104.570 ;
        RECT 8.585 93.840 8.885 104.570 ;
        RECT 9.785 93.840 10.085 104.570 ;
        RECT 10.985 93.840 11.285 104.570 ;
        RECT 12.185 93.840 12.485 104.570 ;
        RECT 13.385 93.840 13.685 104.570 ;
        RECT 14.585 93.840 14.885 104.570 ;
        RECT 15.785 93.840 16.085 104.570 ;
        RECT 16.985 93.840 17.595 104.570 ;
        RECT 6.185 93.510 17.595 93.840 ;
        RECT 19.275 93.840 19.575 104.570 ;
        RECT 20.475 93.840 20.775 104.570 ;
        RECT 21.675 93.840 21.975 104.570 ;
        RECT 22.875 93.840 23.175 104.570 ;
        RECT 24.075 93.840 24.375 104.570 ;
        RECT 25.275 93.840 25.575 104.570 ;
        RECT 26.475 93.840 26.775 104.570 ;
        RECT 27.675 93.840 27.975 104.570 ;
        RECT 28.875 93.840 29.175 104.570 ;
        RECT 30.075 93.840 30.685 104.570 ;
        RECT 19.275 93.510 30.685 93.840 ;
        RECT 32.365 93.860 32.665 104.590 ;
        RECT 33.565 93.860 33.865 104.590 ;
        RECT 34.765 93.860 35.065 104.590 ;
        RECT 35.965 93.860 36.265 104.590 ;
        RECT 37.165 93.860 37.465 104.590 ;
        RECT 38.365 93.860 38.665 104.590 ;
        RECT 39.565 93.860 39.865 104.590 ;
        RECT 40.765 93.860 41.065 104.590 ;
        RECT 41.965 93.860 42.265 104.590 ;
        RECT 43.165 93.860 43.775 104.590 ;
        RECT 32.365 93.530 43.775 93.860 ;
        RECT 45.455 93.860 45.755 104.590 ;
        RECT 46.655 93.860 46.955 104.590 ;
        RECT 47.855 93.860 48.155 104.590 ;
        RECT 49.055 93.860 49.355 104.590 ;
        RECT 50.255 93.860 50.555 104.590 ;
        RECT 51.455 93.860 51.755 104.590 ;
        RECT 52.655 93.860 52.955 104.590 ;
        RECT 53.855 93.860 54.155 104.590 ;
        RECT 55.055 93.860 55.355 104.590 ;
        RECT 56.255 93.860 56.865 104.590 ;
        RECT 45.455 93.530 56.865 93.860 ;
        RECT 58.505 93.860 58.805 104.590 ;
        RECT 59.705 93.860 60.005 104.590 ;
        RECT 60.905 93.860 61.205 104.590 ;
        RECT 62.105 93.860 62.405 104.590 ;
        RECT 63.305 93.860 63.605 104.590 ;
        RECT 64.505 93.860 64.805 104.590 ;
        RECT 65.705 93.860 66.005 104.590 ;
        RECT 66.905 93.860 67.205 104.590 ;
        RECT 68.105 93.860 68.405 104.590 ;
        RECT 69.305 93.860 69.915 104.590 ;
        RECT 58.505 93.530 69.915 93.860 ;
        RECT 71.595 93.860 71.895 104.590 ;
        RECT 72.795 93.860 73.095 104.590 ;
        RECT 73.995 93.860 74.295 104.590 ;
        RECT 75.195 93.860 75.495 104.590 ;
        RECT 76.395 93.860 76.695 104.590 ;
        RECT 77.595 93.860 77.895 104.590 ;
        RECT 78.795 93.860 79.095 104.590 ;
        RECT 79.995 93.860 80.295 104.590 ;
        RECT 81.195 93.860 81.495 104.590 ;
        RECT 82.395 93.860 83.005 104.590 ;
        RECT 71.595 93.530 83.005 93.860 ;
        RECT 84.685 93.880 84.985 104.610 ;
        RECT 85.885 93.880 86.185 104.610 ;
        RECT 87.085 93.880 87.385 104.610 ;
        RECT 88.285 93.880 88.585 104.610 ;
        RECT 89.485 93.880 89.785 104.610 ;
        RECT 90.685 93.880 90.985 104.610 ;
        RECT 91.885 93.880 92.185 104.610 ;
        RECT 93.085 93.880 93.385 104.610 ;
        RECT 94.285 93.880 94.585 104.610 ;
        RECT 95.485 93.880 96.095 104.610 ;
        RECT 84.685 93.550 96.095 93.880 ;
        RECT 97.775 93.880 98.075 104.610 ;
        RECT 98.975 93.880 99.275 104.610 ;
        RECT 100.175 93.880 100.475 104.610 ;
        RECT 101.375 93.880 101.675 104.610 ;
        RECT 102.575 93.880 102.875 104.610 ;
        RECT 103.775 93.880 104.075 104.610 ;
        RECT 104.975 93.880 105.275 104.610 ;
        RECT 106.175 93.880 106.475 104.610 ;
        RECT 107.375 93.880 107.675 104.610 ;
        RECT 108.575 93.880 109.185 104.610 ;
        RECT 97.775 93.550 109.185 93.880 ;
        RECT 110.865 93.880 111.165 104.610 ;
        RECT 112.065 93.880 112.365 104.610 ;
        RECT 113.265 93.880 113.565 104.610 ;
        RECT 114.465 93.880 114.765 104.610 ;
        RECT 115.665 93.880 115.965 104.610 ;
        RECT 116.865 93.880 117.165 104.610 ;
        RECT 118.065 93.880 118.365 104.610 ;
        RECT 119.265 93.880 119.565 104.610 ;
        RECT 120.465 93.880 120.765 104.610 ;
        RECT 121.665 93.880 122.275 104.610 ;
        RECT 110.865 93.550 122.275 93.880 ;
        RECT 123.955 93.880 124.255 104.610 ;
        RECT 125.155 93.880 125.455 104.610 ;
        RECT 126.355 93.880 126.655 104.610 ;
        RECT 127.555 93.880 127.855 104.610 ;
        RECT 128.755 93.880 129.055 104.610 ;
        RECT 129.955 93.880 130.255 104.610 ;
        RECT 131.155 93.880 131.455 104.610 ;
        RECT 132.355 93.880 132.655 104.610 ;
        RECT 133.555 93.880 133.855 104.610 ;
        RECT 134.755 93.880 135.365 104.610 ;
        RECT 123.955 93.550 135.365 93.880 ;
        RECT 137.045 93.900 137.345 104.630 ;
        RECT 138.245 93.900 138.545 104.630 ;
        RECT 139.445 93.900 139.745 104.630 ;
        RECT 140.645 93.900 140.945 104.630 ;
        RECT 141.845 93.900 142.145 104.630 ;
        RECT 143.045 93.900 143.345 104.630 ;
        RECT 144.245 93.900 144.545 104.630 ;
        RECT 145.445 93.900 145.745 104.630 ;
        RECT 146.645 93.900 146.945 104.630 ;
        RECT 147.845 93.900 148.455 104.630 ;
        RECT 137.045 93.570 148.455 93.900 ;
        RECT 150.135 93.900 150.435 104.630 ;
        RECT 151.335 93.900 151.635 104.630 ;
        RECT 152.535 93.900 152.835 104.630 ;
        RECT 153.735 93.900 154.035 104.630 ;
        RECT 154.935 93.900 155.235 104.630 ;
        RECT 156.135 93.900 156.435 104.630 ;
        RECT 157.335 93.900 157.635 104.630 ;
        RECT 158.535 93.900 158.835 104.630 ;
        RECT 159.735 93.900 160.035 104.630 ;
        RECT 160.935 93.900 161.545 104.630 ;
        RECT 150.135 93.570 161.545 93.900 ;
        RECT 167.300 89.440 167.855 89.965 ;
        RECT 1.955 88.320 2.475 88.870 ;
        RECT 1.915 33.160 2.435 33.710 ;
        RECT 166.040 29.885 166.565 30.440 ;
        RECT 6.595 26.640 18.005 26.970 ;
        RECT 6.595 15.910 6.895 26.640 ;
        RECT 7.795 15.910 8.095 26.640 ;
        RECT 8.995 15.910 9.295 26.640 ;
        RECT 10.195 15.910 10.495 26.640 ;
        RECT 11.395 15.910 11.695 26.640 ;
        RECT 12.595 15.910 12.895 26.640 ;
        RECT 13.795 15.910 14.095 26.640 ;
        RECT 14.995 15.910 15.295 26.640 ;
        RECT 16.195 15.910 16.495 26.640 ;
        RECT 17.395 15.910 18.005 26.640 ;
        RECT 19.685 26.640 31.095 26.970 ;
        RECT 19.685 15.910 19.985 26.640 ;
        RECT 20.885 15.910 21.185 26.640 ;
        RECT 22.085 15.910 22.385 26.640 ;
        RECT 23.285 15.910 23.585 26.640 ;
        RECT 24.485 15.910 24.785 26.640 ;
        RECT 25.685 15.910 25.985 26.640 ;
        RECT 26.885 15.910 27.185 26.640 ;
        RECT 28.085 15.910 28.385 26.640 ;
        RECT 29.285 15.910 29.585 26.640 ;
        RECT 30.485 15.910 31.095 26.640 ;
        RECT 32.775 26.620 44.185 26.950 ;
        RECT 32.775 15.890 33.075 26.620 ;
        RECT 33.975 15.890 34.275 26.620 ;
        RECT 35.175 15.890 35.475 26.620 ;
        RECT 36.375 15.890 36.675 26.620 ;
        RECT 37.575 15.890 37.875 26.620 ;
        RECT 38.775 15.890 39.075 26.620 ;
        RECT 39.975 15.890 40.275 26.620 ;
        RECT 41.175 15.890 41.475 26.620 ;
        RECT 42.375 15.890 42.675 26.620 ;
        RECT 43.575 15.890 44.185 26.620 ;
        RECT 45.865 26.620 57.275 26.950 ;
        RECT 45.865 15.890 46.165 26.620 ;
        RECT 47.065 15.890 47.365 26.620 ;
        RECT 48.265 15.890 48.565 26.620 ;
        RECT 49.465 15.890 49.765 26.620 ;
        RECT 50.665 15.890 50.965 26.620 ;
        RECT 51.865 15.890 52.165 26.620 ;
        RECT 53.065 15.890 53.365 26.620 ;
        RECT 54.265 15.890 54.565 26.620 ;
        RECT 55.465 15.890 55.765 26.620 ;
        RECT 56.665 15.890 57.275 26.620 ;
        RECT 58.915 26.620 70.325 26.950 ;
        RECT 58.915 15.890 59.215 26.620 ;
        RECT 60.115 15.890 60.415 26.620 ;
        RECT 61.315 15.890 61.615 26.620 ;
        RECT 62.515 15.890 62.815 26.620 ;
        RECT 63.715 15.890 64.015 26.620 ;
        RECT 64.915 15.890 65.215 26.620 ;
        RECT 66.115 15.890 66.415 26.620 ;
        RECT 67.315 15.890 67.615 26.620 ;
        RECT 68.515 15.890 68.815 26.620 ;
        RECT 69.715 15.890 70.325 26.620 ;
        RECT 72.005 26.620 83.415 26.950 ;
        RECT 72.005 15.890 72.305 26.620 ;
        RECT 73.205 15.890 73.505 26.620 ;
        RECT 74.405 15.890 74.705 26.620 ;
        RECT 75.605 15.890 75.905 26.620 ;
        RECT 76.805 15.890 77.105 26.620 ;
        RECT 78.005 15.890 78.305 26.620 ;
        RECT 79.205 15.890 79.505 26.620 ;
        RECT 80.405 15.890 80.705 26.620 ;
        RECT 81.605 15.890 81.905 26.620 ;
        RECT 82.805 15.890 83.415 26.620 ;
        RECT 85.095 26.600 96.505 26.930 ;
        RECT 85.095 15.870 85.395 26.600 ;
        RECT 86.295 15.870 86.595 26.600 ;
        RECT 87.495 15.870 87.795 26.600 ;
        RECT 88.695 15.870 88.995 26.600 ;
        RECT 89.895 15.870 90.195 26.600 ;
        RECT 91.095 15.870 91.395 26.600 ;
        RECT 92.295 15.870 92.595 26.600 ;
        RECT 93.495 15.870 93.795 26.600 ;
        RECT 94.695 15.870 94.995 26.600 ;
        RECT 95.895 15.870 96.505 26.600 ;
        RECT 98.185 26.600 109.595 26.930 ;
        RECT 98.185 15.870 98.485 26.600 ;
        RECT 99.385 15.870 99.685 26.600 ;
        RECT 100.585 15.870 100.885 26.600 ;
        RECT 101.785 15.870 102.085 26.600 ;
        RECT 102.985 15.870 103.285 26.600 ;
        RECT 104.185 15.870 104.485 26.600 ;
        RECT 105.385 15.870 105.685 26.600 ;
        RECT 106.585 15.870 106.885 26.600 ;
        RECT 107.785 15.870 108.085 26.600 ;
        RECT 108.985 15.870 109.595 26.600 ;
        RECT 111.275 26.600 122.685 26.930 ;
        RECT 111.275 15.870 111.575 26.600 ;
        RECT 112.475 15.870 112.775 26.600 ;
        RECT 113.675 15.870 113.975 26.600 ;
        RECT 114.875 15.870 115.175 26.600 ;
        RECT 116.075 15.870 116.375 26.600 ;
        RECT 117.275 15.870 117.575 26.600 ;
        RECT 118.475 15.870 118.775 26.600 ;
        RECT 119.675 15.870 119.975 26.600 ;
        RECT 120.875 15.870 121.175 26.600 ;
        RECT 122.075 15.870 122.685 26.600 ;
        RECT 124.365 26.600 135.775 26.930 ;
        RECT 124.365 15.870 124.665 26.600 ;
        RECT 125.565 15.870 125.865 26.600 ;
        RECT 126.765 15.870 127.065 26.600 ;
        RECT 127.965 15.870 128.265 26.600 ;
        RECT 129.165 15.870 129.465 26.600 ;
        RECT 130.365 15.870 130.665 26.600 ;
        RECT 131.565 15.870 131.865 26.600 ;
        RECT 132.765 15.870 133.065 26.600 ;
        RECT 133.965 15.870 134.265 26.600 ;
        RECT 135.165 15.870 135.775 26.600 ;
        RECT 137.455 26.580 148.865 26.910 ;
        RECT 137.455 15.850 137.755 26.580 ;
        RECT 138.655 15.850 138.955 26.580 ;
        RECT 139.855 15.850 140.155 26.580 ;
        RECT 141.055 15.850 141.355 26.580 ;
        RECT 142.255 15.850 142.555 26.580 ;
        RECT 143.455 15.850 143.755 26.580 ;
        RECT 144.655 15.850 144.955 26.580 ;
        RECT 145.855 15.850 146.155 26.580 ;
        RECT 147.055 15.850 147.355 26.580 ;
        RECT 148.255 15.850 148.865 26.580 ;
        RECT 150.545 26.580 161.955 26.910 ;
        RECT 150.545 15.850 150.845 26.580 ;
        RECT 151.745 15.850 152.045 26.580 ;
        RECT 152.945 15.850 153.245 26.580 ;
        RECT 154.145 15.850 154.445 26.580 ;
        RECT 155.345 15.850 155.645 26.580 ;
        RECT 156.545 15.850 156.845 26.580 ;
        RECT 157.745 15.850 158.045 26.580 ;
        RECT 158.945 15.850 159.245 26.580 ;
        RECT 160.145 15.850 160.445 26.580 ;
        RECT 161.345 15.850 161.955 26.580 ;
        RECT 6.625 2.200 6.925 12.930 ;
        RECT 7.825 2.200 8.125 12.930 ;
        RECT 9.025 2.200 9.325 12.930 ;
        RECT 10.225 2.200 10.525 12.930 ;
        RECT 11.425 2.200 11.725 12.930 ;
        RECT 12.625 2.200 12.925 12.930 ;
        RECT 13.825 2.200 14.125 12.930 ;
        RECT 15.025 2.200 15.325 12.930 ;
        RECT 16.225 2.200 16.525 12.930 ;
        RECT 17.425 2.200 18.035 12.930 ;
        RECT 6.625 1.870 18.035 2.200 ;
        RECT 19.715 2.200 20.015 12.930 ;
        RECT 20.915 2.200 21.215 12.930 ;
        RECT 22.115 2.200 22.415 12.930 ;
        RECT 23.315 2.200 23.615 12.930 ;
        RECT 24.515 2.200 24.815 12.930 ;
        RECT 25.715 2.200 26.015 12.930 ;
        RECT 26.915 2.200 27.215 12.930 ;
        RECT 28.115 2.200 28.415 12.930 ;
        RECT 29.315 2.200 29.615 12.930 ;
        RECT 30.515 2.200 31.125 12.930 ;
        RECT 19.715 1.870 31.125 2.200 ;
        RECT 32.805 2.220 33.105 12.950 ;
        RECT 34.005 2.220 34.305 12.950 ;
        RECT 35.205 2.220 35.505 12.950 ;
        RECT 36.405 2.220 36.705 12.950 ;
        RECT 37.605 2.220 37.905 12.950 ;
        RECT 38.805 2.220 39.105 12.950 ;
        RECT 40.005 2.220 40.305 12.950 ;
        RECT 41.205 2.220 41.505 12.950 ;
        RECT 42.405 2.220 42.705 12.950 ;
        RECT 43.605 2.220 44.215 12.950 ;
        RECT 32.805 1.890 44.215 2.220 ;
        RECT 45.895 2.220 46.195 12.950 ;
        RECT 47.095 2.220 47.395 12.950 ;
        RECT 48.295 2.220 48.595 12.950 ;
        RECT 49.495 2.220 49.795 12.950 ;
        RECT 50.695 2.220 50.995 12.950 ;
        RECT 51.895 2.220 52.195 12.950 ;
        RECT 53.095 2.220 53.395 12.950 ;
        RECT 54.295 2.220 54.595 12.950 ;
        RECT 55.495 2.220 55.795 12.950 ;
        RECT 56.695 2.220 57.305 12.950 ;
        RECT 45.895 1.890 57.305 2.220 ;
        RECT 58.945 2.220 59.245 12.950 ;
        RECT 60.145 2.220 60.445 12.950 ;
        RECT 61.345 2.220 61.645 12.950 ;
        RECT 62.545 2.220 62.845 12.950 ;
        RECT 63.745 2.220 64.045 12.950 ;
        RECT 64.945 2.220 65.245 12.950 ;
        RECT 66.145 2.220 66.445 12.950 ;
        RECT 67.345 2.220 67.645 12.950 ;
        RECT 68.545 2.220 68.845 12.950 ;
        RECT 69.745 2.220 70.355 12.950 ;
        RECT 58.945 1.890 70.355 2.220 ;
        RECT 72.035 2.220 72.335 12.950 ;
        RECT 73.235 2.220 73.535 12.950 ;
        RECT 74.435 2.220 74.735 12.950 ;
        RECT 75.635 2.220 75.935 12.950 ;
        RECT 76.835 2.220 77.135 12.950 ;
        RECT 78.035 2.220 78.335 12.950 ;
        RECT 79.235 2.220 79.535 12.950 ;
        RECT 80.435 2.220 80.735 12.950 ;
        RECT 81.635 2.220 81.935 12.950 ;
        RECT 82.835 2.220 83.445 12.950 ;
        RECT 72.035 1.890 83.445 2.220 ;
        RECT 85.125 2.240 85.425 12.970 ;
        RECT 86.325 2.240 86.625 12.970 ;
        RECT 87.525 2.240 87.825 12.970 ;
        RECT 88.725 2.240 89.025 12.970 ;
        RECT 89.925 2.240 90.225 12.970 ;
        RECT 91.125 2.240 91.425 12.970 ;
        RECT 92.325 2.240 92.625 12.970 ;
        RECT 93.525 2.240 93.825 12.970 ;
        RECT 94.725 2.240 95.025 12.970 ;
        RECT 95.925 2.240 96.535 12.970 ;
        RECT 85.125 1.910 96.535 2.240 ;
        RECT 98.215 2.240 98.515 12.970 ;
        RECT 99.415 2.240 99.715 12.970 ;
        RECT 100.615 2.240 100.915 12.970 ;
        RECT 101.815 2.240 102.115 12.970 ;
        RECT 103.015 2.240 103.315 12.970 ;
        RECT 104.215 2.240 104.515 12.970 ;
        RECT 105.415 2.240 105.715 12.970 ;
        RECT 106.615 2.240 106.915 12.970 ;
        RECT 107.815 2.240 108.115 12.970 ;
        RECT 109.015 2.240 109.625 12.970 ;
        RECT 98.215 1.910 109.625 2.240 ;
        RECT 111.305 2.240 111.605 12.970 ;
        RECT 112.505 2.240 112.805 12.970 ;
        RECT 113.705 2.240 114.005 12.970 ;
        RECT 114.905 2.240 115.205 12.970 ;
        RECT 116.105 2.240 116.405 12.970 ;
        RECT 117.305 2.240 117.605 12.970 ;
        RECT 118.505 2.240 118.805 12.970 ;
        RECT 119.705 2.240 120.005 12.970 ;
        RECT 120.905 2.240 121.205 12.970 ;
        RECT 122.105 2.240 122.715 12.970 ;
        RECT 111.305 1.910 122.715 2.240 ;
        RECT 124.395 2.240 124.695 12.970 ;
        RECT 125.595 2.240 125.895 12.970 ;
        RECT 126.795 2.240 127.095 12.970 ;
        RECT 127.995 2.240 128.295 12.970 ;
        RECT 129.195 2.240 129.495 12.970 ;
        RECT 130.395 2.240 130.695 12.970 ;
        RECT 131.595 2.240 131.895 12.970 ;
        RECT 132.795 2.240 133.095 12.970 ;
        RECT 133.995 2.240 134.295 12.970 ;
        RECT 135.195 2.240 135.805 12.970 ;
        RECT 124.395 1.910 135.805 2.240 ;
        RECT 137.485 2.260 137.785 12.990 ;
        RECT 138.685 2.260 138.985 12.990 ;
        RECT 139.885 2.260 140.185 12.990 ;
        RECT 141.085 2.260 141.385 12.990 ;
        RECT 142.285 2.260 142.585 12.990 ;
        RECT 143.485 2.260 143.785 12.990 ;
        RECT 144.685 2.260 144.985 12.990 ;
        RECT 145.885 2.260 146.185 12.990 ;
        RECT 147.085 2.260 147.385 12.990 ;
        RECT 148.285 2.260 148.895 12.990 ;
        RECT 137.485 1.930 148.895 2.260 ;
        RECT 150.575 2.260 150.875 12.990 ;
        RECT 151.775 2.260 152.075 12.990 ;
        RECT 152.975 2.260 153.275 12.990 ;
        RECT 154.175 2.260 154.475 12.990 ;
        RECT 155.375 2.260 155.675 12.990 ;
        RECT 156.575 2.260 156.875 12.990 ;
        RECT 157.775 2.260 158.075 12.990 ;
        RECT 158.975 2.260 159.275 12.990 ;
        RECT 160.175 2.260 160.475 12.990 ;
        RECT 161.375 2.260 161.985 12.990 ;
        RECT 150.575 1.930 161.985 2.260 ;
      LAYER via3 ;
        RECT 6.295 118.285 6.615 118.605 ;
        RECT 6.695 118.285 7.015 118.605 ;
        RECT 7.095 118.285 7.415 118.605 ;
        RECT 7.495 118.285 7.815 118.605 ;
        RECT 7.895 118.285 8.215 118.605 ;
        RECT 8.295 118.285 8.615 118.605 ;
        RECT 8.695 118.285 9.015 118.605 ;
        RECT 9.095 118.285 9.415 118.605 ;
        RECT 9.495 118.285 9.815 118.605 ;
        RECT 9.895 118.285 10.215 118.605 ;
        RECT 10.295 118.285 10.615 118.605 ;
        RECT 10.695 118.285 11.015 118.605 ;
        RECT 11.095 118.285 11.415 118.605 ;
        RECT 11.495 118.285 11.815 118.605 ;
        RECT 11.895 118.285 12.215 118.605 ;
        RECT 12.295 118.285 12.615 118.605 ;
        RECT 12.695 118.285 13.015 118.605 ;
        RECT 13.095 118.285 13.415 118.605 ;
        RECT 13.495 118.285 13.815 118.605 ;
        RECT 13.895 118.285 14.215 118.605 ;
        RECT 14.295 118.285 14.615 118.605 ;
        RECT 14.695 118.285 15.015 118.605 ;
        RECT 15.095 118.285 15.415 118.605 ;
        RECT 15.495 118.285 15.815 118.605 ;
        RECT 15.895 118.285 16.215 118.605 ;
        RECT 16.295 118.285 16.615 118.605 ;
        RECT 16.695 118.285 17.015 118.605 ;
        RECT 17.095 118.285 17.415 118.605 ;
        RECT 19.385 118.285 19.705 118.605 ;
        RECT 19.785 118.285 20.105 118.605 ;
        RECT 20.185 118.285 20.505 118.605 ;
        RECT 20.585 118.285 20.905 118.605 ;
        RECT 20.985 118.285 21.305 118.605 ;
        RECT 21.385 118.285 21.705 118.605 ;
        RECT 21.785 118.285 22.105 118.605 ;
        RECT 22.185 118.285 22.505 118.605 ;
        RECT 22.585 118.285 22.905 118.605 ;
        RECT 22.985 118.285 23.305 118.605 ;
        RECT 23.385 118.285 23.705 118.605 ;
        RECT 23.785 118.285 24.105 118.605 ;
        RECT 24.185 118.285 24.505 118.605 ;
        RECT 24.585 118.285 24.905 118.605 ;
        RECT 24.985 118.285 25.305 118.605 ;
        RECT 25.385 118.285 25.705 118.605 ;
        RECT 25.785 118.285 26.105 118.605 ;
        RECT 26.185 118.285 26.505 118.605 ;
        RECT 26.585 118.285 26.905 118.605 ;
        RECT 26.985 118.285 27.305 118.605 ;
        RECT 27.385 118.285 27.705 118.605 ;
        RECT 27.785 118.285 28.105 118.605 ;
        RECT 28.185 118.285 28.505 118.605 ;
        RECT 28.585 118.285 28.905 118.605 ;
        RECT 28.985 118.285 29.305 118.605 ;
        RECT 29.385 118.285 29.705 118.605 ;
        RECT 29.785 118.285 30.105 118.605 ;
        RECT 30.185 118.285 30.505 118.605 ;
        RECT 32.475 118.265 32.795 118.585 ;
        RECT 32.875 118.265 33.195 118.585 ;
        RECT 33.275 118.265 33.595 118.585 ;
        RECT 33.675 118.265 33.995 118.585 ;
        RECT 34.075 118.265 34.395 118.585 ;
        RECT 34.475 118.265 34.795 118.585 ;
        RECT 34.875 118.265 35.195 118.585 ;
        RECT 35.275 118.265 35.595 118.585 ;
        RECT 35.675 118.265 35.995 118.585 ;
        RECT 36.075 118.265 36.395 118.585 ;
        RECT 36.475 118.265 36.795 118.585 ;
        RECT 36.875 118.265 37.195 118.585 ;
        RECT 37.275 118.265 37.595 118.585 ;
        RECT 37.675 118.265 37.995 118.585 ;
        RECT 38.075 118.265 38.395 118.585 ;
        RECT 38.475 118.265 38.795 118.585 ;
        RECT 38.875 118.265 39.195 118.585 ;
        RECT 39.275 118.265 39.595 118.585 ;
        RECT 39.675 118.265 39.995 118.585 ;
        RECT 40.075 118.265 40.395 118.585 ;
        RECT 40.475 118.265 40.795 118.585 ;
        RECT 40.875 118.265 41.195 118.585 ;
        RECT 41.275 118.265 41.595 118.585 ;
        RECT 41.675 118.265 41.995 118.585 ;
        RECT 42.075 118.265 42.395 118.585 ;
        RECT 42.475 118.265 42.795 118.585 ;
        RECT 42.875 118.265 43.195 118.585 ;
        RECT 43.275 118.265 43.595 118.585 ;
        RECT 45.565 118.265 45.885 118.585 ;
        RECT 45.965 118.265 46.285 118.585 ;
        RECT 46.365 118.265 46.685 118.585 ;
        RECT 46.765 118.265 47.085 118.585 ;
        RECT 47.165 118.265 47.485 118.585 ;
        RECT 47.565 118.265 47.885 118.585 ;
        RECT 47.965 118.265 48.285 118.585 ;
        RECT 48.365 118.265 48.685 118.585 ;
        RECT 48.765 118.265 49.085 118.585 ;
        RECT 49.165 118.265 49.485 118.585 ;
        RECT 49.565 118.265 49.885 118.585 ;
        RECT 49.965 118.265 50.285 118.585 ;
        RECT 50.365 118.265 50.685 118.585 ;
        RECT 50.765 118.265 51.085 118.585 ;
        RECT 51.165 118.265 51.485 118.585 ;
        RECT 51.565 118.265 51.885 118.585 ;
        RECT 51.965 118.265 52.285 118.585 ;
        RECT 52.365 118.265 52.685 118.585 ;
        RECT 52.765 118.265 53.085 118.585 ;
        RECT 53.165 118.265 53.485 118.585 ;
        RECT 53.565 118.265 53.885 118.585 ;
        RECT 53.965 118.265 54.285 118.585 ;
        RECT 54.365 118.265 54.685 118.585 ;
        RECT 54.765 118.265 55.085 118.585 ;
        RECT 55.165 118.265 55.485 118.585 ;
        RECT 55.565 118.265 55.885 118.585 ;
        RECT 55.965 118.265 56.285 118.585 ;
        RECT 56.365 118.265 56.685 118.585 ;
        RECT 58.615 118.265 58.935 118.585 ;
        RECT 59.015 118.265 59.335 118.585 ;
        RECT 59.415 118.265 59.735 118.585 ;
        RECT 59.815 118.265 60.135 118.585 ;
        RECT 60.215 118.265 60.535 118.585 ;
        RECT 60.615 118.265 60.935 118.585 ;
        RECT 61.015 118.265 61.335 118.585 ;
        RECT 61.415 118.265 61.735 118.585 ;
        RECT 61.815 118.265 62.135 118.585 ;
        RECT 62.215 118.265 62.535 118.585 ;
        RECT 62.615 118.265 62.935 118.585 ;
        RECT 63.015 118.265 63.335 118.585 ;
        RECT 63.415 118.265 63.735 118.585 ;
        RECT 63.815 118.265 64.135 118.585 ;
        RECT 64.215 118.265 64.535 118.585 ;
        RECT 64.615 118.265 64.935 118.585 ;
        RECT 65.015 118.265 65.335 118.585 ;
        RECT 65.415 118.265 65.735 118.585 ;
        RECT 65.815 118.265 66.135 118.585 ;
        RECT 66.215 118.265 66.535 118.585 ;
        RECT 66.615 118.265 66.935 118.585 ;
        RECT 67.015 118.265 67.335 118.585 ;
        RECT 67.415 118.265 67.735 118.585 ;
        RECT 67.815 118.265 68.135 118.585 ;
        RECT 68.215 118.265 68.535 118.585 ;
        RECT 68.615 118.265 68.935 118.585 ;
        RECT 69.015 118.265 69.335 118.585 ;
        RECT 69.415 118.265 69.735 118.585 ;
        RECT 71.705 118.265 72.025 118.585 ;
        RECT 72.105 118.265 72.425 118.585 ;
        RECT 72.505 118.265 72.825 118.585 ;
        RECT 72.905 118.265 73.225 118.585 ;
        RECT 73.305 118.265 73.625 118.585 ;
        RECT 73.705 118.265 74.025 118.585 ;
        RECT 74.105 118.265 74.425 118.585 ;
        RECT 74.505 118.265 74.825 118.585 ;
        RECT 74.905 118.265 75.225 118.585 ;
        RECT 75.305 118.265 75.625 118.585 ;
        RECT 75.705 118.265 76.025 118.585 ;
        RECT 76.105 118.265 76.425 118.585 ;
        RECT 76.505 118.265 76.825 118.585 ;
        RECT 76.905 118.265 77.225 118.585 ;
        RECT 77.305 118.265 77.625 118.585 ;
        RECT 77.705 118.265 78.025 118.585 ;
        RECT 78.105 118.265 78.425 118.585 ;
        RECT 78.505 118.265 78.825 118.585 ;
        RECT 78.905 118.265 79.225 118.585 ;
        RECT 79.305 118.265 79.625 118.585 ;
        RECT 79.705 118.265 80.025 118.585 ;
        RECT 80.105 118.265 80.425 118.585 ;
        RECT 80.505 118.265 80.825 118.585 ;
        RECT 80.905 118.265 81.225 118.585 ;
        RECT 81.305 118.265 81.625 118.585 ;
        RECT 81.705 118.265 82.025 118.585 ;
        RECT 82.105 118.265 82.425 118.585 ;
        RECT 82.505 118.265 82.825 118.585 ;
        RECT 84.795 118.245 85.115 118.565 ;
        RECT 85.195 118.245 85.515 118.565 ;
        RECT 85.595 118.245 85.915 118.565 ;
        RECT 85.995 118.245 86.315 118.565 ;
        RECT 86.395 118.245 86.715 118.565 ;
        RECT 86.795 118.245 87.115 118.565 ;
        RECT 87.195 118.245 87.515 118.565 ;
        RECT 87.595 118.245 87.915 118.565 ;
        RECT 87.995 118.245 88.315 118.565 ;
        RECT 88.395 118.245 88.715 118.565 ;
        RECT 88.795 118.245 89.115 118.565 ;
        RECT 89.195 118.245 89.515 118.565 ;
        RECT 89.595 118.245 89.915 118.565 ;
        RECT 89.995 118.245 90.315 118.565 ;
        RECT 90.395 118.245 90.715 118.565 ;
        RECT 90.795 118.245 91.115 118.565 ;
        RECT 91.195 118.245 91.515 118.565 ;
        RECT 91.595 118.245 91.915 118.565 ;
        RECT 91.995 118.245 92.315 118.565 ;
        RECT 92.395 118.245 92.715 118.565 ;
        RECT 92.795 118.245 93.115 118.565 ;
        RECT 93.195 118.245 93.515 118.565 ;
        RECT 93.595 118.245 93.915 118.565 ;
        RECT 93.995 118.245 94.315 118.565 ;
        RECT 94.395 118.245 94.715 118.565 ;
        RECT 94.795 118.245 95.115 118.565 ;
        RECT 95.195 118.245 95.515 118.565 ;
        RECT 95.595 118.245 95.915 118.565 ;
        RECT 97.885 118.245 98.205 118.565 ;
        RECT 98.285 118.245 98.605 118.565 ;
        RECT 98.685 118.245 99.005 118.565 ;
        RECT 99.085 118.245 99.405 118.565 ;
        RECT 99.485 118.245 99.805 118.565 ;
        RECT 99.885 118.245 100.205 118.565 ;
        RECT 100.285 118.245 100.605 118.565 ;
        RECT 100.685 118.245 101.005 118.565 ;
        RECT 101.085 118.245 101.405 118.565 ;
        RECT 101.485 118.245 101.805 118.565 ;
        RECT 101.885 118.245 102.205 118.565 ;
        RECT 102.285 118.245 102.605 118.565 ;
        RECT 102.685 118.245 103.005 118.565 ;
        RECT 103.085 118.245 103.405 118.565 ;
        RECT 103.485 118.245 103.805 118.565 ;
        RECT 103.885 118.245 104.205 118.565 ;
        RECT 104.285 118.245 104.605 118.565 ;
        RECT 104.685 118.245 105.005 118.565 ;
        RECT 105.085 118.245 105.405 118.565 ;
        RECT 105.485 118.245 105.805 118.565 ;
        RECT 105.885 118.245 106.205 118.565 ;
        RECT 106.285 118.245 106.605 118.565 ;
        RECT 106.685 118.245 107.005 118.565 ;
        RECT 107.085 118.245 107.405 118.565 ;
        RECT 107.485 118.245 107.805 118.565 ;
        RECT 107.885 118.245 108.205 118.565 ;
        RECT 108.285 118.245 108.605 118.565 ;
        RECT 108.685 118.245 109.005 118.565 ;
        RECT 110.975 118.245 111.295 118.565 ;
        RECT 111.375 118.245 111.695 118.565 ;
        RECT 111.775 118.245 112.095 118.565 ;
        RECT 112.175 118.245 112.495 118.565 ;
        RECT 112.575 118.245 112.895 118.565 ;
        RECT 112.975 118.245 113.295 118.565 ;
        RECT 113.375 118.245 113.695 118.565 ;
        RECT 113.775 118.245 114.095 118.565 ;
        RECT 114.175 118.245 114.495 118.565 ;
        RECT 114.575 118.245 114.895 118.565 ;
        RECT 114.975 118.245 115.295 118.565 ;
        RECT 115.375 118.245 115.695 118.565 ;
        RECT 115.775 118.245 116.095 118.565 ;
        RECT 116.175 118.245 116.495 118.565 ;
        RECT 116.575 118.245 116.895 118.565 ;
        RECT 116.975 118.245 117.295 118.565 ;
        RECT 117.375 118.245 117.695 118.565 ;
        RECT 117.775 118.245 118.095 118.565 ;
        RECT 118.175 118.245 118.495 118.565 ;
        RECT 118.575 118.245 118.895 118.565 ;
        RECT 118.975 118.245 119.295 118.565 ;
        RECT 119.375 118.245 119.695 118.565 ;
        RECT 119.775 118.245 120.095 118.565 ;
        RECT 120.175 118.245 120.495 118.565 ;
        RECT 120.575 118.245 120.895 118.565 ;
        RECT 120.975 118.245 121.295 118.565 ;
        RECT 121.375 118.245 121.695 118.565 ;
        RECT 121.775 118.245 122.095 118.565 ;
        RECT 124.065 118.245 124.385 118.565 ;
        RECT 124.465 118.245 124.785 118.565 ;
        RECT 124.865 118.245 125.185 118.565 ;
        RECT 125.265 118.245 125.585 118.565 ;
        RECT 125.665 118.245 125.985 118.565 ;
        RECT 126.065 118.245 126.385 118.565 ;
        RECT 126.465 118.245 126.785 118.565 ;
        RECT 126.865 118.245 127.185 118.565 ;
        RECT 127.265 118.245 127.585 118.565 ;
        RECT 127.665 118.245 127.985 118.565 ;
        RECT 128.065 118.245 128.385 118.565 ;
        RECT 128.465 118.245 128.785 118.565 ;
        RECT 128.865 118.245 129.185 118.565 ;
        RECT 129.265 118.245 129.585 118.565 ;
        RECT 129.665 118.245 129.985 118.565 ;
        RECT 130.065 118.245 130.385 118.565 ;
        RECT 130.465 118.245 130.785 118.565 ;
        RECT 130.865 118.245 131.185 118.565 ;
        RECT 131.265 118.245 131.585 118.565 ;
        RECT 131.665 118.245 131.985 118.565 ;
        RECT 132.065 118.245 132.385 118.565 ;
        RECT 132.465 118.245 132.785 118.565 ;
        RECT 132.865 118.245 133.185 118.565 ;
        RECT 133.265 118.245 133.585 118.565 ;
        RECT 133.665 118.245 133.985 118.565 ;
        RECT 134.065 118.245 134.385 118.565 ;
        RECT 134.465 118.245 134.785 118.565 ;
        RECT 134.865 118.245 135.185 118.565 ;
        RECT 137.155 118.225 137.475 118.545 ;
        RECT 137.555 118.225 137.875 118.545 ;
        RECT 137.955 118.225 138.275 118.545 ;
        RECT 138.355 118.225 138.675 118.545 ;
        RECT 138.755 118.225 139.075 118.545 ;
        RECT 139.155 118.225 139.475 118.545 ;
        RECT 139.555 118.225 139.875 118.545 ;
        RECT 139.955 118.225 140.275 118.545 ;
        RECT 140.355 118.225 140.675 118.545 ;
        RECT 140.755 118.225 141.075 118.545 ;
        RECT 141.155 118.225 141.475 118.545 ;
        RECT 141.555 118.225 141.875 118.545 ;
        RECT 141.955 118.225 142.275 118.545 ;
        RECT 142.355 118.225 142.675 118.545 ;
        RECT 142.755 118.225 143.075 118.545 ;
        RECT 143.155 118.225 143.475 118.545 ;
        RECT 143.555 118.225 143.875 118.545 ;
        RECT 143.955 118.225 144.275 118.545 ;
        RECT 144.355 118.225 144.675 118.545 ;
        RECT 144.755 118.225 145.075 118.545 ;
        RECT 145.155 118.225 145.475 118.545 ;
        RECT 145.555 118.225 145.875 118.545 ;
        RECT 145.955 118.225 146.275 118.545 ;
        RECT 146.355 118.225 146.675 118.545 ;
        RECT 146.755 118.225 147.075 118.545 ;
        RECT 147.155 118.225 147.475 118.545 ;
        RECT 147.555 118.225 147.875 118.545 ;
        RECT 147.955 118.225 148.275 118.545 ;
        RECT 150.245 118.225 150.565 118.545 ;
        RECT 150.645 118.225 150.965 118.545 ;
        RECT 151.045 118.225 151.365 118.545 ;
        RECT 151.445 118.225 151.765 118.545 ;
        RECT 151.845 118.225 152.165 118.545 ;
        RECT 152.245 118.225 152.565 118.545 ;
        RECT 152.645 118.225 152.965 118.545 ;
        RECT 153.045 118.225 153.365 118.545 ;
        RECT 153.445 118.225 153.765 118.545 ;
        RECT 153.845 118.225 154.165 118.545 ;
        RECT 154.245 118.225 154.565 118.545 ;
        RECT 154.645 118.225 154.965 118.545 ;
        RECT 155.045 118.225 155.365 118.545 ;
        RECT 155.445 118.225 155.765 118.545 ;
        RECT 155.845 118.225 156.165 118.545 ;
        RECT 156.245 118.225 156.565 118.545 ;
        RECT 156.645 118.225 156.965 118.545 ;
        RECT 157.045 118.225 157.365 118.545 ;
        RECT 157.445 118.225 157.765 118.545 ;
        RECT 157.845 118.225 158.165 118.545 ;
        RECT 158.245 118.225 158.565 118.545 ;
        RECT 158.645 118.225 158.965 118.545 ;
        RECT 159.045 118.225 159.365 118.545 ;
        RECT 159.445 118.225 159.765 118.545 ;
        RECT 159.845 118.225 160.165 118.545 ;
        RECT 160.245 118.225 160.565 118.545 ;
        RECT 160.645 118.225 160.965 118.545 ;
        RECT 161.045 118.225 161.365 118.545 ;
        RECT 6.325 93.515 6.645 93.835 ;
        RECT 6.725 93.515 7.045 93.835 ;
        RECT 7.125 93.515 7.445 93.835 ;
        RECT 7.525 93.515 7.845 93.835 ;
        RECT 7.925 93.515 8.245 93.835 ;
        RECT 8.325 93.515 8.645 93.835 ;
        RECT 8.725 93.515 9.045 93.835 ;
        RECT 9.125 93.515 9.445 93.835 ;
        RECT 9.525 93.515 9.845 93.835 ;
        RECT 9.925 93.515 10.245 93.835 ;
        RECT 10.325 93.515 10.645 93.835 ;
        RECT 10.725 93.515 11.045 93.835 ;
        RECT 11.125 93.515 11.445 93.835 ;
        RECT 11.525 93.515 11.845 93.835 ;
        RECT 11.925 93.515 12.245 93.835 ;
        RECT 12.325 93.515 12.645 93.835 ;
        RECT 12.725 93.515 13.045 93.835 ;
        RECT 13.125 93.515 13.445 93.835 ;
        RECT 13.525 93.515 13.845 93.835 ;
        RECT 13.925 93.515 14.245 93.835 ;
        RECT 14.325 93.515 14.645 93.835 ;
        RECT 14.725 93.515 15.045 93.835 ;
        RECT 15.125 93.515 15.445 93.835 ;
        RECT 15.525 93.515 15.845 93.835 ;
        RECT 15.925 93.515 16.245 93.835 ;
        RECT 16.325 93.515 16.645 93.835 ;
        RECT 16.725 93.515 17.045 93.835 ;
        RECT 17.125 93.515 17.445 93.835 ;
        RECT 19.415 93.515 19.735 93.835 ;
        RECT 19.815 93.515 20.135 93.835 ;
        RECT 20.215 93.515 20.535 93.835 ;
        RECT 20.615 93.515 20.935 93.835 ;
        RECT 21.015 93.515 21.335 93.835 ;
        RECT 21.415 93.515 21.735 93.835 ;
        RECT 21.815 93.515 22.135 93.835 ;
        RECT 22.215 93.515 22.535 93.835 ;
        RECT 22.615 93.515 22.935 93.835 ;
        RECT 23.015 93.515 23.335 93.835 ;
        RECT 23.415 93.515 23.735 93.835 ;
        RECT 23.815 93.515 24.135 93.835 ;
        RECT 24.215 93.515 24.535 93.835 ;
        RECT 24.615 93.515 24.935 93.835 ;
        RECT 25.015 93.515 25.335 93.835 ;
        RECT 25.415 93.515 25.735 93.835 ;
        RECT 25.815 93.515 26.135 93.835 ;
        RECT 26.215 93.515 26.535 93.835 ;
        RECT 26.615 93.515 26.935 93.835 ;
        RECT 27.015 93.515 27.335 93.835 ;
        RECT 27.415 93.515 27.735 93.835 ;
        RECT 27.815 93.515 28.135 93.835 ;
        RECT 28.215 93.515 28.535 93.835 ;
        RECT 28.615 93.515 28.935 93.835 ;
        RECT 29.015 93.515 29.335 93.835 ;
        RECT 29.415 93.515 29.735 93.835 ;
        RECT 29.815 93.515 30.135 93.835 ;
        RECT 30.215 93.515 30.535 93.835 ;
        RECT 32.505 93.535 32.825 93.855 ;
        RECT 32.905 93.535 33.225 93.855 ;
        RECT 33.305 93.535 33.625 93.855 ;
        RECT 33.705 93.535 34.025 93.855 ;
        RECT 34.105 93.535 34.425 93.855 ;
        RECT 34.505 93.535 34.825 93.855 ;
        RECT 34.905 93.535 35.225 93.855 ;
        RECT 35.305 93.535 35.625 93.855 ;
        RECT 35.705 93.535 36.025 93.855 ;
        RECT 36.105 93.535 36.425 93.855 ;
        RECT 36.505 93.535 36.825 93.855 ;
        RECT 36.905 93.535 37.225 93.855 ;
        RECT 37.305 93.535 37.625 93.855 ;
        RECT 37.705 93.535 38.025 93.855 ;
        RECT 38.105 93.535 38.425 93.855 ;
        RECT 38.505 93.535 38.825 93.855 ;
        RECT 38.905 93.535 39.225 93.855 ;
        RECT 39.305 93.535 39.625 93.855 ;
        RECT 39.705 93.535 40.025 93.855 ;
        RECT 40.105 93.535 40.425 93.855 ;
        RECT 40.505 93.535 40.825 93.855 ;
        RECT 40.905 93.535 41.225 93.855 ;
        RECT 41.305 93.535 41.625 93.855 ;
        RECT 41.705 93.535 42.025 93.855 ;
        RECT 42.105 93.535 42.425 93.855 ;
        RECT 42.505 93.535 42.825 93.855 ;
        RECT 42.905 93.535 43.225 93.855 ;
        RECT 43.305 93.535 43.625 93.855 ;
        RECT 45.595 93.535 45.915 93.855 ;
        RECT 45.995 93.535 46.315 93.855 ;
        RECT 46.395 93.535 46.715 93.855 ;
        RECT 46.795 93.535 47.115 93.855 ;
        RECT 47.195 93.535 47.515 93.855 ;
        RECT 47.595 93.535 47.915 93.855 ;
        RECT 47.995 93.535 48.315 93.855 ;
        RECT 48.395 93.535 48.715 93.855 ;
        RECT 48.795 93.535 49.115 93.855 ;
        RECT 49.195 93.535 49.515 93.855 ;
        RECT 49.595 93.535 49.915 93.855 ;
        RECT 49.995 93.535 50.315 93.855 ;
        RECT 50.395 93.535 50.715 93.855 ;
        RECT 50.795 93.535 51.115 93.855 ;
        RECT 51.195 93.535 51.515 93.855 ;
        RECT 51.595 93.535 51.915 93.855 ;
        RECT 51.995 93.535 52.315 93.855 ;
        RECT 52.395 93.535 52.715 93.855 ;
        RECT 52.795 93.535 53.115 93.855 ;
        RECT 53.195 93.535 53.515 93.855 ;
        RECT 53.595 93.535 53.915 93.855 ;
        RECT 53.995 93.535 54.315 93.855 ;
        RECT 54.395 93.535 54.715 93.855 ;
        RECT 54.795 93.535 55.115 93.855 ;
        RECT 55.195 93.535 55.515 93.855 ;
        RECT 55.595 93.535 55.915 93.855 ;
        RECT 55.995 93.535 56.315 93.855 ;
        RECT 56.395 93.535 56.715 93.855 ;
        RECT 58.645 93.535 58.965 93.855 ;
        RECT 59.045 93.535 59.365 93.855 ;
        RECT 59.445 93.535 59.765 93.855 ;
        RECT 59.845 93.535 60.165 93.855 ;
        RECT 60.245 93.535 60.565 93.855 ;
        RECT 60.645 93.535 60.965 93.855 ;
        RECT 61.045 93.535 61.365 93.855 ;
        RECT 61.445 93.535 61.765 93.855 ;
        RECT 61.845 93.535 62.165 93.855 ;
        RECT 62.245 93.535 62.565 93.855 ;
        RECT 62.645 93.535 62.965 93.855 ;
        RECT 63.045 93.535 63.365 93.855 ;
        RECT 63.445 93.535 63.765 93.855 ;
        RECT 63.845 93.535 64.165 93.855 ;
        RECT 64.245 93.535 64.565 93.855 ;
        RECT 64.645 93.535 64.965 93.855 ;
        RECT 65.045 93.535 65.365 93.855 ;
        RECT 65.445 93.535 65.765 93.855 ;
        RECT 65.845 93.535 66.165 93.855 ;
        RECT 66.245 93.535 66.565 93.855 ;
        RECT 66.645 93.535 66.965 93.855 ;
        RECT 67.045 93.535 67.365 93.855 ;
        RECT 67.445 93.535 67.765 93.855 ;
        RECT 67.845 93.535 68.165 93.855 ;
        RECT 68.245 93.535 68.565 93.855 ;
        RECT 68.645 93.535 68.965 93.855 ;
        RECT 69.045 93.535 69.365 93.855 ;
        RECT 69.445 93.535 69.765 93.855 ;
        RECT 71.735 93.535 72.055 93.855 ;
        RECT 72.135 93.535 72.455 93.855 ;
        RECT 72.535 93.535 72.855 93.855 ;
        RECT 72.935 93.535 73.255 93.855 ;
        RECT 73.335 93.535 73.655 93.855 ;
        RECT 73.735 93.535 74.055 93.855 ;
        RECT 74.135 93.535 74.455 93.855 ;
        RECT 74.535 93.535 74.855 93.855 ;
        RECT 74.935 93.535 75.255 93.855 ;
        RECT 75.335 93.535 75.655 93.855 ;
        RECT 75.735 93.535 76.055 93.855 ;
        RECT 76.135 93.535 76.455 93.855 ;
        RECT 76.535 93.535 76.855 93.855 ;
        RECT 76.935 93.535 77.255 93.855 ;
        RECT 77.335 93.535 77.655 93.855 ;
        RECT 77.735 93.535 78.055 93.855 ;
        RECT 78.135 93.535 78.455 93.855 ;
        RECT 78.535 93.535 78.855 93.855 ;
        RECT 78.935 93.535 79.255 93.855 ;
        RECT 79.335 93.535 79.655 93.855 ;
        RECT 79.735 93.535 80.055 93.855 ;
        RECT 80.135 93.535 80.455 93.855 ;
        RECT 80.535 93.535 80.855 93.855 ;
        RECT 80.935 93.535 81.255 93.855 ;
        RECT 81.335 93.535 81.655 93.855 ;
        RECT 81.735 93.535 82.055 93.855 ;
        RECT 82.135 93.535 82.455 93.855 ;
        RECT 82.535 93.535 82.855 93.855 ;
        RECT 84.825 93.555 85.145 93.875 ;
        RECT 85.225 93.555 85.545 93.875 ;
        RECT 85.625 93.555 85.945 93.875 ;
        RECT 86.025 93.555 86.345 93.875 ;
        RECT 86.425 93.555 86.745 93.875 ;
        RECT 86.825 93.555 87.145 93.875 ;
        RECT 87.225 93.555 87.545 93.875 ;
        RECT 87.625 93.555 87.945 93.875 ;
        RECT 88.025 93.555 88.345 93.875 ;
        RECT 88.425 93.555 88.745 93.875 ;
        RECT 88.825 93.555 89.145 93.875 ;
        RECT 89.225 93.555 89.545 93.875 ;
        RECT 89.625 93.555 89.945 93.875 ;
        RECT 90.025 93.555 90.345 93.875 ;
        RECT 90.425 93.555 90.745 93.875 ;
        RECT 90.825 93.555 91.145 93.875 ;
        RECT 91.225 93.555 91.545 93.875 ;
        RECT 91.625 93.555 91.945 93.875 ;
        RECT 92.025 93.555 92.345 93.875 ;
        RECT 92.425 93.555 92.745 93.875 ;
        RECT 92.825 93.555 93.145 93.875 ;
        RECT 93.225 93.555 93.545 93.875 ;
        RECT 93.625 93.555 93.945 93.875 ;
        RECT 94.025 93.555 94.345 93.875 ;
        RECT 94.425 93.555 94.745 93.875 ;
        RECT 94.825 93.555 95.145 93.875 ;
        RECT 95.225 93.555 95.545 93.875 ;
        RECT 95.625 93.555 95.945 93.875 ;
        RECT 97.915 93.555 98.235 93.875 ;
        RECT 98.315 93.555 98.635 93.875 ;
        RECT 98.715 93.555 99.035 93.875 ;
        RECT 99.115 93.555 99.435 93.875 ;
        RECT 99.515 93.555 99.835 93.875 ;
        RECT 99.915 93.555 100.235 93.875 ;
        RECT 100.315 93.555 100.635 93.875 ;
        RECT 100.715 93.555 101.035 93.875 ;
        RECT 101.115 93.555 101.435 93.875 ;
        RECT 101.515 93.555 101.835 93.875 ;
        RECT 101.915 93.555 102.235 93.875 ;
        RECT 102.315 93.555 102.635 93.875 ;
        RECT 102.715 93.555 103.035 93.875 ;
        RECT 103.115 93.555 103.435 93.875 ;
        RECT 103.515 93.555 103.835 93.875 ;
        RECT 103.915 93.555 104.235 93.875 ;
        RECT 104.315 93.555 104.635 93.875 ;
        RECT 104.715 93.555 105.035 93.875 ;
        RECT 105.115 93.555 105.435 93.875 ;
        RECT 105.515 93.555 105.835 93.875 ;
        RECT 105.915 93.555 106.235 93.875 ;
        RECT 106.315 93.555 106.635 93.875 ;
        RECT 106.715 93.555 107.035 93.875 ;
        RECT 107.115 93.555 107.435 93.875 ;
        RECT 107.515 93.555 107.835 93.875 ;
        RECT 107.915 93.555 108.235 93.875 ;
        RECT 108.315 93.555 108.635 93.875 ;
        RECT 108.715 93.555 109.035 93.875 ;
        RECT 111.005 93.555 111.325 93.875 ;
        RECT 111.405 93.555 111.725 93.875 ;
        RECT 111.805 93.555 112.125 93.875 ;
        RECT 112.205 93.555 112.525 93.875 ;
        RECT 112.605 93.555 112.925 93.875 ;
        RECT 113.005 93.555 113.325 93.875 ;
        RECT 113.405 93.555 113.725 93.875 ;
        RECT 113.805 93.555 114.125 93.875 ;
        RECT 114.205 93.555 114.525 93.875 ;
        RECT 114.605 93.555 114.925 93.875 ;
        RECT 115.005 93.555 115.325 93.875 ;
        RECT 115.405 93.555 115.725 93.875 ;
        RECT 115.805 93.555 116.125 93.875 ;
        RECT 116.205 93.555 116.525 93.875 ;
        RECT 116.605 93.555 116.925 93.875 ;
        RECT 117.005 93.555 117.325 93.875 ;
        RECT 117.405 93.555 117.725 93.875 ;
        RECT 117.805 93.555 118.125 93.875 ;
        RECT 118.205 93.555 118.525 93.875 ;
        RECT 118.605 93.555 118.925 93.875 ;
        RECT 119.005 93.555 119.325 93.875 ;
        RECT 119.405 93.555 119.725 93.875 ;
        RECT 119.805 93.555 120.125 93.875 ;
        RECT 120.205 93.555 120.525 93.875 ;
        RECT 120.605 93.555 120.925 93.875 ;
        RECT 121.005 93.555 121.325 93.875 ;
        RECT 121.405 93.555 121.725 93.875 ;
        RECT 121.805 93.555 122.125 93.875 ;
        RECT 124.095 93.555 124.415 93.875 ;
        RECT 124.495 93.555 124.815 93.875 ;
        RECT 124.895 93.555 125.215 93.875 ;
        RECT 125.295 93.555 125.615 93.875 ;
        RECT 125.695 93.555 126.015 93.875 ;
        RECT 126.095 93.555 126.415 93.875 ;
        RECT 126.495 93.555 126.815 93.875 ;
        RECT 126.895 93.555 127.215 93.875 ;
        RECT 127.295 93.555 127.615 93.875 ;
        RECT 127.695 93.555 128.015 93.875 ;
        RECT 128.095 93.555 128.415 93.875 ;
        RECT 128.495 93.555 128.815 93.875 ;
        RECT 128.895 93.555 129.215 93.875 ;
        RECT 129.295 93.555 129.615 93.875 ;
        RECT 129.695 93.555 130.015 93.875 ;
        RECT 130.095 93.555 130.415 93.875 ;
        RECT 130.495 93.555 130.815 93.875 ;
        RECT 130.895 93.555 131.215 93.875 ;
        RECT 131.295 93.555 131.615 93.875 ;
        RECT 131.695 93.555 132.015 93.875 ;
        RECT 132.095 93.555 132.415 93.875 ;
        RECT 132.495 93.555 132.815 93.875 ;
        RECT 132.895 93.555 133.215 93.875 ;
        RECT 133.295 93.555 133.615 93.875 ;
        RECT 133.695 93.555 134.015 93.875 ;
        RECT 134.095 93.555 134.415 93.875 ;
        RECT 134.495 93.555 134.815 93.875 ;
        RECT 134.895 93.555 135.215 93.875 ;
        RECT 137.185 93.575 137.505 93.895 ;
        RECT 137.585 93.575 137.905 93.895 ;
        RECT 137.985 93.575 138.305 93.895 ;
        RECT 138.385 93.575 138.705 93.895 ;
        RECT 138.785 93.575 139.105 93.895 ;
        RECT 139.185 93.575 139.505 93.895 ;
        RECT 139.585 93.575 139.905 93.895 ;
        RECT 139.985 93.575 140.305 93.895 ;
        RECT 140.385 93.575 140.705 93.895 ;
        RECT 140.785 93.575 141.105 93.895 ;
        RECT 141.185 93.575 141.505 93.895 ;
        RECT 141.585 93.575 141.905 93.895 ;
        RECT 141.985 93.575 142.305 93.895 ;
        RECT 142.385 93.575 142.705 93.895 ;
        RECT 142.785 93.575 143.105 93.895 ;
        RECT 143.185 93.575 143.505 93.895 ;
        RECT 143.585 93.575 143.905 93.895 ;
        RECT 143.985 93.575 144.305 93.895 ;
        RECT 144.385 93.575 144.705 93.895 ;
        RECT 144.785 93.575 145.105 93.895 ;
        RECT 145.185 93.575 145.505 93.895 ;
        RECT 145.585 93.575 145.905 93.895 ;
        RECT 145.985 93.575 146.305 93.895 ;
        RECT 146.385 93.575 146.705 93.895 ;
        RECT 146.785 93.575 147.105 93.895 ;
        RECT 147.185 93.575 147.505 93.895 ;
        RECT 147.585 93.575 147.905 93.895 ;
        RECT 147.985 93.575 148.305 93.895 ;
        RECT 150.275 93.575 150.595 93.895 ;
        RECT 150.675 93.575 150.995 93.895 ;
        RECT 151.075 93.575 151.395 93.895 ;
        RECT 151.475 93.575 151.795 93.895 ;
        RECT 151.875 93.575 152.195 93.895 ;
        RECT 152.275 93.575 152.595 93.895 ;
        RECT 152.675 93.575 152.995 93.895 ;
        RECT 153.075 93.575 153.395 93.895 ;
        RECT 153.475 93.575 153.795 93.895 ;
        RECT 153.875 93.575 154.195 93.895 ;
        RECT 154.275 93.575 154.595 93.895 ;
        RECT 154.675 93.575 154.995 93.895 ;
        RECT 155.075 93.575 155.395 93.895 ;
        RECT 155.475 93.575 155.795 93.895 ;
        RECT 155.875 93.575 156.195 93.895 ;
        RECT 156.275 93.575 156.595 93.895 ;
        RECT 156.675 93.575 156.995 93.895 ;
        RECT 157.075 93.575 157.395 93.895 ;
        RECT 157.475 93.575 157.795 93.895 ;
        RECT 157.875 93.575 158.195 93.895 ;
        RECT 158.275 93.575 158.595 93.895 ;
        RECT 158.675 93.575 158.995 93.895 ;
        RECT 159.075 93.575 159.395 93.895 ;
        RECT 159.475 93.575 159.795 93.895 ;
        RECT 159.875 93.575 160.195 93.895 ;
        RECT 160.275 93.575 160.595 93.895 ;
        RECT 160.675 93.575 160.995 93.895 ;
        RECT 161.075 93.575 161.395 93.895 ;
        RECT 167.350 89.440 167.825 89.965 ;
        RECT 1.955 88.370 2.475 88.840 ;
        RECT 1.915 33.190 2.435 33.660 ;
        RECT 166.040 29.935 166.565 30.410 ;
        RECT 6.735 26.645 7.055 26.965 ;
        RECT 7.135 26.645 7.455 26.965 ;
        RECT 7.535 26.645 7.855 26.965 ;
        RECT 7.935 26.645 8.255 26.965 ;
        RECT 8.335 26.645 8.655 26.965 ;
        RECT 8.735 26.645 9.055 26.965 ;
        RECT 9.135 26.645 9.455 26.965 ;
        RECT 9.535 26.645 9.855 26.965 ;
        RECT 9.935 26.645 10.255 26.965 ;
        RECT 10.335 26.645 10.655 26.965 ;
        RECT 10.735 26.645 11.055 26.965 ;
        RECT 11.135 26.645 11.455 26.965 ;
        RECT 11.535 26.645 11.855 26.965 ;
        RECT 11.935 26.645 12.255 26.965 ;
        RECT 12.335 26.645 12.655 26.965 ;
        RECT 12.735 26.645 13.055 26.965 ;
        RECT 13.135 26.645 13.455 26.965 ;
        RECT 13.535 26.645 13.855 26.965 ;
        RECT 13.935 26.645 14.255 26.965 ;
        RECT 14.335 26.645 14.655 26.965 ;
        RECT 14.735 26.645 15.055 26.965 ;
        RECT 15.135 26.645 15.455 26.965 ;
        RECT 15.535 26.645 15.855 26.965 ;
        RECT 15.935 26.645 16.255 26.965 ;
        RECT 16.335 26.645 16.655 26.965 ;
        RECT 16.735 26.645 17.055 26.965 ;
        RECT 17.135 26.645 17.455 26.965 ;
        RECT 17.535 26.645 17.855 26.965 ;
        RECT 19.825 26.645 20.145 26.965 ;
        RECT 20.225 26.645 20.545 26.965 ;
        RECT 20.625 26.645 20.945 26.965 ;
        RECT 21.025 26.645 21.345 26.965 ;
        RECT 21.425 26.645 21.745 26.965 ;
        RECT 21.825 26.645 22.145 26.965 ;
        RECT 22.225 26.645 22.545 26.965 ;
        RECT 22.625 26.645 22.945 26.965 ;
        RECT 23.025 26.645 23.345 26.965 ;
        RECT 23.425 26.645 23.745 26.965 ;
        RECT 23.825 26.645 24.145 26.965 ;
        RECT 24.225 26.645 24.545 26.965 ;
        RECT 24.625 26.645 24.945 26.965 ;
        RECT 25.025 26.645 25.345 26.965 ;
        RECT 25.425 26.645 25.745 26.965 ;
        RECT 25.825 26.645 26.145 26.965 ;
        RECT 26.225 26.645 26.545 26.965 ;
        RECT 26.625 26.645 26.945 26.965 ;
        RECT 27.025 26.645 27.345 26.965 ;
        RECT 27.425 26.645 27.745 26.965 ;
        RECT 27.825 26.645 28.145 26.965 ;
        RECT 28.225 26.645 28.545 26.965 ;
        RECT 28.625 26.645 28.945 26.965 ;
        RECT 29.025 26.645 29.345 26.965 ;
        RECT 29.425 26.645 29.745 26.965 ;
        RECT 29.825 26.645 30.145 26.965 ;
        RECT 30.225 26.645 30.545 26.965 ;
        RECT 30.625 26.645 30.945 26.965 ;
        RECT 32.915 26.625 33.235 26.945 ;
        RECT 33.315 26.625 33.635 26.945 ;
        RECT 33.715 26.625 34.035 26.945 ;
        RECT 34.115 26.625 34.435 26.945 ;
        RECT 34.515 26.625 34.835 26.945 ;
        RECT 34.915 26.625 35.235 26.945 ;
        RECT 35.315 26.625 35.635 26.945 ;
        RECT 35.715 26.625 36.035 26.945 ;
        RECT 36.115 26.625 36.435 26.945 ;
        RECT 36.515 26.625 36.835 26.945 ;
        RECT 36.915 26.625 37.235 26.945 ;
        RECT 37.315 26.625 37.635 26.945 ;
        RECT 37.715 26.625 38.035 26.945 ;
        RECT 38.115 26.625 38.435 26.945 ;
        RECT 38.515 26.625 38.835 26.945 ;
        RECT 38.915 26.625 39.235 26.945 ;
        RECT 39.315 26.625 39.635 26.945 ;
        RECT 39.715 26.625 40.035 26.945 ;
        RECT 40.115 26.625 40.435 26.945 ;
        RECT 40.515 26.625 40.835 26.945 ;
        RECT 40.915 26.625 41.235 26.945 ;
        RECT 41.315 26.625 41.635 26.945 ;
        RECT 41.715 26.625 42.035 26.945 ;
        RECT 42.115 26.625 42.435 26.945 ;
        RECT 42.515 26.625 42.835 26.945 ;
        RECT 42.915 26.625 43.235 26.945 ;
        RECT 43.315 26.625 43.635 26.945 ;
        RECT 43.715 26.625 44.035 26.945 ;
        RECT 46.005 26.625 46.325 26.945 ;
        RECT 46.405 26.625 46.725 26.945 ;
        RECT 46.805 26.625 47.125 26.945 ;
        RECT 47.205 26.625 47.525 26.945 ;
        RECT 47.605 26.625 47.925 26.945 ;
        RECT 48.005 26.625 48.325 26.945 ;
        RECT 48.405 26.625 48.725 26.945 ;
        RECT 48.805 26.625 49.125 26.945 ;
        RECT 49.205 26.625 49.525 26.945 ;
        RECT 49.605 26.625 49.925 26.945 ;
        RECT 50.005 26.625 50.325 26.945 ;
        RECT 50.405 26.625 50.725 26.945 ;
        RECT 50.805 26.625 51.125 26.945 ;
        RECT 51.205 26.625 51.525 26.945 ;
        RECT 51.605 26.625 51.925 26.945 ;
        RECT 52.005 26.625 52.325 26.945 ;
        RECT 52.405 26.625 52.725 26.945 ;
        RECT 52.805 26.625 53.125 26.945 ;
        RECT 53.205 26.625 53.525 26.945 ;
        RECT 53.605 26.625 53.925 26.945 ;
        RECT 54.005 26.625 54.325 26.945 ;
        RECT 54.405 26.625 54.725 26.945 ;
        RECT 54.805 26.625 55.125 26.945 ;
        RECT 55.205 26.625 55.525 26.945 ;
        RECT 55.605 26.625 55.925 26.945 ;
        RECT 56.005 26.625 56.325 26.945 ;
        RECT 56.405 26.625 56.725 26.945 ;
        RECT 56.805 26.625 57.125 26.945 ;
        RECT 59.055 26.625 59.375 26.945 ;
        RECT 59.455 26.625 59.775 26.945 ;
        RECT 59.855 26.625 60.175 26.945 ;
        RECT 60.255 26.625 60.575 26.945 ;
        RECT 60.655 26.625 60.975 26.945 ;
        RECT 61.055 26.625 61.375 26.945 ;
        RECT 61.455 26.625 61.775 26.945 ;
        RECT 61.855 26.625 62.175 26.945 ;
        RECT 62.255 26.625 62.575 26.945 ;
        RECT 62.655 26.625 62.975 26.945 ;
        RECT 63.055 26.625 63.375 26.945 ;
        RECT 63.455 26.625 63.775 26.945 ;
        RECT 63.855 26.625 64.175 26.945 ;
        RECT 64.255 26.625 64.575 26.945 ;
        RECT 64.655 26.625 64.975 26.945 ;
        RECT 65.055 26.625 65.375 26.945 ;
        RECT 65.455 26.625 65.775 26.945 ;
        RECT 65.855 26.625 66.175 26.945 ;
        RECT 66.255 26.625 66.575 26.945 ;
        RECT 66.655 26.625 66.975 26.945 ;
        RECT 67.055 26.625 67.375 26.945 ;
        RECT 67.455 26.625 67.775 26.945 ;
        RECT 67.855 26.625 68.175 26.945 ;
        RECT 68.255 26.625 68.575 26.945 ;
        RECT 68.655 26.625 68.975 26.945 ;
        RECT 69.055 26.625 69.375 26.945 ;
        RECT 69.455 26.625 69.775 26.945 ;
        RECT 69.855 26.625 70.175 26.945 ;
        RECT 72.145 26.625 72.465 26.945 ;
        RECT 72.545 26.625 72.865 26.945 ;
        RECT 72.945 26.625 73.265 26.945 ;
        RECT 73.345 26.625 73.665 26.945 ;
        RECT 73.745 26.625 74.065 26.945 ;
        RECT 74.145 26.625 74.465 26.945 ;
        RECT 74.545 26.625 74.865 26.945 ;
        RECT 74.945 26.625 75.265 26.945 ;
        RECT 75.345 26.625 75.665 26.945 ;
        RECT 75.745 26.625 76.065 26.945 ;
        RECT 76.145 26.625 76.465 26.945 ;
        RECT 76.545 26.625 76.865 26.945 ;
        RECT 76.945 26.625 77.265 26.945 ;
        RECT 77.345 26.625 77.665 26.945 ;
        RECT 77.745 26.625 78.065 26.945 ;
        RECT 78.145 26.625 78.465 26.945 ;
        RECT 78.545 26.625 78.865 26.945 ;
        RECT 78.945 26.625 79.265 26.945 ;
        RECT 79.345 26.625 79.665 26.945 ;
        RECT 79.745 26.625 80.065 26.945 ;
        RECT 80.145 26.625 80.465 26.945 ;
        RECT 80.545 26.625 80.865 26.945 ;
        RECT 80.945 26.625 81.265 26.945 ;
        RECT 81.345 26.625 81.665 26.945 ;
        RECT 81.745 26.625 82.065 26.945 ;
        RECT 82.145 26.625 82.465 26.945 ;
        RECT 82.545 26.625 82.865 26.945 ;
        RECT 82.945 26.625 83.265 26.945 ;
        RECT 85.235 26.605 85.555 26.925 ;
        RECT 85.635 26.605 85.955 26.925 ;
        RECT 86.035 26.605 86.355 26.925 ;
        RECT 86.435 26.605 86.755 26.925 ;
        RECT 86.835 26.605 87.155 26.925 ;
        RECT 87.235 26.605 87.555 26.925 ;
        RECT 87.635 26.605 87.955 26.925 ;
        RECT 88.035 26.605 88.355 26.925 ;
        RECT 88.435 26.605 88.755 26.925 ;
        RECT 88.835 26.605 89.155 26.925 ;
        RECT 89.235 26.605 89.555 26.925 ;
        RECT 89.635 26.605 89.955 26.925 ;
        RECT 90.035 26.605 90.355 26.925 ;
        RECT 90.435 26.605 90.755 26.925 ;
        RECT 90.835 26.605 91.155 26.925 ;
        RECT 91.235 26.605 91.555 26.925 ;
        RECT 91.635 26.605 91.955 26.925 ;
        RECT 92.035 26.605 92.355 26.925 ;
        RECT 92.435 26.605 92.755 26.925 ;
        RECT 92.835 26.605 93.155 26.925 ;
        RECT 93.235 26.605 93.555 26.925 ;
        RECT 93.635 26.605 93.955 26.925 ;
        RECT 94.035 26.605 94.355 26.925 ;
        RECT 94.435 26.605 94.755 26.925 ;
        RECT 94.835 26.605 95.155 26.925 ;
        RECT 95.235 26.605 95.555 26.925 ;
        RECT 95.635 26.605 95.955 26.925 ;
        RECT 96.035 26.605 96.355 26.925 ;
        RECT 98.325 26.605 98.645 26.925 ;
        RECT 98.725 26.605 99.045 26.925 ;
        RECT 99.125 26.605 99.445 26.925 ;
        RECT 99.525 26.605 99.845 26.925 ;
        RECT 99.925 26.605 100.245 26.925 ;
        RECT 100.325 26.605 100.645 26.925 ;
        RECT 100.725 26.605 101.045 26.925 ;
        RECT 101.125 26.605 101.445 26.925 ;
        RECT 101.525 26.605 101.845 26.925 ;
        RECT 101.925 26.605 102.245 26.925 ;
        RECT 102.325 26.605 102.645 26.925 ;
        RECT 102.725 26.605 103.045 26.925 ;
        RECT 103.125 26.605 103.445 26.925 ;
        RECT 103.525 26.605 103.845 26.925 ;
        RECT 103.925 26.605 104.245 26.925 ;
        RECT 104.325 26.605 104.645 26.925 ;
        RECT 104.725 26.605 105.045 26.925 ;
        RECT 105.125 26.605 105.445 26.925 ;
        RECT 105.525 26.605 105.845 26.925 ;
        RECT 105.925 26.605 106.245 26.925 ;
        RECT 106.325 26.605 106.645 26.925 ;
        RECT 106.725 26.605 107.045 26.925 ;
        RECT 107.125 26.605 107.445 26.925 ;
        RECT 107.525 26.605 107.845 26.925 ;
        RECT 107.925 26.605 108.245 26.925 ;
        RECT 108.325 26.605 108.645 26.925 ;
        RECT 108.725 26.605 109.045 26.925 ;
        RECT 109.125 26.605 109.445 26.925 ;
        RECT 111.415 26.605 111.735 26.925 ;
        RECT 111.815 26.605 112.135 26.925 ;
        RECT 112.215 26.605 112.535 26.925 ;
        RECT 112.615 26.605 112.935 26.925 ;
        RECT 113.015 26.605 113.335 26.925 ;
        RECT 113.415 26.605 113.735 26.925 ;
        RECT 113.815 26.605 114.135 26.925 ;
        RECT 114.215 26.605 114.535 26.925 ;
        RECT 114.615 26.605 114.935 26.925 ;
        RECT 115.015 26.605 115.335 26.925 ;
        RECT 115.415 26.605 115.735 26.925 ;
        RECT 115.815 26.605 116.135 26.925 ;
        RECT 116.215 26.605 116.535 26.925 ;
        RECT 116.615 26.605 116.935 26.925 ;
        RECT 117.015 26.605 117.335 26.925 ;
        RECT 117.415 26.605 117.735 26.925 ;
        RECT 117.815 26.605 118.135 26.925 ;
        RECT 118.215 26.605 118.535 26.925 ;
        RECT 118.615 26.605 118.935 26.925 ;
        RECT 119.015 26.605 119.335 26.925 ;
        RECT 119.415 26.605 119.735 26.925 ;
        RECT 119.815 26.605 120.135 26.925 ;
        RECT 120.215 26.605 120.535 26.925 ;
        RECT 120.615 26.605 120.935 26.925 ;
        RECT 121.015 26.605 121.335 26.925 ;
        RECT 121.415 26.605 121.735 26.925 ;
        RECT 121.815 26.605 122.135 26.925 ;
        RECT 122.215 26.605 122.535 26.925 ;
        RECT 124.505 26.605 124.825 26.925 ;
        RECT 124.905 26.605 125.225 26.925 ;
        RECT 125.305 26.605 125.625 26.925 ;
        RECT 125.705 26.605 126.025 26.925 ;
        RECT 126.105 26.605 126.425 26.925 ;
        RECT 126.505 26.605 126.825 26.925 ;
        RECT 126.905 26.605 127.225 26.925 ;
        RECT 127.305 26.605 127.625 26.925 ;
        RECT 127.705 26.605 128.025 26.925 ;
        RECT 128.105 26.605 128.425 26.925 ;
        RECT 128.505 26.605 128.825 26.925 ;
        RECT 128.905 26.605 129.225 26.925 ;
        RECT 129.305 26.605 129.625 26.925 ;
        RECT 129.705 26.605 130.025 26.925 ;
        RECT 130.105 26.605 130.425 26.925 ;
        RECT 130.505 26.605 130.825 26.925 ;
        RECT 130.905 26.605 131.225 26.925 ;
        RECT 131.305 26.605 131.625 26.925 ;
        RECT 131.705 26.605 132.025 26.925 ;
        RECT 132.105 26.605 132.425 26.925 ;
        RECT 132.505 26.605 132.825 26.925 ;
        RECT 132.905 26.605 133.225 26.925 ;
        RECT 133.305 26.605 133.625 26.925 ;
        RECT 133.705 26.605 134.025 26.925 ;
        RECT 134.105 26.605 134.425 26.925 ;
        RECT 134.505 26.605 134.825 26.925 ;
        RECT 134.905 26.605 135.225 26.925 ;
        RECT 135.305 26.605 135.625 26.925 ;
        RECT 137.595 26.585 137.915 26.905 ;
        RECT 137.995 26.585 138.315 26.905 ;
        RECT 138.395 26.585 138.715 26.905 ;
        RECT 138.795 26.585 139.115 26.905 ;
        RECT 139.195 26.585 139.515 26.905 ;
        RECT 139.595 26.585 139.915 26.905 ;
        RECT 139.995 26.585 140.315 26.905 ;
        RECT 140.395 26.585 140.715 26.905 ;
        RECT 140.795 26.585 141.115 26.905 ;
        RECT 141.195 26.585 141.515 26.905 ;
        RECT 141.595 26.585 141.915 26.905 ;
        RECT 141.995 26.585 142.315 26.905 ;
        RECT 142.395 26.585 142.715 26.905 ;
        RECT 142.795 26.585 143.115 26.905 ;
        RECT 143.195 26.585 143.515 26.905 ;
        RECT 143.595 26.585 143.915 26.905 ;
        RECT 143.995 26.585 144.315 26.905 ;
        RECT 144.395 26.585 144.715 26.905 ;
        RECT 144.795 26.585 145.115 26.905 ;
        RECT 145.195 26.585 145.515 26.905 ;
        RECT 145.595 26.585 145.915 26.905 ;
        RECT 145.995 26.585 146.315 26.905 ;
        RECT 146.395 26.585 146.715 26.905 ;
        RECT 146.795 26.585 147.115 26.905 ;
        RECT 147.195 26.585 147.515 26.905 ;
        RECT 147.595 26.585 147.915 26.905 ;
        RECT 147.995 26.585 148.315 26.905 ;
        RECT 148.395 26.585 148.715 26.905 ;
        RECT 150.685 26.585 151.005 26.905 ;
        RECT 151.085 26.585 151.405 26.905 ;
        RECT 151.485 26.585 151.805 26.905 ;
        RECT 151.885 26.585 152.205 26.905 ;
        RECT 152.285 26.585 152.605 26.905 ;
        RECT 152.685 26.585 153.005 26.905 ;
        RECT 153.085 26.585 153.405 26.905 ;
        RECT 153.485 26.585 153.805 26.905 ;
        RECT 153.885 26.585 154.205 26.905 ;
        RECT 154.285 26.585 154.605 26.905 ;
        RECT 154.685 26.585 155.005 26.905 ;
        RECT 155.085 26.585 155.405 26.905 ;
        RECT 155.485 26.585 155.805 26.905 ;
        RECT 155.885 26.585 156.205 26.905 ;
        RECT 156.285 26.585 156.605 26.905 ;
        RECT 156.685 26.585 157.005 26.905 ;
        RECT 157.085 26.585 157.405 26.905 ;
        RECT 157.485 26.585 157.805 26.905 ;
        RECT 157.885 26.585 158.205 26.905 ;
        RECT 158.285 26.585 158.605 26.905 ;
        RECT 158.685 26.585 159.005 26.905 ;
        RECT 159.085 26.585 159.405 26.905 ;
        RECT 159.485 26.585 159.805 26.905 ;
        RECT 159.885 26.585 160.205 26.905 ;
        RECT 160.285 26.585 160.605 26.905 ;
        RECT 160.685 26.585 161.005 26.905 ;
        RECT 161.085 26.585 161.405 26.905 ;
        RECT 161.485 26.585 161.805 26.905 ;
        RECT 6.765 1.875 7.085 2.195 ;
        RECT 7.165 1.875 7.485 2.195 ;
        RECT 7.565 1.875 7.885 2.195 ;
        RECT 7.965 1.875 8.285 2.195 ;
        RECT 8.365 1.875 8.685 2.195 ;
        RECT 8.765 1.875 9.085 2.195 ;
        RECT 9.165 1.875 9.485 2.195 ;
        RECT 9.565 1.875 9.885 2.195 ;
        RECT 9.965 1.875 10.285 2.195 ;
        RECT 10.365 1.875 10.685 2.195 ;
        RECT 10.765 1.875 11.085 2.195 ;
        RECT 11.165 1.875 11.485 2.195 ;
        RECT 11.565 1.875 11.885 2.195 ;
        RECT 11.965 1.875 12.285 2.195 ;
        RECT 12.365 1.875 12.685 2.195 ;
        RECT 12.765 1.875 13.085 2.195 ;
        RECT 13.165 1.875 13.485 2.195 ;
        RECT 13.565 1.875 13.885 2.195 ;
        RECT 13.965 1.875 14.285 2.195 ;
        RECT 14.365 1.875 14.685 2.195 ;
        RECT 14.765 1.875 15.085 2.195 ;
        RECT 15.165 1.875 15.485 2.195 ;
        RECT 15.565 1.875 15.885 2.195 ;
        RECT 15.965 1.875 16.285 2.195 ;
        RECT 16.365 1.875 16.685 2.195 ;
        RECT 16.765 1.875 17.085 2.195 ;
        RECT 17.165 1.875 17.485 2.195 ;
        RECT 17.565 1.875 17.885 2.195 ;
        RECT 19.855 1.875 20.175 2.195 ;
        RECT 20.255 1.875 20.575 2.195 ;
        RECT 20.655 1.875 20.975 2.195 ;
        RECT 21.055 1.875 21.375 2.195 ;
        RECT 21.455 1.875 21.775 2.195 ;
        RECT 21.855 1.875 22.175 2.195 ;
        RECT 22.255 1.875 22.575 2.195 ;
        RECT 22.655 1.875 22.975 2.195 ;
        RECT 23.055 1.875 23.375 2.195 ;
        RECT 23.455 1.875 23.775 2.195 ;
        RECT 23.855 1.875 24.175 2.195 ;
        RECT 24.255 1.875 24.575 2.195 ;
        RECT 24.655 1.875 24.975 2.195 ;
        RECT 25.055 1.875 25.375 2.195 ;
        RECT 25.455 1.875 25.775 2.195 ;
        RECT 25.855 1.875 26.175 2.195 ;
        RECT 26.255 1.875 26.575 2.195 ;
        RECT 26.655 1.875 26.975 2.195 ;
        RECT 27.055 1.875 27.375 2.195 ;
        RECT 27.455 1.875 27.775 2.195 ;
        RECT 27.855 1.875 28.175 2.195 ;
        RECT 28.255 1.875 28.575 2.195 ;
        RECT 28.655 1.875 28.975 2.195 ;
        RECT 29.055 1.875 29.375 2.195 ;
        RECT 29.455 1.875 29.775 2.195 ;
        RECT 29.855 1.875 30.175 2.195 ;
        RECT 30.255 1.875 30.575 2.195 ;
        RECT 30.655 1.875 30.975 2.195 ;
        RECT 32.945 1.895 33.265 2.215 ;
        RECT 33.345 1.895 33.665 2.215 ;
        RECT 33.745 1.895 34.065 2.215 ;
        RECT 34.145 1.895 34.465 2.215 ;
        RECT 34.545 1.895 34.865 2.215 ;
        RECT 34.945 1.895 35.265 2.215 ;
        RECT 35.345 1.895 35.665 2.215 ;
        RECT 35.745 1.895 36.065 2.215 ;
        RECT 36.145 1.895 36.465 2.215 ;
        RECT 36.545 1.895 36.865 2.215 ;
        RECT 36.945 1.895 37.265 2.215 ;
        RECT 37.345 1.895 37.665 2.215 ;
        RECT 37.745 1.895 38.065 2.215 ;
        RECT 38.145 1.895 38.465 2.215 ;
        RECT 38.545 1.895 38.865 2.215 ;
        RECT 38.945 1.895 39.265 2.215 ;
        RECT 39.345 1.895 39.665 2.215 ;
        RECT 39.745 1.895 40.065 2.215 ;
        RECT 40.145 1.895 40.465 2.215 ;
        RECT 40.545 1.895 40.865 2.215 ;
        RECT 40.945 1.895 41.265 2.215 ;
        RECT 41.345 1.895 41.665 2.215 ;
        RECT 41.745 1.895 42.065 2.215 ;
        RECT 42.145 1.895 42.465 2.215 ;
        RECT 42.545 1.895 42.865 2.215 ;
        RECT 42.945 1.895 43.265 2.215 ;
        RECT 43.345 1.895 43.665 2.215 ;
        RECT 43.745 1.895 44.065 2.215 ;
        RECT 46.035 1.895 46.355 2.215 ;
        RECT 46.435 1.895 46.755 2.215 ;
        RECT 46.835 1.895 47.155 2.215 ;
        RECT 47.235 1.895 47.555 2.215 ;
        RECT 47.635 1.895 47.955 2.215 ;
        RECT 48.035 1.895 48.355 2.215 ;
        RECT 48.435 1.895 48.755 2.215 ;
        RECT 48.835 1.895 49.155 2.215 ;
        RECT 49.235 1.895 49.555 2.215 ;
        RECT 49.635 1.895 49.955 2.215 ;
        RECT 50.035 1.895 50.355 2.215 ;
        RECT 50.435 1.895 50.755 2.215 ;
        RECT 50.835 1.895 51.155 2.215 ;
        RECT 51.235 1.895 51.555 2.215 ;
        RECT 51.635 1.895 51.955 2.215 ;
        RECT 52.035 1.895 52.355 2.215 ;
        RECT 52.435 1.895 52.755 2.215 ;
        RECT 52.835 1.895 53.155 2.215 ;
        RECT 53.235 1.895 53.555 2.215 ;
        RECT 53.635 1.895 53.955 2.215 ;
        RECT 54.035 1.895 54.355 2.215 ;
        RECT 54.435 1.895 54.755 2.215 ;
        RECT 54.835 1.895 55.155 2.215 ;
        RECT 55.235 1.895 55.555 2.215 ;
        RECT 55.635 1.895 55.955 2.215 ;
        RECT 56.035 1.895 56.355 2.215 ;
        RECT 56.435 1.895 56.755 2.215 ;
        RECT 56.835 1.895 57.155 2.215 ;
        RECT 59.085 1.895 59.405 2.215 ;
        RECT 59.485 1.895 59.805 2.215 ;
        RECT 59.885 1.895 60.205 2.215 ;
        RECT 60.285 1.895 60.605 2.215 ;
        RECT 60.685 1.895 61.005 2.215 ;
        RECT 61.085 1.895 61.405 2.215 ;
        RECT 61.485 1.895 61.805 2.215 ;
        RECT 61.885 1.895 62.205 2.215 ;
        RECT 62.285 1.895 62.605 2.215 ;
        RECT 62.685 1.895 63.005 2.215 ;
        RECT 63.085 1.895 63.405 2.215 ;
        RECT 63.485 1.895 63.805 2.215 ;
        RECT 63.885 1.895 64.205 2.215 ;
        RECT 64.285 1.895 64.605 2.215 ;
        RECT 64.685 1.895 65.005 2.215 ;
        RECT 65.085 1.895 65.405 2.215 ;
        RECT 65.485 1.895 65.805 2.215 ;
        RECT 65.885 1.895 66.205 2.215 ;
        RECT 66.285 1.895 66.605 2.215 ;
        RECT 66.685 1.895 67.005 2.215 ;
        RECT 67.085 1.895 67.405 2.215 ;
        RECT 67.485 1.895 67.805 2.215 ;
        RECT 67.885 1.895 68.205 2.215 ;
        RECT 68.285 1.895 68.605 2.215 ;
        RECT 68.685 1.895 69.005 2.215 ;
        RECT 69.085 1.895 69.405 2.215 ;
        RECT 69.485 1.895 69.805 2.215 ;
        RECT 69.885 1.895 70.205 2.215 ;
        RECT 72.175 1.895 72.495 2.215 ;
        RECT 72.575 1.895 72.895 2.215 ;
        RECT 72.975 1.895 73.295 2.215 ;
        RECT 73.375 1.895 73.695 2.215 ;
        RECT 73.775 1.895 74.095 2.215 ;
        RECT 74.175 1.895 74.495 2.215 ;
        RECT 74.575 1.895 74.895 2.215 ;
        RECT 74.975 1.895 75.295 2.215 ;
        RECT 75.375 1.895 75.695 2.215 ;
        RECT 75.775 1.895 76.095 2.215 ;
        RECT 76.175 1.895 76.495 2.215 ;
        RECT 76.575 1.895 76.895 2.215 ;
        RECT 76.975 1.895 77.295 2.215 ;
        RECT 77.375 1.895 77.695 2.215 ;
        RECT 77.775 1.895 78.095 2.215 ;
        RECT 78.175 1.895 78.495 2.215 ;
        RECT 78.575 1.895 78.895 2.215 ;
        RECT 78.975 1.895 79.295 2.215 ;
        RECT 79.375 1.895 79.695 2.215 ;
        RECT 79.775 1.895 80.095 2.215 ;
        RECT 80.175 1.895 80.495 2.215 ;
        RECT 80.575 1.895 80.895 2.215 ;
        RECT 80.975 1.895 81.295 2.215 ;
        RECT 81.375 1.895 81.695 2.215 ;
        RECT 81.775 1.895 82.095 2.215 ;
        RECT 82.175 1.895 82.495 2.215 ;
        RECT 82.575 1.895 82.895 2.215 ;
        RECT 82.975 1.895 83.295 2.215 ;
        RECT 85.265 1.915 85.585 2.235 ;
        RECT 85.665 1.915 85.985 2.235 ;
        RECT 86.065 1.915 86.385 2.235 ;
        RECT 86.465 1.915 86.785 2.235 ;
        RECT 86.865 1.915 87.185 2.235 ;
        RECT 87.265 1.915 87.585 2.235 ;
        RECT 87.665 1.915 87.985 2.235 ;
        RECT 88.065 1.915 88.385 2.235 ;
        RECT 88.465 1.915 88.785 2.235 ;
        RECT 88.865 1.915 89.185 2.235 ;
        RECT 89.265 1.915 89.585 2.235 ;
        RECT 89.665 1.915 89.985 2.235 ;
        RECT 90.065 1.915 90.385 2.235 ;
        RECT 90.465 1.915 90.785 2.235 ;
        RECT 90.865 1.915 91.185 2.235 ;
        RECT 91.265 1.915 91.585 2.235 ;
        RECT 91.665 1.915 91.985 2.235 ;
        RECT 92.065 1.915 92.385 2.235 ;
        RECT 92.465 1.915 92.785 2.235 ;
        RECT 92.865 1.915 93.185 2.235 ;
        RECT 93.265 1.915 93.585 2.235 ;
        RECT 93.665 1.915 93.985 2.235 ;
        RECT 94.065 1.915 94.385 2.235 ;
        RECT 94.465 1.915 94.785 2.235 ;
        RECT 94.865 1.915 95.185 2.235 ;
        RECT 95.265 1.915 95.585 2.235 ;
        RECT 95.665 1.915 95.985 2.235 ;
        RECT 96.065 1.915 96.385 2.235 ;
        RECT 98.355 1.915 98.675 2.235 ;
        RECT 98.755 1.915 99.075 2.235 ;
        RECT 99.155 1.915 99.475 2.235 ;
        RECT 99.555 1.915 99.875 2.235 ;
        RECT 99.955 1.915 100.275 2.235 ;
        RECT 100.355 1.915 100.675 2.235 ;
        RECT 100.755 1.915 101.075 2.235 ;
        RECT 101.155 1.915 101.475 2.235 ;
        RECT 101.555 1.915 101.875 2.235 ;
        RECT 101.955 1.915 102.275 2.235 ;
        RECT 102.355 1.915 102.675 2.235 ;
        RECT 102.755 1.915 103.075 2.235 ;
        RECT 103.155 1.915 103.475 2.235 ;
        RECT 103.555 1.915 103.875 2.235 ;
        RECT 103.955 1.915 104.275 2.235 ;
        RECT 104.355 1.915 104.675 2.235 ;
        RECT 104.755 1.915 105.075 2.235 ;
        RECT 105.155 1.915 105.475 2.235 ;
        RECT 105.555 1.915 105.875 2.235 ;
        RECT 105.955 1.915 106.275 2.235 ;
        RECT 106.355 1.915 106.675 2.235 ;
        RECT 106.755 1.915 107.075 2.235 ;
        RECT 107.155 1.915 107.475 2.235 ;
        RECT 107.555 1.915 107.875 2.235 ;
        RECT 107.955 1.915 108.275 2.235 ;
        RECT 108.355 1.915 108.675 2.235 ;
        RECT 108.755 1.915 109.075 2.235 ;
        RECT 109.155 1.915 109.475 2.235 ;
        RECT 111.445 1.915 111.765 2.235 ;
        RECT 111.845 1.915 112.165 2.235 ;
        RECT 112.245 1.915 112.565 2.235 ;
        RECT 112.645 1.915 112.965 2.235 ;
        RECT 113.045 1.915 113.365 2.235 ;
        RECT 113.445 1.915 113.765 2.235 ;
        RECT 113.845 1.915 114.165 2.235 ;
        RECT 114.245 1.915 114.565 2.235 ;
        RECT 114.645 1.915 114.965 2.235 ;
        RECT 115.045 1.915 115.365 2.235 ;
        RECT 115.445 1.915 115.765 2.235 ;
        RECT 115.845 1.915 116.165 2.235 ;
        RECT 116.245 1.915 116.565 2.235 ;
        RECT 116.645 1.915 116.965 2.235 ;
        RECT 117.045 1.915 117.365 2.235 ;
        RECT 117.445 1.915 117.765 2.235 ;
        RECT 117.845 1.915 118.165 2.235 ;
        RECT 118.245 1.915 118.565 2.235 ;
        RECT 118.645 1.915 118.965 2.235 ;
        RECT 119.045 1.915 119.365 2.235 ;
        RECT 119.445 1.915 119.765 2.235 ;
        RECT 119.845 1.915 120.165 2.235 ;
        RECT 120.245 1.915 120.565 2.235 ;
        RECT 120.645 1.915 120.965 2.235 ;
        RECT 121.045 1.915 121.365 2.235 ;
        RECT 121.445 1.915 121.765 2.235 ;
        RECT 121.845 1.915 122.165 2.235 ;
        RECT 122.245 1.915 122.565 2.235 ;
        RECT 124.535 1.915 124.855 2.235 ;
        RECT 124.935 1.915 125.255 2.235 ;
        RECT 125.335 1.915 125.655 2.235 ;
        RECT 125.735 1.915 126.055 2.235 ;
        RECT 126.135 1.915 126.455 2.235 ;
        RECT 126.535 1.915 126.855 2.235 ;
        RECT 126.935 1.915 127.255 2.235 ;
        RECT 127.335 1.915 127.655 2.235 ;
        RECT 127.735 1.915 128.055 2.235 ;
        RECT 128.135 1.915 128.455 2.235 ;
        RECT 128.535 1.915 128.855 2.235 ;
        RECT 128.935 1.915 129.255 2.235 ;
        RECT 129.335 1.915 129.655 2.235 ;
        RECT 129.735 1.915 130.055 2.235 ;
        RECT 130.135 1.915 130.455 2.235 ;
        RECT 130.535 1.915 130.855 2.235 ;
        RECT 130.935 1.915 131.255 2.235 ;
        RECT 131.335 1.915 131.655 2.235 ;
        RECT 131.735 1.915 132.055 2.235 ;
        RECT 132.135 1.915 132.455 2.235 ;
        RECT 132.535 1.915 132.855 2.235 ;
        RECT 132.935 1.915 133.255 2.235 ;
        RECT 133.335 1.915 133.655 2.235 ;
        RECT 133.735 1.915 134.055 2.235 ;
        RECT 134.135 1.915 134.455 2.235 ;
        RECT 134.535 1.915 134.855 2.235 ;
        RECT 134.935 1.915 135.255 2.235 ;
        RECT 135.335 1.915 135.655 2.235 ;
        RECT 137.625 1.935 137.945 2.255 ;
        RECT 138.025 1.935 138.345 2.255 ;
        RECT 138.425 1.935 138.745 2.255 ;
        RECT 138.825 1.935 139.145 2.255 ;
        RECT 139.225 1.935 139.545 2.255 ;
        RECT 139.625 1.935 139.945 2.255 ;
        RECT 140.025 1.935 140.345 2.255 ;
        RECT 140.425 1.935 140.745 2.255 ;
        RECT 140.825 1.935 141.145 2.255 ;
        RECT 141.225 1.935 141.545 2.255 ;
        RECT 141.625 1.935 141.945 2.255 ;
        RECT 142.025 1.935 142.345 2.255 ;
        RECT 142.425 1.935 142.745 2.255 ;
        RECT 142.825 1.935 143.145 2.255 ;
        RECT 143.225 1.935 143.545 2.255 ;
        RECT 143.625 1.935 143.945 2.255 ;
        RECT 144.025 1.935 144.345 2.255 ;
        RECT 144.425 1.935 144.745 2.255 ;
        RECT 144.825 1.935 145.145 2.255 ;
        RECT 145.225 1.935 145.545 2.255 ;
        RECT 145.625 1.935 145.945 2.255 ;
        RECT 146.025 1.935 146.345 2.255 ;
        RECT 146.425 1.935 146.745 2.255 ;
        RECT 146.825 1.935 147.145 2.255 ;
        RECT 147.225 1.935 147.545 2.255 ;
        RECT 147.625 1.935 147.945 2.255 ;
        RECT 148.025 1.935 148.345 2.255 ;
        RECT 148.425 1.935 148.745 2.255 ;
        RECT 150.715 1.935 151.035 2.255 ;
        RECT 151.115 1.935 151.435 2.255 ;
        RECT 151.515 1.935 151.835 2.255 ;
        RECT 151.915 1.935 152.235 2.255 ;
        RECT 152.315 1.935 152.635 2.255 ;
        RECT 152.715 1.935 153.035 2.255 ;
        RECT 153.115 1.935 153.435 2.255 ;
        RECT 153.515 1.935 153.835 2.255 ;
        RECT 153.915 1.935 154.235 2.255 ;
        RECT 154.315 1.935 154.635 2.255 ;
        RECT 154.715 1.935 155.035 2.255 ;
        RECT 155.115 1.935 155.435 2.255 ;
        RECT 155.515 1.935 155.835 2.255 ;
        RECT 155.915 1.935 156.235 2.255 ;
        RECT 156.315 1.935 156.635 2.255 ;
        RECT 156.715 1.935 157.035 2.255 ;
        RECT 157.115 1.935 157.435 2.255 ;
        RECT 157.515 1.935 157.835 2.255 ;
        RECT 157.915 1.935 158.235 2.255 ;
        RECT 158.315 1.935 158.635 2.255 ;
        RECT 158.715 1.935 159.035 2.255 ;
        RECT 159.115 1.935 159.435 2.255 ;
        RECT 159.515 1.935 159.835 2.255 ;
        RECT 159.915 1.935 160.235 2.255 ;
        RECT 160.315 1.935 160.635 2.255 ;
        RECT 160.715 1.935 161.035 2.255 ;
        RECT 161.115 1.935 161.435 2.255 ;
        RECT 161.515 1.935 161.835 2.255 ;
      LAYER met4 ;
        RECT 1.415 118.260 3.015 119.860 ;
        RECT 6.155 118.280 17.565 118.610 ;
        RECT 19.245 118.280 30.655 118.610 ;
        RECT 1.615 93.440 2.815 118.260 ;
        RECT 6.755 117.055 8.255 118.280 ;
        RECT 6.755 107.550 7.055 117.055 ;
        RECT 7.955 108.775 8.255 117.055 ;
        RECT 9.155 107.550 9.455 118.280 ;
        RECT 10.355 107.550 10.655 118.280 ;
        RECT 11.555 107.550 11.855 118.280 ;
        RECT 12.755 107.550 13.055 118.280 ;
        RECT 13.955 117.055 15.455 118.280 ;
        RECT 13.955 107.550 14.255 117.055 ;
        RECT 15.155 108.775 15.455 117.055 ;
        RECT 16.355 107.550 16.655 118.280 ;
        RECT 19.845 117.055 21.345 118.280 ;
        RECT 19.845 107.550 20.145 117.055 ;
        RECT 21.045 108.775 21.345 117.055 ;
        RECT 22.245 107.550 22.545 118.280 ;
        RECT 23.445 107.550 23.745 118.280 ;
        RECT 24.645 107.550 24.945 118.280 ;
        RECT 25.845 107.550 26.145 118.280 ;
        RECT 27.045 117.055 28.545 118.280 ;
        RECT 27.045 107.550 27.345 117.055 ;
        RECT 28.245 108.775 28.545 117.055 ;
        RECT 29.445 107.550 29.745 118.280 ;
        RECT 32.335 118.260 43.745 118.590 ;
        RECT 45.425 118.260 56.835 118.590 ;
        RECT 58.475 118.260 69.885 118.590 ;
        RECT 71.565 118.260 82.975 118.590 ;
        RECT 32.935 117.035 34.435 118.260 ;
        RECT 32.935 107.530 33.235 117.035 ;
        RECT 34.135 108.755 34.435 117.035 ;
        RECT 35.335 107.530 35.635 118.260 ;
        RECT 36.535 107.530 36.835 118.260 ;
        RECT 37.735 107.530 38.035 118.260 ;
        RECT 38.935 107.530 39.235 118.260 ;
        RECT 40.135 117.035 41.635 118.260 ;
        RECT 40.135 107.530 40.435 117.035 ;
        RECT 41.335 108.755 41.635 117.035 ;
        RECT 42.535 107.530 42.835 118.260 ;
        RECT 46.025 117.035 47.525 118.260 ;
        RECT 46.025 107.530 46.325 117.035 ;
        RECT 47.225 108.755 47.525 117.035 ;
        RECT 48.425 107.530 48.725 118.260 ;
        RECT 49.625 107.530 49.925 118.260 ;
        RECT 50.825 107.530 51.125 118.260 ;
        RECT 52.025 107.530 52.325 118.260 ;
        RECT 53.225 117.035 54.725 118.260 ;
        RECT 53.225 107.530 53.525 117.035 ;
        RECT 54.425 108.755 54.725 117.035 ;
        RECT 55.625 107.530 55.925 118.260 ;
        RECT 59.075 117.035 60.575 118.260 ;
        RECT 59.075 107.530 59.375 117.035 ;
        RECT 60.275 108.755 60.575 117.035 ;
        RECT 61.475 107.530 61.775 118.260 ;
        RECT 62.675 107.530 62.975 118.260 ;
        RECT 63.875 107.530 64.175 118.260 ;
        RECT 65.075 107.530 65.375 118.260 ;
        RECT 66.275 117.035 67.775 118.260 ;
        RECT 66.275 107.530 66.575 117.035 ;
        RECT 67.475 108.755 67.775 117.035 ;
        RECT 68.675 107.530 68.975 118.260 ;
        RECT 72.165 117.035 73.665 118.260 ;
        RECT 72.165 107.530 72.465 117.035 ;
        RECT 73.365 108.755 73.665 117.035 ;
        RECT 74.565 107.530 74.865 118.260 ;
        RECT 75.765 107.530 76.065 118.260 ;
        RECT 76.965 107.530 77.265 118.260 ;
        RECT 78.165 107.530 78.465 118.260 ;
        RECT 79.365 117.035 80.865 118.260 ;
        RECT 79.365 107.530 79.665 117.035 ;
        RECT 80.565 108.755 80.865 117.035 ;
        RECT 81.765 107.530 82.065 118.260 ;
        RECT 84.655 118.240 96.065 118.570 ;
        RECT 97.745 118.240 109.155 118.570 ;
        RECT 110.835 118.240 122.245 118.570 ;
        RECT 123.925 118.240 135.335 118.570 ;
        RECT 85.255 117.015 86.755 118.240 ;
        RECT 85.255 107.510 85.555 117.015 ;
        RECT 86.455 108.735 86.755 117.015 ;
        RECT 87.655 107.510 87.955 118.240 ;
        RECT 88.855 107.510 89.155 118.240 ;
        RECT 90.055 107.510 90.355 118.240 ;
        RECT 91.255 107.510 91.555 118.240 ;
        RECT 92.455 117.015 93.955 118.240 ;
        RECT 92.455 107.510 92.755 117.015 ;
        RECT 93.655 108.735 93.955 117.015 ;
        RECT 94.855 107.510 95.155 118.240 ;
        RECT 98.345 117.015 99.845 118.240 ;
        RECT 98.345 107.510 98.645 117.015 ;
        RECT 99.545 108.735 99.845 117.015 ;
        RECT 100.745 107.510 101.045 118.240 ;
        RECT 101.945 107.510 102.245 118.240 ;
        RECT 103.145 107.510 103.445 118.240 ;
        RECT 104.345 107.510 104.645 118.240 ;
        RECT 105.545 117.015 107.045 118.240 ;
        RECT 105.545 107.510 105.845 117.015 ;
        RECT 106.745 108.735 107.045 117.015 ;
        RECT 107.945 107.510 108.245 118.240 ;
        RECT 111.435 117.015 112.935 118.240 ;
        RECT 111.435 107.510 111.735 117.015 ;
        RECT 112.635 108.735 112.935 117.015 ;
        RECT 113.835 107.510 114.135 118.240 ;
        RECT 115.035 107.510 115.335 118.240 ;
        RECT 116.235 107.510 116.535 118.240 ;
        RECT 117.435 107.510 117.735 118.240 ;
        RECT 118.635 117.015 120.135 118.240 ;
        RECT 118.635 107.510 118.935 117.015 ;
        RECT 119.835 108.735 120.135 117.015 ;
        RECT 121.035 107.510 121.335 118.240 ;
        RECT 124.525 117.015 126.025 118.240 ;
        RECT 124.525 107.510 124.825 117.015 ;
        RECT 125.725 108.735 126.025 117.015 ;
        RECT 126.925 107.510 127.225 118.240 ;
        RECT 128.125 107.510 128.425 118.240 ;
        RECT 129.325 107.510 129.625 118.240 ;
        RECT 130.525 107.510 130.825 118.240 ;
        RECT 131.725 117.015 133.225 118.240 ;
        RECT 131.725 107.510 132.025 117.015 ;
        RECT 132.925 108.735 133.225 117.015 ;
        RECT 134.125 107.510 134.425 118.240 ;
        RECT 137.015 118.220 148.425 118.550 ;
        RECT 150.105 118.220 161.515 118.550 ;
        RECT 137.615 116.995 139.115 118.220 ;
        RECT 137.615 107.490 137.915 116.995 ;
        RECT 138.815 108.715 139.115 116.995 ;
        RECT 140.015 107.490 140.315 118.220 ;
        RECT 141.215 107.490 141.515 118.220 ;
        RECT 142.415 107.490 142.715 118.220 ;
        RECT 143.615 107.490 143.915 118.220 ;
        RECT 144.815 116.995 146.315 118.220 ;
        RECT 144.815 107.490 145.115 116.995 ;
        RECT 146.015 108.715 146.315 116.995 ;
        RECT 147.215 107.490 147.515 118.220 ;
        RECT 150.705 116.995 152.205 118.220 ;
        RECT 150.705 107.490 151.005 116.995 ;
        RECT 151.905 108.715 152.205 116.995 ;
        RECT 153.105 107.490 153.405 118.220 ;
        RECT 154.305 107.490 154.605 118.220 ;
        RECT 155.505 107.490 155.805 118.220 ;
        RECT 156.705 107.490 157.005 118.220 ;
        RECT 157.905 116.995 159.405 118.220 ;
        RECT 157.905 107.490 158.205 116.995 ;
        RECT 159.105 108.715 159.405 116.995 ;
        RECT 160.305 107.490 160.605 118.220 ;
        RECT 166.775 118.210 168.375 119.810 ;
        RECT 6.785 95.065 7.085 104.570 ;
        RECT 7.985 95.065 8.285 103.345 ;
        RECT 6.785 93.840 8.285 95.065 ;
        RECT 9.185 93.840 9.485 104.570 ;
        RECT 10.385 93.840 10.685 104.570 ;
        RECT 11.585 93.840 11.885 104.570 ;
        RECT 12.785 93.840 13.085 104.570 ;
        RECT 13.985 95.065 14.285 104.570 ;
        RECT 15.185 95.065 15.485 103.345 ;
        RECT 13.985 93.840 15.485 95.065 ;
        RECT 16.385 93.840 16.685 104.570 ;
        RECT 19.875 95.065 20.175 104.570 ;
        RECT 21.075 95.065 21.375 103.345 ;
        RECT 19.875 93.840 21.375 95.065 ;
        RECT 22.275 93.840 22.575 104.570 ;
        RECT 23.475 93.840 23.775 104.570 ;
        RECT 24.675 93.840 24.975 104.570 ;
        RECT 25.875 93.840 26.175 104.570 ;
        RECT 27.075 95.065 27.375 104.570 ;
        RECT 28.275 95.065 28.575 103.345 ;
        RECT 27.075 93.840 28.575 95.065 ;
        RECT 29.475 93.840 29.775 104.570 ;
        RECT 32.965 95.085 33.265 104.590 ;
        RECT 34.165 95.085 34.465 103.365 ;
        RECT 32.965 93.860 34.465 95.085 ;
        RECT 35.365 93.860 35.665 104.590 ;
        RECT 36.565 93.860 36.865 104.590 ;
        RECT 37.765 93.860 38.065 104.590 ;
        RECT 38.965 93.860 39.265 104.590 ;
        RECT 40.165 95.085 40.465 104.590 ;
        RECT 41.365 95.085 41.665 103.365 ;
        RECT 40.165 93.860 41.665 95.085 ;
        RECT 42.565 93.860 42.865 104.590 ;
        RECT 46.055 95.085 46.355 104.590 ;
        RECT 47.255 95.085 47.555 103.365 ;
        RECT 46.055 93.860 47.555 95.085 ;
        RECT 48.455 93.860 48.755 104.590 ;
        RECT 49.655 93.860 49.955 104.590 ;
        RECT 50.855 93.860 51.155 104.590 ;
        RECT 52.055 93.860 52.355 104.590 ;
        RECT 53.255 95.085 53.555 104.590 ;
        RECT 54.455 95.085 54.755 103.365 ;
        RECT 53.255 93.860 54.755 95.085 ;
        RECT 55.655 93.860 55.955 104.590 ;
        RECT 59.105 95.085 59.405 104.590 ;
        RECT 60.305 95.085 60.605 103.365 ;
        RECT 59.105 93.860 60.605 95.085 ;
        RECT 61.505 93.860 61.805 104.590 ;
        RECT 62.705 93.860 63.005 104.590 ;
        RECT 63.905 93.860 64.205 104.590 ;
        RECT 65.105 93.860 65.405 104.590 ;
        RECT 66.305 95.085 66.605 104.590 ;
        RECT 67.505 95.085 67.805 103.365 ;
        RECT 66.305 93.860 67.805 95.085 ;
        RECT 68.705 93.860 69.005 104.590 ;
        RECT 72.195 95.085 72.495 104.590 ;
        RECT 73.395 95.085 73.695 103.365 ;
        RECT 72.195 93.860 73.695 95.085 ;
        RECT 74.595 93.860 74.895 104.590 ;
        RECT 75.795 93.860 76.095 104.590 ;
        RECT 76.995 93.860 77.295 104.590 ;
        RECT 78.195 93.860 78.495 104.590 ;
        RECT 79.395 95.085 79.695 104.590 ;
        RECT 80.595 95.085 80.895 103.365 ;
        RECT 79.395 93.860 80.895 95.085 ;
        RECT 81.795 93.860 82.095 104.590 ;
        RECT 85.285 95.105 85.585 104.610 ;
        RECT 86.485 95.105 86.785 103.385 ;
        RECT 85.285 93.880 86.785 95.105 ;
        RECT 87.685 93.880 87.985 104.610 ;
        RECT 88.885 93.880 89.185 104.610 ;
        RECT 90.085 93.880 90.385 104.610 ;
        RECT 91.285 93.880 91.585 104.610 ;
        RECT 92.485 95.105 92.785 104.610 ;
        RECT 93.685 95.105 93.985 103.385 ;
        RECT 92.485 93.880 93.985 95.105 ;
        RECT 94.885 93.880 95.185 104.610 ;
        RECT 98.375 95.105 98.675 104.610 ;
        RECT 99.575 95.105 99.875 103.385 ;
        RECT 98.375 93.880 99.875 95.105 ;
        RECT 100.775 93.880 101.075 104.610 ;
        RECT 101.975 93.880 102.275 104.610 ;
        RECT 103.175 93.880 103.475 104.610 ;
        RECT 104.375 93.880 104.675 104.610 ;
        RECT 105.575 95.105 105.875 104.610 ;
        RECT 106.775 95.105 107.075 103.385 ;
        RECT 105.575 93.880 107.075 95.105 ;
        RECT 107.975 93.880 108.275 104.610 ;
        RECT 111.465 95.105 111.765 104.610 ;
        RECT 112.665 95.105 112.965 103.385 ;
        RECT 111.465 93.880 112.965 95.105 ;
        RECT 113.865 93.880 114.165 104.610 ;
        RECT 115.065 93.880 115.365 104.610 ;
        RECT 116.265 93.880 116.565 104.610 ;
        RECT 117.465 93.880 117.765 104.610 ;
        RECT 118.665 95.105 118.965 104.610 ;
        RECT 119.865 95.105 120.165 103.385 ;
        RECT 118.665 93.880 120.165 95.105 ;
        RECT 121.065 93.880 121.365 104.610 ;
        RECT 124.555 95.105 124.855 104.610 ;
        RECT 125.755 95.105 126.055 103.385 ;
        RECT 124.555 93.880 126.055 95.105 ;
        RECT 126.955 93.880 127.255 104.610 ;
        RECT 128.155 93.880 128.455 104.610 ;
        RECT 129.355 93.880 129.655 104.610 ;
        RECT 130.555 93.880 130.855 104.610 ;
        RECT 131.755 95.105 132.055 104.610 ;
        RECT 132.955 95.105 133.255 103.385 ;
        RECT 131.755 93.880 133.255 95.105 ;
        RECT 134.155 93.880 134.455 104.610 ;
        RECT 137.645 95.125 137.945 104.630 ;
        RECT 138.845 95.125 139.145 103.405 ;
        RECT 137.645 93.900 139.145 95.125 ;
        RECT 140.045 93.900 140.345 104.630 ;
        RECT 141.245 93.900 141.545 104.630 ;
        RECT 142.445 93.900 142.745 104.630 ;
        RECT 143.645 93.900 143.945 104.630 ;
        RECT 144.845 95.125 145.145 104.630 ;
        RECT 146.045 95.125 146.345 103.405 ;
        RECT 144.845 93.900 146.345 95.125 ;
        RECT 147.245 93.900 147.545 104.630 ;
        RECT 150.735 95.125 151.035 104.630 ;
        RECT 151.935 95.125 152.235 103.405 ;
        RECT 150.735 93.900 152.235 95.125 ;
        RECT 153.135 93.900 153.435 104.630 ;
        RECT 154.335 93.900 154.635 104.630 ;
        RECT 155.535 93.900 155.835 104.630 ;
        RECT 156.735 93.900 157.035 104.630 ;
        RECT 157.935 95.125 158.235 104.630 ;
        RECT 159.135 95.125 159.435 103.405 ;
        RECT 157.935 93.900 159.435 95.125 ;
        RECT 160.335 93.900 160.635 104.630 ;
        RECT 6.185 93.510 17.595 93.840 ;
        RECT 19.275 93.510 30.685 93.840 ;
        RECT 32.365 93.530 43.775 93.860 ;
        RECT 45.455 93.530 56.865 93.860 ;
        RECT 58.505 93.530 69.915 93.860 ;
        RECT 71.595 93.530 83.005 93.860 ;
        RECT 84.685 93.550 96.095 93.880 ;
        RECT 97.775 93.550 109.185 93.880 ;
        RECT 110.865 93.550 122.275 93.880 ;
        RECT 123.955 93.550 135.365 93.880 ;
        RECT 137.045 93.570 148.455 93.900 ;
        RECT 150.135 93.570 161.545 93.900 ;
        RECT 166.975 93.630 168.175 118.210 ;
        RECT 1.415 91.840 3.015 93.440 ;
        RECT 166.775 92.030 168.375 93.630 ;
        RECT 1.615 28.310 2.815 91.840 ;
        RECT 166.975 89.160 168.175 92.030 ;
        RECT 1.415 1.000 3.015 28.310 ;
        RECT 165.735 28.070 166.935 30.790 ;
        RECT 6.595 26.640 18.005 26.970 ;
        RECT 19.685 26.640 31.095 26.970 ;
        RECT 7.195 25.415 8.695 26.640 ;
        RECT 7.195 15.910 7.495 25.415 ;
        RECT 8.395 17.135 8.695 25.415 ;
        RECT 9.595 15.910 9.895 26.640 ;
        RECT 10.795 15.910 11.095 26.640 ;
        RECT 11.995 15.910 12.295 26.640 ;
        RECT 13.195 15.910 13.495 26.640 ;
        RECT 14.395 25.415 15.895 26.640 ;
        RECT 14.395 15.910 14.695 25.415 ;
        RECT 15.595 17.135 15.895 25.415 ;
        RECT 16.795 15.910 17.095 26.640 ;
        RECT 20.285 25.415 21.785 26.640 ;
        RECT 20.285 15.910 20.585 25.415 ;
        RECT 21.485 17.135 21.785 25.415 ;
        RECT 22.685 15.910 22.985 26.640 ;
        RECT 23.885 15.910 24.185 26.640 ;
        RECT 25.085 15.910 25.385 26.640 ;
        RECT 26.285 15.910 26.585 26.640 ;
        RECT 27.485 25.415 28.985 26.640 ;
        RECT 27.485 15.910 27.785 25.415 ;
        RECT 28.685 17.135 28.985 25.415 ;
        RECT 29.885 15.910 30.185 26.640 ;
        RECT 32.775 26.620 44.185 26.950 ;
        RECT 45.865 26.620 57.275 26.950 ;
        RECT 58.915 26.620 70.325 26.950 ;
        RECT 72.005 26.620 83.415 26.950 ;
        RECT 33.375 25.395 34.875 26.620 ;
        RECT 33.375 15.890 33.675 25.395 ;
        RECT 34.575 17.115 34.875 25.395 ;
        RECT 35.775 15.890 36.075 26.620 ;
        RECT 36.975 15.890 37.275 26.620 ;
        RECT 38.175 15.890 38.475 26.620 ;
        RECT 39.375 15.890 39.675 26.620 ;
        RECT 40.575 25.395 42.075 26.620 ;
        RECT 40.575 15.890 40.875 25.395 ;
        RECT 41.775 17.115 42.075 25.395 ;
        RECT 42.975 15.890 43.275 26.620 ;
        RECT 46.465 25.395 47.965 26.620 ;
        RECT 46.465 15.890 46.765 25.395 ;
        RECT 47.665 17.115 47.965 25.395 ;
        RECT 48.865 15.890 49.165 26.620 ;
        RECT 50.065 15.890 50.365 26.620 ;
        RECT 51.265 15.890 51.565 26.620 ;
        RECT 52.465 15.890 52.765 26.620 ;
        RECT 53.665 25.395 55.165 26.620 ;
        RECT 53.665 15.890 53.965 25.395 ;
        RECT 54.865 17.115 55.165 25.395 ;
        RECT 56.065 15.890 56.365 26.620 ;
        RECT 59.515 25.395 61.015 26.620 ;
        RECT 59.515 15.890 59.815 25.395 ;
        RECT 60.715 17.115 61.015 25.395 ;
        RECT 61.915 15.890 62.215 26.620 ;
        RECT 63.115 15.890 63.415 26.620 ;
        RECT 64.315 15.890 64.615 26.620 ;
        RECT 65.515 15.890 65.815 26.620 ;
        RECT 66.715 25.395 68.215 26.620 ;
        RECT 66.715 15.890 67.015 25.395 ;
        RECT 67.915 17.115 68.215 25.395 ;
        RECT 69.115 15.890 69.415 26.620 ;
        RECT 72.605 25.395 74.105 26.620 ;
        RECT 72.605 15.890 72.905 25.395 ;
        RECT 73.805 17.115 74.105 25.395 ;
        RECT 75.005 15.890 75.305 26.620 ;
        RECT 76.205 15.890 76.505 26.620 ;
        RECT 77.405 15.890 77.705 26.620 ;
        RECT 78.605 15.890 78.905 26.620 ;
        RECT 79.805 25.395 81.305 26.620 ;
        RECT 79.805 15.890 80.105 25.395 ;
        RECT 81.005 17.115 81.305 25.395 ;
        RECT 82.205 15.890 82.505 26.620 ;
        RECT 85.095 26.600 96.505 26.930 ;
        RECT 98.185 26.600 109.595 26.930 ;
        RECT 111.275 26.600 122.685 26.930 ;
        RECT 124.365 26.600 135.775 26.930 ;
        RECT 85.695 25.375 87.195 26.600 ;
        RECT 85.695 15.870 85.995 25.375 ;
        RECT 86.895 17.095 87.195 25.375 ;
        RECT 88.095 15.870 88.395 26.600 ;
        RECT 89.295 15.870 89.595 26.600 ;
        RECT 90.495 15.870 90.795 26.600 ;
        RECT 91.695 15.870 91.995 26.600 ;
        RECT 92.895 25.375 94.395 26.600 ;
        RECT 92.895 15.870 93.195 25.375 ;
        RECT 94.095 17.095 94.395 25.375 ;
        RECT 95.295 15.870 95.595 26.600 ;
        RECT 98.785 25.375 100.285 26.600 ;
        RECT 98.785 15.870 99.085 25.375 ;
        RECT 99.985 17.095 100.285 25.375 ;
        RECT 101.185 15.870 101.485 26.600 ;
        RECT 102.385 15.870 102.685 26.600 ;
        RECT 103.585 15.870 103.885 26.600 ;
        RECT 104.785 15.870 105.085 26.600 ;
        RECT 105.985 25.375 107.485 26.600 ;
        RECT 105.985 15.870 106.285 25.375 ;
        RECT 107.185 17.095 107.485 25.375 ;
        RECT 108.385 15.870 108.685 26.600 ;
        RECT 111.875 25.375 113.375 26.600 ;
        RECT 111.875 15.870 112.175 25.375 ;
        RECT 113.075 17.095 113.375 25.375 ;
        RECT 114.275 15.870 114.575 26.600 ;
        RECT 115.475 15.870 115.775 26.600 ;
        RECT 116.675 15.870 116.975 26.600 ;
        RECT 117.875 15.870 118.175 26.600 ;
        RECT 119.075 25.375 120.575 26.600 ;
        RECT 119.075 15.870 119.375 25.375 ;
        RECT 120.275 17.095 120.575 25.375 ;
        RECT 121.475 15.870 121.775 26.600 ;
        RECT 124.965 25.375 126.465 26.600 ;
        RECT 124.965 15.870 125.265 25.375 ;
        RECT 126.165 17.095 126.465 25.375 ;
        RECT 127.365 15.870 127.665 26.600 ;
        RECT 128.565 15.870 128.865 26.600 ;
        RECT 129.765 15.870 130.065 26.600 ;
        RECT 130.965 15.870 131.265 26.600 ;
        RECT 132.165 25.375 133.665 26.600 ;
        RECT 132.165 15.870 132.465 25.375 ;
        RECT 133.365 17.095 133.665 25.375 ;
        RECT 134.565 15.870 134.865 26.600 ;
        RECT 137.455 26.580 148.865 26.910 ;
        RECT 150.545 26.580 161.955 26.910 ;
        RECT 138.055 25.355 139.555 26.580 ;
        RECT 138.055 15.850 138.355 25.355 ;
        RECT 139.255 17.075 139.555 25.355 ;
        RECT 140.455 15.850 140.755 26.580 ;
        RECT 141.655 15.850 141.955 26.580 ;
        RECT 142.855 15.850 143.155 26.580 ;
        RECT 144.055 15.850 144.355 26.580 ;
        RECT 145.255 25.355 146.755 26.580 ;
        RECT 145.255 15.850 145.555 25.355 ;
        RECT 146.455 17.075 146.755 25.355 ;
        RECT 147.655 15.850 147.955 26.580 ;
        RECT 151.145 25.355 152.645 26.580 ;
        RECT 151.145 15.850 151.445 25.355 ;
        RECT 152.345 17.075 152.645 25.355 ;
        RECT 153.545 15.850 153.845 26.580 ;
        RECT 154.745 15.850 155.045 26.580 ;
        RECT 155.945 15.850 156.245 26.580 ;
        RECT 157.145 15.850 157.445 26.580 ;
        RECT 158.345 25.355 159.845 26.580 ;
        RECT 158.345 15.850 158.645 25.355 ;
        RECT 159.545 17.075 159.845 25.355 ;
        RECT 160.745 15.850 161.045 26.580 ;
        RECT 165.535 26.470 167.135 28.070 ;
        RECT 7.225 3.425 7.525 12.930 ;
        RECT 8.425 3.425 8.725 11.705 ;
        RECT 7.225 2.200 8.725 3.425 ;
        RECT 9.625 2.200 9.925 12.930 ;
        RECT 10.825 2.200 11.125 12.930 ;
        RECT 12.025 2.200 12.325 12.930 ;
        RECT 13.225 2.200 13.525 12.930 ;
        RECT 14.425 3.425 14.725 12.930 ;
        RECT 15.625 3.425 15.925 11.705 ;
        RECT 14.425 2.200 15.925 3.425 ;
        RECT 16.825 2.200 17.125 12.930 ;
        RECT 20.315 3.425 20.615 12.930 ;
        RECT 21.515 3.425 21.815 11.705 ;
        RECT 20.315 2.200 21.815 3.425 ;
        RECT 22.715 2.200 23.015 12.930 ;
        RECT 23.915 2.200 24.215 12.930 ;
        RECT 25.115 2.200 25.415 12.930 ;
        RECT 26.315 2.200 26.615 12.930 ;
        RECT 27.515 3.425 27.815 12.930 ;
        RECT 28.715 3.425 29.015 11.705 ;
        RECT 27.515 2.200 29.015 3.425 ;
        RECT 29.915 2.200 30.215 12.930 ;
        RECT 33.405 3.445 33.705 12.950 ;
        RECT 34.605 3.445 34.905 11.725 ;
        RECT 33.405 2.220 34.905 3.445 ;
        RECT 35.805 2.220 36.105 12.950 ;
        RECT 37.005 2.220 37.305 12.950 ;
        RECT 38.205 2.220 38.505 12.950 ;
        RECT 39.405 2.220 39.705 12.950 ;
        RECT 40.605 3.445 40.905 12.950 ;
        RECT 41.805 3.445 42.105 11.725 ;
        RECT 40.605 2.220 42.105 3.445 ;
        RECT 43.005 2.220 43.305 12.950 ;
        RECT 46.495 3.445 46.795 12.950 ;
        RECT 47.695 3.445 47.995 11.725 ;
        RECT 46.495 2.220 47.995 3.445 ;
        RECT 48.895 2.220 49.195 12.950 ;
        RECT 50.095 2.220 50.395 12.950 ;
        RECT 51.295 2.220 51.595 12.950 ;
        RECT 52.495 2.220 52.795 12.950 ;
        RECT 53.695 3.445 53.995 12.950 ;
        RECT 54.895 3.445 55.195 11.725 ;
        RECT 53.695 2.220 55.195 3.445 ;
        RECT 56.095 2.220 56.395 12.950 ;
        RECT 59.545 3.445 59.845 12.950 ;
        RECT 60.745 3.445 61.045 11.725 ;
        RECT 59.545 2.220 61.045 3.445 ;
        RECT 61.945 2.220 62.245 12.950 ;
        RECT 63.145 2.220 63.445 12.950 ;
        RECT 64.345 2.220 64.645 12.950 ;
        RECT 65.545 2.220 65.845 12.950 ;
        RECT 66.745 3.445 67.045 12.950 ;
        RECT 67.945 3.445 68.245 11.725 ;
        RECT 66.745 2.220 68.245 3.445 ;
        RECT 69.145 2.220 69.445 12.950 ;
        RECT 72.635 3.445 72.935 12.950 ;
        RECT 73.835 3.445 74.135 11.725 ;
        RECT 72.635 2.220 74.135 3.445 ;
        RECT 75.035 2.220 75.335 12.950 ;
        RECT 76.235 2.220 76.535 12.950 ;
        RECT 77.435 2.220 77.735 12.950 ;
        RECT 78.635 2.220 78.935 12.950 ;
        RECT 79.835 3.445 80.135 12.950 ;
        RECT 81.035 3.445 81.335 11.725 ;
        RECT 79.835 2.220 81.335 3.445 ;
        RECT 82.235 2.220 82.535 12.950 ;
        RECT 85.725 3.465 86.025 12.970 ;
        RECT 86.925 3.465 87.225 11.745 ;
        RECT 85.725 2.240 87.225 3.465 ;
        RECT 88.125 2.240 88.425 12.970 ;
        RECT 89.325 2.240 89.625 12.970 ;
        RECT 90.525 2.240 90.825 12.970 ;
        RECT 91.725 2.240 92.025 12.970 ;
        RECT 92.925 3.465 93.225 12.970 ;
        RECT 94.125 3.465 94.425 11.745 ;
        RECT 92.925 2.240 94.425 3.465 ;
        RECT 95.325 2.240 95.625 12.970 ;
        RECT 98.815 3.465 99.115 12.970 ;
        RECT 100.015 3.465 100.315 11.745 ;
        RECT 98.815 2.240 100.315 3.465 ;
        RECT 101.215 2.240 101.515 12.970 ;
        RECT 102.415 2.240 102.715 12.970 ;
        RECT 103.615 2.240 103.915 12.970 ;
        RECT 104.815 2.240 105.115 12.970 ;
        RECT 106.015 3.465 106.315 12.970 ;
        RECT 107.215 3.465 107.515 11.745 ;
        RECT 106.015 2.240 107.515 3.465 ;
        RECT 108.415 2.240 108.715 12.970 ;
        RECT 111.905 3.465 112.205 12.970 ;
        RECT 113.105 3.465 113.405 11.745 ;
        RECT 111.905 2.240 113.405 3.465 ;
        RECT 114.305 2.240 114.605 12.970 ;
        RECT 115.505 2.240 115.805 12.970 ;
        RECT 116.705 2.240 117.005 12.970 ;
        RECT 117.905 2.240 118.205 12.970 ;
        RECT 119.105 3.465 119.405 12.970 ;
        RECT 120.305 3.465 120.605 11.745 ;
        RECT 119.105 2.240 120.605 3.465 ;
        RECT 121.505 2.240 121.805 12.970 ;
        RECT 124.995 3.465 125.295 12.970 ;
        RECT 126.195 3.465 126.495 11.745 ;
        RECT 124.995 2.240 126.495 3.465 ;
        RECT 127.395 2.240 127.695 12.970 ;
        RECT 128.595 2.240 128.895 12.970 ;
        RECT 129.795 2.240 130.095 12.970 ;
        RECT 130.995 2.240 131.295 12.970 ;
        RECT 132.195 3.465 132.495 12.970 ;
        RECT 133.395 3.465 133.695 11.745 ;
        RECT 132.195 2.240 133.695 3.465 ;
        RECT 134.595 2.240 134.895 12.970 ;
        RECT 138.085 3.485 138.385 12.990 ;
        RECT 139.285 3.485 139.585 11.765 ;
        RECT 138.085 2.260 139.585 3.485 ;
        RECT 140.485 2.260 140.785 12.990 ;
        RECT 141.685 2.260 141.985 12.990 ;
        RECT 142.885 2.260 143.185 12.990 ;
        RECT 144.085 2.260 144.385 12.990 ;
        RECT 145.285 3.485 145.585 12.990 ;
        RECT 146.485 3.485 146.785 11.765 ;
        RECT 145.285 2.260 146.785 3.485 ;
        RECT 147.685 2.260 147.985 12.990 ;
        RECT 151.175 3.485 151.475 12.990 ;
        RECT 152.375 3.485 152.675 11.765 ;
        RECT 151.175 2.260 152.675 3.485 ;
        RECT 153.575 2.260 153.875 12.990 ;
        RECT 154.775 2.260 155.075 12.990 ;
        RECT 155.975 2.260 156.275 12.990 ;
        RECT 157.175 2.260 157.475 12.990 ;
        RECT 158.375 3.485 158.675 12.990 ;
        RECT 159.575 3.485 159.875 11.765 ;
        RECT 158.375 2.260 159.875 3.485 ;
        RECT 160.775 2.260 161.075 12.990 ;
        RECT 6.625 1.870 18.035 2.200 ;
        RECT 19.715 1.870 31.125 2.200 ;
        RECT 32.805 1.890 44.215 2.220 ;
        RECT 45.895 1.890 57.305 2.220 ;
        RECT 58.945 1.890 70.355 2.220 ;
        RECT 72.035 1.890 83.445 2.220 ;
        RECT 85.125 1.910 96.535 2.240 ;
        RECT 98.215 1.910 109.625 2.240 ;
        RECT 111.305 1.910 122.715 2.240 ;
        RECT 124.395 1.910 135.805 2.240 ;
        RECT 137.485 1.930 148.895 2.260 ;
        RECT 150.575 1.930 161.985 2.260 ;
        RECT 165.735 2.250 166.935 26.470 ;
        RECT 165.535 0.650 167.135 2.250 ;
      LAYER via4 ;
        RECT 6.915 117.055 8.095 118.235 ;
        RECT 14.115 117.055 15.295 118.235 ;
        RECT 20.005 117.055 21.185 118.235 ;
        RECT 27.205 117.055 28.385 118.235 ;
        RECT 33.095 117.035 34.275 118.215 ;
        RECT 40.295 117.035 41.475 118.215 ;
        RECT 46.185 117.035 47.365 118.215 ;
        RECT 53.385 117.035 54.565 118.215 ;
        RECT 59.235 117.035 60.415 118.215 ;
        RECT 66.435 117.035 67.615 118.215 ;
        RECT 72.325 117.035 73.505 118.215 ;
        RECT 79.525 117.035 80.705 118.215 ;
        RECT 85.415 117.015 86.595 118.195 ;
        RECT 92.615 117.015 93.795 118.195 ;
        RECT 98.505 117.015 99.685 118.195 ;
        RECT 105.705 117.015 106.885 118.195 ;
        RECT 111.595 117.015 112.775 118.195 ;
        RECT 118.795 117.015 119.975 118.195 ;
        RECT 124.685 117.015 125.865 118.195 ;
        RECT 131.885 117.015 133.065 118.195 ;
        RECT 137.775 116.995 138.955 118.175 ;
        RECT 144.975 116.995 146.155 118.175 ;
        RECT 150.865 116.995 152.045 118.175 ;
        RECT 158.065 116.995 159.245 118.175 ;
        RECT 6.945 93.885 8.125 95.065 ;
        RECT 14.145 93.885 15.325 95.065 ;
        RECT 20.035 93.885 21.215 95.065 ;
        RECT 27.235 93.885 28.415 95.065 ;
        RECT 33.125 93.905 34.305 95.085 ;
        RECT 40.325 93.905 41.505 95.085 ;
        RECT 46.215 93.905 47.395 95.085 ;
        RECT 53.415 93.905 54.595 95.085 ;
        RECT 59.265 93.905 60.445 95.085 ;
        RECT 66.465 93.905 67.645 95.085 ;
        RECT 72.355 93.905 73.535 95.085 ;
        RECT 79.555 93.905 80.735 95.085 ;
        RECT 85.445 93.925 86.625 95.105 ;
        RECT 92.645 93.925 93.825 95.105 ;
        RECT 98.535 93.925 99.715 95.105 ;
        RECT 105.735 93.925 106.915 95.105 ;
        RECT 111.625 93.925 112.805 95.105 ;
        RECT 118.825 93.925 120.005 95.105 ;
        RECT 124.715 93.925 125.895 95.105 ;
        RECT 131.915 93.925 133.095 95.105 ;
        RECT 137.805 93.945 138.985 95.125 ;
        RECT 145.005 93.945 146.185 95.125 ;
        RECT 150.895 93.945 152.075 95.125 ;
        RECT 158.095 93.945 159.275 95.125 ;
        RECT 1.415 26.710 3.015 28.310 ;
        RECT 7.355 25.415 8.535 26.595 ;
        RECT 14.555 25.415 15.735 26.595 ;
        RECT 20.445 25.415 21.625 26.595 ;
        RECT 27.645 25.415 28.825 26.595 ;
        RECT 33.535 25.395 34.715 26.575 ;
        RECT 40.735 25.395 41.915 26.575 ;
        RECT 46.625 25.395 47.805 26.575 ;
        RECT 53.825 25.395 55.005 26.575 ;
        RECT 59.675 25.395 60.855 26.575 ;
        RECT 66.875 25.395 68.055 26.575 ;
        RECT 72.765 25.395 73.945 26.575 ;
        RECT 79.965 25.395 81.145 26.575 ;
        RECT 85.855 25.375 87.035 26.555 ;
        RECT 93.055 25.375 94.235 26.555 ;
        RECT 98.945 25.375 100.125 26.555 ;
        RECT 106.145 25.375 107.325 26.555 ;
        RECT 112.035 25.375 113.215 26.555 ;
        RECT 119.235 25.375 120.415 26.555 ;
        RECT 125.125 25.375 126.305 26.555 ;
        RECT 132.325 25.375 133.505 26.555 ;
        RECT 138.215 25.355 139.395 26.535 ;
        RECT 145.415 25.355 146.595 26.535 ;
        RECT 151.305 25.355 152.485 26.535 ;
        RECT 158.505 25.355 159.685 26.535 ;
        RECT 7.385 2.245 8.565 3.425 ;
        RECT 14.585 2.245 15.765 3.425 ;
        RECT 20.475 2.245 21.655 3.425 ;
        RECT 27.675 2.245 28.855 3.425 ;
        RECT 33.565 2.265 34.745 3.445 ;
        RECT 40.765 2.265 41.945 3.445 ;
        RECT 46.655 2.265 47.835 3.445 ;
        RECT 53.855 2.265 55.035 3.445 ;
        RECT 59.705 2.265 60.885 3.445 ;
        RECT 66.905 2.265 68.085 3.445 ;
        RECT 72.795 2.265 73.975 3.445 ;
        RECT 79.995 2.265 81.175 3.445 ;
        RECT 85.885 2.285 87.065 3.465 ;
        RECT 93.085 2.285 94.265 3.465 ;
        RECT 98.975 2.285 100.155 3.465 ;
        RECT 106.175 2.285 107.355 3.465 ;
        RECT 112.065 2.285 113.245 3.465 ;
        RECT 119.265 2.285 120.445 3.465 ;
        RECT 125.155 2.285 126.335 3.465 ;
        RECT 132.355 2.285 133.535 3.465 ;
        RECT 138.245 2.305 139.425 3.485 ;
        RECT 145.445 2.305 146.625 3.485 ;
        RECT 151.335 2.305 152.515 3.485 ;
        RECT 158.535 2.305 159.715 3.485 ;
      LAYER met5 ;
        RECT 0.000 117.500 169.120 120.810 ;
        RECT 6.155 116.935 17.565 117.500 ;
        RECT 19.245 116.935 30.655 117.500 ;
        RECT 6.155 110.195 7.755 116.935 ;
        RECT 12.555 110.195 14.155 116.935 ;
        RECT 19.245 110.195 20.845 116.935 ;
        RECT 25.645 110.195 27.245 116.935 ;
        RECT 32.335 116.915 43.745 117.500 ;
        RECT 45.425 116.915 56.835 117.500 ;
        RECT 58.475 116.915 69.885 117.500 ;
        RECT 71.565 116.915 82.975 117.500 ;
        RECT 32.335 110.175 33.935 116.915 ;
        RECT 38.735 110.175 40.335 116.915 ;
        RECT 45.425 110.175 47.025 116.915 ;
        RECT 51.825 110.175 53.425 116.915 ;
        RECT 58.475 110.175 60.075 116.915 ;
        RECT 64.875 110.175 66.475 116.915 ;
        RECT 71.565 110.175 73.165 116.915 ;
        RECT 77.965 110.175 79.565 116.915 ;
        RECT 84.655 116.895 96.065 117.500 ;
        RECT 97.745 116.895 109.155 117.500 ;
        RECT 110.835 116.895 122.245 117.500 ;
        RECT 123.925 116.895 135.335 117.500 ;
        RECT 84.655 110.155 86.255 116.895 ;
        RECT 91.055 110.155 92.655 116.895 ;
        RECT 97.745 110.155 99.345 116.895 ;
        RECT 104.145 110.155 105.745 116.895 ;
        RECT 110.835 110.155 112.435 116.895 ;
        RECT 117.235 110.155 118.835 116.895 ;
        RECT 123.925 110.155 125.525 116.895 ;
        RECT 130.325 110.155 131.925 116.895 ;
        RECT 137.015 116.875 148.425 117.500 ;
        RECT 150.105 116.875 161.515 117.500 ;
        RECT 137.015 110.135 138.615 116.875 ;
        RECT 143.415 110.135 145.015 116.875 ;
        RECT 150.105 110.135 151.705 116.875 ;
        RECT 156.505 110.135 158.105 116.875 ;
        RECT 6.185 95.185 7.785 101.925 ;
        RECT 12.585 95.185 14.185 101.925 ;
        RECT 19.275 95.185 20.875 101.925 ;
        RECT 25.675 95.185 27.275 101.925 ;
        RECT 32.365 95.205 33.965 101.945 ;
        RECT 38.765 95.205 40.365 101.945 ;
        RECT 45.455 95.205 47.055 101.945 ;
        RECT 51.855 95.205 53.455 101.945 ;
        RECT 58.505 95.205 60.105 101.945 ;
        RECT 64.905 95.205 66.505 101.945 ;
        RECT 71.595 95.205 73.195 101.945 ;
        RECT 77.995 95.205 79.595 101.945 ;
        RECT 84.685 95.225 86.285 101.965 ;
        RECT 91.085 95.225 92.685 101.965 ;
        RECT 97.775 95.225 99.375 101.965 ;
        RECT 104.175 95.225 105.775 101.965 ;
        RECT 110.865 95.225 112.465 101.965 ;
        RECT 117.265 95.225 118.865 101.965 ;
        RECT 123.955 95.225 125.555 101.965 ;
        RECT 130.355 95.225 131.955 101.965 ;
        RECT 137.045 95.245 138.645 101.985 ;
        RECT 143.445 95.245 145.045 101.985 ;
        RECT 150.135 95.245 151.735 101.985 ;
        RECT 156.535 95.245 158.135 101.985 ;
        RECT 6.185 94.550 17.595 95.185 ;
        RECT 19.275 94.550 30.685 95.185 ;
        RECT 32.365 94.550 43.775 95.205 ;
        RECT 45.455 94.550 56.865 95.205 ;
        RECT 58.505 94.550 69.915 95.205 ;
        RECT 71.595 94.550 83.005 95.205 ;
        RECT 84.685 94.550 96.095 95.225 ;
        RECT 97.775 94.550 109.185 95.225 ;
        RECT 110.865 94.550 122.275 95.225 ;
        RECT 123.955 94.550 135.365 95.225 ;
        RECT 137.045 94.550 148.455 95.245 ;
        RECT 150.135 94.550 161.545 95.245 ;
        RECT 0.570 91.240 169.320 94.550 ;
        RECT 0.800 25.690 167.540 29.000 ;
        RECT 6.595 25.295 18.005 25.690 ;
        RECT 19.685 25.295 31.095 25.690 ;
        RECT 6.595 18.555 8.195 25.295 ;
        RECT 12.995 18.555 14.595 25.295 ;
        RECT 19.685 18.555 21.285 25.295 ;
        RECT 26.085 18.555 27.685 25.295 ;
        RECT 32.775 25.275 44.185 25.690 ;
        RECT 45.865 25.275 57.275 25.690 ;
        RECT 58.915 25.275 70.325 25.690 ;
        RECT 72.005 25.275 83.415 25.690 ;
        RECT 32.775 18.535 34.375 25.275 ;
        RECT 39.175 18.535 40.775 25.275 ;
        RECT 45.865 18.535 47.465 25.275 ;
        RECT 52.265 18.535 53.865 25.275 ;
        RECT 58.915 18.535 60.515 25.275 ;
        RECT 65.315 18.535 66.915 25.275 ;
        RECT 72.005 18.535 73.605 25.275 ;
        RECT 78.405 18.535 80.005 25.275 ;
        RECT 85.095 25.255 96.505 25.690 ;
        RECT 98.185 25.255 109.595 25.690 ;
        RECT 111.275 25.255 122.685 25.690 ;
        RECT 124.365 25.255 135.775 25.690 ;
        RECT 85.095 18.515 86.695 25.255 ;
        RECT 91.495 18.515 93.095 25.255 ;
        RECT 98.185 18.515 99.785 25.255 ;
        RECT 104.585 18.515 106.185 25.255 ;
        RECT 111.275 18.515 112.875 25.255 ;
        RECT 117.675 18.515 119.275 25.255 ;
        RECT 124.365 18.515 125.965 25.255 ;
        RECT 130.765 18.515 132.365 25.255 ;
        RECT 137.455 25.235 148.865 25.690 ;
        RECT 150.545 25.235 161.955 25.690 ;
        RECT 137.455 18.495 139.055 25.235 ;
        RECT 143.855 18.495 145.455 25.235 ;
        RECT 150.545 18.495 152.145 25.235 ;
        RECT 156.945 18.495 158.545 25.235 ;
        RECT 6.625 3.545 8.225 10.285 ;
        RECT 13.025 3.545 14.625 10.285 ;
        RECT 19.715 3.545 21.315 10.285 ;
        RECT 26.115 3.545 27.715 10.285 ;
        RECT 32.805 3.565 34.405 10.305 ;
        RECT 39.205 3.565 40.805 10.305 ;
        RECT 45.895 3.565 47.495 10.305 ;
        RECT 52.295 3.565 53.895 10.305 ;
        RECT 58.945 3.565 60.545 10.305 ;
        RECT 65.345 3.565 66.945 10.305 ;
        RECT 72.035 3.565 73.635 10.305 ;
        RECT 78.435 3.565 80.035 10.305 ;
        RECT 85.125 3.585 86.725 10.325 ;
        RECT 91.525 3.585 93.125 10.325 ;
        RECT 98.215 3.585 99.815 10.325 ;
        RECT 104.615 3.585 106.215 10.325 ;
        RECT 111.305 3.585 112.905 10.325 ;
        RECT 117.705 3.585 119.305 10.325 ;
        RECT 124.395 3.585 125.995 10.325 ;
        RECT 130.795 3.585 132.395 10.325 ;
        RECT 137.485 3.605 139.085 10.345 ;
        RECT 143.885 3.605 145.485 10.345 ;
        RECT 150.575 3.605 152.175 10.345 ;
        RECT 156.975 3.605 158.575 10.345 ;
        RECT 6.625 3.310 18.035 3.545 ;
        RECT 19.715 3.310 31.125 3.545 ;
        RECT 32.805 3.310 44.215 3.565 ;
        RECT 45.895 3.310 57.305 3.565 ;
        RECT 58.945 3.310 70.355 3.565 ;
        RECT 72.035 3.310 83.445 3.565 ;
        RECT 85.125 3.310 96.535 3.585 ;
        RECT 98.215 3.310 109.625 3.585 ;
        RECT 111.305 3.310 122.715 3.585 ;
        RECT 124.395 3.310 135.805 3.585 ;
        RECT 137.485 3.310 148.895 3.605 ;
        RECT 150.575 3.310 161.985 3.605 ;
        RECT 0.590 0.000 167.850 3.310 ;
    END
  END avdd
  PIN avss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 11.435 75.560 19.005 78.350 ;
        RECT 21.050 75.560 28.620 78.350 ;
        RECT 30.665 75.560 38.235 78.350 ;
        RECT 40.280 75.560 47.850 78.350 ;
        RECT 149.840 67.215 156.230 70.005 ;
        RECT 157.830 67.215 161.860 70.005 ;
        RECT 162.735 67.215 165.585 70.005 ;
        RECT 165.855 67.545 168.645 69.805 ;
        RECT 168.650 67.610 171.440 69.870 ;
        RECT 171.635 66.040 174.905 66.470 ;
        RECT 152.955 61.235 155.215 62.385 ;
        RECT 155.245 61.235 157.505 62.410 ;
        RECT 152.955 61.055 157.505 61.235 ;
        RECT 152.955 57.815 155.215 61.055 ;
        RECT 155.245 57.840 157.505 61.055 ;
        RECT 157.545 57.855 159.805 62.425 ;
        RECT 171.635 55.470 172.065 66.040 ;
        RECT 174.475 55.470 174.905 66.040 ;
        RECT 171.635 55.040 174.905 55.470 ;
        RECT 149.955 49.975 156.345 52.765 ;
        RECT 157.945 49.975 161.975 52.765 ;
        RECT 162.850 49.975 165.700 52.765 ;
        RECT 165.970 50.175 168.760 52.435 ;
        RECT 168.765 50.110 171.555 52.370 ;
        RECT 11.435 41.500 19.005 44.290 ;
        RECT 21.050 41.500 28.620 44.290 ;
        RECT 30.665 41.500 38.235 44.290 ;
        RECT 40.280 41.500 47.850 44.290 ;
      LAYER li1 ;
        RECT 147.625 88.460 147.795 89.490 ;
        RECT 147.625 88.230 148.615 88.460 ;
        RECT 147.625 87.560 147.795 88.230 ;
        RECT 147.625 87.350 148.615 87.560 ;
        RECT 147.625 87.085 147.795 87.350 ;
        RECT 147.625 86.855 148.615 87.085 ;
        RECT 147.625 86.185 147.795 86.855 ;
        RECT 147.625 85.975 148.615 86.185 ;
        RECT 147.625 85.715 147.795 85.975 ;
        RECT 147.625 85.485 148.615 85.715 ;
        RECT 147.625 84.815 147.795 85.485 ;
        RECT 147.625 84.605 148.615 84.815 ;
        RECT 147.625 84.340 147.795 84.605 ;
        RECT 147.625 84.110 148.615 84.340 ;
        RECT 147.625 83.440 147.795 84.110 ;
        RECT 147.625 83.230 148.615 83.440 ;
        RECT 147.625 82.960 147.795 83.230 ;
        RECT 147.625 82.730 148.615 82.960 ;
        RECT 147.625 82.060 147.795 82.730 ;
        RECT 147.625 81.850 148.615 82.060 ;
        RECT 9.825 81.665 50.125 81.835 ;
        RECT 10.830 80.895 14.340 81.665 ;
        RECT 14.545 81.205 14.810 81.665 ;
        RECT 15.480 81.205 15.650 81.665 ;
        RECT 16.320 81.200 16.570 81.665 ;
        RECT 16.810 81.205 17.075 81.665 ;
        RECT 17.745 81.205 17.915 81.665 ;
        RECT 18.585 81.200 18.835 81.665 ;
        RECT 19.065 80.915 20.275 81.665 ;
        RECT 10.830 80.375 12.480 80.895 ;
        RECT 19.065 80.375 19.585 80.915 ;
        RECT 20.445 80.895 23.955 81.665 ;
        RECT 24.160 81.205 24.425 81.665 ;
        RECT 25.095 81.205 25.265 81.665 ;
        RECT 25.935 81.200 26.185 81.665 ;
        RECT 26.425 81.205 26.690 81.665 ;
        RECT 27.360 81.205 27.530 81.665 ;
        RECT 28.200 81.200 28.450 81.665 ;
        RECT 28.680 80.915 29.890 81.665 ;
        RECT 20.445 80.375 22.095 80.895 ;
        RECT 28.680 80.375 29.200 80.915 ;
        RECT 30.060 80.895 33.570 81.665 ;
        RECT 33.775 81.205 34.040 81.665 ;
        RECT 34.710 81.205 34.880 81.665 ;
        RECT 35.550 81.200 35.800 81.665 ;
        RECT 36.040 81.205 36.305 81.665 ;
        RECT 36.975 81.205 37.145 81.665 ;
        RECT 37.815 81.200 38.065 81.665 ;
        RECT 38.295 80.915 39.505 81.665 ;
        RECT 30.060 80.375 31.710 80.895 ;
        RECT 38.295 80.375 38.815 80.915 ;
        RECT 39.675 80.895 43.185 81.665 ;
        RECT 43.390 81.205 43.655 81.665 ;
        RECT 44.325 81.205 44.495 81.665 ;
        RECT 45.165 81.200 45.415 81.665 ;
        RECT 45.655 81.205 45.920 81.665 ;
        RECT 46.590 81.205 46.760 81.665 ;
        RECT 47.430 81.200 47.680 81.665 ;
        RECT 47.910 80.915 49.120 81.665 ;
        RECT 147.625 81.585 147.795 81.850 ;
        RECT 147.625 81.355 148.615 81.585 ;
        RECT 39.675 80.375 41.325 80.895 ;
        RECT 47.910 80.375 48.430 80.915 ;
        RECT 147.625 80.685 147.795 81.355 ;
        RECT 147.625 80.475 148.615 80.685 ;
        RECT 147.625 80.210 147.795 80.475 ;
        RECT 147.625 79.980 148.615 80.210 ;
        RECT 147.625 79.310 147.795 79.980 ;
        RECT 147.625 79.100 148.615 79.310 ;
        RECT 147.625 78.840 147.795 79.100 ;
        RECT 147.625 78.610 148.615 78.840 ;
        RECT 12.640 78.000 17.800 78.170 ;
        RECT 22.255 78.000 27.415 78.170 ;
        RECT 31.870 78.000 37.030 78.170 ;
        RECT 41.485 78.000 46.645 78.170 ;
        RECT 147.625 77.940 147.795 78.610 ;
        RECT 147.625 77.730 148.615 77.940 ;
        RECT 11.615 76.285 11.785 77.625 ;
        RECT 18.655 76.995 18.825 77.625 ;
        RECT 18.655 76.590 18.830 76.995 ;
        RECT 18.640 76.390 18.840 76.590 ;
        RECT 18.655 76.285 18.825 76.390 ;
        RECT 21.230 76.285 21.400 77.625 ;
        RECT 28.270 76.995 28.440 77.625 ;
        RECT 28.270 76.590 28.445 76.995 ;
        RECT 28.255 76.390 28.455 76.590 ;
        RECT 28.270 76.285 28.440 76.390 ;
        RECT 30.845 76.285 31.015 77.625 ;
        RECT 37.885 76.995 38.055 77.625 ;
        RECT 37.885 76.590 38.060 76.995 ;
        RECT 37.870 76.390 38.070 76.590 ;
        RECT 37.885 76.285 38.055 76.390 ;
        RECT 40.460 76.285 40.630 77.625 ;
        RECT 47.500 76.995 47.670 77.625 ;
        RECT 147.625 77.465 147.795 77.730 ;
        RECT 147.625 77.235 148.615 77.465 ;
        RECT 47.500 76.590 47.675 76.995 ;
        RECT 47.485 76.390 47.685 76.590 ;
        RECT 147.625 76.565 147.795 77.235 ;
        RECT 47.500 76.285 47.670 76.390 ;
        RECT 147.625 76.355 148.615 76.565 ;
        RECT 147.625 75.305 147.795 76.355 ;
        RECT 151.180 67.620 151.350 68.885 ;
        RECT 152.360 68.255 152.530 68.885 ;
        RECT 153.540 68.290 153.710 68.885 ;
        RECT 152.360 68.025 152.535 68.255 ;
        RECT 152.365 67.620 152.535 68.025 ;
        RECT 151.180 67.605 152.535 67.620 ;
        RECT 153.530 68.025 153.710 68.290 ;
        RECT 154.720 68.280 154.890 68.885 ;
        RECT 154.720 68.025 154.905 68.280 ;
        RECT 159.170 68.190 159.340 68.885 ;
        RECT 160.350 68.205 160.520 68.885 ;
        RECT 153.530 67.605 153.700 68.025 ;
        RECT 154.735 67.605 154.905 68.025 ;
        RECT 147.125 67.565 147.340 67.580 ;
        RECT 151.180 67.565 154.905 67.605 ;
        RECT 159.165 67.565 159.340 68.190 ;
        RECT 160.345 67.565 160.520 68.205 ;
        RECT 164.075 68.225 164.245 68.885 ;
        RECT 166.035 68.465 166.205 69.130 ;
        RECT 168.830 68.635 169.000 69.195 ;
        RECT 168.825 68.530 169.000 68.635 ;
        RECT 166.035 68.295 167.525 68.465 ;
        RECT 168.825 68.360 170.320 68.530 ;
        RECT 164.075 67.565 164.250 68.225 ;
        RECT 166.035 67.565 166.205 68.295 ;
        RECT 147.015 67.550 166.205 67.565 ;
        RECT 168.825 68.285 169.000 68.360 ;
        RECT 168.825 67.550 168.995 68.285 ;
        RECT 147.015 67.395 168.995 67.550 ;
        RECT 147.125 58.200 147.340 67.395 ;
        RECT 166.035 67.380 168.995 67.395 ;
        RECT 171.765 66.170 174.775 66.340 ;
        RECT 153.705 60.965 153.875 61.615 ;
        RECT 153.130 60.755 153.875 60.965 ;
        RECT 153.130 60.750 153.845 60.755 ;
        RECT 153.130 58.870 153.345 60.750 ;
        RECT 153.705 58.870 153.875 59.485 ;
        RECT 153.130 58.655 153.875 58.870 ;
        RECT 153.130 58.200 153.345 58.655 ;
        RECT 153.705 58.625 153.875 58.655 ;
        RECT 158.220 58.200 159.130 58.205 ;
        RECT 147.125 58.035 159.130 58.200 ;
        RECT 147.125 57.985 158.520 58.035 ;
        RECT 147.125 52.585 147.340 57.985 ;
        RECT 171.765 55.340 171.935 66.170 ;
        RECT 172.895 65.335 173.935 65.505 ;
        RECT 172.895 63.765 173.935 63.935 ;
        RECT 172.895 62.195 173.935 62.365 ;
        RECT 172.895 59.145 173.935 59.315 ;
        RECT 172.895 57.575 173.935 57.745 ;
        RECT 172.895 56.005 173.935 56.175 ;
        RECT 174.605 55.340 174.775 66.170 ;
        RECT 171.765 55.170 174.775 55.340 ;
        RECT 166.150 52.585 169.110 52.600 ;
        RECT 147.020 52.540 169.110 52.585 ;
        RECT 172.010 52.540 172.180 55.170 ;
        RECT 147.020 52.430 172.180 52.540 ;
        RECT 147.020 52.415 166.320 52.430 ;
        RECT 147.020 52.390 147.340 52.415 ;
        RECT 147.020 44.395 147.190 52.390 ;
        RECT 151.295 52.375 155.020 52.415 ;
        RECT 151.295 52.360 152.650 52.375 ;
        RECT 151.295 51.095 151.465 52.360 ;
        RECT 152.480 51.955 152.650 52.360 ;
        RECT 152.475 51.725 152.650 51.955 ;
        RECT 153.645 51.955 153.815 52.375 ;
        RECT 154.850 51.955 155.020 52.375 ;
        RECT 152.475 51.095 152.645 51.725 ;
        RECT 153.645 51.690 153.825 51.955 ;
        RECT 153.655 51.095 153.825 51.690 ;
        RECT 154.835 51.700 155.020 51.955 ;
        RECT 159.280 51.790 159.455 52.415 ;
        RECT 154.835 51.095 155.005 51.700 ;
        RECT 159.285 51.095 159.455 51.790 ;
        RECT 160.460 51.775 160.635 52.415 ;
        RECT 160.465 51.095 160.635 51.775 ;
        RECT 164.190 51.755 164.365 52.415 ;
        RECT 164.190 51.095 164.360 51.755 ;
        RECT 166.150 51.685 166.320 52.415 ;
        RECT 168.790 52.370 172.180 52.430 ;
        RECT 168.940 51.695 169.110 52.370 ;
        RECT 166.150 51.515 167.640 51.685 ;
        RECT 168.940 51.620 169.115 51.695 ;
        RECT 166.150 50.850 166.320 51.515 ;
        RECT 168.940 51.450 170.435 51.620 ;
        RECT 168.940 51.345 169.115 51.450 ;
        RECT 168.945 50.785 169.115 51.345 ;
        RECT 147.625 44.395 147.795 44.545 ;
        RECT 147.020 44.225 147.795 44.395 ;
        RECT 11.615 42.225 11.785 43.565 ;
        RECT 18.655 43.460 18.825 43.565 ;
        RECT 18.640 43.260 18.840 43.460 ;
        RECT 18.655 42.855 18.830 43.260 ;
        RECT 18.655 42.225 18.825 42.855 ;
        RECT 21.230 42.225 21.400 43.565 ;
        RECT 28.270 43.460 28.440 43.565 ;
        RECT 28.255 43.260 28.455 43.460 ;
        RECT 28.270 42.855 28.445 43.260 ;
        RECT 28.270 42.225 28.440 42.855 ;
        RECT 30.845 42.225 31.015 43.565 ;
        RECT 37.885 43.460 38.055 43.565 ;
        RECT 37.870 43.260 38.070 43.460 ;
        RECT 37.885 42.855 38.060 43.260 ;
        RECT 37.885 42.225 38.055 42.855 ;
        RECT 40.460 42.225 40.630 43.565 ;
        RECT 47.500 43.460 47.670 43.565 ;
        RECT 147.625 43.495 147.795 44.225 ;
        RECT 47.485 43.260 47.685 43.460 ;
        RECT 147.625 43.285 148.615 43.495 ;
        RECT 47.500 42.855 47.675 43.260 ;
        RECT 47.500 42.225 47.670 42.855 ;
        RECT 147.625 42.615 147.795 43.285 ;
        RECT 147.625 42.385 148.615 42.615 ;
        RECT 147.625 42.120 147.795 42.385 ;
        RECT 147.625 41.910 148.615 42.120 ;
        RECT 12.640 41.680 17.800 41.850 ;
        RECT 22.255 41.680 27.415 41.850 ;
        RECT 31.870 41.680 37.030 41.850 ;
        RECT 41.485 41.680 46.645 41.850 ;
        RECT 147.625 41.240 147.795 41.910 ;
        RECT 147.625 41.010 148.615 41.240 ;
        RECT 147.625 40.750 147.795 41.010 ;
        RECT 147.625 40.540 148.615 40.750 ;
        RECT 147.625 39.870 147.795 40.540 ;
        RECT 147.625 39.640 148.615 39.870 ;
        RECT 10.830 38.955 12.480 39.475 ;
        RECT 10.830 38.185 14.340 38.955 ;
        RECT 19.065 38.935 19.585 39.475 ;
        RECT 20.445 38.955 22.095 39.475 ;
        RECT 14.545 38.185 14.810 38.645 ;
        RECT 15.480 38.185 15.650 38.645 ;
        RECT 16.320 38.185 16.570 38.650 ;
        RECT 16.810 38.185 17.075 38.645 ;
        RECT 17.745 38.185 17.915 38.645 ;
        RECT 18.585 38.185 18.835 38.650 ;
        RECT 19.065 38.185 20.275 38.935 ;
        RECT 20.445 38.185 23.955 38.955 ;
        RECT 28.680 38.935 29.200 39.475 ;
        RECT 30.060 38.955 31.710 39.475 ;
        RECT 24.160 38.185 24.425 38.645 ;
        RECT 25.095 38.185 25.265 38.645 ;
        RECT 25.935 38.185 26.185 38.650 ;
        RECT 26.425 38.185 26.690 38.645 ;
        RECT 27.360 38.185 27.530 38.645 ;
        RECT 28.200 38.185 28.450 38.650 ;
        RECT 28.680 38.185 29.890 38.935 ;
        RECT 30.060 38.185 33.570 38.955 ;
        RECT 38.295 38.935 38.815 39.475 ;
        RECT 39.675 38.955 41.325 39.475 ;
        RECT 33.775 38.185 34.040 38.645 ;
        RECT 34.710 38.185 34.880 38.645 ;
        RECT 35.550 38.185 35.800 38.650 ;
        RECT 36.040 38.185 36.305 38.645 ;
        RECT 36.975 38.185 37.145 38.645 ;
        RECT 37.815 38.185 38.065 38.650 ;
        RECT 38.295 38.185 39.505 38.935 ;
        RECT 39.675 38.185 43.185 38.955 ;
        RECT 47.910 38.935 48.430 39.475 ;
        RECT 147.625 39.375 147.795 39.640 ;
        RECT 147.625 39.165 148.615 39.375 ;
        RECT 43.390 38.185 43.655 38.645 ;
        RECT 44.325 38.185 44.495 38.645 ;
        RECT 45.165 38.185 45.415 38.650 ;
        RECT 45.655 38.185 45.920 38.645 ;
        RECT 46.590 38.185 46.760 38.645 ;
        RECT 47.430 38.185 47.680 38.650 ;
        RECT 47.910 38.185 49.120 38.935 ;
        RECT 147.625 38.495 147.795 39.165 ;
        RECT 147.625 38.265 148.615 38.495 ;
        RECT 9.825 38.015 50.125 38.185 ;
        RECT 147.625 38.000 147.795 38.265 ;
        RECT 147.625 37.790 148.615 38.000 ;
        RECT 147.625 37.120 147.795 37.790 ;
        RECT 147.625 36.890 148.615 37.120 ;
        RECT 147.625 36.620 147.795 36.890 ;
        RECT 147.625 36.410 148.615 36.620 ;
        RECT 147.625 35.740 147.795 36.410 ;
        RECT 147.625 35.510 148.615 35.740 ;
        RECT 147.625 35.245 147.795 35.510 ;
        RECT 147.625 35.035 148.615 35.245 ;
        RECT 147.625 34.365 147.795 35.035 ;
        RECT 147.625 34.135 148.615 34.365 ;
        RECT 147.625 33.875 147.795 34.135 ;
        RECT 147.625 33.665 148.615 33.875 ;
        RECT 147.625 32.995 147.795 33.665 ;
        RECT 147.625 32.765 148.615 32.995 ;
        RECT 147.625 32.500 147.795 32.765 ;
        RECT 147.625 32.290 148.615 32.500 ;
        RECT 147.625 31.620 147.795 32.290 ;
        RECT 147.625 31.390 148.615 31.620 ;
        RECT 147.625 30.360 147.795 31.390 ;
        RECT 148.785 31.370 149.035 31.700 ;
      LAYER mcon ;
        RECT 147.625 89.175 147.795 89.345 ;
        RECT 147.625 88.715 147.795 88.885 ;
        RECT 147.625 88.270 147.795 88.440 ;
        RECT 147.625 87.810 147.795 87.980 ;
        RECT 147.625 86.895 147.795 87.065 ;
        RECT 147.625 86.435 147.795 86.605 ;
        RECT 147.625 85.525 147.795 85.695 ;
        RECT 147.625 85.065 147.795 85.235 ;
        RECT 147.625 84.150 147.795 84.320 ;
        RECT 147.625 83.690 147.795 83.860 ;
        RECT 147.625 82.770 147.795 82.940 ;
        RECT 147.625 82.310 147.795 82.480 ;
        RECT 9.970 81.665 10.140 81.835 ;
        RECT 10.430 81.665 10.600 81.835 ;
        RECT 10.890 81.665 11.060 81.835 ;
        RECT 11.350 81.665 11.520 81.835 ;
        RECT 11.810 81.665 11.980 81.835 ;
        RECT 12.270 81.665 12.440 81.835 ;
        RECT 12.730 81.665 12.900 81.835 ;
        RECT 13.190 81.665 13.360 81.835 ;
        RECT 13.650 81.665 13.820 81.835 ;
        RECT 14.110 81.665 14.280 81.835 ;
        RECT 14.560 81.665 14.730 81.835 ;
        RECT 15.020 81.665 15.190 81.835 ;
        RECT 15.480 81.665 15.650 81.835 ;
        RECT 15.940 81.665 16.110 81.835 ;
        RECT 16.400 81.665 16.570 81.835 ;
        RECT 16.825 81.665 16.995 81.835 ;
        RECT 17.285 81.665 17.455 81.835 ;
        RECT 17.745 81.665 17.915 81.835 ;
        RECT 18.205 81.665 18.375 81.835 ;
        RECT 18.665 81.665 18.835 81.835 ;
        RECT 19.125 81.665 19.295 81.835 ;
        RECT 19.585 81.665 19.755 81.835 ;
        RECT 20.045 81.665 20.215 81.835 ;
        RECT 20.505 81.665 20.675 81.835 ;
        RECT 20.965 81.665 21.135 81.835 ;
        RECT 21.425 81.665 21.595 81.835 ;
        RECT 21.885 81.665 22.055 81.835 ;
        RECT 22.345 81.665 22.515 81.835 ;
        RECT 22.805 81.665 22.975 81.835 ;
        RECT 23.265 81.665 23.435 81.835 ;
        RECT 23.725 81.665 23.895 81.835 ;
        RECT 24.175 81.665 24.345 81.835 ;
        RECT 24.635 81.665 24.805 81.835 ;
        RECT 25.095 81.665 25.265 81.835 ;
        RECT 25.555 81.665 25.725 81.835 ;
        RECT 26.015 81.665 26.185 81.835 ;
        RECT 26.440 81.665 26.610 81.835 ;
        RECT 26.900 81.665 27.070 81.835 ;
        RECT 27.360 81.665 27.530 81.835 ;
        RECT 27.820 81.665 27.990 81.835 ;
        RECT 28.280 81.665 28.450 81.835 ;
        RECT 28.740 81.665 28.910 81.835 ;
        RECT 29.200 81.665 29.370 81.835 ;
        RECT 29.660 81.665 29.830 81.835 ;
        RECT 30.120 81.665 30.290 81.835 ;
        RECT 30.580 81.665 30.750 81.835 ;
        RECT 31.040 81.665 31.210 81.835 ;
        RECT 31.500 81.665 31.670 81.835 ;
        RECT 31.960 81.665 32.130 81.835 ;
        RECT 32.420 81.665 32.590 81.835 ;
        RECT 32.880 81.665 33.050 81.835 ;
        RECT 33.340 81.665 33.510 81.835 ;
        RECT 33.790 81.665 33.960 81.835 ;
        RECT 34.250 81.665 34.420 81.835 ;
        RECT 34.710 81.665 34.880 81.835 ;
        RECT 35.170 81.665 35.340 81.835 ;
        RECT 35.630 81.665 35.800 81.835 ;
        RECT 36.055 81.665 36.225 81.835 ;
        RECT 36.515 81.665 36.685 81.835 ;
        RECT 36.975 81.665 37.145 81.835 ;
        RECT 37.435 81.665 37.605 81.835 ;
        RECT 37.895 81.665 38.065 81.835 ;
        RECT 38.355 81.665 38.525 81.835 ;
        RECT 38.815 81.665 38.985 81.835 ;
        RECT 39.275 81.665 39.445 81.835 ;
        RECT 39.735 81.665 39.905 81.835 ;
        RECT 40.195 81.665 40.365 81.835 ;
        RECT 40.655 81.665 40.825 81.835 ;
        RECT 41.115 81.665 41.285 81.835 ;
        RECT 41.575 81.665 41.745 81.835 ;
        RECT 42.035 81.665 42.205 81.835 ;
        RECT 42.495 81.665 42.665 81.835 ;
        RECT 42.955 81.665 43.125 81.835 ;
        RECT 43.405 81.665 43.575 81.835 ;
        RECT 43.865 81.665 44.035 81.835 ;
        RECT 44.325 81.665 44.495 81.835 ;
        RECT 44.785 81.665 44.955 81.835 ;
        RECT 45.245 81.665 45.415 81.835 ;
        RECT 45.670 81.665 45.840 81.835 ;
        RECT 46.130 81.665 46.300 81.835 ;
        RECT 46.590 81.665 46.760 81.835 ;
        RECT 47.050 81.665 47.220 81.835 ;
        RECT 47.510 81.665 47.680 81.835 ;
        RECT 47.970 81.665 48.140 81.835 ;
        RECT 48.430 81.665 48.600 81.835 ;
        RECT 48.890 81.665 49.060 81.835 ;
        RECT 49.350 81.665 49.520 81.835 ;
        RECT 49.810 81.665 49.980 81.835 ;
        RECT 147.625 81.395 147.795 81.565 ;
        RECT 147.625 80.935 147.795 81.105 ;
        RECT 147.625 80.020 147.795 80.190 ;
        RECT 147.625 79.560 147.795 79.730 ;
        RECT 147.625 78.650 147.795 78.820 ;
        RECT 147.625 78.190 147.795 78.360 ;
        RECT 18.640 76.390 18.840 76.590 ;
        RECT 28.255 76.390 28.455 76.590 ;
        RECT 37.870 76.390 38.070 76.590 ;
        RECT 147.625 77.275 147.795 77.445 ;
        RECT 147.625 76.815 147.795 76.985 ;
        RECT 47.485 76.390 47.685 76.590 ;
        RECT 147.625 75.910 147.795 76.080 ;
        RECT 147.625 75.450 147.795 75.620 ;
        RECT 151.180 68.190 151.350 68.720 ;
        RECT 152.360 68.190 152.530 68.720 ;
        RECT 153.540 68.190 153.710 68.720 ;
        RECT 154.720 68.190 154.890 68.720 ;
        RECT 160.350 68.190 160.520 68.720 ;
        RECT 164.075 68.190 164.245 68.720 ;
        RECT 166.830 68.295 167.360 68.465 ;
        RECT 169.625 68.360 170.155 68.530 ;
        RECT 173.150 65.335 173.320 65.505 ;
        RECT 173.510 65.335 173.680 65.505 ;
        RECT 171.765 64.080 171.935 64.250 ;
        RECT 171.765 63.720 171.935 63.890 ;
        RECT 173.150 63.765 173.320 63.935 ;
        RECT 173.510 63.765 173.680 63.935 ;
        RECT 171.765 63.080 171.935 63.250 ;
        RECT 171.765 62.720 171.935 62.890 ;
        RECT 171.765 62.080 171.935 62.250 ;
        RECT 173.150 62.195 173.320 62.365 ;
        RECT 173.510 62.195 173.680 62.365 ;
        RECT 171.765 61.720 171.935 61.890 ;
        RECT 153.705 60.920 153.875 61.450 ;
        RECT 171.765 61.080 171.935 61.250 ;
        RECT 171.765 60.720 171.935 60.890 ;
        RECT 171.765 60.080 171.935 60.250 ;
        RECT 171.765 59.720 171.935 59.890 ;
        RECT 153.705 58.790 153.875 59.320 ;
        RECT 171.765 59.080 171.935 59.250 ;
        RECT 173.150 59.145 173.320 59.315 ;
        RECT 173.510 59.145 173.680 59.315 ;
        RECT 171.765 58.720 171.935 58.890 ;
        RECT 171.765 58.080 171.935 58.250 ;
        RECT 171.765 57.720 171.935 57.890 ;
        RECT 173.150 57.575 173.320 57.745 ;
        RECT 173.510 57.575 173.680 57.745 ;
        RECT 173.150 56.005 173.320 56.175 ;
        RECT 173.510 56.005 173.680 56.175 ;
        RECT 151.295 51.260 151.465 51.790 ;
        RECT 152.475 51.260 152.645 51.790 ;
        RECT 153.655 51.260 153.825 51.790 ;
        RECT 154.835 51.260 155.005 51.790 ;
        RECT 159.285 51.260 159.455 51.790 ;
        RECT 160.465 51.260 160.635 51.790 ;
        RECT 164.190 51.260 164.360 51.790 ;
        RECT 166.945 51.515 167.475 51.685 ;
        RECT 169.740 51.450 170.270 51.620 ;
        RECT 147.625 44.230 147.795 44.400 ;
        RECT 147.625 43.770 147.795 43.940 ;
        RECT 18.640 43.260 18.840 43.460 ;
        RECT 28.255 43.260 28.455 43.460 ;
        RECT 37.870 43.260 38.070 43.460 ;
        RECT 47.485 43.260 47.685 43.460 ;
        RECT 147.625 43.325 147.795 43.495 ;
        RECT 147.625 42.865 147.795 43.035 ;
        RECT 147.625 42.405 147.795 42.575 ;
        RECT 147.625 41.950 147.795 42.120 ;
        RECT 147.625 41.490 147.795 41.660 ;
        RECT 147.625 41.030 147.795 41.200 ;
        RECT 147.625 40.580 147.795 40.750 ;
        RECT 147.625 40.120 147.795 40.290 ;
        RECT 147.625 39.660 147.795 39.830 ;
        RECT 147.625 39.205 147.795 39.375 ;
        RECT 147.625 38.745 147.795 38.915 ;
        RECT 147.625 38.285 147.795 38.455 ;
        RECT 9.970 38.015 10.140 38.185 ;
        RECT 10.430 38.015 10.600 38.185 ;
        RECT 10.890 38.015 11.060 38.185 ;
        RECT 11.350 38.015 11.520 38.185 ;
        RECT 11.810 38.015 11.980 38.185 ;
        RECT 12.270 38.015 12.440 38.185 ;
        RECT 12.730 38.015 12.900 38.185 ;
        RECT 13.190 38.015 13.360 38.185 ;
        RECT 13.650 38.015 13.820 38.185 ;
        RECT 14.110 38.015 14.280 38.185 ;
        RECT 14.560 38.015 14.730 38.185 ;
        RECT 15.020 38.015 15.190 38.185 ;
        RECT 15.480 38.015 15.650 38.185 ;
        RECT 15.940 38.015 16.110 38.185 ;
        RECT 16.400 38.015 16.570 38.185 ;
        RECT 16.825 38.015 16.995 38.185 ;
        RECT 17.285 38.015 17.455 38.185 ;
        RECT 17.745 38.015 17.915 38.185 ;
        RECT 18.205 38.015 18.375 38.185 ;
        RECT 18.665 38.015 18.835 38.185 ;
        RECT 19.125 38.015 19.295 38.185 ;
        RECT 19.585 38.015 19.755 38.185 ;
        RECT 20.045 38.015 20.215 38.185 ;
        RECT 20.505 38.015 20.675 38.185 ;
        RECT 20.965 38.015 21.135 38.185 ;
        RECT 21.425 38.015 21.595 38.185 ;
        RECT 21.885 38.015 22.055 38.185 ;
        RECT 22.345 38.015 22.515 38.185 ;
        RECT 22.805 38.015 22.975 38.185 ;
        RECT 23.265 38.015 23.435 38.185 ;
        RECT 23.725 38.015 23.895 38.185 ;
        RECT 24.175 38.015 24.345 38.185 ;
        RECT 24.635 38.015 24.805 38.185 ;
        RECT 25.095 38.015 25.265 38.185 ;
        RECT 25.555 38.015 25.725 38.185 ;
        RECT 26.015 38.015 26.185 38.185 ;
        RECT 26.440 38.015 26.610 38.185 ;
        RECT 26.900 38.015 27.070 38.185 ;
        RECT 27.360 38.015 27.530 38.185 ;
        RECT 27.820 38.015 27.990 38.185 ;
        RECT 28.280 38.015 28.450 38.185 ;
        RECT 28.740 38.015 28.910 38.185 ;
        RECT 29.200 38.015 29.370 38.185 ;
        RECT 29.660 38.015 29.830 38.185 ;
        RECT 30.120 38.015 30.290 38.185 ;
        RECT 30.580 38.015 30.750 38.185 ;
        RECT 31.040 38.015 31.210 38.185 ;
        RECT 31.500 38.015 31.670 38.185 ;
        RECT 31.960 38.015 32.130 38.185 ;
        RECT 32.420 38.015 32.590 38.185 ;
        RECT 32.880 38.015 33.050 38.185 ;
        RECT 33.340 38.015 33.510 38.185 ;
        RECT 33.790 38.015 33.960 38.185 ;
        RECT 34.250 38.015 34.420 38.185 ;
        RECT 34.710 38.015 34.880 38.185 ;
        RECT 35.170 38.015 35.340 38.185 ;
        RECT 35.630 38.015 35.800 38.185 ;
        RECT 36.055 38.015 36.225 38.185 ;
        RECT 36.515 38.015 36.685 38.185 ;
        RECT 36.975 38.015 37.145 38.185 ;
        RECT 37.435 38.015 37.605 38.185 ;
        RECT 37.895 38.015 38.065 38.185 ;
        RECT 38.355 38.015 38.525 38.185 ;
        RECT 38.815 38.015 38.985 38.185 ;
        RECT 39.275 38.015 39.445 38.185 ;
        RECT 39.735 38.015 39.905 38.185 ;
        RECT 40.195 38.015 40.365 38.185 ;
        RECT 40.655 38.015 40.825 38.185 ;
        RECT 41.115 38.015 41.285 38.185 ;
        RECT 41.575 38.015 41.745 38.185 ;
        RECT 42.035 38.015 42.205 38.185 ;
        RECT 42.495 38.015 42.665 38.185 ;
        RECT 42.955 38.015 43.125 38.185 ;
        RECT 43.405 38.015 43.575 38.185 ;
        RECT 43.865 38.015 44.035 38.185 ;
        RECT 44.325 38.015 44.495 38.185 ;
        RECT 44.785 38.015 44.955 38.185 ;
        RECT 45.245 38.015 45.415 38.185 ;
        RECT 45.670 38.015 45.840 38.185 ;
        RECT 46.130 38.015 46.300 38.185 ;
        RECT 46.590 38.015 46.760 38.185 ;
        RECT 47.050 38.015 47.220 38.185 ;
        RECT 47.510 38.015 47.680 38.185 ;
        RECT 47.970 38.015 48.140 38.185 ;
        RECT 48.430 38.015 48.600 38.185 ;
        RECT 48.890 38.015 49.060 38.185 ;
        RECT 49.350 38.015 49.520 38.185 ;
        RECT 49.810 38.015 49.980 38.185 ;
        RECT 147.625 37.830 147.795 38.000 ;
        RECT 147.625 37.370 147.795 37.540 ;
        RECT 147.625 36.910 147.795 37.080 ;
        RECT 147.625 36.450 147.795 36.620 ;
        RECT 147.625 35.990 147.795 36.160 ;
        RECT 147.625 35.530 147.795 35.700 ;
        RECT 147.625 35.075 147.795 35.245 ;
        RECT 147.625 34.615 147.795 34.785 ;
        RECT 147.625 34.155 147.795 34.325 ;
        RECT 147.625 33.705 147.795 33.875 ;
        RECT 147.625 33.245 147.795 33.415 ;
        RECT 147.625 32.785 147.795 32.955 ;
        RECT 147.625 32.330 147.795 32.500 ;
        RECT 147.625 31.870 147.795 32.040 ;
        RECT 147.625 31.410 147.795 31.580 ;
        RECT 148.810 31.390 149.010 31.590 ;
        RECT 147.625 30.965 147.795 31.135 ;
        RECT 147.625 30.505 147.795 30.675 ;
      LAYER met1 ;
        RECT 6.435 107.250 6.575 118.140 ;
        RECT 6.995 107.250 7.135 118.140 ;
        RECT 7.555 107.250 7.695 118.140 ;
        RECT 8.115 107.250 8.255 118.140 ;
        RECT 8.675 107.250 8.815 118.140 ;
        RECT 9.235 107.250 9.375 118.140 ;
        RECT 9.795 107.250 9.935 118.140 ;
        RECT 10.355 107.250 10.495 118.140 ;
        RECT 10.915 107.250 11.055 118.140 ;
        RECT 11.475 107.250 11.615 118.140 ;
        RECT 12.035 107.250 12.175 118.140 ;
        RECT 12.595 107.250 12.735 118.140 ;
        RECT 13.155 107.250 13.295 118.140 ;
        RECT 13.715 107.250 13.855 118.140 ;
        RECT 14.275 107.250 14.415 118.140 ;
        RECT 14.835 107.250 14.975 118.140 ;
        RECT 15.395 107.250 15.535 118.140 ;
        RECT 15.955 107.250 16.095 118.140 ;
        RECT 16.515 107.250 16.655 118.140 ;
        RECT 17.075 107.250 17.215 118.140 ;
        RECT 19.525 107.250 19.665 118.140 ;
        RECT 20.085 107.250 20.225 118.140 ;
        RECT 20.645 107.250 20.785 118.140 ;
        RECT 21.205 107.250 21.345 118.140 ;
        RECT 21.765 107.250 21.905 118.140 ;
        RECT 22.325 107.250 22.465 118.140 ;
        RECT 22.885 107.250 23.025 118.140 ;
        RECT 23.445 107.250 23.585 118.140 ;
        RECT 24.005 107.250 24.145 118.140 ;
        RECT 24.565 107.250 24.705 118.140 ;
        RECT 25.125 107.250 25.265 118.140 ;
        RECT 25.685 107.250 25.825 118.140 ;
        RECT 26.245 107.250 26.385 118.140 ;
        RECT 26.805 107.250 26.945 118.140 ;
        RECT 27.365 107.250 27.505 118.140 ;
        RECT 27.925 107.250 28.065 118.140 ;
        RECT 28.485 107.250 28.625 118.140 ;
        RECT 29.045 107.250 29.185 118.140 ;
        RECT 29.605 107.250 29.745 118.140 ;
        RECT 30.165 107.250 30.305 118.140 ;
        RECT 6.155 106.920 17.565 107.250 ;
        RECT 19.245 106.920 30.655 107.250 ;
        RECT 32.615 107.230 32.755 118.120 ;
        RECT 33.175 107.230 33.315 118.120 ;
        RECT 33.735 107.230 33.875 118.120 ;
        RECT 34.295 107.230 34.435 118.120 ;
        RECT 34.855 107.230 34.995 118.120 ;
        RECT 35.415 107.230 35.555 118.120 ;
        RECT 35.975 107.230 36.115 118.120 ;
        RECT 36.535 107.230 36.675 118.120 ;
        RECT 37.095 107.230 37.235 118.120 ;
        RECT 37.655 107.230 37.795 118.120 ;
        RECT 38.215 107.230 38.355 118.120 ;
        RECT 38.775 107.230 38.915 118.120 ;
        RECT 39.335 107.230 39.475 118.120 ;
        RECT 39.895 107.230 40.035 118.120 ;
        RECT 40.455 107.230 40.595 118.120 ;
        RECT 41.015 107.230 41.155 118.120 ;
        RECT 41.575 107.230 41.715 118.120 ;
        RECT 42.135 107.230 42.275 118.120 ;
        RECT 42.695 107.230 42.835 118.120 ;
        RECT 43.255 107.230 43.395 118.120 ;
        RECT 45.705 107.230 45.845 118.120 ;
        RECT 46.265 107.230 46.405 118.120 ;
        RECT 46.825 107.230 46.965 118.120 ;
        RECT 47.385 107.230 47.525 118.120 ;
        RECT 47.945 107.230 48.085 118.120 ;
        RECT 48.505 107.230 48.645 118.120 ;
        RECT 49.065 107.230 49.205 118.120 ;
        RECT 49.625 107.230 49.765 118.120 ;
        RECT 50.185 107.230 50.325 118.120 ;
        RECT 50.745 107.230 50.885 118.120 ;
        RECT 51.305 107.230 51.445 118.120 ;
        RECT 51.865 107.230 52.005 118.120 ;
        RECT 52.425 107.230 52.565 118.120 ;
        RECT 52.985 107.230 53.125 118.120 ;
        RECT 53.545 107.230 53.685 118.120 ;
        RECT 54.105 107.230 54.245 118.120 ;
        RECT 54.665 107.230 54.805 118.120 ;
        RECT 55.225 107.230 55.365 118.120 ;
        RECT 55.785 107.230 55.925 118.120 ;
        RECT 56.345 107.230 56.485 118.120 ;
        RECT 58.755 107.230 58.895 118.120 ;
        RECT 59.315 107.230 59.455 118.120 ;
        RECT 59.875 107.230 60.015 118.120 ;
        RECT 60.435 107.230 60.575 118.120 ;
        RECT 60.995 107.230 61.135 118.120 ;
        RECT 61.555 107.230 61.695 118.120 ;
        RECT 62.115 107.230 62.255 118.120 ;
        RECT 62.675 107.230 62.815 118.120 ;
        RECT 63.235 107.230 63.375 118.120 ;
        RECT 63.795 107.230 63.935 118.120 ;
        RECT 64.355 107.230 64.495 118.120 ;
        RECT 64.915 107.230 65.055 118.120 ;
        RECT 65.475 107.230 65.615 118.120 ;
        RECT 66.035 107.230 66.175 118.120 ;
        RECT 66.595 107.230 66.735 118.120 ;
        RECT 67.155 107.230 67.295 118.120 ;
        RECT 67.715 107.230 67.855 118.120 ;
        RECT 68.275 107.230 68.415 118.120 ;
        RECT 68.835 107.230 68.975 118.120 ;
        RECT 69.395 107.230 69.535 118.120 ;
        RECT 71.845 107.230 71.985 118.120 ;
        RECT 72.405 107.230 72.545 118.120 ;
        RECT 72.965 107.230 73.105 118.120 ;
        RECT 73.525 107.230 73.665 118.120 ;
        RECT 74.085 107.230 74.225 118.120 ;
        RECT 74.645 107.230 74.785 118.120 ;
        RECT 75.205 107.230 75.345 118.120 ;
        RECT 75.765 107.230 75.905 118.120 ;
        RECT 76.325 107.230 76.465 118.120 ;
        RECT 76.885 107.230 77.025 118.120 ;
        RECT 77.445 107.230 77.585 118.120 ;
        RECT 78.005 107.230 78.145 118.120 ;
        RECT 78.565 107.230 78.705 118.120 ;
        RECT 79.125 107.230 79.265 118.120 ;
        RECT 79.685 107.230 79.825 118.120 ;
        RECT 80.245 107.230 80.385 118.120 ;
        RECT 80.805 107.230 80.945 118.120 ;
        RECT 81.365 107.230 81.505 118.120 ;
        RECT 81.925 107.230 82.065 118.120 ;
        RECT 82.485 107.230 82.625 118.120 ;
        RECT 32.335 106.900 43.745 107.230 ;
        RECT 45.425 106.900 56.835 107.230 ;
        RECT 58.475 106.900 69.885 107.230 ;
        RECT 71.565 106.900 82.975 107.230 ;
        RECT 84.935 107.210 85.075 118.100 ;
        RECT 85.495 107.210 85.635 118.100 ;
        RECT 86.055 107.210 86.195 118.100 ;
        RECT 86.615 107.210 86.755 118.100 ;
        RECT 87.175 107.210 87.315 118.100 ;
        RECT 87.735 107.210 87.875 118.100 ;
        RECT 88.295 107.210 88.435 118.100 ;
        RECT 88.855 107.210 88.995 118.100 ;
        RECT 89.415 107.210 89.555 118.100 ;
        RECT 89.975 107.210 90.115 118.100 ;
        RECT 90.535 107.210 90.675 118.100 ;
        RECT 91.095 107.210 91.235 118.100 ;
        RECT 91.655 107.210 91.795 118.100 ;
        RECT 92.215 107.210 92.355 118.100 ;
        RECT 92.775 107.210 92.915 118.100 ;
        RECT 93.335 107.210 93.475 118.100 ;
        RECT 93.895 107.210 94.035 118.100 ;
        RECT 94.455 107.210 94.595 118.100 ;
        RECT 95.015 107.210 95.155 118.100 ;
        RECT 95.575 107.210 95.715 118.100 ;
        RECT 98.025 107.210 98.165 118.100 ;
        RECT 98.585 107.210 98.725 118.100 ;
        RECT 99.145 107.210 99.285 118.100 ;
        RECT 99.705 107.210 99.845 118.100 ;
        RECT 100.265 107.210 100.405 118.100 ;
        RECT 100.825 107.210 100.965 118.100 ;
        RECT 101.385 107.210 101.525 118.100 ;
        RECT 101.945 107.210 102.085 118.100 ;
        RECT 102.505 107.210 102.645 118.100 ;
        RECT 103.065 107.210 103.205 118.100 ;
        RECT 103.625 107.210 103.765 118.100 ;
        RECT 104.185 107.210 104.325 118.100 ;
        RECT 104.745 107.210 104.885 118.100 ;
        RECT 105.305 107.210 105.445 118.100 ;
        RECT 105.865 107.210 106.005 118.100 ;
        RECT 106.425 107.210 106.565 118.100 ;
        RECT 106.985 107.210 107.125 118.100 ;
        RECT 107.545 107.210 107.685 118.100 ;
        RECT 108.105 107.210 108.245 118.100 ;
        RECT 108.665 107.210 108.805 118.100 ;
        RECT 111.115 107.210 111.255 118.100 ;
        RECT 111.675 107.210 111.815 118.100 ;
        RECT 112.235 107.210 112.375 118.100 ;
        RECT 112.795 107.210 112.935 118.100 ;
        RECT 113.355 107.210 113.495 118.100 ;
        RECT 113.915 107.210 114.055 118.100 ;
        RECT 114.475 107.210 114.615 118.100 ;
        RECT 115.035 107.210 115.175 118.100 ;
        RECT 115.595 107.210 115.735 118.100 ;
        RECT 116.155 107.210 116.295 118.100 ;
        RECT 116.715 107.210 116.855 118.100 ;
        RECT 117.275 107.210 117.415 118.100 ;
        RECT 117.835 107.210 117.975 118.100 ;
        RECT 118.395 107.210 118.535 118.100 ;
        RECT 118.955 107.210 119.095 118.100 ;
        RECT 119.515 107.210 119.655 118.100 ;
        RECT 120.075 107.210 120.215 118.100 ;
        RECT 120.635 107.210 120.775 118.100 ;
        RECT 121.195 107.210 121.335 118.100 ;
        RECT 121.755 107.210 121.895 118.100 ;
        RECT 124.205 107.210 124.345 118.100 ;
        RECT 124.765 107.210 124.905 118.100 ;
        RECT 125.325 107.210 125.465 118.100 ;
        RECT 125.885 107.210 126.025 118.100 ;
        RECT 126.445 107.210 126.585 118.100 ;
        RECT 127.005 107.210 127.145 118.100 ;
        RECT 127.565 107.210 127.705 118.100 ;
        RECT 128.125 107.210 128.265 118.100 ;
        RECT 128.685 107.210 128.825 118.100 ;
        RECT 129.245 107.210 129.385 118.100 ;
        RECT 129.805 107.210 129.945 118.100 ;
        RECT 130.365 107.210 130.505 118.100 ;
        RECT 130.925 107.210 131.065 118.100 ;
        RECT 131.485 107.210 131.625 118.100 ;
        RECT 132.045 107.210 132.185 118.100 ;
        RECT 132.605 107.210 132.745 118.100 ;
        RECT 133.165 107.210 133.305 118.100 ;
        RECT 133.725 107.210 133.865 118.100 ;
        RECT 134.285 107.210 134.425 118.100 ;
        RECT 134.845 107.210 134.985 118.100 ;
        RECT 84.655 106.880 96.065 107.210 ;
        RECT 97.745 106.880 109.155 107.210 ;
        RECT 110.835 106.880 122.245 107.210 ;
        RECT 123.925 106.880 135.335 107.210 ;
        RECT 137.295 107.190 137.435 118.080 ;
        RECT 137.855 107.190 137.995 118.080 ;
        RECT 138.415 107.190 138.555 118.080 ;
        RECT 138.975 107.190 139.115 118.080 ;
        RECT 139.535 107.190 139.675 118.080 ;
        RECT 140.095 107.190 140.235 118.080 ;
        RECT 140.655 107.190 140.795 118.080 ;
        RECT 141.215 107.190 141.355 118.080 ;
        RECT 141.775 107.190 141.915 118.080 ;
        RECT 142.335 107.190 142.475 118.080 ;
        RECT 142.895 107.190 143.035 118.080 ;
        RECT 143.455 107.190 143.595 118.080 ;
        RECT 144.015 107.190 144.155 118.080 ;
        RECT 144.575 107.190 144.715 118.080 ;
        RECT 145.135 107.190 145.275 118.080 ;
        RECT 145.695 107.190 145.835 118.080 ;
        RECT 146.255 107.190 146.395 118.080 ;
        RECT 146.815 107.190 146.955 118.080 ;
        RECT 147.375 107.190 147.515 118.080 ;
        RECT 147.935 107.190 148.075 118.080 ;
        RECT 150.385 107.190 150.525 118.080 ;
        RECT 150.945 107.190 151.085 118.080 ;
        RECT 151.505 107.190 151.645 118.080 ;
        RECT 152.065 107.190 152.205 118.080 ;
        RECT 152.625 107.190 152.765 118.080 ;
        RECT 153.185 107.190 153.325 118.080 ;
        RECT 153.745 107.190 153.885 118.080 ;
        RECT 154.305 107.190 154.445 118.080 ;
        RECT 154.865 107.190 155.005 118.080 ;
        RECT 155.425 107.190 155.565 118.080 ;
        RECT 155.985 107.190 156.125 118.080 ;
        RECT 156.545 107.190 156.685 118.080 ;
        RECT 157.105 107.190 157.245 118.080 ;
        RECT 157.665 107.190 157.805 118.080 ;
        RECT 158.225 107.190 158.365 118.080 ;
        RECT 158.785 107.190 158.925 118.080 ;
        RECT 159.345 107.190 159.485 118.080 ;
        RECT 159.905 107.190 160.045 118.080 ;
        RECT 160.465 107.190 160.605 118.080 ;
        RECT 161.025 107.190 161.165 118.080 ;
        RECT 137.015 106.860 148.425 107.190 ;
        RECT 150.105 106.860 161.515 107.190 ;
        RECT 6.185 104.870 17.595 105.200 ;
        RECT 19.275 104.870 30.685 105.200 ;
        RECT 32.365 104.890 43.775 105.220 ;
        RECT 45.455 104.890 56.865 105.220 ;
        RECT 58.505 104.890 69.915 105.220 ;
        RECT 71.595 104.890 83.005 105.220 ;
        RECT 84.685 104.910 96.095 105.240 ;
        RECT 97.775 104.910 109.185 105.240 ;
        RECT 110.865 104.910 122.275 105.240 ;
        RECT 123.955 104.910 135.365 105.240 ;
        RECT 137.045 104.930 148.455 105.260 ;
        RECT 150.135 104.930 161.545 105.260 ;
        RECT 6.465 93.980 6.605 104.870 ;
        RECT 7.025 93.980 7.165 104.870 ;
        RECT 7.585 93.980 7.725 104.870 ;
        RECT 8.145 93.980 8.285 104.870 ;
        RECT 8.705 93.980 8.845 104.870 ;
        RECT 9.265 93.980 9.405 104.870 ;
        RECT 9.825 93.980 9.965 104.870 ;
        RECT 10.385 93.980 10.525 104.870 ;
        RECT 10.945 93.980 11.085 104.870 ;
        RECT 11.505 93.980 11.645 104.870 ;
        RECT 12.065 93.980 12.205 104.870 ;
        RECT 12.625 93.980 12.765 104.870 ;
        RECT 13.185 93.980 13.325 104.870 ;
        RECT 13.745 93.980 13.885 104.870 ;
        RECT 14.305 93.980 14.445 104.870 ;
        RECT 14.865 93.980 15.005 104.870 ;
        RECT 15.425 93.980 15.565 104.870 ;
        RECT 15.985 93.980 16.125 104.870 ;
        RECT 16.545 93.980 16.685 104.870 ;
        RECT 17.105 93.980 17.245 104.870 ;
        RECT 19.555 93.980 19.695 104.870 ;
        RECT 20.115 93.980 20.255 104.870 ;
        RECT 20.675 93.980 20.815 104.870 ;
        RECT 21.235 93.980 21.375 104.870 ;
        RECT 21.795 93.980 21.935 104.870 ;
        RECT 22.355 93.980 22.495 104.870 ;
        RECT 22.915 93.980 23.055 104.870 ;
        RECT 23.475 93.980 23.615 104.870 ;
        RECT 24.035 93.980 24.175 104.870 ;
        RECT 24.595 93.980 24.735 104.870 ;
        RECT 25.155 93.980 25.295 104.870 ;
        RECT 25.715 93.980 25.855 104.870 ;
        RECT 26.275 93.980 26.415 104.870 ;
        RECT 26.835 93.980 26.975 104.870 ;
        RECT 27.395 93.980 27.535 104.870 ;
        RECT 27.955 93.980 28.095 104.870 ;
        RECT 28.515 93.980 28.655 104.870 ;
        RECT 29.075 93.980 29.215 104.870 ;
        RECT 29.635 93.980 29.775 104.870 ;
        RECT 30.195 93.980 30.335 104.870 ;
        RECT 32.645 94.000 32.785 104.890 ;
        RECT 33.205 94.000 33.345 104.890 ;
        RECT 33.765 94.000 33.905 104.890 ;
        RECT 34.325 94.000 34.465 104.890 ;
        RECT 34.885 94.000 35.025 104.890 ;
        RECT 35.445 94.000 35.585 104.890 ;
        RECT 36.005 94.000 36.145 104.890 ;
        RECT 36.565 94.000 36.705 104.890 ;
        RECT 37.125 94.000 37.265 104.890 ;
        RECT 37.685 94.000 37.825 104.890 ;
        RECT 38.245 94.000 38.385 104.890 ;
        RECT 38.805 94.000 38.945 104.890 ;
        RECT 39.365 94.000 39.505 104.890 ;
        RECT 39.925 94.000 40.065 104.890 ;
        RECT 40.485 94.000 40.625 104.890 ;
        RECT 41.045 94.000 41.185 104.890 ;
        RECT 41.605 94.000 41.745 104.890 ;
        RECT 42.165 94.000 42.305 104.890 ;
        RECT 42.725 94.000 42.865 104.890 ;
        RECT 43.285 94.000 43.425 104.890 ;
        RECT 45.735 94.000 45.875 104.890 ;
        RECT 46.295 94.000 46.435 104.890 ;
        RECT 46.855 94.000 46.995 104.890 ;
        RECT 47.415 94.000 47.555 104.890 ;
        RECT 47.975 94.000 48.115 104.890 ;
        RECT 48.535 94.000 48.675 104.890 ;
        RECT 49.095 94.000 49.235 104.890 ;
        RECT 49.655 94.000 49.795 104.890 ;
        RECT 50.215 94.000 50.355 104.890 ;
        RECT 50.775 94.000 50.915 104.890 ;
        RECT 51.335 94.000 51.475 104.890 ;
        RECT 51.895 94.000 52.035 104.890 ;
        RECT 52.455 94.000 52.595 104.890 ;
        RECT 53.015 94.000 53.155 104.890 ;
        RECT 53.575 94.000 53.715 104.890 ;
        RECT 54.135 94.000 54.275 104.890 ;
        RECT 54.695 94.000 54.835 104.890 ;
        RECT 55.255 94.000 55.395 104.890 ;
        RECT 55.815 94.000 55.955 104.890 ;
        RECT 56.375 94.000 56.515 104.890 ;
        RECT 58.785 94.000 58.925 104.890 ;
        RECT 59.345 94.000 59.485 104.890 ;
        RECT 59.905 94.000 60.045 104.890 ;
        RECT 60.465 94.000 60.605 104.890 ;
        RECT 61.025 94.000 61.165 104.890 ;
        RECT 61.585 94.000 61.725 104.890 ;
        RECT 62.145 94.000 62.285 104.890 ;
        RECT 62.705 94.000 62.845 104.890 ;
        RECT 63.265 94.000 63.405 104.890 ;
        RECT 63.825 94.000 63.965 104.890 ;
        RECT 64.385 94.000 64.525 104.890 ;
        RECT 64.945 94.000 65.085 104.890 ;
        RECT 65.505 94.000 65.645 104.890 ;
        RECT 66.065 94.000 66.205 104.890 ;
        RECT 66.625 94.000 66.765 104.890 ;
        RECT 67.185 94.000 67.325 104.890 ;
        RECT 67.745 94.000 67.885 104.890 ;
        RECT 68.305 94.000 68.445 104.890 ;
        RECT 68.865 94.000 69.005 104.890 ;
        RECT 69.425 94.000 69.565 104.890 ;
        RECT 71.875 94.000 72.015 104.890 ;
        RECT 72.435 94.000 72.575 104.890 ;
        RECT 72.995 94.000 73.135 104.890 ;
        RECT 73.555 94.000 73.695 104.890 ;
        RECT 74.115 94.000 74.255 104.890 ;
        RECT 74.675 94.000 74.815 104.890 ;
        RECT 75.235 94.000 75.375 104.890 ;
        RECT 75.795 94.000 75.935 104.890 ;
        RECT 76.355 94.000 76.495 104.890 ;
        RECT 76.915 94.000 77.055 104.890 ;
        RECT 77.475 94.000 77.615 104.890 ;
        RECT 78.035 94.000 78.175 104.890 ;
        RECT 78.595 94.000 78.735 104.890 ;
        RECT 79.155 94.000 79.295 104.890 ;
        RECT 79.715 94.000 79.855 104.890 ;
        RECT 80.275 94.000 80.415 104.890 ;
        RECT 80.835 94.000 80.975 104.890 ;
        RECT 81.395 94.000 81.535 104.890 ;
        RECT 81.955 94.000 82.095 104.890 ;
        RECT 82.515 94.000 82.655 104.890 ;
        RECT 84.965 94.020 85.105 104.910 ;
        RECT 85.525 94.020 85.665 104.910 ;
        RECT 86.085 94.020 86.225 104.910 ;
        RECT 86.645 94.020 86.785 104.910 ;
        RECT 87.205 94.020 87.345 104.910 ;
        RECT 87.765 94.020 87.905 104.910 ;
        RECT 88.325 94.020 88.465 104.910 ;
        RECT 88.885 94.020 89.025 104.910 ;
        RECT 89.445 94.020 89.585 104.910 ;
        RECT 90.005 94.020 90.145 104.910 ;
        RECT 90.565 94.020 90.705 104.910 ;
        RECT 91.125 94.020 91.265 104.910 ;
        RECT 91.685 94.020 91.825 104.910 ;
        RECT 92.245 94.020 92.385 104.910 ;
        RECT 92.805 94.020 92.945 104.910 ;
        RECT 93.365 94.020 93.505 104.910 ;
        RECT 93.925 94.020 94.065 104.910 ;
        RECT 94.485 94.020 94.625 104.910 ;
        RECT 95.045 94.020 95.185 104.910 ;
        RECT 95.605 94.020 95.745 104.910 ;
        RECT 98.055 94.020 98.195 104.910 ;
        RECT 98.615 94.020 98.755 104.910 ;
        RECT 99.175 94.020 99.315 104.910 ;
        RECT 99.735 94.020 99.875 104.910 ;
        RECT 100.295 94.020 100.435 104.910 ;
        RECT 100.855 94.020 100.995 104.910 ;
        RECT 101.415 94.020 101.555 104.910 ;
        RECT 101.975 94.020 102.115 104.910 ;
        RECT 102.535 94.020 102.675 104.910 ;
        RECT 103.095 94.020 103.235 104.910 ;
        RECT 103.655 94.020 103.795 104.910 ;
        RECT 104.215 94.020 104.355 104.910 ;
        RECT 104.775 94.020 104.915 104.910 ;
        RECT 105.335 94.020 105.475 104.910 ;
        RECT 105.895 94.020 106.035 104.910 ;
        RECT 106.455 94.020 106.595 104.910 ;
        RECT 107.015 94.020 107.155 104.910 ;
        RECT 107.575 94.020 107.715 104.910 ;
        RECT 108.135 94.020 108.275 104.910 ;
        RECT 108.695 94.020 108.835 104.910 ;
        RECT 111.145 94.020 111.285 104.910 ;
        RECT 111.705 94.020 111.845 104.910 ;
        RECT 112.265 94.020 112.405 104.910 ;
        RECT 112.825 94.020 112.965 104.910 ;
        RECT 113.385 94.020 113.525 104.910 ;
        RECT 113.945 94.020 114.085 104.910 ;
        RECT 114.505 94.020 114.645 104.910 ;
        RECT 115.065 94.020 115.205 104.910 ;
        RECT 115.625 94.020 115.765 104.910 ;
        RECT 116.185 94.020 116.325 104.910 ;
        RECT 116.745 94.020 116.885 104.910 ;
        RECT 117.305 94.020 117.445 104.910 ;
        RECT 117.865 94.020 118.005 104.910 ;
        RECT 118.425 94.020 118.565 104.910 ;
        RECT 118.985 94.020 119.125 104.910 ;
        RECT 119.545 94.020 119.685 104.910 ;
        RECT 120.105 94.020 120.245 104.910 ;
        RECT 120.665 94.020 120.805 104.910 ;
        RECT 121.225 94.020 121.365 104.910 ;
        RECT 121.785 94.020 121.925 104.910 ;
        RECT 124.235 94.020 124.375 104.910 ;
        RECT 124.795 94.020 124.935 104.910 ;
        RECT 125.355 94.020 125.495 104.910 ;
        RECT 125.915 94.020 126.055 104.910 ;
        RECT 126.475 94.020 126.615 104.910 ;
        RECT 127.035 94.020 127.175 104.910 ;
        RECT 127.595 94.020 127.735 104.910 ;
        RECT 128.155 94.020 128.295 104.910 ;
        RECT 128.715 94.020 128.855 104.910 ;
        RECT 129.275 94.020 129.415 104.910 ;
        RECT 129.835 94.020 129.975 104.910 ;
        RECT 130.395 94.020 130.535 104.910 ;
        RECT 130.955 94.020 131.095 104.910 ;
        RECT 131.515 94.020 131.655 104.910 ;
        RECT 132.075 94.020 132.215 104.910 ;
        RECT 132.635 94.020 132.775 104.910 ;
        RECT 133.195 94.020 133.335 104.910 ;
        RECT 133.755 94.020 133.895 104.910 ;
        RECT 134.315 94.020 134.455 104.910 ;
        RECT 134.875 94.020 135.015 104.910 ;
        RECT 137.325 94.040 137.465 104.930 ;
        RECT 137.885 94.040 138.025 104.930 ;
        RECT 138.445 94.040 138.585 104.930 ;
        RECT 139.005 94.040 139.145 104.930 ;
        RECT 139.565 94.040 139.705 104.930 ;
        RECT 140.125 94.040 140.265 104.930 ;
        RECT 140.685 94.040 140.825 104.930 ;
        RECT 141.245 94.040 141.385 104.930 ;
        RECT 141.805 94.040 141.945 104.930 ;
        RECT 142.365 94.040 142.505 104.930 ;
        RECT 142.925 94.040 143.065 104.930 ;
        RECT 143.485 94.040 143.625 104.930 ;
        RECT 144.045 94.040 144.185 104.930 ;
        RECT 144.605 94.040 144.745 104.930 ;
        RECT 145.165 94.040 145.305 104.930 ;
        RECT 145.725 94.040 145.865 104.930 ;
        RECT 146.285 94.040 146.425 104.930 ;
        RECT 146.845 94.040 146.985 104.930 ;
        RECT 147.405 94.040 147.545 104.930 ;
        RECT 147.965 94.040 148.105 104.930 ;
        RECT 150.415 94.040 150.555 104.930 ;
        RECT 150.975 94.040 151.115 104.930 ;
        RECT 151.535 94.040 151.675 104.930 ;
        RECT 152.095 94.040 152.235 104.930 ;
        RECT 152.655 94.040 152.795 104.930 ;
        RECT 153.215 94.040 153.355 104.930 ;
        RECT 153.775 94.040 153.915 104.930 ;
        RECT 154.335 94.040 154.475 104.930 ;
        RECT 154.895 94.040 155.035 104.930 ;
        RECT 155.455 94.040 155.595 104.930 ;
        RECT 156.015 94.040 156.155 104.930 ;
        RECT 156.575 94.040 156.715 104.930 ;
        RECT 157.135 94.040 157.275 104.930 ;
        RECT 157.695 94.040 157.835 104.930 ;
        RECT 158.255 94.040 158.395 104.930 ;
        RECT 158.815 94.040 158.955 104.930 ;
        RECT 159.375 94.040 159.515 104.930 ;
        RECT 159.935 94.040 160.075 104.930 ;
        RECT 160.495 94.040 160.635 104.930 ;
        RECT 161.055 94.040 161.195 104.930 ;
        RECT 147.460 90.270 163.380 90.745 ;
        RECT 147.460 89.490 147.935 90.270 ;
        RECT 147.460 89.180 147.950 89.490 ;
        RECT 4.760 81.970 5.230 89.175 ;
        RECT 9.825 81.970 50.125 81.990 ;
        RECT 4.760 81.510 50.125 81.970 ;
        RECT 4.760 81.500 10.575 81.510 ;
        RECT 18.610 76.330 18.870 76.650 ;
        RECT 28.225 76.330 28.485 76.650 ;
        RECT 37.840 76.330 38.100 76.650 ;
        RECT 47.455 76.330 47.715 76.650 ;
        RECT 147.470 75.305 147.950 89.180 ;
        RECT 151.150 68.130 151.380 68.780 ;
        RECT 152.330 68.130 152.560 68.780 ;
        RECT 153.510 68.130 153.740 68.780 ;
        RECT 154.690 68.130 154.920 68.780 ;
        RECT 159.140 68.130 159.370 68.780 ;
        RECT 160.320 68.130 160.550 68.780 ;
        RECT 164.045 68.130 164.275 68.780 ;
        RECT 166.770 68.265 167.420 68.495 ;
        RECT 169.565 68.330 170.215 68.560 ;
        RECT 171.700 65.535 172.000 65.770 ;
        RECT 171.700 65.305 173.915 65.535 ;
        RECT 171.700 63.965 172.000 65.305 ;
        RECT 171.700 63.735 173.915 63.965 ;
        RECT 171.700 62.395 172.000 63.735 ;
        RECT 171.700 62.165 173.915 62.395 ;
        RECT 153.675 60.860 153.905 61.510 ;
        RECT 153.675 58.730 153.905 59.380 ;
        RECT 171.700 59.345 172.000 62.165 ;
        RECT 171.700 59.115 173.915 59.345 ;
        RECT 171.700 57.775 172.000 59.115 ;
        RECT 171.700 57.545 173.915 57.775 ;
        RECT 171.700 56.205 172.000 57.545 ;
        RECT 171.700 55.975 173.915 56.205 ;
        RECT 171.700 55.740 172.000 55.975 ;
        RECT 151.265 51.200 151.495 51.850 ;
        RECT 152.445 51.200 152.675 51.850 ;
        RECT 153.625 51.200 153.855 51.850 ;
        RECT 154.805 51.200 155.035 51.850 ;
        RECT 159.255 51.200 159.485 51.850 ;
        RECT 160.435 51.200 160.665 51.850 ;
        RECT 164.160 51.200 164.390 51.850 ;
        RECT 166.885 51.485 167.535 51.715 ;
        RECT 169.680 51.420 170.330 51.650 ;
        RECT 18.610 43.200 18.870 43.520 ;
        RECT 28.225 43.200 28.485 43.520 ;
        RECT 37.840 43.200 38.100 43.520 ;
        RECT 47.455 43.200 47.715 43.520 ;
        RECT 4.750 38.340 10.575 38.350 ;
        RECT 4.750 37.880 50.125 38.340 ;
        RECT 4.750 33.185 5.220 37.880 ;
        RECT 9.825 37.860 50.125 37.880 ;
        RECT 147.470 30.670 147.950 44.545 ;
        RECT 148.780 31.330 149.040 31.650 ;
        RECT 147.460 30.360 147.950 30.670 ;
        RECT 147.460 29.690 147.935 30.360 ;
        RECT 163.275 29.690 163.750 29.720 ;
        RECT 147.460 29.215 163.750 29.690 ;
        RECT 163.275 29.185 163.750 29.215 ;
        RECT 6.875 15.610 7.015 26.500 ;
        RECT 7.435 15.610 7.575 26.500 ;
        RECT 7.995 15.610 8.135 26.500 ;
        RECT 8.555 15.610 8.695 26.500 ;
        RECT 9.115 15.610 9.255 26.500 ;
        RECT 9.675 15.610 9.815 26.500 ;
        RECT 10.235 15.610 10.375 26.500 ;
        RECT 10.795 15.610 10.935 26.500 ;
        RECT 11.355 15.610 11.495 26.500 ;
        RECT 11.915 15.610 12.055 26.500 ;
        RECT 12.475 15.610 12.615 26.500 ;
        RECT 13.035 15.610 13.175 26.500 ;
        RECT 13.595 15.610 13.735 26.500 ;
        RECT 14.155 15.610 14.295 26.500 ;
        RECT 14.715 15.610 14.855 26.500 ;
        RECT 15.275 15.610 15.415 26.500 ;
        RECT 15.835 15.610 15.975 26.500 ;
        RECT 16.395 15.610 16.535 26.500 ;
        RECT 16.955 15.610 17.095 26.500 ;
        RECT 17.515 15.610 17.655 26.500 ;
        RECT 19.965 15.610 20.105 26.500 ;
        RECT 20.525 15.610 20.665 26.500 ;
        RECT 21.085 15.610 21.225 26.500 ;
        RECT 21.645 15.610 21.785 26.500 ;
        RECT 22.205 15.610 22.345 26.500 ;
        RECT 22.765 15.610 22.905 26.500 ;
        RECT 23.325 15.610 23.465 26.500 ;
        RECT 23.885 15.610 24.025 26.500 ;
        RECT 24.445 15.610 24.585 26.500 ;
        RECT 25.005 15.610 25.145 26.500 ;
        RECT 25.565 15.610 25.705 26.500 ;
        RECT 26.125 15.610 26.265 26.500 ;
        RECT 26.685 15.610 26.825 26.500 ;
        RECT 27.245 15.610 27.385 26.500 ;
        RECT 27.805 15.610 27.945 26.500 ;
        RECT 28.365 15.610 28.505 26.500 ;
        RECT 28.925 15.610 29.065 26.500 ;
        RECT 29.485 15.610 29.625 26.500 ;
        RECT 30.045 15.610 30.185 26.500 ;
        RECT 30.605 15.610 30.745 26.500 ;
        RECT 6.595 15.280 18.005 15.610 ;
        RECT 19.685 15.280 31.095 15.610 ;
        RECT 33.055 15.590 33.195 26.480 ;
        RECT 33.615 15.590 33.755 26.480 ;
        RECT 34.175 15.590 34.315 26.480 ;
        RECT 34.735 15.590 34.875 26.480 ;
        RECT 35.295 15.590 35.435 26.480 ;
        RECT 35.855 15.590 35.995 26.480 ;
        RECT 36.415 15.590 36.555 26.480 ;
        RECT 36.975 15.590 37.115 26.480 ;
        RECT 37.535 15.590 37.675 26.480 ;
        RECT 38.095 15.590 38.235 26.480 ;
        RECT 38.655 15.590 38.795 26.480 ;
        RECT 39.215 15.590 39.355 26.480 ;
        RECT 39.775 15.590 39.915 26.480 ;
        RECT 40.335 15.590 40.475 26.480 ;
        RECT 40.895 15.590 41.035 26.480 ;
        RECT 41.455 15.590 41.595 26.480 ;
        RECT 42.015 15.590 42.155 26.480 ;
        RECT 42.575 15.590 42.715 26.480 ;
        RECT 43.135 15.590 43.275 26.480 ;
        RECT 43.695 15.590 43.835 26.480 ;
        RECT 46.145 15.590 46.285 26.480 ;
        RECT 46.705 15.590 46.845 26.480 ;
        RECT 47.265 15.590 47.405 26.480 ;
        RECT 47.825 15.590 47.965 26.480 ;
        RECT 48.385 15.590 48.525 26.480 ;
        RECT 48.945 15.590 49.085 26.480 ;
        RECT 49.505 15.590 49.645 26.480 ;
        RECT 50.065 15.590 50.205 26.480 ;
        RECT 50.625 15.590 50.765 26.480 ;
        RECT 51.185 15.590 51.325 26.480 ;
        RECT 51.745 15.590 51.885 26.480 ;
        RECT 52.305 15.590 52.445 26.480 ;
        RECT 52.865 15.590 53.005 26.480 ;
        RECT 53.425 15.590 53.565 26.480 ;
        RECT 53.985 15.590 54.125 26.480 ;
        RECT 54.545 15.590 54.685 26.480 ;
        RECT 55.105 15.590 55.245 26.480 ;
        RECT 55.665 15.590 55.805 26.480 ;
        RECT 56.225 15.590 56.365 26.480 ;
        RECT 56.785 15.590 56.925 26.480 ;
        RECT 59.195 15.590 59.335 26.480 ;
        RECT 59.755 15.590 59.895 26.480 ;
        RECT 60.315 15.590 60.455 26.480 ;
        RECT 60.875 15.590 61.015 26.480 ;
        RECT 61.435 15.590 61.575 26.480 ;
        RECT 61.995 15.590 62.135 26.480 ;
        RECT 62.555 15.590 62.695 26.480 ;
        RECT 63.115 15.590 63.255 26.480 ;
        RECT 63.675 15.590 63.815 26.480 ;
        RECT 64.235 15.590 64.375 26.480 ;
        RECT 64.795 15.590 64.935 26.480 ;
        RECT 65.355 15.590 65.495 26.480 ;
        RECT 65.915 15.590 66.055 26.480 ;
        RECT 66.475 15.590 66.615 26.480 ;
        RECT 67.035 15.590 67.175 26.480 ;
        RECT 67.595 15.590 67.735 26.480 ;
        RECT 68.155 15.590 68.295 26.480 ;
        RECT 68.715 15.590 68.855 26.480 ;
        RECT 69.275 15.590 69.415 26.480 ;
        RECT 69.835 15.590 69.975 26.480 ;
        RECT 72.285 15.590 72.425 26.480 ;
        RECT 72.845 15.590 72.985 26.480 ;
        RECT 73.405 15.590 73.545 26.480 ;
        RECT 73.965 15.590 74.105 26.480 ;
        RECT 74.525 15.590 74.665 26.480 ;
        RECT 75.085 15.590 75.225 26.480 ;
        RECT 75.645 15.590 75.785 26.480 ;
        RECT 76.205 15.590 76.345 26.480 ;
        RECT 76.765 15.590 76.905 26.480 ;
        RECT 77.325 15.590 77.465 26.480 ;
        RECT 77.885 15.590 78.025 26.480 ;
        RECT 78.445 15.590 78.585 26.480 ;
        RECT 79.005 15.590 79.145 26.480 ;
        RECT 79.565 15.590 79.705 26.480 ;
        RECT 80.125 15.590 80.265 26.480 ;
        RECT 80.685 15.590 80.825 26.480 ;
        RECT 81.245 15.590 81.385 26.480 ;
        RECT 81.805 15.590 81.945 26.480 ;
        RECT 82.365 15.590 82.505 26.480 ;
        RECT 82.925 15.590 83.065 26.480 ;
        RECT 32.775 15.260 44.185 15.590 ;
        RECT 45.865 15.260 57.275 15.590 ;
        RECT 58.915 15.260 70.325 15.590 ;
        RECT 72.005 15.260 83.415 15.590 ;
        RECT 85.375 15.570 85.515 26.460 ;
        RECT 85.935 15.570 86.075 26.460 ;
        RECT 86.495 15.570 86.635 26.460 ;
        RECT 87.055 15.570 87.195 26.460 ;
        RECT 87.615 15.570 87.755 26.460 ;
        RECT 88.175 15.570 88.315 26.460 ;
        RECT 88.735 15.570 88.875 26.460 ;
        RECT 89.295 15.570 89.435 26.460 ;
        RECT 89.855 15.570 89.995 26.460 ;
        RECT 90.415 15.570 90.555 26.460 ;
        RECT 90.975 15.570 91.115 26.460 ;
        RECT 91.535 15.570 91.675 26.460 ;
        RECT 92.095 15.570 92.235 26.460 ;
        RECT 92.655 15.570 92.795 26.460 ;
        RECT 93.215 15.570 93.355 26.460 ;
        RECT 93.775 15.570 93.915 26.460 ;
        RECT 94.335 15.570 94.475 26.460 ;
        RECT 94.895 15.570 95.035 26.460 ;
        RECT 95.455 15.570 95.595 26.460 ;
        RECT 96.015 15.570 96.155 26.460 ;
        RECT 98.465 15.570 98.605 26.460 ;
        RECT 99.025 15.570 99.165 26.460 ;
        RECT 99.585 15.570 99.725 26.460 ;
        RECT 100.145 15.570 100.285 26.460 ;
        RECT 100.705 15.570 100.845 26.460 ;
        RECT 101.265 15.570 101.405 26.460 ;
        RECT 101.825 15.570 101.965 26.460 ;
        RECT 102.385 15.570 102.525 26.460 ;
        RECT 102.945 15.570 103.085 26.460 ;
        RECT 103.505 15.570 103.645 26.460 ;
        RECT 104.065 15.570 104.205 26.460 ;
        RECT 104.625 15.570 104.765 26.460 ;
        RECT 105.185 15.570 105.325 26.460 ;
        RECT 105.745 15.570 105.885 26.460 ;
        RECT 106.305 15.570 106.445 26.460 ;
        RECT 106.865 15.570 107.005 26.460 ;
        RECT 107.425 15.570 107.565 26.460 ;
        RECT 107.985 15.570 108.125 26.460 ;
        RECT 108.545 15.570 108.685 26.460 ;
        RECT 109.105 15.570 109.245 26.460 ;
        RECT 111.555 15.570 111.695 26.460 ;
        RECT 112.115 15.570 112.255 26.460 ;
        RECT 112.675 15.570 112.815 26.460 ;
        RECT 113.235 15.570 113.375 26.460 ;
        RECT 113.795 15.570 113.935 26.460 ;
        RECT 114.355 15.570 114.495 26.460 ;
        RECT 114.915 15.570 115.055 26.460 ;
        RECT 115.475 15.570 115.615 26.460 ;
        RECT 116.035 15.570 116.175 26.460 ;
        RECT 116.595 15.570 116.735 26.460 ;
        RECT 117.155 15.570 117.295 26.460 ;
        RECT 117.715 15.570 117.855 26.460 ;
        RECT 118.275 15.570 118.415 26.460 ;
        RECT 118.835 15.570 118.975 26.460 ;
        RECT 119.395 15.570 119.535 26.460 ;
        RECT 119.955 15.570 120.095 26.460 ;
        RECT 120.515 15.570 120.655 26.460 ;
        RECT 121.075 15.570 121.215 26.460 ;
        RECT 121.635 15.570 121.775 26.460 ;
        RECT 122.195 15.570 122.335 26.460 ;
        RECT 124.645 15.570 124.785 26.460 ;
        RECT 125.205 15.570 125.345 26.460 ;
        RECT 125.765 15.570 125.905 26.460 ;
        RECT 126.325 15.570 126.465 26.460 ;
        RECT 126.885 15.570 127.025 26.460 ;
        RECT 127.445 15.570 127.585 26.460 ;
        RECT 128.005 15.570 128.145 26.460 ;
        RECT 128.565 15.570 128.705 26.460 ;
        RECT 129.125 15.570 129.265 26.460 ;
        RECT 129.685 15.570 129.825 26.460 ;
        RECT 130.245 15.570 130.385 26.460 ;
        RECT 130.805 15.570 130.945 26.460 ;
        RECT 131.365 15.570 131.505 26.460 ;
        RECT 131.925 15.570 132.065 26.460 ;
        RECT 132.485 15.570 132.625 26.460 ;
        RECT 133.045 15.570 133.185 26.460 ;
        RECT 133.605 15.570 133.745 26.460 ;
        RECT 134.165 15.570 134.305 26.460 ;
        RECT 134.725 15.570 134.865 26.460 ;
        RECT 135.285 15.570 135.425 26.460 ;
        RECT 85.095 15.240 96.505 15.570 ;
        RECT 98.185 15.240 109.595 15.570 ;
        RECT 111.275 15.240 122.685 15.570 ;
        RECT 124.365 15.240 135.775 15.570 ;
        RECT 137.735 15.550 137.875 26.440 ;
        RECT 138.295 15.550 138.435 26.440 ;
        RECT 138.855 15.550 138.995 26.440 ;
        RECT 139.415 15.550 139.555 26.440 ;
        RECT 139.975 15.550 140.115 26.440 ;
        RECT 140.535 15.550 140.675 26.440 ;
        RECT 141.095 15.550 141.235 26.440 ;
        RECT 141.655 15.550 141.795 26.440 ;
        RECT 142.215 15.550 142.355 26.440 ;
        RECT 142.775 15.550 142.915 26.440 ;
        RECT 143.335 15.550 143.475 26.440 ;
        RECT 143.895 15.550 144.035 26.440 ;
        RECT 144.455 15.550 144.595 26.440 ;
        RECT 145.015 15.550 145.155 26.440 ;
        RECT 145.575 15.550 145.715 26.440 ;
        RECT 146.135 15.550 146.275 26.440 ;
        RECT 146.695 15.550 146.835 26.440 ;
        RECT 147.255 15.550 147.395 26.440 ;
        RECT 147.815 15.550 147.955 26.440 ;
        RECT 148.375 15.550 148.515 26.440 ;
        RECT 150.825 15.550 150.965 26.440 ;
        RECT 151.385 15.550 151.525 26.440 ;
        RECT 151.945 15.550 152.085 26.440 ;
        RECT 152.505 15.550 152.645 26.440 ;
        RECT 153.065 15.550 153.205 26.440 ;
        RECT 153.625 15.550 153.765 26.440 ;
        RECT 154.185 15.550 154.325 26.440 ;
        RECT 154.745 15.550 154.885 26.440 ;
        RECT 155.305 15.550 155.445 26.440 ;
        RECT 155.865 15.550 156.005 26.440 ;
        RECT 156.425 15.550 156.565 26.440 ;
        RECT 156.985 15.550 157.125 26.440 ;
        RECT 157.545 15.550 157.685 26.440 ;
        RECT 158.105 15.550 158.245 26.440 ;
        RECT 158.665 15.550 158.805 26.440 ;
        RECT 159.225 15.550 159.365 26.440 ;
        RECT 159.785 15.550 159.925 26.440 ;
        RECT 160.345 15.550 160.485 26.440 ;
        RECT 160.905 15.550 161.045 26.440 ;
        RECT 161.465 15.550 161.605 26.440 ;
        RECT 137.455 15.220 148.865 15.550 ;
        RECT 150.545 15.220 161.955 15.550 ;
        RECT 6.625 13.230 18.035 13.560 ;
        RECT 19.715 13.230 31.125 13.560 ;
        RECT 32.805 13.250 44.215 13.580 ;
        RECT 45.895 13.250 57.305 13.580 ;
        RECT 58.945 13.250 70.355 13.580 ;
        RECT 72.035 13.250 83.445 13.580 ;
        RECT 85.125 13.270 96.535 13.600 ;
        RECT 98.215 13.270 109.625 13.600 ;
        RECT 111.305 13.270 122.715 13.600 ;
        RECT 124.395 13.270 135.805 13.600 ;
        RECT 137.485 13.290 148.895 13.620 ;
        RECT 150.575 13.290 161.985 13.620 ;
        RECT 6.905 2.340 7.045 13.230 ;
        RECT 7.465 2.340 7.605 13.230 ;
        RECT 8.025 2.340 8.165 13.230 ;
        RECT 8.585 2.340 8.725 13.230 ;
        RECT 9.145 2.340 9.285 13.230 ;
        RECT 9.705 2.340 9.845 13.230 ;
        RECT 10.265 2.340 10.405 13.230 ;
        RECT 10.825 2.340 10.965 13.230 ;
        RECT 11.385 2.340 11.525 13.230 ;
        RECT 11.945 2.340 12.085 13.230 ;
        RECT 12.505 2.340 12.645 13.230 ;
        RECT 13.065 2.340 13.205 13.230 ;
        RECT 13.625 2.340 13.765 13.230 ;
        RECT 14.185 2.340 14.325 13.230 ;
        RECT 14.745 2.340 14.885 13.230 ;
        RECT 15.305 2.340 15.445 13.230 ;
        RECT 15.865 2.340 16.005 13.230 ;
        RECT 16.425 2.340 16.565 13.230 ;
        RECT 16.985 2.340 17.125 13.230 ;
        RECT 17.545 2.340 17.685 13.230 ;
        RECT 19.995 2.340 20.135 13.230 ;
        RECT 20.555 2.340 20.695 13.230 ;
        RECT 21.115 2.340 21.255 13.230 ;
        RECT 21.675 2.340 21.815 13.230 ;
        RECT 22.235 2.340 22.375 13.230 ;
        RECT 22.795 2.340 22.935 13.230 ;
        RECT 23.355 2.340 23.495 13.230 ;
        RECT 23.915 2.340 24.055 13.230 ;
        RECT 24.475 2.340 24.615 13.230 ;
        RECT 25.035 2.340 25.175 13.230 ;
        RECT 25.595 2.340 25.735 13.230 ;
        RECT 26.155 2.340 26.295 13.230 ;
        RECT 26.715 2.340 26.855 13.230 ;
        RECT 27.275 2.340 27.415 13.230 ;
        RECT 27.835 2.340 27.975 13.230 ;
        RECT 28.395 2.340 28.535 13.230 ;
        RECT 28.955 2.340 29.095 13.230 ;
        RECT 29.515 2.340 29.655 13.230 ;
        RECT 30.075 2.340 30.215 13.230 ;
        RECT 30.635 2.340 30.775 13.230 ;
        RECT 33.085 2.360 33.225 13.250 ;
        RECT 33.645 2.360 33.785 13.250 ;
        RECT 34.205 2.360 34.345 13.250 ;
        RECT 34.765 2.360 34.905 13.250 ;
        RECT 35.325 2.360 35.465 13.250 ;
        RECT 35.885 2.360 36.025 13.250 ;
        RECT 36.445 2.360 36.585 13.250 ;
        RECT 37.005 2.360 37.145 13.250 ;
        RECT 37.565 2.360 37.705 13.250 ;
        RECT 38.125 2.360 38.265 13.250 ;
        RECT 38.685 2.360 38.825 13.250 ;
        RECT 39.245 2.360 39.385 13.250 ;
        RECT 39.805 2.360 39.945 13.250 ;
        RECT 40.365 2.360 40.505 13.250 ;
        RECT 40.925 2.360 41.065 13.250 ;
        RECT 41.485 2.360 41.625 13.250 ;
        RECT 42.045 2.360 42.185 13.250 ;
        RECT 42.605 2.360 42.745 13.250 ;
        RECT 43.165 2.360 43.305 13.250 ;
        RECT 43.725 2.360 43.865 13.250 ;
        RECT 46.175 2.360 46.315 13.250 ;
        RECT 46.735 2.360 46.875 13.250 ;
        RECT 47.295 2.360 47.435 13.250 ;
        RECT 47.855 2.360 47.995 13.250 ;
        RECT 48.415 2.360 48.555 13.250 ;
        RECT 48.975 2.360 49.115 13.250 ;
        RECT 49.535 2.360 49.675 13.250 ;
        RECT 50.095 2.360 50.235 13.250 ;
        RECT 50.655 2.360 50.795 13.250 ;
        RECT 51.215 2.360 51.355 13.250 ;
        RECT 51.775 2.360 51.915 13.250 ;
        RECT 52.335 2.360 52.475 13.250 ;
        RECT 52.895 2.360 53.035 13.250 ;
        RECT 53.455 2.360 53.595 13.250 ;
        RECT 54.015 2.360 54.155 13.250 ;
        RECT 54.575 2.360 54.715 13.250 ;
        RECT 55.135 2.360 55.275 13.250 ;
        RECT 55.695 2.360 55.835 13.250 ;
        RECT 56.255 2.360 56.395 13.250 ;
        RECT 56.815 2.360 56.955 13.250 ;
        RECT 59.225 2.360 59.365 13.250 ;
        RECT 59.785 2.360 59.925 13.250 ;
        RECT 60.345 2.360 60.485 13.250 ;
        RECT 60.905 2.360 61.045 13.250 ;
        RECT 61.465 2.360 61.605 13.250 ;
        RECT 62.025 2.360 62.165 13.250 ;
        RECT 62.585 2.360 62.725 13.250 ;
        RECT 63.145 2.360 63.285 13.250 ;
        RECT 63.705 2.360 63.845 13.250 ;
        RECT 64.265 2.360 64.405 13.250 ;
        RECT 64.825 2.360 64.965 13.250 ;
        RECT 65.385 2.360 65.525 13.250 ;
        RECT 65.945 2.360 66.085 13.250 ;
        RECT 66.505 2.360 66.645 13.250 ;
        RECT 67.065 2.360 67.205 13.250 ;
        RECT 67.625 2.360 67.765 13.250 ;
        RECT 68.185 2.360 68.325 13.250 ;
        RECT 68.745 2.360 68.885 13.250 ;
        RECT 69.305 2.360 69.445 13.250 ;
        RECT 69.865 2.360 70.005 13.250 ;
        RECT 72.315 2.360 72.455 13.250 ;
        RECT 72.875 2.360 73.015 13.250 ;
        RECT 73.435 2.360 73.575 13.250 ;
        RECT 73.995 2.360 74.135 13.250 ;
        RECT 74.555 2.360 74.695 13.250 ;
        RECT 75.115 2.360 75.255 13.250 ;
        RECT 75.675 2.360 75.815 13.250 ;
        RECT 76.235 2.360 76.375 13.250 ;
        RECT 76.795 2.360 76.935 13.250 ;
        RECT 77.355 2.360 77.495 13.250 ;
        RECT 77.915 2.360 78.055 13.250 ;
        RECT 78.475 2.360 78.615 13.250 ;
        RECT 79.035 2.360 79.175 13.250 ;
        RECT 79.595 2.360 79.735 13.250 ;
        RECT 80.155 2.360 80.295 13.250 ;
        RECT 80.715 2.360 80.855 13.250 ;
        RECT 81.275 2.360 81.415 13.250 ;
        RECT 81.835 2.360 81.975 13.250 ;
        RECT 82.395 2.360 82.535 13.250 ;
        RECT 82.955 2.360 83.095 13.250 ;
        RECT 85.405 2.380 85.545 13.270 ;
        RECT 85.965 2.380 86.105 13.270 ;
        RECT 86.525 2.380 86.665 13.270 ;
        RECT 87.085 2.380 87.225 13.270 ;
        RECT 87.645 2.380 87.785 13.270 ;
        RECT 88.205 2.380 88.345 13.270 ;
        RECT 88.765 2.380 88.905 13.270 ;
        RECT 89.325 2.380 89.465 13.270 ;
        RECT 89.885 2.380 90.025 13.270 ;
        RECT 90.445 2.380 90.585 13.270 ;
        RECT 91.005 2.380 91.145 13.270 ;
        RECT 91.565 2.380 91.705 13.270 ;
        RECT 92.125 2.380 92.265 13.270 ;
        RECT 92.685 2.380 92.825 13.270 ;
        RECT 93.245 2.380 93.385 13.270 ;
        RECT 93.805 2.380 93.945 13.270 ;
        RECT 94.365 2.380 94.505 13.270 ;
        RECT 94.925 2.380 95.065 13.270 ;
        RECT 95.485 2.380 95.625 13.270 ;
        RECT 96.045 2.380 96.185 13.270 ;
        RECT 98.495 2.380 98.635 13.270 ;
        RECT 99.055 2.380 99.195 13.270 ;
        RECT 99.615 2.380 99.755 13.270 ;
        RECT 100.175 2.380 100.315 13.270 ;
        RECT 100.735 2.380 100.875 13.270 ;
        RECT 101.295 2.380 101.435 13.270 ;
        RECT 101.855 2.380 101.995 13.270 ;
        RECT 102.415 2.380 102.555 13.270 ;
        RECT 102.975 2.380 103.115 13.270 ;
        RECT 103.535 2.380 103.675 13.270 ;
        RECT 104.095 2.380 104.235 13.270 ;
        RECT 104.655 2.380 104.795 13.270 ;
        RECT 105.215 2.380 105.355 13.270 ;
        RECT 105.775 2.380 105.915 13.270 ;
        RECT 106.335 2.380 106.475 13.270 ;
        RECT 106.895 2.380 107.035 13.270 ;
        RECT 107.455 2.380 107.595 13.270 ;
        RECT 108.015 2.380 108.155 13.270 ;
        RECT 108.575 2.380 108.715 13.270 ;
        RECT 109.135 2.380 109.275 13.270 ;
        RECT 111.585 2.380 111.725 13.270 ;
        RECT 112.145 2.380 112.285 13.270 ;
        RECT 112.705 2.380 112.845 13.270 ;
        RECT 113.265 2.380 113.405 13.270 ;
        RECT 113.825 2.380 113.965 13.270 ;
        RECT 114.385 2.380 114.525 13.270 ;
        RECT 114.945 2.380 115.085 13.270 ;
        RECT 115.505 2.380 115.645 13.270 ;
        RECT 116.065 2.380 116.205 13.270 ;
        RECT 116.625 2.380 116.765 13.270 ;
        RECT 117.185 2.380 117.325 13.270 ;
        RECT 117.745 2.380 117.885 13.270 ;
        RECT 118.305 2.380 118.445 13.270 ;
        RECT 118.865 2.380 119.005 13.270 ;
        RECT 119.425 2.380 119.565 13.270 ;
        RECT 119.985 2.380 120.125 13.270 ;
        RECT 120.545 2.380 120.685 13.270 ;
        RECT 121.105 2.380 121.245 13.270 ;
        RECT 121.665 2.380 121.805 13.270 ;
        RECT 122.225 2.380 122.365 13.270 ;
        RECT 124.675 2.380 124.815 13.270 ;
        RECT 125.235 2.380 125.375 13.270 ;
        RECT 125.795 2.380 125.935 13.270 ;
        RECT 126.355 2.380 126.495 13.270 ;
        RECT 126.915 2.380 127.055 13.270 ;
        RECT 127.475 2.380 127.615 13.270 ;
        RECT 128.035 2.380 128.175 13.270 ;
        RECT 128.595 2.380 128.735 13.270 ;
        RECT 129.155 2.380 129.295 13.270 ;
        RECT 129.715 2.380 129.855 13.270 ;
        RECT 130.275 2.380 130.415 13.270 ;
        RECT 130.835 2.380 130.975 13.270 ;
        RECT 131.395 2.380 131.535 13.270 ;
        RECT 131.955 2.380 132.095 13.270 ;
        RECT 132.515 2.380 132.655 13.270 ;
        RECT 133.075 2.380 133.215 13.270 ;
        RECT 133.635 2.380 133.775 13.270 ;
        RECT 134.195 2.380 134.335 13.270 ;
        RECT 134.755 2.380 134.895 13.270 ;
        RECT 135.315 2.380 135.455 13.270 ;
        RECT 137.765 2.400 137.905 13.290 ;
        RECT 138.325 2.400 138.465 13.290 ;
        RECT 138.885 2.400 139.025 13.290 ;
        RECT 139.445 2.400 139.585 13.290 ;
        RECT 140.005 2.400 140.145 13.290 ;
        RECT 140.565 2.400 140.705 13.290 ;
        RECT 141.125 2.400 141.265 13.290 ;
        RECT 141.685 2.400 141.825 13.290 ;
        RECT 142.245 2.400 142.385 13.290 ;
        RECT 142.805 2.400 142.945 13.290 ;
        RECT 143.365 2.400 143.505 13.290 ;
        RECT 143.925 2.400 144.065 13.290 ;
        RECT 144.485 2.400 144.625 13.290 ;
        RECT 145.045 2.400 145.185 13.290 ;
        RECT 145.605 2.400 145.745 13.290 ;
        RECT 146.165 2.400 146.305 13.290 ;
        RECT 146.725 2.400 146.865 13.290 ;
        RECT 147.285 2.400 147.425 13.290 ;
        RECT 147.845 2.400 147.985 13.290 ;
        RECT 148.405 2.400 148.545 13.290 ;
        RECT 150.855 2.400 150.995 13.290 ;
        RECT 151.415 2.400 151.555 13.290 ;
        RECT 151.975 2.400 152.115 13.290 ;
        RECT 152.535 2.400 152.675 13.290 ;
        RECT 153.095 2.400 153.235 13.290 ;
        RECT 153.655 2.400 153.795 13.290 ;
        RECT 154.215 2.400 154.355 13.290 ;
        RECT 154.775 2.400 154.915 13.290 ;
        RECT 155.335 2.400 155.475 13.290 ;
        RECT 155.895 2.400 156.035 13.290 ;
        RECT 156.455 2.400 156.595 13.290 ;
        RECT 157.015 2.400 157.155 13.290 ;
        RECT 157.575 2.400 157.715 13.290 ;
        RECT 158.135 2.400 158.275 13.290 ;
        RECT 158.695 2.400 158.835 13.290 ;
        RECT 159.255 2.400 159.395 13.290 ;
        RECT 159.815 2.400 159.955 13.290 ;
        RECT 160.375 2.400 160.515 13.290 ;
        RECT 160.935 2.400 161.075 13.290 ;
        RECT 161.495 2.400 161.635 13.290 ;
      LAYER via ;
        RECT 6.275 106.955 6.535 107.215 ;
        RECT 6.595 106.955 6.855 107.215 ;
        RECT 7.335 106.955 7.595 107.215 ;
        RECT 7.655 106.955 7.915 107.215 ;
        RECT 8.455 106.955 8.715 107.215 ;
        RECT 8.775 106.955 9.035 107.215 ;
        RECT 9.575 106.955 9.835 107.215 ;
        RECT 9.895 106.955 10.155 107.215 ;
        RECT 10.695 106.955 10.955 107.215 ;
        RECT 11.015 106.955 11.275 107.215 ;
        RECT 11.815 106.955 12.075 107.215 ;
        RECT 12.135 106.955 12.395 107.215 ;
        RECT 12.935 106.955 13.195 107.215 ;
        RECT 13.255 106.955 13.515 107.215 ;
        RECT 14.055 106.955 14.315 107.215 ;
        RECT 14.375 106.955 14.635 107.215 ;
        RECT 15.175 106.955 15.435 107.215 ;
        RECT 15.495 106.955 15.755 107.215 ;
        RECT 16.295 106.955 16.555 107.215 ;
        RECT 16.615 106.955 16.875 107.215 ;
        RECT 19.365 106.955 19.625 107.215 ;
        RECT 19.685 106.955 19.945 107.215 ;
        RECT 20.425 106.955 20.685 107.215 ;
        RECT 20.745 106.955 21.005 107.215 ;
        RECT 21.545 106.955 21.805 107.215 ;
        RECT 21.865 106.955 22.125 107.215 ;
        RECT 22.665 106.955 22.925 107.215 ;
        RECT 22.985 106.955 23.245 107.215 ;
        RECT 23.785 106.955 24.045 107.215 ;
        RECT 24.105 106.955 24.365 107.215 ;
        RECT 24.905 106.955 25.165 107.215 ;
        RECT 25.225 106.955 25.485 107.215 ;
        RECT 26.025 106.955 26.285 107.215 ;
        RECT 26.345 106.955 26.605 107.215 ;
        RECT 27.145 106.955 27.405 107.215 ;
        RECT 27.465 106.955 27.725 107.215 ;
        RECT 28.265 106.955 28.525 107.215 ;
        RECT 28.585 106.955 28.845 107.215 ;
        RECT 29.385 106.955 29.645 107.215 ;
        RECT 29.705 106.955 29.965 107.215 ;
        RECT 32.455 106.935 32.715 107.195 ;
        RECT 32.775 106.935 33.035 107.195 ;
        RECT 33.515 106.935 33.775 107.195 ;
        RECT 33.835 106.935 34.095 107.195 ;
        RECT 34.635 106.935 34.895 107.195 ;
        RECT 34.955 106.935 35.215 107.195 ;
        RECT 35.755 106.935 36.015 107.195 ;
        RECT 36.075 106.935 36.335 107.195 ;
        RECT 36.875 106.935 37.135 107.195 ;
        RECT 37.195 106.935 37.455 107.195 ;
        RECT 37.995 106.935 38.255 107.195 ;
        RECT 38.315 106.935 38.575 107.195 ;
        RECT 39.115 106.935 39.375 107.195 ;
        RECT 39.435 106.935 39.695 107.195 ;
        RECT 40.235 106.935 40.495 107.195 ;
        RECT 40.555 106.935 40.815 107.195 ;
        RECT 41.355 106.935 41.615 107.195 ;
        RECT 41.675 106.935 41.935 107.195 ;
        RECT 42.475 106.935 42.735 107.195 ;
        RECT 42.795 106.935 43.055 107.195 ;
        RECT 45.545 106.935 45.805 107.195 ;
        RECT 45.865 106.935 46.125 107.195 ;
        RECT 46.605 106.935 46.865 107.195 ;
        RECT 46.925 106.935 47.185 107.195 ;
        RECT 47.725 106.935 47.985 107.195 ;
        RECT 48.045 106.935 48.305 107.195 ;
        RECT 48.845 106.935 49.105 107.195 ;
        RECT 49.165 106.935 49.425 107.195 ;
        RECT 49.965 106.935 50.225 107.195 ;
        RECT 50.285 106.935 50.545 107.195 ;
        RECT 51.085 106.935 51.345 107.195 ;
        RECT 51.405 106.935 51.665 107.195 ;
        RECT 52.205 106.935 52.465 107.195 ;
        RECT 52.525 106.935 52.785 107.195 ;
        RECT 53.325 106.935 53.585 107.195 ;
        RECT 53.645 106.935 53.905 107.195 ;
        RECT 54.445 106.935 54.705 107.195 ;
        RECT 54.765 106.935 55.025 107.195 ;
        RECT 55.565 106.935 55.825 107.195 ;
        RECT 55.885 106.935 56.145 107.195 ;
        RECT 58.595 106.935 58.855 107.195 ;
        RECT 58.915 106.935 59.175 107.195 ;
        RECT 59.655 106.935 59.915 107.195 ;
        RECT 59.975 106.935 60.235 107.195 ;
        RECT 60.775 106.935 61.035 107.195 ;
        RECT 61.095 106.935 61.355 107.195 ;
        RECT 61.895 106.935 62.155 107.195 ;
        RECT 62.215 106.935 62.475 107.195 ;
        RECT 63.015 106.935 63.275 107.195 ;
        RECT 63.335 106.935 63.595 107.195 ;
        RECT 64.135 106.935 64.395 107.195 ;
        RECT 64.455 106.935 64.715 107.195 ;
        RECT 65.255 106.935 65.515 107.195 ;
        RECT 65.575 106.935 65.835 107.195 ;
        RECT 66.375 106.935 66.635 107.195 ;
        RECT 66.695 106.935 66.955 107.195 ;
        RECT 67.495 106.935 67.755 107.195 ;
        RECT 67.815 106.935 68.075 107.195 ;
        RECT 68.615 106.935 68.875 107.195 ;
        RECT 68.935 106.935 69.195 107.195 ;
        RECT 71.685 106.935 71.945 107.195 ;
        RECT 72.005 106.935 72.265 107.195 ;
        RECT 72.745 106.935 73.005 107.195 ;
        RECT 73.065 106.935 73.325 107.195 ;
        RECT 73.865 106.935 74.125 107.195 ;
        RECT 74.185 106.935 74.445 107.195 ;
        RECT 74.985 106.935 75.245 107.195 ;
        RECT 75.305 106.935 75.565 107.195 ;
        RECT 76.105 106.935 76.365 107.195 ;
        RECT 76.425 106.935 76.685 107.195 ;
        RECT 77.225 106.935 77.485 107.195 ;
        RECT 77.545 106.935 77.805 107.195 ;
        RECT 78.345 106.935 78.605 107.195 ;
        RECT 78.665 106.935 78.925 107.195 ;
        RECT 79.465 106.935 79.725 107.195 ;
        RECT 79.785 106.935 80.045 107.195 ;
        RECT 80.585 106.935 80.845 107.195 ;
        RECT 80.905 106.935 81.165 107.195 ;
        RECT 81.705 106.935 81.965 107.195 ;
        RECT 82.025 106.935 82.285 107.195 ;
        RECT 84.775 106.915 85.035 107.175 ;
        RECT 85.095 106.915 85.355 107.175 ;
        RECT 85.835 106.915 86.095 107.175 ;
        RECT 86.155 106.915 86.415 107.175 ;
        RECT 86.955 106.915 87.215 107.175 ;
        RECT 87.275 106.915 87.535 107.175 ;
        RECT 88.075 106.915 88.335 107.175 ;
        RECT 88.395 106.915 88.655 107.175 ;
        RECT 89.195 106.915 89.455 107.175 ;
        RECT 89.515 106.915 89.775 107.175 ;
        RECT 90.315 106.915 90.575 107.175 ;
        RECT 90.635 106.915 90.895 107.175 ;
        RECT 91.435 106.915 91.695 107.175 ;
        RECT 91.755 106.915 92.015 107.175 ;
        RECT 92.555 106.915 92.815 107.175 ;
        RECT 92.875 106.915 93.135 107.175 ;
        RECT 93.675 106.915 93.935 107.175 ;
        RECT 93.995 106.915 94.255 107.175 ;
        RECT 94.795 106.915 95.055 107.175 ;
        RECT 95.115 106.915 95.375 107.175 ;
        RECT 97.865 106.915 98.125 107.175 ;
        RECT 98.185 106.915 98.445 107.175 ;
        RECT 98.925 106.915 99.185 107.175 ;
        RECT 99.245 106.915 99.505 107.175 ;
        RECT 100.045 106.915 100.305 107.175 ;
        RECT 100.365 106.915 100.625 107.175 ;
        RECT 101.165 106.915 101.425 107.175 ;
        RECT 101.485 106.915 101.745 107.175 ;
        RECT 102.285 106.915 102.545 107.175 ;
        RECT 102.605 106.915 102.865 107.175 ;
        RECT 103.405 106.915 103.665 107.175 ;
        RECT 103.725 106.915 103.985 107.175 ;
        RECT 104.525 106.915 104.785 107.175 ;
        RECT 104.845 106.915 105.105 107.175 ;
        RECT 105.645 106.915 105.905 107.175 ;
        RECT 105.965 106.915 106.225 107.175 ;
        RECT 106.765 106.915 107.025 107.175 ;
        RECT 107.085 106.915 107.345 107.175 ;
        RECT 107.885 106.915 108.145 107.175 ;
        RECT 108.205 106.915 108.465 107.175 ;
        RECT 110.955 106.915 111.215 107.175 ;
        RECT 111.275 106.915 111.535 107.175 ;
        RECT 112.015 106.915 112.275 107.175 ;
        RECT 112.335 106.915 112.595 107.175 ;
        RECT 113.135 106.915 113.395 107.175 ;
        RECT 113.455 106.915 113.715 107.175 ;
        RECT 114.255 106.915 114.515 107.175 ;
        RECT 114.575 106.915 114.835 107.175 ;
        RECT 115.375 106.915 115.635 107.175 ;
        RECT 115.695 106.915 115.955 107.175 ;
        RECT 116.495 106.915 116.755 107.175 ;
        RECT 116.815 106.915 117.075 107.175 ;
        RECT 117.615 106.915 117.875 107.175 ;
        RECT 117.935 106.915 118.195 107.175 ;
        RECT 118.735 106.915 118.995 107.175 ;
        RECT 119.055 106.915 119.315 107.175 ;
        RECT 119.855 106.915 120.115 107.175 ;
        RECT 120.175 106.915 120.435 107.175 ;
        RECT 120.975 106.915 121.235 107.175 ;
        RECT 121.295 106.915 121.555 107.175 ;
        RECT 124.045 106.915 124.305 107.175 ;
        RECT 124.365 106.915 124.625 107.175 ;
        RECT 125.105 106.915 125.365 107.175 ;
        RECT 125.425 106.915 125.685 107.175 ;
        RECT 126.225 106.915 126.485 107.175 ;
        RECT 126.545 106.915 126.805 107.175 ;
        RECT 127.345 106.915 127.605 107.175 ;
        RECT 127.665 106.915 127.925 107.175 ;
        RECT 128.465 106.915 128.725 107.175 ;
        RECT 128.785 106.915 129.045 107.175 ;
        RECT 129.585 106.915 129.845 107.175 ;
        RECT 129.905 106.915 130.165 107.175 ;
        RECT 130.705 106.915 130.965 107.175 ;
        RECT 131.025 106.915 131.285 107.175 ;
        RECT 131.825 106.915 132.085 107.175 ;
        RECT 132.145 106.915 132.405 107.175 ;
        RECT 132.945 106.915 133.205 107.175 ;
        RECT 133.265 106.915 133.525 107.175 ;
        RECT 134.065 106.915 134.325 107.175 ;
        RECT 134.385 106.915 134.645 107.175 ;
        RECT 137.135 106.895 137.395 107.155 ;
        RECT 137.455 106.895 137.715 107.155 ;
        RECT 138.195 106.895 138.455 107.155 ;
        RECT 138.515 106.895 138.775 107.155 ;
        RECT 139.315 106.895 139.575 107.155 ;
        RECT 139.635 106.895 139.895 107.155 ;
        RECT 140.435 106.895 140.695 107.155 ;
        RECT 140.755 106.895 141.015 107.155 ;
        RECT 141.555 106.895 141.815 107.155 ;
        RECT 141.875 106.895 142.135 107.155 ;
        RECT 142.675 106.895 142.935 107.155 ;
        RECT 142.995 106.895 143.255 107.155 ;
        RECT 143.795 106.895 144.055 107.155 ;
        RECT 144.115 106.895 144.375 107.155 ;
        RECT 144.915 106.895 145.175 107.155 ;
        RECT 145.235 106.895 145.495 107.155 ;
        RECT 146.035 106.895 146.295 107.155 ;
        RECT 146.355 106.895 146.615 107.155 ;
        RECT 147.155 106.895 147.415 107.155 ;
        RECT 147.475 106.895 147.735 107.155 ;
        RECT 150.225 106.895 150.485 107.155 ;
        RECT 150.545 106.895 150.805 107.155 ;
        RECT 151.285 106.895 151.545 107.155 ;
        RECT 151.605 106.895 151.865 107.155 ;
        RECT 152.405 106.895 152.665 107.155 ;
        RECT 152.725 106.895 152.985 107.155 ;
        RECT 153.525 106.895 153.785 107.155 ;
        RECT 153.845 106.895 154.105 107.155 ;
        RECT 154.645 106.895 154.905 107.155 ;
        RECT 154.965 106.895 155.225 107.155 ;
        RECT 155.765 106.895 156.025 107.155 ;
        RECT 156.085 106.895 156.345 107.155 ;
        RECT 156.885 106.895 157.145 107.155 ;
        RECT 157.205 106.895 157.465 107.155 ;
        RECT 158.005 106.895 158.265 107.155 ;
        RECT 158.325 106.895 158.585 107.155 ;
        RECT 159.125 106.895 159.385 107.155 ;
        RECT 159.445 106.895 159.705 107.155 ;
        RECT 160.245 106.895 160.505 107.155 ;
        RECT 160.565 106.895 160.825 107.155 ;
        RECT 6.305 104.905 6.565 105.165 ;
        RECT 6.625 104.905 6.885 105.165 ;
        RECT 7.365 104.905 7.625 105.165 ;
        RECT 7.685 104.905 7.945 105.165 ;
        RECT 8.485 104.905 8.745 105.165 ;
        RECT 8.805 104.905 9.065 105.165 ;
        RECT 9.605 104.905 9.865 105.165 ;
        RECT 9.925 104.905 10.185 105.165 ;
        RECT 10.725 104.905 10.985 105.165 ;
        RECT 11.045 104.905 11.305 105.165 ;
        RECT 11.845 104.905 12.105 105.165 ;
        RECT 12.165 104.905 12.425 105.165 ;
        RECT 12.965 104.905 13.225 105.165 ;
        RECT 13.285 104.905 13.545 105.165 ;
        RECT 14.085 104.905 14.345 105.165 ;
        RECT 14.405 104.905 14.665 105.165 ;
        RECT 15.205 104.905 15.465 105.165 ;
        RECT 15.525 104.905 15.785 105.165 ;
        RECT 16.325 104.905 16.585 105.165 ;
        RECT 16.645 104.905 16.905 105.165 ;
        RECT 19.395 104.905 19.655 105.165 ;
        RECT 19.715 104.905 19.975 105.165 ;
        RECT 20.455 104.905 20.715 105.165 ;
        RECT 20.775 104.905 21.035 105.165 ;
        RECT 21.575 104.905 21.835 105.165 ;
        RECT 21.895 104.905 22.155 105.165 ;
        RECT 22.695 104.905 22.955 105.165 ;
        RECT 23.015 104.905 23.275 105.165 ;
        RECT 23.815 104.905 24.075 105.165 ;
        RECT 24.135 104.905 24.395 105.165 ;
        RECT 24.935 104.905 25.195 105.165 ;
        RECT 25.255 104.905 25.515 105.165 ;
        RECT 26.055 104.905 26.315 105.165 ;
        RECT 26.375 104.905 26.635 105.165 ;
        RECT 27.175 104.905 27.435 105.165 ;
        RECT 27.495 104.905 27.755 105.165 ;
        RECT 28.295 104.905 28.555 105.165 ;
        RECT 28.615 104.905 28.875 105.165 ;
        RECT 29.415 104.905 29.675 105.165 ;
        RECT 29.735 104.905 29.995 105.165 ;
        RECT 32.485 104.925 32.745 105.185 ;
        RECT 32.805 104.925 33.065 105.185 ;
        RECT 33.545 104.925 33.805 105.185 ;
        RECT 33.865 104.925 34.125 105.185 ;
        RECT 34.665 104.925 34.925 105.185 ;
        RECT 34.985 104.925 35.245 105.185 ;
        RECT 35.785 104.925 36.045 105.185 ;
        RECT 36.105 104.925 36.365 105.185 ;
        RECT 36.905 104.925 37.165 105.185 ;
        RECT 37.225 104.925 37.485 105.185 ;
        RECT 38.025 104.925 38.285 105.185 ;
        RECT 38.345 104.925 38.605 105.185 ;
        RECT 39.145 104.925 39.405 105.185 ;
        RECT 39.465 104.925 39.725 105.185 ;
        RECT 40.265 104.925 40.525 105.185 ;
        RECT 40.585 104.925 40.845 105.185 ;
        RECT 41.385 104.925 41.645 105.185 ;
        RECT 41.705 104.925 41.965 105.185 ;
        RECT 42.505 104.925 42.765 105.185 ;
        RECT 42.825 104.925 43.085 105.185 ;
        RECT 45.575 104.925 45.835 105.185 ;
        RECT 45.895 104.925 46.155 105.185 ;
        RECT 46.635 104.925 46.895 105.185 ;
        RECT 46.955 104.925 47.215 105.185 ;
        RECT 47.755 104.925 48.015 105.185 ;
        RECT 48.075 104.925 48.335 105.185 ;
        RECT 48.875 104.925 49.135 105.185 ;
        RECT 49.195 104.925 49.455 105.185 ;
        RECT 49.995 104.925 50.255 105.185 ;
        RECT 50.315 104.925 50.575 105.185 ;
        RECT 51.115 104.925 51.375 105.185 ;
        RECT 51.435 104.925 51.695 105.185 ;
        RECT 52.235 104.925 52.495 105.185 ;
        RECT 52.555 104.925 52.815 105.185 ;
        RECT 53.355 104.925 53.615 105.185 ;
        RECT 53.675 104.925 53.935 105.185 ;
        RECT 54.475 104.925 54.735 105.185 ;
        RECT 54.795 104.925 55.055 105.185 ;
        RECT 55.595 104.925 55.855 105.185 ;
        RECT 55.915 104.925 56.175 105.185 ;
        RECT 58.625 104.925 58.885 105.185 ;
        RECT 58.945 104.925 59.205 105.185 ;
        RECT 59.685 104.925 59.945 105.185 ;
        RECT 60.005 104.925 60.265 105.185 ;
        RECT 60.805 104.925 61.065 105.185 ;
        RECT 61.125 104.925 61.385 105.185 ;
        RECT 61.925 104.925 62.185 105.185 ;
        RECT 62.245 104.925 62.505 105.185 ;
        RECT 63.045 104.925 63.305 105.185 ;
        RECT 63.365 104.925 63.625 105.185 ;
        RECT 64.165 104.925 64.425 105.185 ;
        RECT 64.485 104.925 64.745 105.185 ;
        RECT 65.285 104.925 65.545 105.185 ;
        RECT 65.605 104.925 65.865 105.185 ;
        RECT 66.405 104.925 66.665 105.185 ;
        RECT 66.725 104.925 66.985 105.185 ;
        RECT 67.525 104.925 67.785 105.185 ;
        RECT 67.845 104.925 68.105 105.185 ;
        RECT 68.645 104.925 68.905 105.185 ;
        RECT 68.965 104.925 69.225 105.185 ;
        RECT 71.715 104.925 71.975 105.185 ;
        RECT 72.035 104.925 72.295 105.185 ;
        RECT 72.775 104.925 73.035 105.185 ;
        RECT 73.095 104.925 73.355 105.185 ;
        RECT 73.895 104.925 74.155 105.185 ;
        RECT 74.215 104.925 74.475 105.185 ;
        RECT 75.015 104.925 75.275 105.185 ;
        RECT 75.335 104.925 75.595 105.185 ;
        RECT 76.135 104.925 76.395 105.185 ;
        RECT 76.455 104.925 76.715 105.185 ;
        RECT 77.255 104.925 77.515 105.185 ;
        RECT 77.575 104.925 77.835 105.185 ;
        RECT 78.375 104.925 78.635 105.185 ;
        RECT 78.695 104.925 78.955 105.185 ;
        RECT 79.495 104.925 79.755 105.185 ;
        RECT 79.815 104.925 80.075 105.185 ;
        RECT 80.615 104.925 80.875 105.185 ;
        RECT 80.935 104.925 81.195 105.185 ;
        RECT 81.735 104.925 81.995 105.185 ;
        RECT 82.055 104.925 82.315 105.185 ;
        RECT 84.805 104.945 85.065 105.205 ;
        RECT 85.125 104.945 85.385 105.205 ;
        RECT 85.865 104.945 86.125 105.205 ;
        RECT 86.185 104.945 86.445 105.205 ;
        RECT 86.985 104.945 87.245 105.205 ;
        RECT 87.305 104.945 87.565 105.205 ;
        RECT 88.105 104.945 88.365 105.205 ;
        RECT 88.425 104.945 88.685 105.205 ;
        RECT 89.225 104.945 89.485 105.205 ;
        RECT 89.545 104.945 89.805 105.205 ;
        RECT 90.345 104.945 90.605 105.205 ;
        RECT 90.665 104.945 90.925 105.205 ;
        RECT 91.465 104.945 91.725 105.205 ;
        RECT 91.785 104.945 92.045 105.205 ;
        RECT 92.585 104.945 92.845 105.205 ;
        RECT 92.905 104.945 93.165 105.205 ;
        RECT 93.705 104.945 93.965 105.205 ;
        RECT 94.025 104.945 94.285 105.205 ;
        RECT 94.825 104.945 95.085 105.205 ;
        RECT 95.145 104.945 95.405 105.205 ;
        RECT 97.895 104.945 98.155 105.205 ;
        RECT 98.215 104.945 98.475 105.205 ;
        RECT 98.955 104.945 99.215 105.205 ;
        RECT 99.275 104.945 99.535 105.205 ;
        RECT 100.075 104.945 100.335 105.205 ;
        RECT 100.395 104.945 100.655 105.205 ;
        RECT 101.195 104.945 101.455 105.205 ;
        RECT 101.515 104.945 101.775 105.205 ;
        RECT 102.315 104.945 102.575 105.205 ;
        RECT 102.635 104.945 102.895 105.205 ;
        RECT 103.435 104.945 103.695 105.205 ;
        RECT 103.755 104.945 104.015 105.205 ;
        RECT 104.555 104.945 104.815 105.205 ;
        RECT 104.875 104.945 105.135 105.205 ;
        RECT 105.675 104.945 105.935 105.205 ;
        RECT 105.995 104.945 106.255 105.205 ;
        RECT 106.795 104.945 107.055 105.205 ;
        RECT 107.115 104.945 107.375 105.205 ;
        RECT 107.915 104.945 108.175 105.205 ;
        RECT 108.235 104.945 108.495 105.205 ;
        RECT 110.985 104.945 111.245 105.205 ;
        RECT 111.305 104.945 111.565 105.205 ;
        RECT 112.045 104.945 112.305 105.205 ;
        RECT 112.365 104.945 112.625 105.205 ;
        RECT 113.165 104.945 113.425 105.205 ;
        RECT 113.485 104.945 113.745 105.205 ;
        RECT 114.285 104.945 114.545 105.205 ;
        RECT 114.605 104.945 114.865 105.205 ;
        RECT 115.405 104.945 115.665 105.205 ;
        RECT 115.725 104.945 115.985 105.205 ;
        RECT 116.525 104.945 116.785 105.205 ;
        RECT 116.845 104.945 117.105 105.205 ;
        RECT 117.645 104.945 117.905 105.205 ;
        RECT 117.965 104.945 118.225 105.205 ;
        RECT 118.765 104.945 119.025 105.205 ;
        RECT 119.085 104.945 119.345 105.205 ;
        RECT 119.885 104.945 120.145 105.205 ;
        RECT 120.205 104.945 120.465 105.205 ;
        RECT 121.005 104.945 121.265 105.205 ;
        RECT 121.325 104.945 121.585 105.205 ;
        RECT 124.075 104.945 124.335 105.205 ;
        RECT 124.395 104.945 124.655 105.205 ;
        RECT 125.135 104.945 125.395 105.205 ;
        RECT 125.455 104.945 125.715 105.205 ;
        RECT 126.255 104.945 126.515 105.205 ;
        RECT 126.575 104.945 126.835 105.205 ;
        RECT 127.375 104.945 127.635 105.205 ;
        RECT 127.695 104.945 127.955 105.205 ;
        RECT 128.495 104.945 128.755 105.205 ;
        RECT 128.815 104.945 129.075 105.205 ;
        RECT 129.615 104.945 129.875 105.205 ;
        RECT 129.935 104.945 130.195 105.205 ;
        RECT 130.735 104.945 130.995 105.205 ;
        RECT 131.055 104.945 131.315 105.205 ;
        RECT 131.855 104.945 132.115 105.205 ;
        RECT 132.175 104.945 132.435 105.205 ;
        RECT 132.975 104.945 133.235 105.205 ;
        RECT 133.295 104.945 133.555 105.205 ;
        RECT 134.095 104.945 134.355 105.205 ;
        RECT 134.415 104.945 134.675 105.205 ;
        RECT 137.165 104.965 137.425 105.225 ;
        RECT 137.485 104.965 137.745 105.225 ;
        RECT 138.225 104.965 138.485 105.225 ;
        RECT 138.545 104.965 138.805 105.225 ;
        RECT 139.345 104.965 139.605 105.225 ;
        RECT 139.665 104.965 139.925 105.225 ;
        RECT 140.465 104.965 140.725 105.225 ;
        RECT 140.785 104.965 141.045 105.225 ;
        RECT 141.585 104.965 141.845 105.225 ;
        RECT 141.905 104.965 142.165 105.225 ;
        RECT 142.705 104.965 142.965 105.225 ;
        RECT 143.025 104.965 143.285 105.225 ;
        RECT 143.825 104.965 144.085 105.225 ;
        RECT 144.145 104.965 144.405 105.225 ;
        RECT 144.945 104.965 145.205 105.225 ;
        RECT 145.265 104.965 145.525 105.225 ;
        RECT 146.065 104.965 146.325 105.225 ;
        RECT 146.385 104.965 146.645 105.225 ;
        RECT 147.185 104.965 147.445 105.225 ;
        RECT 147.505 104.965 147.765 105.225 ;
        RECT 150.255 104.965 150.515 105.225 ;
        RECT 150.575 104.965 150.835 105.225 ;
        RECT 151.315 104.965 151.575 105.225 ;
        RECT 151.635 104.965 151.895 105.225 ;
        RECT 152.435 104.965 152.695 105.225 ;
        RECT 152.755 104.965 153.015 105.225 ;
        RECT 153.555 104.965 153.815 105.225 ;
        RECT 153.875 104.965 154.135 105.225 ;
        RECT 154.675 104.965 154.935 105.225 ;
        RECT 154.995 104.965 155.255 105.225 ;
        RECT 155.795 104.965 156.055 105.225 ;
        RECT 156.115 104.965 156.375 105.225 ;
        RECT 156.915 104.965 157.175 105.225 ;
        RECT 157.235 104.965 157.495 105.225 ;
        RECT 158.035 104.965 158.295 105.225 ;
        RECT 158.355 104.965 158.615 105.225 ;
        RECT 159.155 104.965 159.415 105.225 ;
        RECT 159.475 104.965 159.735 105.225 ;
        RECT 160.275 104.965 160.535 105.225 ;
        RECT 160.595 104.965 160.855 105.225 ;
        RECT 162.875 90.270 163.350 90.745 ;
        RECT 4.760 88.675 5.230 89.145 ;
        RECT 19.725 81.625 19.985 81.885 ;
        RECT 29.340 81.625 29.600 81.885 ;
        RECT 38.955 81.625 39.215 81.885 ;
        RECT 48.570 81.625 48.830 81.885 ;
        RECT 18.610 76.360 18.870 76.620 ;
        RECT 28.225 76.360 28.485 76.620 ;
        RECT 37.840 76.360 38.100 76.620 ;
        RECT 47.455 76.360 47.715 76.620 ;
        RECT 171.720 65.450 171.980 65.710 ;
        RECT 171.720 65.130 171.980 65.390 ;
        RECT 171.720 63.880 171.980 64.140 ;
        RECT 171.720 63.560 171.980 63.820 ;
        RECT 171.720 62.310 171.980 62.570 ;
        RECT 171.720 61.990 171.980 62.250 ;
        RECT 171.720 59.260 171.980 59.520 ;
        RECT 171.720 58.940 171.980 59.200 ;
        RECT 171.720 57.690 171.980 57.950 ;
        RECT 171.720 57.370 171.980 57.630 ;
        RECT 171.720 56.120 171.980 56.380 ;
        RECT 171.720 55.800 171.980 56.060 ;
        RECT 18.610 43.230 18.870 43.490 ;
        RECT 28.225 43.230 28.485 43.490 ;
        RECT 37.840 43.230 38.100 43.490 ;
        RECT 47.455 43.230 47.715 43.490 ;
        RECT 19.725 37.965 19.985 38.225 ;
        RECT 29.340 37.965 29.600 38.225 ;
        RECT 38.955 37.965 39.215 38.225 ;
        RECT 48.570 37.965 48.830 38.225 ;
        RECT 4.750 33.215 5.220 33.685 ;
        RECT 148.780 31.360 149.040 31.620 ;
        RECT 150.975 29.300 151.235 29.560 ;
        RECT 163.275 29.215 163.750 29.690 ;
        RECT 6.715 15.315 6.975 15.575 ;
        RECT 7.035 15.315 7.295 15.575 ;
        RECT 7.775 15.315 8.035 15.575 ;
        RECT 8.095 15.315 8.355 15.575 ;
        RECT 8.895 15.315 9.155 15.575 ;
        RECT 9.215 15.315 9.475 15.575 ;
        RECT 10.015 15.315 10.275 15.575 ;
        RECT 10.335 15.315 10.595 15.575 ;
        RECT 11.135 15.315 11.395 15.575 ;
        RECT 11.455 15.315 11.715 15.575 ;
        RECT 12.255 15.315 12.515 15.575 ;
        RECT 12.575 15.315 12.835 15.575 ;
        RECT 13.375 15.315 13.635 15.575 ;
        RECT 13.695 15.315 13.955 15.575 ;
        RECT 14.495 15.315 14.755 15.575 ;
        RECT 14.815 15.315 15.075 15.575 ;
        RECT 15.615 15.315 15.875 15.575 ;
        RECT 15.935 15.315 16.195 15.575 ;
        RECT 16.735 15.315 16.995 15.575 ;
        RECT 17.055 15.315 17.315 15.575 ;
        RECT 19.805 15.315 20.065 15.575 ;
        RECT 20.125 15.315 20.385 15.575 ;
        RECT 20.865 15.315 21.125 15.575 ;
        RECT 21.185 15.315 21.445 15.575 ;
        RECT 21.985 15.315 22.245 15.575 ;
        RECT 22.305 15.315 22.565 15.575 ;
        RECT 23.105 15.315 23.365 15.575 ;
        RECT 23.425 15.315 23.685 15.575 ;
        RECT 24.225 15.315 24.485 15.575 ;
        RECT 24.545 15.315 24.805 15.575 ;
        RECT 25.345 15.315 25.605 15.575 ;
        RECT 25.665 15.315 25.925 15.575 ;
        RECT 26.465 15.315 26.725 15.575 ;
        RECT 26.785 15.315 27.045 15.575 ;
        RECT 27.585 15.315 27.845 15.575 ;
        RECT 27.905 15.315 28.165 15.575 ;
        RECT 28.705 15.315 28.965 15.575 ;
        RECT 29.025 15.315 29.285 15.575 ;
        RECT 29.825 15.315 30.085 15.575 ;
        RECT 30.145 15.315 30.405 15.575 ;
        RECT 32.895 15.295 33.155 15.555 ;
        RECT 33.215 15.295 33.475 15.555 ;
        RECT 33.955 15.295 34.215 15.555 ;
        RECT 34.275 15.295 34.535 15.555 ;
        RECT 35.075 15.295 35.335 15.555 ;
        RECT 35.395 15.295 35.655 15.555 ;
        RECT 36.195 15.295 36.455 15.555 ;
        RECT 36.515 15.295 36.775 15.555 ;
        RECT 37.315 15.295 37.575 15.555 ;
        RECT 37.635 15.295 37.895 15.555 ;
        RECT 38.435 15.295 38.695 15.555 ;
        RECT 38.755 15.295 39.015 15.555 ;
        RECT 39.555 15.295 39.815 15.555 ;
        RECT 39.875 15.295 40.135 15.555 ;
        RECT 40.675 15.295 40.935 15.555 ;
        RECT 40.995 15.295 41.255 15.555 ;
        RECT 41.795 15.295 42.055 15.555 ;
        RECT 42.115 15.295 42.375 15.555 ;
        RECT 42.915 15.295 43.175 15.555 ;
        RECT 43.235 15.295 43.495 15.555 ;
        RECT 45.985 15.295 46.245 15.555 ;
        RECT 46.305 15.295 46.565 15.555 ;
        RECT 47.045 15.295 47.305 15.555 ;
        RECT 47.365 15.295 47.625 15.555 ;
        RECT 48.165 15.295 48.425 15.555 ;
        RECT 48.485 15.295 48.745 15.555 ;
        RECT 49.285 15.295 49.545 15.555 ;
        RECT 49.605 15.295 49.865 15.555 ;
        RECT 50.405 15.295 50.665 15.555 ;
        RECT 50.725 15.295 50.985 15.555 ;
        RECT 51.525 15.295 51.785 15.555 ;
        RECT 51.845 15.295 52.105 15.555 ;
        RECT 52.645 15.295 52.905 15.555 ;
        RECT 52.965 15.295 53.225 15.555 ;
        RECT 53.765 15.295 54.025 15.555 ;
        RECT 54.085 15.295 54.345 15.555 ;
        RECT 54.885 15.295 55.145 15.555 ;
        RECT 55.205 15.295 55.465 15.555 ;
        RECT 56.005 15.295 56.265 15.555 ;
        RECT 56.325 15.295 56.585 15.555 ;
        RECT 59.035 15.295 59.295 15.555 ;
        RECT 59.355 15.295 59.615 15.555 ;
        RECT 60.095 15.295 60.355 15.555 ;
        RECT 60.415 15.295 60.675 15.555 ;
        RECT 61.215 15.295 61.475 15.555 ;
        RECT 61.535 15.295 61.795 15.555 ;
        RECT 62.335 15.295 62.595 15.555 ;
        RECT 62.655 15.295 62.915 15.555 ;
        RECT 63.455 15.295 63.715 15.555 ;
        RECT 63.775 15.295 64.035 15.555 ;
        RECT 64.575 15.295 64.835 15.555 ;
        RECT 64.895 15.295 65.155 15.555 ;
        RECT 65.695 15.295 65.955 15.555 ;
        RECT 66.015 15.295 66.275 15.555 ;
        RECT 66.815 15.295 67.075 15.555 ;
        RECT 67.135 15.295 67.395 15.555 ;
        RECT 67.935 15.295 68.195 15.555 ;
        RECT 68.255 15.295 68.515 15.555 ;
        RECT 69.055 15.295 69.315 15.555 ;
        RECT 69.375 15.295 69.635 15.555 ;
        RECT 72.125 15.295 72.385 15.555 ;
        RECT 72.445 15.295 72.705 15.555 ;
        RECT 73.185 15.295 73.445 15.555 ;
        RECT 73.505 15.295 73.765 15.555 ;
        RECT 74.305 15.295 74.565 15.555 ;
        RECT 74.625 15.295 74.885 15.555 ;
        RECT 75.425 15.295 75.685 15.555 ;
        RECT 75.745 15.295 76.005 15.555 ;
        RECT 76.545 15.295 76.805 15.555 ;
        RECT 76.865 15.295 77.125 15.555 ;
        RECT 77.665 15.295 77.925 15.555 ;
        RECT 77.985 15.295 78.245 15.555 ;
        RECT 78.785 15.295 79.045 15.555 ;
        RECT 79.105 15.295 79.365 15.555 ;
        RECT 79.905 15.295 80.165 15.555 ;
        RECT 80.225 15.295 80.485 15.555 ;
        RECT 81.025 15.295 81.285 15.555 ;
        RECT 81.345 15.295 81.605 15.555 ;
        RECT 82.145 15.295 82.405 15.555 ;
        RECT 82.465 15.295 82.725 15.555 ;
        RECT 85.215 15.275 85.475 15.535 ;
        RECT 85.535 15.275 85.795 15.535 ;
        RECT 86.275 15.275 86.535 15.535 ;
        RECT 86.595 15.275 86.855 15.535 ;
        RECT 87.395 15.275 87.655 15.535 ;
        RECT 87.715 15.275 87.975 15.535 ;
        RECT 88.515 15.275 88.775 15.535 ;
        RECT 88.835 15.275 89.095 15.535 ;
        RECT 89.635 15.275 89.895 15.535 ;
        RECT 89.955 15.275 90.215 15.535 ;
        RECT 90.755 15.275 91.015 15.535 ;
        RECT 91.075 15.275 91.335 15.535 ;
        RECT 91.875 15.275 92.135 15.535 ;
        RECT 92.195 15.275 92.455 15.535 ;
        RECT 92.995 15.275 93.255 15.535 ;
        RECT 93.315 15.275 93.575 15.535 ;
        RECT 94.115 15.275 94.375 15.535 ;
        RECT 94.435 15.275 94.695 15.535 ;
        RECT 95.235 15.275 95.495 15.535 ;
        RECT 95.555 15.275 95.815 15.535 ;
        RECT 98.305 15.275 98.565 15.535 ;
        RECT 98.625 15.275 98.885 15.535 ;
        RECT 99.365 15.275 99.625 15.535 ;
        RECT 99.685 15.275 99.945 15.535 ;
        RECT 100.485 15.275 100.745 15.535 ;
        RECT 100.805 15.275 101.065 15.535 ;
        RECT 101.605 15.275 101.865 15.535 ;
        RECT 101.925 15.275 102.185 15.535 ;
        RECT 102.725 15.275 102.985 15.535 ;
        RECT 103.045 15.275 103.305 15.535 ;
        RECT 103.845 15.275 104.105 15.535 ;
        RECT 104.165 15.275 104.425 15.535 ;
        RECT 104.965 15.275 105.225 15.535 ;
        RECT 105.285 15.275 105.545 15.535 ;
        RECT 106.085 15.275 106.345 15.535 ;
        RECT 106.405 15.275 106.665 15.535 ;
        RECT 107.205 15.275 107.465 15.535 ;
        RECT 107.525 15.275 107.785 15.535 ;
        RECT 108.325 15.275 108.585 15.535 ;
        RECT 108.645 15.275 108.905 15.535 ;
        RECT 111.395 15.275 111.655 15.535 ;
        RECT 111.715 15.275 111.975 15.535 ;
        RECT 112.455 15.275 112.715 15.535 ;
        RECT 112.775 15.275 113.035 15.535 ;
        RECT 113.575 15.275 113.835 15.535 ;
        RECT 113.895 15.275 114.155 15.535 ;
        RECT 114.695 15.275 114.955 15.535 ;
        RECT 115.015 15.275 115.275 15.535 ;
        RECT 115.815 15.275 116.075 15.535 ;
        RECT 116.135 15.275 116.395 15.535 ;
        RECT 116.935 15.275 117.195 15.535 ;
        RECT 117.255 15.275 117.515 15.535 ;
        RECT 118.055 15.275 118.315 15.535 ;
        RECT 118.375 15.275 118.635 15.535 ;
        RECT 119.175 15.275 119.435 15.535 ;
        RECT 119.495 15.275 119.755 15.535 ;
        RECT 120.295 15.275 120.555 15.535 ;
        RECT 120.615 15.275 120.875 15.535 ;
        RECT 121.415 15.275 121.675 15.535 ;
        RECT 121.735 15.275 121.995 15.535 ;
        RECT 124.485 15.275 124.745 15.535 ;
        RECT 124.805 15.275 125.065 15.535 ;
        RECT 125.545 15.275 125.805 15.535 ;
        RECT 125.865 15.275 126.125 15.535 ;
        RECT 126.665 15.275 126.925 15.535 ;
        RECT 126.985 15.275 127.245 15.535 ;
        RECT 127.785 15.275 128.045 15.535 ;
        RECT 128.105 15.275 128.365 15.535 ;
        RECT 128.905 15.275 129.165 15.535 ;
        RECT 129.225 15.275 129.485 15.535 ;
        RECT 130.025 15.275 130.285 15.535 ;
        RECT 130.345 15.275 130.605 15.535 ;
        RECT 131.145 15.275 131.405 15.535 ;
        RECT 131.465 15.275 131.725 15.535 ;
        RECT 132.265 15.275 132.525 15.535 ;
        RECT 132.585 15.275 132.845 15.535 ;
        RECT 133.385 15.275 133.645 15.535 ;
        RECT 133.705 15.275 133.965 15.535 ;
        RECT 134.505 15.275 134.765 15.535 ;
        RECT 134.825 15.275 135.085 15.535 ;
        RECT 137.575 15.255 137.835 15.515 ;
        RECT 137.895 15.255 138.155 15.515 ;
        RECT 138.635 15.255 138.895 15.515 ;
        RECT 138.955 15.255 139.215 15.515 ;
        RECT 139.755 15.255 140.015 15.515 ;
        RECT 140.075 15.255 140.335 15.515 ;
        RECT 140.875 15.255 141.135 15.515 ;
        RECT 141.195 15.255 141.455 15.515 ;
        RECT 141.995 15.255 142.255 15.515 ;
        RECT 142.315 15.255 142.575 15.515 ;
        RECT 143.115 15.255 143.375 15.515 ;
        RECT 143.435 15.255 143.695 15.515 ;
        RECT 144.235 15.255 144.495 15.515 ;
        RECT 144.555 15.255 144.815 15.515 ;
        RECT 145.355 15.255 145.615 15.515 ;
        RECT 145.675 15.255 145.935 15.515 ;
        RECT 146.475 15.255 146.735 15.515 ;
        RECT 146.795 15.255 147.055 15.515 ;
        RECT 147.595 15.255 147.855 15.515 ;
        RECT 147.915 15.255 148.175 15.515 ;
        RECT 150.665 15.255 150.925 15.515 ;
        RECT 150.985 15.255 151.245 15.515 ;
        RECT 151.725 15.255 151.985 15.515 ;
        RECT 152.045 15.255 152.305 15.515 ;
        RECT 152.845 15.255 153.105 15.515 ;
        RECT 153.165 15.255 153.425 15.515 ;
        RECT 153.965 15.255 154.225 15.515 ;
        RECT 154.285 15.255 154.545 15.515 ;
        RECT 155.085 15.255 155.345 15.515 ;
        RECT 155.405 15.255 155.665 15.515 ;
        RECT 156.205 15.255 156.465 15.515 ;
        RECT 156.525 15.255 156.785 15.515 ;
        RECT 157.325 15.255 157.585 15.515 ;
        RECT 157.645 15.255 157.905 15.515 ;
        RECT 158.445 15.255 158.705 15.515 ;
        RECT 158.765 15.255 159.025 15.515 ;
        RECT 159.565 15.255 159.825 15.515 ;
        RECT 159.885 15.255 160.145 15.515 ;
        RECT 160.685 15.255 160.945 15.515 ;
        RECT 161.005 15.255 161.265 15.515 ;
        RECT 6.745 13.265 7.005 13.525 ;
        RECT 7.065 13.265 7.325 13.525 ;
        RECT 7.805 13.265 8.065 13.525 ;
        RECT 8.125 13.265 8.385 13.525 ;
        RECT 8.925 13.265 9.185 13.525 ;
        RECT 9.245 13.265 9.505 13.525 ;
        RECT 10.045 13.265 10.305 13.525 ;
        RECT 10.365 13.265 10.625 13.525 ;
        RECT 11.165 13.265 11.425 13.525 ;
        RECT 11.485 13.265 11.745 13.525 ;
        RECT 12.285 13.265 12.545 13.525 ;
        RECT 12.605 13.265 12.865 13.525 ;
        RECT 13.405 13.265 13.665 13.525 ;
        RECT 13.725 13.265 13.985 13.525 ;
        RECT 14.525 13.265 14.785 13.525 ;
        RECT 14.845 13.265 15.105 13.525 ;
        RECT 15.645 13.265 15.905 13.525 ;
        RECT 15.965 13.265 16.225 13.525 ;
        RECT 16.765 13.265 17.025 13.525 ;
        RECT 17.085 13.265 17.345 13.525 ;
        RECT 19.835 13.265 20.095 13.525 ;
        RECT 20.155 13.265 20.415 13.525 ;
        RECT 20.895 13.265 21.155 13.525 ;
        RECT 21.215 13.265 21.475 13.525 ;
        RECT 22.015 13.265 22.275 13.525 ;
        RECT 22.335 13.265 22.595 13.525 ;
        RECT 23.135 13.265 23.395 13.525 ;
        RECT 23.455 13.265 23.715 13.525 ;
        RECT 24.255 13.265 24.515 13.525 ;
        RECT 24.575 13.265 24.835 13.525 ;
        RECT 25.375 13.265 25.635 13.525 ;
        RECT 25.695 13.265 25.955 13.525 ;
        RECT 26.495 13.265 26.755 13.525 ;
        RECT 26.815 13.265 27.075 13.525 ;
        RECT 27.615 13.265 27.875 13.525 ;
        RECT 27.935 13.265 28.195 13.525 ;
        RECT 28.735 13.265 28.995 13.525 ;
        RECT 29.055 13.265 29.315 13.525 ;
        RECT 29.855 13.265 30.115 13.525 ;
        RECT 30.175 13.265 30.435 13.525 ;
        RECT 32.925 13.285 33.185 13.545 ;
        RECT 33.245 13.285 33.505 13.545 ;
        RECT 33.985 13.285 34.245 13.545 ;
        RECT 34.305 13.285 34.565 13.545 ;
        RECT 35.105 13.285 35.365 13.545 ;
        RECT 35.425 13.285 35.685 13.545 ;
        RECT 36.225 13.285 36.485 13.545 ;
        RECT 36.545 13.285 36.805 13.545 ;
        RECT 37.345 13.285 37.605 13.545 ;
        RECT 37.665 13.285 37.925 13.545 ;
        RECT 38.465 13.285 38.725 13.545 ;
        RECT 38.785 13.285 39.045 13.545 ;
        RECT 39.585 13.285 39.845 13.545 ;
        RECT 39.905 13.285 40.165 13.545 ;
        RECT 40.705 13.285 40.965 13.545 ;
        RECT 41.025 13.285 41.285 13.545 ;
        RECT 41.825 13.285 42.085 13.545 ;
        RECT 42.145 13.285 42.405 13.545 ;
        RECT 42.945 13.285 43.205 13.545 ;
        RECT 43.265 13.285 43.525 13.545 ;
        RECT 46.015 13.285 46.275 13.545 ;
        RECT 46.335 13.285 46.595 13.545 ;
        RECT 47.075 13.285 47.335 13.545 ;
        RECT 47.395 13.285 47.655 13.545 ;
        RECT 48.195 13.285 48.455 13.545 ;
        RECT 48.515 13.285 48.775 13.545 ;
        RECT 49.315 13.285 49.575 13.545 ;
        RECT 49.635 13.285 49.895 13.545 ;
        RECT 50.435 13.285 50.695 13.545 ;
        RECT 50.755 13.285 51.015 13.545 ;
        RECT 51.555 13.285 51.815 13.545 ;
        RECT 51.875 13.285 52.135 13.545 ;
        RECT 52.675 13.285 52.935 13.545 ;
        RECT 52.995 13.285 53.255 13.545 ;
        RECT 53.795 13.285 54.055 13.545 ;
        RECT 54.115 13.285 54.375 13.545 ;
        RECT 54.915 13.285 55.175 13.545 ;
        RECT 55.235 13.285 55.495 13.545 ;
        RECT 56.035 13.285 56.295 13.545 ;
        RECT 56.355 13.285 56.615 13.545 ;
        RECT 59.065 13.285 59.325 13.545 ;
        RECT 59.385 13.285 59.645 13.545 ;
        RECT 60.125 13.285 60.385 13.545 ;
        RECT 60.445 13.285 60.705 13.545 ;
        RECT 61.245 13.285 61.505 13.545 ;
        RECT 61.565 13.285 61.825 13.545 ;
        RECT 62.365 13.285 62.625 13.545 ;
        RECT 62.685 13.285 62.945 13.545 ;
        RECT 63.485 13.285 63.745 13.545 ;
        RECT 63.805 13.285 64.065 13.545 ;
        RECT 64.605 13.285 64.865 13.545 ;
        RECT 64.925 13.285 65.185 13.545 ;
        RECT 65.725 13.285 65.985 13.545 ;
        RECT 66.045 13.285 66.305 13.545 ;
        RECT 66.845 13.285 67.105 13.545 ;
        RECT 67.165 13.285 67.425 13.545 ;
        RECT 67.965 13.285 68.225 13.545 ;
        RECT 68.285 13.285 68.545 13.545 ;
        RECT 69.085 13.285 69.345 13.545 ;
        RECT 69.405 13.285 69.665 13.545 ;
        RECT 72.155 13.285 72.415 13.545 ;
        RECT 72.475 13.285 72.735 13.545 ;
        RECT 73.215 13.285 73.475 13.545 ;
        RECT 73.535 13.285 73.795 13.545 ;
        RECT 74.335 13.285 74.595 13.545 ;
        RECT 74.655 13.285 74.915 13.545 ;
        RECT 75.455 13.285 75.715 13.545 ;
        RECT 75.775 13.285 76.035 13.545 ;
        RECT 76.575 13.285 76.835 13.545 ;
        RECT 76.895 13.285 77.155 13.545 ;
        RECT 77.695 13.285 77.955 13.545 ;
        RECT 78.015 13.285 78.275 13.545 ;
        RECT 78.815 13.285 79.075 13.545 ;
        RECT 79.135 13.285 79.395 13.545 ;
        RECT 79.935 13.285 80.195 13.545 ;
        RECT 80.255 13.285 80.515 13.545 ;
        RECT 81.055 13.285 81.315 13.545 ;
        RECT 81.375 13.285 81.635 13.545 ;
        RECT 82.175 13.285 82.435 13.545 ;
        RECT 82.495 13.285 82.755 13.545 ;
        RECT 85.245 13.305 85.505 13.565 ;
        RECT 85.565 13.305 85.825 13.565 ;
        RECT 86.305 13.305 86.565 13.565 ;
        RECT 86.625 13.305 86.885 13.565 ;
        RECT 87.425 13.305 87.685 13.565 ;
        RECT 87.745 13.305 88.005 13.565 ;
        RECT 88.545 13.305 88.805 13.565 ;
        RECT 88.865 13.305 89.125 13.565 ;
        RECT 89.665 13.305 89.925 13.565 ;
        RECT 89.985 13.305 90.245 13.565 ;
        RECT 90.785 13.305 91.045 13.565 ;
        RECT 91.105 13.305 91.365 13.565 ;
        RECT 91.905 13.305 92.165 13.565 ;
        RECT 92.225 13.305 92.485 13.565 ;
        RECT 93.025 13.305 93.285 13.565 ;
        RECT 93.345 13.305 93.605 13.565 ;
        RECT 94.145 13.305 94.405 13.565 ;
        RECT 94.465 13.305 94.725 13.565 ;
        RECT 95.265 13.305 95.525 13.565 ;
        RECT 95.585 13.305 95.845 13.565 ;
        RECT 98.335 13.305 98.595 13.565 ;
        RECT 98.655 13.305 98.915 13.565 ;
        RECT 99.395 13.305 99.655 13.565 ;
        RECT 99.715 13.305 99.975 13.565 ;
        RECT 100.515 13.305 100.775 13.565 ;
        RECT 100.835 13.305 101.095 13.565 ;
        RECT 101.635 13.305 101.895 13.565 ;
        RECT 101.955 13.305 102.215 13.565 ;
        RECT 102.755 13.305 103.015 13.565 ;
        RECT 103.075 13.305 103.335 13.565 ;
        RECT 103.875 13.305 104.135 13.565 ;
        RECT 104.195 13.305 104.455 13.565 ;
        RECT 104.995 13.305 105.255 13.565 ;
        RECT 105.315 13.305 105.575 13.565 ;
        RECT 106.115 13.305 106.375 13.565 ;
        RECT 106.435 13.305 106.695 13.565 ;
        RECT 107.235 13.305 107.495 13.565 ;
        RECT 107.555 13.305 107.815 13.565 ;
        RECT 108.355 13.305 108.615 13.565 ;
        RECT 108.675 13.305 108.935 13.565 ;
        RECT 111.425 13.305 111.685 13.565 ;
        RECT 111.745 13.305 112.005 13.565 ;
        RECT 112.485 13.305 112.745 13.565 ;
        RECT 112.805 13.305 113.065 13.565 ;
        RECT 113.605 13.305 113.865 13.565 ;
        RECT 113.925 13.305 114.185 13.565 ;
        RECT 114.725 13.305 114.985 13.565 ;
        RECT 115.045 13.305 115.305 13.565 ;
        RECT 115.845 13.305 116.105 13.565 ;
        RECT 116.165 13.305 116.425 13.565 ;
        RECT 116.965 13.305 117.225 13.565 ;
        RECT 117.285 13.305 117.545 13.565 ;
        RECT 118.085 13.305 118.345 13.565 ;
        RECT 118.405 13.305 118.665 13.565 ;
        RECT 119.205 13.305 119.465 13.565 ;
        RECT 119.525 13.305 119.785 13.565 ;
        RECT 120.325 13.305 120.585 13.565 ;
        RECT 120.645 13.305 120.905 13.565 ;
        RECT 121.445 13.305 121.705 13.565 ;
        RECT 121.765 13.305 122.025 13.565 ;
        RECT 124.515 13.305 124.775 13.565 ;
        RECT 124.835 13.305 125.095 13.565 ;
        RECT 125.575 13.305 125.835 13.565 ;
        RECT 125.895 13.305 126.155 13.565 ;
        RECT 126.695 13.305 126.955 13.565 ;
        RECT 127.015 13.305 127.275 13.565 ;
        RECT 127.815 13.305 128.075 13.565 ;
        RECT 128.135 13.305 128.395 13.565 ;
        RECT 128.935 13.305 129.195 13.565 ;
        RECT 129.255 13.305 129.515 13.565 ;
        RECT 130.055 13.305 130.315 13.565 ;
        RECT 130.375 13.305 130.635 13.565 ;
        RECT 131.175 13.305 131.435 13.565 ;
        RECT 131.495 13.305 131.755 13.565 ;
        RECT 132.295 13.305 132.555 13.565 ;
        RECT 132.615 13.305 132.875 13.565 ;
        RECT 133.415 13.305 133.675 13.565 ;
        RECT 133.735 13.305 133.995 13.565 ;
        RECT 134.535 13.305 134.795 13.565 ;
        RECT 134.855 13.305 135.115 13.565 ;
        RECT 137.605 13.325 137.865 13.585 ;
        RECT 137.925 13.325 138.185 13.585 ;
        RECT 138.665 13.325 138.925 13.585 ;
        RECT 138.985 13.325 139.245 13.585 ;
        RECT 139.785 13.325 140.045 13.585 ;
        RECT 140.105 13.325 140.365 13.585 ;
        RECT 140.905 13.325 141.165 13.585 ;
        RECT 141.225 13.325 141.485 13.585 ;
        RECT 142.025 13.325 142.285 13.585 ;
        RECT 142.345 13.325 142.605 13.585 ;
        RECT 143.145 13.325 143.405 13.585 ;
        RECT 143.465 13.325 143.725 13.585 ;
        RECT 144.265 13.325 144.525 13.585 ;
        RECT 144.585 13.325 144.845 13.585 ;
        RECT 145.385 13.325 145.645 13.585 ;
        RECT 145.705 13.325 145.965 13.585 ;
        RECT 146.505 13.325 146.765 13.585 ;
        RECT 146.825 13.325 147.085 13.585 ;
        RECT 147.625 13.325 147.885 13.585 ;
        RECT 147.945 13.325 148.205 13.585 ;
        RECT 150.695 13.325 150.955 13.585 ;
        RECT 151.015 13.325 151.275 13.585 ;
        RECT 151.755 13.325 152.015 13.585 ;
        RECT 152.075 13.325 152.335 13.585 ;
        RECT 152.875 13.325 153.135 13.585 ;
        RECT 153.195 13.325 153.455 13.585 ;
        RECT 153.995 13.325 154.255 13.585 ;
        RECT 154.315 13.325 154.575 13.585 ;
        RECT 155.115 13.325 155.375 13.585 ;
        RECT 155.435 13.325 155.695 13.585 ;
        RECT 156.235 13.325 156.495 13.585 ;
        RECT 156.555 13.325 156.815 13.585 ;
        RECT 157.355 13.325 157.615 13.585 ;
        RECT 157.675 13.325 157.935 13.585 ;
        RECT 158.475 13.325 158.735 13.585 ;
        RECT 158.795 13.325 159.055 13.585 ;
        RECT 159.595 13.325 159.855 13.585 ;
        RECT 159.915 13.325 160.175 13.585 ;
        RECT 160.715 13.325 160.975 13.585 ;
        RECT 161.035 13.325 161.295 13.585 ;
      LAYER met2 ;
        RECT 6.155 107.250 6.295 118.610 ;
        RECT 6.715 107.250 6.855 118.140 ;
        RECT 6.155 106.920 6.855 107.250 ;
        RECT 7.275 107.250 7.415 118.610 ;
        RECT 7.835 107.250 7.975 118.140 ;
        RECT 7.275 106.920 7.975 107.250 ;
        RECT 8.395 107.250 8.535 118.610 ;
        RECT 8.955 107.250 9.095 118.140 ;
        RECT 8.395 106.920 9.095 107.250 ;
        RECT 9.515 107.250 9.655 118.610 ;
        RECT 10.075 107.250 10.215 118.140 ;
        RECT 9.515 106.920 10.215 107.250 ;
        RECT 10.635 107.250 10.775 118.610 ;
        RECT 11.195 107.250 11.335 118.140 ;
        RECT 10.635 106.920 11.335 107.250 ;
        RECT 11.755 107.250 11.895 118.610 ;
        RECT 12.315 107.250 12.455 118.140 ;
        RECT 11.755 106.920 12.455 107.250 ;
        RECT 12.875 107.250 13.015 118.610 ;
        RECT 13.435 107.250 13.575 118.140 ;
        RECT 12.875 106.920 13.575 107.250 ;
        RECT 13.995 107.250 14.135 118.610 ;
        RECT 14.555 107.250 14.695 118.140 ;
        RECT 13.995 106.920 14.695 107.250 ;
        RECT 15.115 107.250 15.255 118.610 ;
        RECT 15.675 107.250 15.815 118.140 ;
        RECT 15.115 106.920 15.815 107.250 ;
        RECT 16.235 107.250 16.375 118.140 ;
        RECT 16.795 107.250 16.935 118.140 ;
        RECT 17.355 107.250 17.565 118.140 ;
        RECT 16.235 106.920 17.565 107.250 ;
        RECT 19.245 107.250 19.385 118.610 ;
        RECT 19.805 107.250 19.945 118.140 ;
        RECT 19.245 106.920 19.945 107.250 ;
        RECT 20.365 107.250 20.505 118.610 ;
        RECT 20.925 107.250 21.065 118.140 ;
        RECT 20.365 106.920 21.065 107.250 ;
        RECT 21.485 107.250 21.625 118.610 ;
        RECT 22.045 107.250 22.185 118.140 ;
        RECT 21.485 106.920 22.185 107.250 ;
        RECT 22.605 107.250 22.745 118.610 ;
        RECT 23.165 107.250 23.305 118.140 ;
        RECT 22.605 106.920 23.305 107.250 ;
        RECT 23.725 107.250 23.865 118.610 ;
        RECT 24.285 107.250 24.425 118.140 ;
        RECT 23.725 106.920 24.425 107.250 ;
        RECT 24.845 107.250 24.985 118.610 ;
        RECT 25.405 107.250 25.545 118.140 ;
        RECT 24.845 106.920 25.545 107.250 ;
        RECT 25.965 107.250 26.105 118.610 ;
        RECT 26.525 107.250 26.665 118.140 ;
        RECT 25.965 106.920 26.665 107.250 ;
        RECT 27.085 107.250 27.225 118.610 ;
        RECT 27.645 107.250 27.785 118.140 ;
        RECT 27.085 106.920 27.785 107.250 ;
        RECT 28.205 107.250 28.345 118.610 ;
        RECT 28.765 107.250 28.905 118.140 ;
        RECT 28.205 106.920 28.905 107.250 ;
        RECT 29.325 107.250 29.465 118.140 ;
        RECT 29.885 107.250 30.025 118.140 ;
        RECT 30.445 107.250 30.655 118.140 ;
        RECT 29.325 106.920 30.655 107.250 ;
        RECT 32.335 107.230 32.475 118.590 ;
        RECT 32.895 107.230 33.035 118.120 ;
        RECT 32.335 106.900 33.035 107.230 ;
        RECT 33.455 107.230 33.595 118.590 ;
        RECT 34.015 107.230 34.155 118.120 ;
        RECT 33.455 106.900 34.155 107.230 ;
        RECT 34.575 107.230 34.715 118.590 ;
        RECT 35.135 107.230 35.275 118.120 ;
        RECT 34.575 106.900 35.275 107.230 ;
        RECT 35.695 107.230 35.835 118.590 ;
        RECT 36.255 107.230 36.395 118.120 ;
        RECT 35.695 106.900 36.395 107.230 ;
        RECT 36.815 107.230 36.955 118.590 ;
        RECT 37.375 107.230 37.515 118.120 ;
        RECT 36.815 106.900 37.515 107.230 ;
        RECT 37.935 107.230 38.075 118.590 ;
        RECT 38.495 107.230 38.635 118.120 ;
        RECT 37.935 106.900 38.635 107.230 ;
        RECT 39.055 107.230 39.195 118.590 ;
        RECT 39.615 107.230 39.755 118.120 ;
        RECT 39.055 106.900 39.755 107.230 ;
        RECT 40.175 107.230 40.315 118.590 ;
        RECT 40.735 107.230 40.875 118.120 ;
        RECT 40.175 106.900 40.875 107.230 ;
        RECT 41.295 107.230 41.435 118.590 ;
        RECT 41.855 107.230 41.995 118.120 ;
        RECT 41.295 106.900 41.995 107.230 ;
        RECT 42.415 107.230 42.555 118.120 ;
        RECT 42.975 107.230 43.115 118.120 ;
        RECT 43.535 107.230 43.745 118.120 ;
        RECT 42.415 106.900 43.745 107.230 ;
        RECT 45.425 107.230 45.565 118.590 ;
        RECT 45.985 107.230 46.125 118.120 ;
        RECT 45.425 106.900 46.125 107.230 ;
        RECT 46.545 107.230 46.685 118.590 ;
        RECT 47.105 107.230 47.245 118.120 ;
        RECT 46.545 106.900 47.245 107.230 ;
        RECT 47.665 107.230 47.805 118.590 ;
        RECT 48.225 107.230 48.365 118.120 ;
        RECT 47.665 106.900 48.365 107.230 ;
        RECT 48.785 107.230 48.925 118.590 ;
        RECT 49.345 107.230 49.485 118.120 ;
        RECT 48.785 106.900 49.485 107.230 ;
        RECT 49.905 107.230 50.045 118.590 ;
        RECT 50.465 107.230 50.605 118.120 ;
        RECT 49.905 106.900 50.605 107.230 ;
        RECT 51.025 107.230 51.165 118.590 ;
        RECT 51.585 107.230 51.725 118.120 ;
        RECT 51.025 106.900 51.725 107.230 ;
        RECT 52.145 107.230 52.285 118.590 ;
        RECT 52.705 107.230 52.845 118.120 ;
        RECT 52.145 106.900 52.845 107.230 ;
        RECT 53.265 107.230 53.405 118.590 ;
        RECT 53.825 107.230 53.965 118.120 ;
        RECT 53.265 106.900 53.965 107.230 ;
        RECT 54.385 107.230 54.525 118.590 ;
        RECT 54.945 107.230 55.085 118.120 ;
        RECT 54.385 106.900 55.085 107.230 ;
        RECT 55.505 107.230 55.645 118.120 ;
        RECT 56.065 107.230 56.205 118.120 ;
        RECT 56.625 107.230 56.835 118.120 ;
        RECT 55.505 106.900 56.835 107.230 ;
        RECT 58.475 107.230 58.615 118.590 ;
        RECT 59.035 107.230 59.175 118.120 ;
        RECT 58.475 106.900 59.175 107.230 ;
        RECT 59.595 107.230 59.735 118.590 ;
        RECT 60.155 107.230 60.295 118.120 ;
        RECT 59.595 106.900 60.295 107.230 ;
        RECT 60.715 107.230 60.855 118.590 ;
        RECT 61.275 107.230 61.415 118.120 ;
        RECT 60.715 106.900 61.415 107.230 ;
        RECT 61.835 107.230 61.975 118.590 ;
        RECT 62.395 107.230 62.535 118.120 ;
        RECT 61.835 106.900 62.535 107.230 ;
        RECT 62.955 107.230 63.095 118.590 ;
        RECT 63.515 107.230 63.655 118.120 ;
        RECT 62.955 106.900 63.655 107.230 ;
        RECT 64.075 107.230 64.215 118.590 ;
        RECT 64.635 107.230 64.775 118.120 ;
        RECT 64.075 106.900 64.775 107.230 ;
        RECT 65.195 107.230 65.335 118.590 ;
        RECT 65.755 107.230 65.895 118.120 ;
        RECT 65.195 106.900 65.895 107.230 ;
        RECT 66.315 107.230 66.455 118.590 ;
        RECT 66.875 107.230 67.015 118.120 ;
        RECT 66.315 106.900 67.015 107.230 ;
        RECT 67.435 107.230 67.575 118.590 ;
        RECT 67.995 107.230 68.135 118.120 ;
        RECT 67.435 106.900 68.135 107.230 ;
        RECT 68.555 107.230 68.695 118.120 ;
        RECT 69.115 107.230 69.255 118.120 ;
        RECT 69.675 107.230 69.885 118.120 ;
        RECT 68.555 106.900 69.885 107.230 ;
        RECT 71.565 107.230 71.705 118.590 ;
        RECT 72.125 107.230 72.265 118.120 ;
        RECT 71.565 106.900 72.265 107.230 ;
        RECT 72.685 107.230 72.825 118.590 ;
        RECT 73.245 107.230 73.385 118.120 ;
        RECT 72.685 106.900 73.385 107.230 ;
        RECT 73.805 107.230 73.945 118.590 ;
        RECT 74.365 107.230 74.505 118.120 ;
        RECT 73.805 106.900 74.505 107.230 ;
        RECT 74.925 107.230 75.065 118.590 ;
        RECT 75.485 107.230 75.625 118.120 ;
        RECT 74.925 106.900 75.625 107.230 ;
        RECT 76.045 107.230 76.185 118.590 ;
        RECT 76.605 107.230 76.745 118.120 ;
        RECT 76.045 106.900 76.745 107.230 ;
        RECT 77.165 107.230 77.305 118.590 ;
        RECT 77.725 107.230 77.865 118.120 ;
        RECT 77.165 106.900 77.865 107.230 ;
        RECT 78.285 107.230 78.425 118.590 ;
        RECT 78.845 107.230 78.985 118.120 ;
        RECT 78.285 106.900 78.985 107.230 ;
        RECT 79.405 107.230 79.545 118.590 ;
        RECT 79.965 107.230 80.105 118.120 ;
        RECT 79.405 106.900 80.105 107.230 ;
        RECT 80.525 107.230 80.665 118.590 ;
        RECT 81.085 107.230 81.225 118.120 ;
        RECT 80.525 106.900 81.225 107.230 ;
        RECT 81.645 107.230 81.785 118.120 ;
        RECT 82.205 107.230 82.345 118.120 ;
        RECT 82.765 107.230 82.975 118.120 ;
        RECT 81.645 106.900 82.975 107.230 ;
        RECT 84.655 107.210 84.795 118.570 ;
        RECT 85.215 107.210 85.355 118.100 ;
        RECT 84.655 106.880 85.355 107.210 ;
        RECT 85.775 107.210 85.915 118.570 ;
        RECT 86.335 107.210 86.475 118.100 ;
        RECT 85.775 106.880 86.475 107.210 ;
        RECT 86.895 107.210 87.035 118.570 ;
        RECT 87.455 107.210 87.595 118.100 ;
        RECT 86.895 106.880 87.595 107.210 ;
        RECT 88.015 107.210 88.155 118.570 ;
        RECT 88.575 107.210 88.715 118.100 ;
        RECT 88.015 106.880 88.715 107.210 ;
        RECT 89.135 107.210 89.275 118.570 ;
        RECT 89.695 107.210 89.835 118.100 ;
        RECT 89.135 106.880 89.835 107.210 ;
        RECT 90.255 107.210 90.395 118.570 ;
        RECT 90.815 107.210 90.955 118.100 ;
        RECT 90.255 106.880 90.955 107.210 ;
        RECT 91.375 107.210 91.515 118.570 ;
        RECT 91.935 107.210 92.075 118.100 ;
        RECT 91.375 106.880 92.075 107.210 ;
        RECT 92.495 107.210 92.635 118.570 ;
        RECT 93.055 107.210 93.195 118.100 ;
        RECT 92.495 106.880 93.195 107.210 ;
        RECT 93.615 107.210 93.755 118.570 ;
        RECT 94.175 107.210 94.315 118.100 ;
        RECT 93.615 106.880 94.315 107.210 ;
        RECT 94.735 107.210 94.875 118.100 ;
        RECT 95.295 107.210 95.435 118.100 ;
        RECT 95.855 107.210 96.065 118.100 ;
        RECT 94.735 106.880 96.065 107.210 ;
        RECT 97.745 107.210 97.885 118.570 ;
        RECT 98.305 107.210 98.445 118.100 ;
        RECT 97.745 106.880 98.445 107.210 ;
        RECT 98.865 107.210 99.005 118.570 ;
        RECT 99.425 107.210 99.565 118.100 ;
        RECT 98.865 106.880 99.565 107.210 ;
        RECT 99.985 107.210 100.125 118.570 ;
        RECT 100.545 107.210 100.685 118.100 ;
        RECT 99.985 106.880 100.685 107.210 ;
        RECT 101.105 107.210 101.245 118.570 ;
        RECT 101.665 107.210 101.805 118.100 ;
        RECT 101.105 106.880 101.805 107.210 ;
        RECT 102.225 107.210 102.365 118.570 ;
        RECT 102.785 107.210 102.925 118.100 ;
        RECT 102.225 106.880 102.925 107.210 ;
        RECT 103.345 107.210 103.485 118.570 ;
        RECT 103.905 107.210 104.045 118.100 ;
        RECT 103.345 106.880 104.045 107.210 ;
        RECT 104.465 107.210 104.605 118.570 ;
        RECT 105.025 107.210 105.165 118.100 ;
        RECT 104.465 106.880 105.165 107.210 ;
        RECT 105.585 107.210 105.725 118.570 ;
        RECT 106.145 107.210 106.285 118.100 ;
        RECT 105.585 106.880 106.285 107.210 ;
        RECT 106.705 107.210 106.845 118.570 ;
        RECT 107.265 107.210 107.405 118.100 ;
        RECT 106.705 106.880 107.405 107.210 ;
        RECT 107.825 107.210 107.965 118.100 ;
        RECT 108.385 107.210 108.525 118.100 ;
        RECT 108.945 107.210 109.155 118.100 ;
        RECT 107.825 106.880 109.155 107.210 ;
        RECT 110.835 107.210 110.975 118.570 ;
        RECT 111.395 107.210 111.535 118.100 ;
        RECT 110.835 106.880 111.535 107.210 ;
        RECT 111.955 107.210 112.095 118.570 ;
        RECT 112.515 107.210 112.655 118.100 ;
        RECT 111.955 106.880 112.655 107.210 ;
        RECT 113.075 107.210 113.215 118.570 ;
        RECT 113.635 107.210 113.775 118.100 ;
        RECT 113.075 106.880 113.775 107.210 ;
        RECT 114.195 107.210 114.335 118.570 ;
        RECT 114.755 107.210 114.895 118.100 ;
        RECT 114.195 106.880 114.895 107.210 ;
        RECT 115.315 107.210 115.455 118.570 ;
        RECT 115.875 107.210 116.015 118.100 ;
        RECT 115.315 106.880 116.015 107.210 ;
        RECT 116.435 107.210 116.575 118.570 ;
        RECT 116.995 107.210 117.135 118.100 ;
        RECT 116.435 106.880 117.135 107.210 ;
        RECT 117.555 107.210 117.695 118.570 ;
        RECT 118.115 107.210 118.255 118.100 ;
        RECT 117.555 106.880 118.255 107.210 ;
        RECT 118.675 107.210 118.815 118.570 ;
        RECT 119.235 107.210 119.375 118.100 ;
        RECT 118.675 106.880 119.375 107.210 ;
        RECT 119.795 107.210 119.935 118.570 ;
        RECT 120.355 107.210 120.495 118.100 ;
        RECT 119.795 106.880 120.495 107.210 ;
        RECT 120.915 107.210 121.055 118.100 ;
        RECT 121.475 107.210 121.615 118.100 ;
        RECT 122.035 107.210 122.245 118.100 ;
        RECT 120.915 106.880 122.245 107.210 ;
        RECT 123.925 107.210 124.065 118.570 ;
        RECT 124.485 107.210 124.625 118.100 ;
        RECT 123.925 106.880 124.625 107.210 ;
        RECT 125.045 107.210 125.185 118.570 ;
        RECT 125.605 107.210 125.745 118.100 ;
        RECT 125.045 106.880 125.745 107.210 ;
        RECT 126.165 107.210 126.305 118.570 ;
        RECT 126.725 107.210 126.865 118.100 ;
        RECT 126.165 106.880 126.865 107.210 ;
        RECT 127.285 107.210 127.425 118.570 ;
        RECT 127.845 107.210 127.985 118.100 ;
        RECT 127.285 106.880 127.985 107.210 ;
        RECT 128.405 107.210 128.545 118.570 ;
        RECT 128.965 107.210 129.105 118.100 ;
        RECT 128.405 106.880 129.105 107.210 ;
        RECT 129.525 107.210 129.665 118.570 ;
        RECT 130.085 107.210 130.225 118.100 ;
        RECT 129.525 106.880 130.225 107.210 ;
        RECT 130.645 107.210 130.785 118.570 ;
        RECT 131.205 107.210 131.345 118.100 ;
        RECT 130.645 106.880 131.345 107.210 ;
        RECT 131.765 107.210 131.905 118.570 ;
        RECT 132.325 107.210 132.465 118.100 ;
        RECT 131.765 106.880 132.465 107.210 ;
        RECT 132.885 107.210 133.025 118.570 ;
        RECT 133.445 107.210 133.585 118.100 ;
        RECT 132.885 106.880 133.585 107.210 ;
        RECT 134.005 107.210 134.145 118.100 ;
        RECT 134.565 107.210 134.705 118.100 ;
        RECT 135.125 107.210 135.335 118.100 ;
        RECT 134.005 106.880 135.335 107.210 ;
        RECT 137.015 107.190 137.155 118.550 ;
        RECT 137.575 107.190 137.715 118.080 ;
        RECT 137.015 106.860 137.715 107.190 ;
        RECT 138.135 107.190 138.275 118.550 ;
        RECT 138.695 107.190 138.835 118.080 ;
        RECT 138.135 106.860 138.835 107.190 ;
        RECT 139.255 107.190 139.395 118.550 ;
        RECT 139.815 107.190 139.955 118.080 ;
        RECT 139.255 106.860 139.955 107.190 ;
        RECT 140.375 107.190 140.515 118.550 ;
        RECT 140.935 107.190 141.075 118.080 ;
        RECT 140.375 106.860 141.075 107.190 ;
        RECT 141.495 107.190 141.635 118.550 ;
        RECT 142.055 107.190 142.195 118.080 ;
        RECT 141.495 106.860 142.195 107.190 ;
        RECT 142.615 107.190 142.755 118.550 ;
        RECT 143.175 107.190 143.315 118.080 ;
        RECT 142.615 106.860 143.315 107.190 ;
        RECT 143.735 107.190 143.875 118.550 ;
        RECT 144.295 107.190 144.435 118.080 ;
        RECT 143.735 106.860 144.435 107.190 ;
        RECT 144.855 107.190 144.995 118.550 ;
        RECT 145.415 107.190 145.555 118.080 ;
        RECT 144.855 106.860 145.555 107.190 ;
        RECT 145.975 107.190 146.115 118.550 ;
        RECT 146.535 107.190 146.675 118.080 ;
        RECT 145.975 106.860 146.675 107.190 ;
        RECT 147.095 107.190 147.235 118.080 ;
        RECT 147.655 107.190 147.795 118.080 ;
        RECT 148.215 107.190 148.425 118.080 ;
        RECT 147.095 106.860 148.425 107.190 ;
        RECT 150.105 107.190 150.245 118.550 ;
        RECT 150.665 107.190 150.805 118.080 ;
        RECT 150.105 106.860 150.805 107.190 ;
        RECT 151.225 107.190 151.365 118.550 ;
        RECT 151.785 107.190 151.925 118.080 ;
        RECT 151.225 106.860 151.925 107.190 ;
        RECT 152.345 107.190 152.485 118.550 ;
        RECT 152.905 107.190 153.045 118.080 ;
        RECT 152.345 106.860 153.045 107.190 ;
        RECT 153.465 107.190 153.605 118.550 ;
        RECT 154.025 107.190 154.165 118.080 ;
        RECT 153.465 106.860 154.165 107.190 ;
        RECT 154.585 107.190 154.725 118.550 ;
        RECT 155.145 107.190 155.285 118.080 ;
        RECT 154.585 106.860 155.285 107.190 ;
        RECT 155.705 107.190 155.845 118.550 ;
        RECT 156.265 107.190 156.405 118.080 ;
        RECT 155.705 106.860 156.405 107.190 ;
        RECT 156.825 107.190 156.965 118.550 ;
        RECT 157.385 107.190 157.525 118.080 ;
        RECT 156.825 106.860 157.525 107.190 ;
        RECT 157.945 107.190 158.085 118.550 ;
        RECT 158.505 107.190 158.645 118.080 ;
        RECT 157.945 106.860 158.645 107.190 ;
        RECT 159.065 107.190 159.205 118.550 ;
        RECT 159.625 107.190 159.765 118.080 ;
        RECT 159.065 106.860 159.765 107.190 ;
        RECT 160.185 107.190 160.325 118.080 ;
        RECT 160.745 107.190 160.885 118.080 ;
        RECT 161.305 107.190 161.515 118.080 ;
        RECT 160.185 106.860 161.515 107.190 ;
        RECT 6.185 104.870 6.885 105.200 ;
        RECT 6.185 93.510 6.325 104.870 ;
        RECT 6.745 93.980 6.885 104.870 ;
        RECT 7.305 104.870 8.005 105.200 ;
        RECT 7.305 93.510 7.445 104.870 ;
        RECT 7.865 93.980 8.005 104.870 ;
        RECT 8.425 104.870 9.125 105.200 ;
        RECT 8.425 93.510 8.565 104.870 ;
        RECT 8.985 93.980 9.125 104.870 ;
        RECT 9.545 104.870 10.245 105.200 ;
        RECT 9.545 93.510 9.685 104.870 ;
        RECT 10.105 93.980 10.245 104.870 ;
        RECT 10.665 104.870 11.365 105.200 ;
        RECT 10.665 93.510 10.805 104.870 ;
        RECT 11.225 93.980 11.365 104.870 ;
        RECT 11.785 104.870 12.485 105.200 ;
        RECT 11.785 93.510 11.925 104.870 ;
        RECT 12.345 93.980 12.485 104.870 ;
        RECT 12.905 104.870 13.605 105.200 ;
        RECT 12.905 93.510 13.045 104.870 ;
        RECT 13.465 93.980 13.605 104.870 ;
        RECT 14.025 104.870 14.725 105.200 ;
        RECT 14.025 93.510 14.165 104.870 ;
        RECT 14.585 93.980 14.725 104.870 ;
        RECT 15.145 104.870 15.845 105.200 ;
        RECT 15.145 93.510 15.285 104.870 ;
        RECT 15.705 93.980 15.845 104.870 ;
        RECT 16.265 104.870 17.595 105.200 ;
        RECT 16.265 93.980 16.405 104.870 ;
        RECT 16.825 93.980 16.965 104.870 ;
        RECT 17.385 93.980 17.595 104.870 ;
        RECT 19.275 104.870 19.975 105.200 ;
        RECT 19.275 93.510 19.415 104.870 ;
        RECT 19.835 93.980 19.975 104.870 ;
        RECT 20.395 104.870 21.095 105.200 ;
        RECT 20.395 93.510 20.535 104.870 ;
        RECT 20.955 93.980 21.095 104.870 ;
        RECT 21.515 104.870 22.215 105.200 ;
        RECT 21.515 93.510 21.655 104.870 ;
        RECT 22.075 93.980 22.215 104.870 ;
        RECT 22.635 104.870 23.335 105.200 ;
        RECT 22.635 93.510 22.775 104.870 ;
        RECT 23.195 93.980 23.335 104.870 ;
        RECT 23.755 104.870 24.455 105.200 ;
        RECT 23.755 93.510 23.895 104.870 ;
        RECT 24.315 93.980 24.455 104.870 ;
        RECT 24.875 104.870 25.575 105.200 ;
        RECT 24.875 93.510 25.015 104.870 ;
        RECT 25.435 93.980 25.575 104.870 ;
        RECT 25.995 104.870 26.695 105.200 ;
        RECT 25.995 93.510 26.135 104.870 ;
        RECT 26.555 93.980 26.695 104.870 ;
        RECT 27.115 104.870 27.815 105.200 ;
        RECT 27.115 93.510 27.255 104.870 ;
        RECT 27.675 93.980 27.815 104.870 ;
        RECT 28.235 104.870 28.935 105.200 ;
        RECT 28.235 93.510 28.375 104.870 ;
        RECT 28.795 93.980 28.935 104.870 ;
        RECT 29.355 104.870 30.685 105.200 ;
        RECT 29.355 93.980 29.495 104.870 ;
        RECT 29.915 93.980 30.055 104.870 ;
        RECT 30.475 93.980 30.685 104.870 ;
        RECT 32.365 104.890 33.065 105.220 ;
        RECT 32.365 93.530 32.505 104.890 ;
        RECT 32.925 94.000 33.065 104.890 ;
        RECT 33.485 104.890 34.185 105.220 ;
        RECT 33.485 93.530 33.625 104.890 ;
        RECT 34.045 94.000 34.185 104.890 ;
        RECT 34.605 104.890 35.305 105.220 ;
        RECT 34.605 93.530 34.745 104.890 ;
        RECT 35.165 94.000 35.305 104.890 ;
        RECT 35.725 104.890 36.425 105.220 ;
        RECT 35.725 93.530 35.865 104.890 ;
        RECT 36.285 94.000 36.425 104.890 ;
        RECT 36.845 104.890 37.545 105.220 ;
        RECT 36.845 93.530 36.985 104.890 ;
        RECT 37.405 94.000 37.545 104.890 ;
        RECT 37.965 104.890 38.665 105.220 ;
        RECT 37.965 93.530 38.105 104.890 ;
        RECT 38.525 94.000 38.665 104.890 ;
        RECT 39.085 104.890 39.785 105.220 ;
        RECT 39.085 93.530 39.225 104.890 ;
        RECT 39.645 94.000 39.785 104.890 ;
        RECT 40.205 104.890 40.905 105.220 ;
        RECT 40.205 93.530 40.345 104.890 ;
        RECT 40.765 94.000 40.905 104.890 ;
        RECT 41.325 104.890 42.025 105.220 ;
        RECT 41.325 93.530 41.465 104.890 ;
        RECT 41.885 94.000 42.025 104.890 ;
        RECT 42.445 104.890 43.775 105.220 ;
        RECT 42.445 94.000 42.585 104.890 ;
        RECT 43.005 94.000 43.145 104.890 ;
        RECT 43.565 94.000 43.775 104.890 ;
        RECT 45.455 104.890 46.155 105.220 ;
        RECT 45.455 93.530 45.595 104.890 ;
        RECT 46.015 94.000 46.155 104.890 ;
        RECT 46.575 104.890 47.275 105.220 ;
        RECT 46.575 93.530 46.715 104.890 ;
        RECT 47.135 94.000 47.275 104.890 ;
        RECT 47.695 104.890 48.395 105.220 ;
        RECT 47.695 93.530 47.835 104.890 ;
        RECT 48.255 94.000 48.395 104.890 ;
        RECT 48.815 104.890 49.515 105.220 ;
        RECT 48.815 93.530 48.955 104.890 ;
        RECT 49.375 94.000 49.515 104.890 ;
        RECT 49.935 104.890 50.635 105.220 ;
        RECT 49.935 93.530 50.075 104.890 ;
        RECT 50.495 94.000 50.635 104.890 ;
        RECT 51.055 104.890 51.755 105.220 ;
        RECT 51.055 93.530 51.195 104.890 ;
        RECT 51.615 94.000 51.755 104.890 ;
        RECT 52.175 104.890 52.875 105.220 ;
        RECT 52.175 93.530 52.315 104.890 ;
        RECT 52.735 94.000 52.875 104.890 ;
        RECT 53.295 104.890 53.995 105.220 ;
        RECT 53.295 93.530 53.435 104.890 ;
        RECT 53.855 94.000 53.995 104.890 ;
        RECT 54.415 104.890 55.115 105.220 ;
        RECT 54.415 93.530 54.555 104.890 ;
        RECT 54.975 94.000 55.115 104.890 ;
        RECT 55.535 104.890 56.865 105.220 ;
        RECT 55.535 94.000 55.675 104.890 ;
        RECT 56.095 94.000 56.235 104.890 ;
        RECT 56.655 94.000 56.865 104.890 ;
        RECT 58.505 104.890 59.205 105.220 ;
        RECT 58.505 93.530 58.645 104.890 ;
        RECT 59.065 94.000 59.205 104.890 ;
        RECT 59.625 104.890 60.325 105.220 ;
        RECT 59.625 93.530 59.765 104.890 ;
        RECT 60.185 94.000 60.325 104.890 ;
        RECT 60.745 104.890 61.445 105.220 ;
        RECT 60.745 93.530 60.885 104.890 ;
        RECT 61.305 94.000 61.445 104.890 ;
        RECT 61.865 104.890 62.565 105.220 ;
        RECT 61.865 93.530 62.005 104.890 ;
        RECT 62.425 94.000 62.565 104.890 ;
        RECT 62.985 104.890 63.685 105.220 ;
        RECT 62.985 93.530 63.125 104.890 ;
        RECT 63.545 94.000 63.685 104.890 ;
        RECT 64.105 104.890 64.805 105.220 ;
        RECT 64.105 93.530 64.245 104.890 ;
        RECT 64.665 94.000 64.805 104.890 ;
        RECT 65.225 104.890 65.925 105.220 ;
        RECT 65.225 93.530 65.365 104.890 ;
        RECT 65.785 94.000 65.925 104.890 ;
        RECT 66.345 104.890 67.045 105.220 ;
        RECT 66.345 93.530 66.485 104.890 ;
        RECT 66.905 94.000 67.045 104.890 ;
        RECT 67.465 104.890 68.165 105.220 ;
        RECT 67.465 93.530 67.605 104.890 ;
        RECT 68.025 94.000 68.165 104.890 ;
        RECT 68.585 104.890 69.915 105.220 ;
        RECT 68.585 94.000 68.725 104.890 ;
        RECT 69.145 94.000 69.285 104.890 ;
        RECT 69.705 94.000 69.915 104.890 ;
        RECT 71.595 104.890 72.295 105.220 ;
        RECT 71.595 93.530 71.735 104.890 ;
        RECT 72.155 94.000 72.295 104.890 ;
        RECT 72.715 104.890 73.415 105.220 ;
        RECT 72.715 93.530 72.855 104.890 ;
        RECT 73.275 94.000 73.415 104.890 ;
        RECT 73.835 104.890 74.535 105.220 ;
        RECT 73.835 93.530 73.975 104.890 ;
        RECT 74.395 94.000 74.535 104.890 ;
        RECT 74.955 104.890 75.655 105.220 ;
        RECT 74.955 93.530 75.095 104.890 ;
        RECT 75.515 94.000 75.655 104.890 ;
        RECT 76.075 104.890 76.775 105.220 ;
        RECT 76.075 93.530 76.215 104.890 ;
        RECT 76.635 94.000 76.775 104.890 ;
        RECT 77.195 104.890 77.895 105.220 ;
        RECT 77.195 93.530 77.335 104.890 ;
        RECT 77.755 94.000 77.895 104.890 ;
        RECT 78.315 104.890 79.015 105.220 ;
        RECT 78.315 93.530 78.455 104.890 ;
        RECT 78.875 94.000 79.015 104.890 ;
        RECT 79.435 104.890 80.135 105.220 ;
        RECT 79.435 93.530 79.575 104.890 ;
        RECT 79.995 94.000 80.135 104.890 ;
        RECT 80.555 104.890 81.255 105.220 ;
        RECT 80.555 93.530 80.695 104.890 ;
        RECT 81.115 94.000 81.255 104.890 ;
        RECT 81.675 104.890 83.005 105.220 ;
        RECT 81.675 94.000 81.815 104.890 ;
        RECT 82.235 94.000 82.375 104.890 ;
        RECT 82.795 94.000 83.005 104.890 ;
        RECT 84.685 104.910 85.385 105.240 ;
        RECT 84.685 93.550 84.825 104.910 ;
        RECT 85.245 94.020 85.385 104.910 ;
        RECT 85.805 104.910 86.505 105.240 ;
        RECT 85.805 93.550 85.945 104.910 ;
        RECT 86.365 94.020 86.505 104.910 ;
        RECT 86.925 104.910 87.625 105.240 ;
        RECT 86.925 93.550 87.065 104.910 ;
        RECT 87.485 94.020 87.625 104.910 ;
        RECT 88.045 104.910 88.745 105.240 ;
        RECT 88.045 93.550 88.185 104.910 ;
        RECT 88.605 94.020 88.745 104.910 ;
        RECT 89.165 104.910 89.865 105.240 ;
        RECT 89.165 93.550 89.305 104.910 ;
        RECT 89.725 94.020 89.865 104.910 ;
        RECT 90.285 104.910 90.985 105.240 ;
        RECT 90.285 93.550 90.425 104.910 ;
        RECT 90.845 94.020 90.985 104.910 ;
        RECT 91.405 104.910 92.105 105.240 ;
        RECT 91.405 93.550 91.545 104.910 ;
        RECT 91.965 94.020 92.105 104.910 ;
        RECT 92.525 104.910 93.225 105.240 ;
        RECT 92.525 93.550 92.665 104.910 ;
        RECT 93.085 94.020 93.225 104.910 ;
        RECT 93.645 104.910 94.345 105.240 ;
        RECT 93.645 93.550 93.785 104.910 ;
        RECT 94.205 94.020 94.345 104.910 ;
        RECT 94.765 104.910 96.095 105.240 ;
        RECT 94.765 94.020 94.905 104.910 ;
        RECT 95.325 94.020 95.465 104.910 ;
        RECT 95.885 94.020 96.095 104.910 ;
        RECT 97.775 104.910 98.475 105.240 ;
        RECT 97.775 93.550 97.915 104.910 ;
        RECT 98.335 94.020 98.475 104.910 ;
        RECT 98.895 104.910 99.595 105.240 ;
        RECT 98.895 93.550 99.035 104.910 ;
        RECT 99.455 94.020 99.595 104.910 ;
        RECT 100.015 104.910 100.715 105.240 ;
        RECT 100.015 93.550 100.155 104.910 ;
        RECT 100.575 94.020 100.715 104.910 ;
        RECT 101.135 104.910 101.835 105.240 ;
        RECT 101.135 93.550 101.275 104.910 ;
        RECT 101.695 94.020 101.835 104.910 ;
        RECT 102.255 104.910 102.955 105.240 ;
        RECT 102.255 93.550 102.395 104.910 ;
        RECT 102.815 94.020 102.955 104.910 ;
        RECT 103.375 104.910 104.075 105.240 ;
        RECT 103.375 93.550 103.515 104.910 ;
        RECT 103.935 94.020 104.075 104.910 ;
        RECT 104.495 104.910 105.195 105.240 ;
        RECT 104.495 93.550 104.635 104.910 ;
        RECT 105.055 94.020 105.195 104.910 ;
        RECT 105.615 104.910 106.315 105.240 ;
        RECT 105.615 93.550 105.755 104.910 ;
        RECT 106.175 94.020 106.315 104.910 ;
        RECT 106.735 104.910 107.435 105.240 ;
        RECT 106.735 93.550 106.875 104.910 ;
        RECT 107.295 94.020 107.435 104.910 ;
        RECT 107.855 104.910 109.185 105.240 ;
        RECT 107.855 94.020 107.995 104.910 ;
        RECT 108.415 94.020 108.555 104.910 ;
        RECT 108.975 94.020 109.185 104.910 ;
        RECT 110.865 104.910 111.565 105.240 ;
        RECT 110.865 93.550 111.005 104.910 ;
        RECT 111.425 94.020 111.565 104.910 ;
        RECT 111.985 104.910 112.685 105.240 ;
        RECT 111.985 93.550 112.125 104.910 ;
        RECT 112.545 94.020 112.685 104.910 ;
        RECT 113.105 104.910 113.805 105.240 ;
        RECT 113.105 93.550 113.245 104.910 ;
        RECT 113.665 94.020 113.805 104.910 ;
        RECT 114.225 104.910 114.925 105.240 ;
        RECT 114.225 93.550 114.365 104.910 ;
        RECT 114.785 94.020 114.925 104.910 ;
        RECT 115.345 104.910 116.045 105.240 ;
        RECT 115.345 93.550 115.485 104.910 ;
        RECT 115.905 94.020 116.045 104.910 ;
        RECT 116.465 104.910 117.165 105.240 ;
        RECT 116.465 93.550 116.605 104.910 ;
        RECT 117.025 94.020 117.165 104.910 ;
        RECT 117.585 104.910 118.285 105.240 ;
        RECT 117.585 93.550 117.725 104.910 ;
        RECT 118.145 94.020 118.285 104.910 ;
        RECT 118.705 104.910 119.405 105.240 ;
        RECT 118.705 93.550 118.845 104.910 ;
        RECT 119.265 94.020 119.405 104.910 ;
        RECT 119.825 104.910 120.525 105.240 ;
        RECT 119.825 93.550 119.965 104.910 ;
        RECT 120.385 94.020 120.525 104.910 ;
        RECT 120.945 104.910 122.275 105.240 ;
        RECT 120.945 94.020 121.085 104.910 ;
        RECT 121.505 94.020 121.645 104.910 ;
        RECT 122.065 94.020 122.275 104.910 ;
        RECT 123.955 104.910 124.655 105.240 ;
        RECT 123.955 93.550 124.095 104.910 ;
        RECT 124.515 94.020 124.655 104.910 ;
        RECT 125.075 104.910 125.775 105.240 ;
        RECT 125.075 93.550 125.215 104.910 ;
        RECT 125.635 94.020 125.775 104.910 ;
        RECT 126.195 104.910 126.895 105.240 ;
        RECT 126.195 93.550 126.335 104.910 ;
        RECT 126.755 94.020 126.895 104.910 ;
        RECT 127.315 104.910 128.015 105.240 ;
        RECT 127.315 93.550 127.455 104.910 ;
        RECT 127.875 94.020 128.015 104.910 ;
        RECT 128.435 104.910 129.135 105.240 ;
        RECT 128.435 93.550 128.575 104.910 ;
        RECT 128.995 94.020 129.135 104.910 ;
        RECT 129.555 104.910 130.255 105.240 ;
        RECT 129.555 93.550 129.695 104.910 ;
        RECT 130.115 94.020 130.255 104.910 ;
        RECT 130.675 104.910 131.375 105.240 ;
        RECT 130.675 93.550 130.815 104.910 ;
        RECT 131.235 94.020 131.375 104.910 ;
        RECT 131.795 104.910 132.495 105.240 ;
        RECT 131.795 93.550 131.935 104.910 ;
        RECT 132.355 94.020 132.495 104.910 ;
        RECT 132.915 104.910 133.615 105.240 ;
        RECT 132.915 93.550 133.055 104.910 ;
        RECT 133.475 94.020 133.615 104.910 ;
        RECT 134.035 104.910 135.365 105.240 ;
        RECT 134.035 94.020 134.175 104.910 ;
        RECT 134.595 94.020 134.735 104.910 ;
        RECT 135.155 94.020 135.365 104.910 ;
        RECT 137.045 104.930 137.745 105.260 ;
        RECT 137.045 93.570 137.185 104.930 ;
        RECT 137.605 94.040 137.745 104.930 ;
        RECT 138.165 104.930 138.865 105.260 ;
        RECT 138.165 93.570 138.305 104.930 ;
        RECT 138.725 94.040 138.865 104.930 ;
        RECT 139.285 104.930 139.985 105.260 ;
        RECT 139.285 93.570 139.425 104.930 ;
        RECT 139.845 94.040 139.985 104.930 ;
        RECT 140.405 104.930 141.105 105.260 ;
        RECT 140.405 93.570 140.545 104.930 ;
        RECT 140.965 94.040 141.105 104.930 ;
        RECT 141.525 104.930 142.225 105.260 ;
        RECT 141.525 93.570 141.665 104.930 ;
        RECT 142.085 94.040 142.225 104.930 ;
        RECT 142.645 104.930 143.345 105.260 ;
        RECT 142.645 93.570 142.785 104.930 ;
        RECT 143.205 94.040 143.345 104.930 ;
        RECT 143.765 104.930 144.465 105.260 ;
        RECT 143.765 93.570 143.905 104.930 ;
        RECT 144.325 94.040 144.465 104.930 ;
        RECT 144.885 104.930 145.585 105.260 ;
        RECT 144.885 93.570 145.025 104.930 ;
        RECT 145.445 94.040 145.585 104.930 ;
        RECT 146.005 104.930 146.705 105.260 ;
        RECT 146.005 93.570 146.145 104.930 ;
        RECT 146.565 94.040 146.705 104.930 ;
        RECT 147.125 104.930 148.455 105.260 ;
        RECT 147.125 94.040 147.265 104.930 ;
        RECT 147.685 94.040 147.825 104.930 ;
        RECT 148.245 94.040 148.455 104.930 ;
        RECT 150.135 104.930 150.835 105.260 ;
        RECT 150.135 93.570 150.275 104.930 ;
        RECT 150.695 94.040 150.835 104.930 ;
        RECT 151.255 104.930 151.955 105.260 ;
        RECT 151.255 93.570 151.395 104.930 ;
        RECT 151.815 94.040 151.955 104.930 ;
        RECT 152.375 104.930 153.075 105.260 ;
        RECT 152.375 93.570 152.515 104.930 ;
        RECT 152.935 94.040 153.075 104.930 ;
        RECT 153.495 104.930 154.195 105.260 ;
        RECT 153.495 93.570 153.635 104.930 ;
        RECT 154.055 94.040 154.195 104.930 ;
        RECT 154.615 104.930 155.315 105.260 ;
        RECT 154.615 93.570 154.755 104.930 ;
        RECT 155.175 94.040 155.315 104.930 ;
        RECT 155.735 104.930 156.435 105.260 ;
        RECT 155.735 93.570 155.875 104.930 ;
        RECT 156.295 94.040 156.435 104.930 ;
        RECT 156.855 104.930 157.555 105.260 ;
        RECT 156.855 93.570 156.995 104.930 ;
        RECT 157.415 94.040 157.555 104.930 ;
        RECT 157.975 104.930 158.675 105.260 ;
        RECT 157.975 93.570 158.115 104.930 ;
        RECT 158.535 94.040 158.675 104.930 ;
        RECT 159.095 104.930 159.795 105.260 ;
        RECT 159.095 93.570 159.235 104.930 ;
        RECT 159.655 94.040 159.795 104.930 ;
        RECT 160.215 104.930 161.545 105.260 ;
        RECT 160.215 94.040 160.355 104.930 ;
        RECT 160.775 94.040 160.915 104.930 ;
        RECT 161.335 94.040 161.545 104.930 ;
        RECT 162.875 90.745 163.350 90.775 ;
        RECT 162.830 90.270 163.395 90.745 ;
        RECT 162.875 90.240 163.350 90.270 ;
        RECT 4.760 89.145 5.230 89.190 ;
        RECT 4.730 88.675 5.260 89.145 ;
        RECT 4.760 88.630 5.230 88.675 ;
        RECT 19.725 81.595 19.985 81.915 ;
        RECT 29.340 81.595 29.600 81.915 ;
        RECT 38.955 81.595 39.215 81.915 ;
        RECT 48.570 81.595 48.830 81.915 ;
        RECT 18.580 76.580 18.900 76.620 ;
        RECT 19.765 76.580 19.940 81.595 ;
        RECT 18.580 76.405 19.940 76.580 ;
        RECT 28.195 76.580 28.515 76.620 ;
        RECT 29.380 76.580 29.555 81.595 ;
        RECT 28.195 76.405 29.555 76.580 ;
        RECT 37.810 76.580 38.130 76.620 ;
        RECT 38.995 76.580 39.170 81.595 ;
        RECT 37.810 76.405 39.170 76.580 ;
        RECT 47.425 76.580 47.745 76.620 ;
        RECT 48.610 76.580 48.785 81.595 ;
        RECT 47.425 76.405 48.785 76.580 ;
        RECT 18.580 76.360 18.900 76.405 ;
        RECT 28.195 76.360 28.515 76.405 ;
        RECT 37.810 76.360 38.130 76.405 ;
        RECT 47.425 76.360 47.745 76.405 ;
        RECT 171.650 55.790 172.050 65.720 ;
        RECT 18.580 43.445 18.900 43.490 ;
        RECT 28.195 43.445 28.515 43.490 ;
        RECT 37.810 43.445 38.130 43.490 ;
        RECT 47.425 43.445 47.745 43.490 ;
        RECT 18.580 43.270 19.940 43.445 ;
        RECT 18.580 43.230 18.900 43.270 ;
        RECT 19.765 38.255 19.940 43.270 ;
        RECT 28.195 43.270 29.555 43.445 ;
        RECT 28.195 43.230 28.515 43.270 ;
        RECT 29.380 38.255 29.555 43.270 ;
        RECT 37.810 43.270 39.170 43.445 ;
        RECT 37.810 43.230 38.130 43.270 ;
        RECT 38.995 38.255 39.170 43.270 ;
        RECT 47.425 43.270 48.785 43.445 ;
        RECT 47.425 43.230 47.745 43.270 ;
        RECT 48.610 38.255 48.785 43.270 ;
        RECT 19.725 37.935 19.985 38.255 ;
        RECT 29.340 37.935 29.600 38.255 ;
        RECT 38.955 37.935 39.215 38.255 ;
        RECT 48.570 37.935 48.830 38.255 ;
        RECT 4.750 33.685 5.220 33.730 ;
        RECT 4.720 33.215 5.250 33.685 ;
        RECT 4.750 33.170 5.220 33.215 ;
        RECT 148.750 31.575 149.070 31.620 ;
        RECT 148.750 31.405 151.205 31.575 ;
        RECT 148.750 31.360 149.070 31.405 ;
        RECT 151.020 29.590 151.190 31.405 ;
        RECT 163.275 29.690 163.750 29.735 ;
        RECT 150.975 29.270 151.235 29.590 ;
        RECT 163.245 29.215 163.780 29.690 ;
        RECT 163.275 29.170 163.750 29.215 ;
        RECT 6.595 15.610 6.735 26.970 ;
        RECT 7.155 15.610 7.295 26.500 ;
        RECT 6.595 15.280 7.295 15.610 ;
        RECT 7.715 15.610 7.855 26.970 ;
        RECT 8.275 15.610 8.415 26.500 ;
        RECT 7.715 15.280 8.415 15.610 ;
        RECT 8.835 15.610 8.975 26.970 ;
        RECT 9.395 15.610 9.535 26.500 ;
        RECT 8.835 15.280 9.535 15.610 ;
        RECT 9.955 15.610 10.095 26.970 ;
        RECT 10.515 15.610 10.655 26.500 ;
        RECT 9.955 15.280 10.655 15.610 ;
        RECT 11.075 15.610 11.215 26.970 ;
        RECT 11.635 15.610 11.775 26.500 ;
        RECT 11.075 15.280 11.775 15.610 ;
        RECT 12.195 15.610 12.335 26.970 ;
        RECT 12.755 15.610 12.895 26.500 ;
        RECT 12.195 15.280 12.895 15.610 ;
        RECT 13.315 15.610 13.455 26.970 ;
        RECT 13.875 15.610 14.015 26.500 ;
        RECT 13.315 15.280 14.015 15.610 ;
        RECT 14.435 15.610 14.575 26.970 ;
        RECT 14.995 15.610 15.135 26.500 ;
        RECT 14.435 15.280 15.135 15.610 ;
        RECT 15.555 15.610 15.695 26.970 ;
        RECT 16.115 15.610 16.255 26.500 ;
        RECT 15.555 15.280 16.255 15.610 ;
        RECT 16.675 15.610 16.815 26.500 ;
        RECT 17.235 15.610 17.375 26.500 ;
        RECT 17.795 15.610 18.005 26.500 ;
        RECT 16.675 15.280 18.005 15.610 ;
        RECT 19.685 15.610 19.825 26.970 ;
        RECT 20.245 15.610 20.385 26.500 ;
        RECT 19.685 15.280 20.385 15.610 ;
        RECT 20.805 15.610 20.945 26.970 ;
        RECT 21.365 15.610 21.505 26.500 ;
        RECT 20.805 15.280 21.505 15.610 ;
        RECT 21.925 15.610 22.065 26.970 ;
        RECT 22.485 15.610 22.625 26.500 ;
        RECT 21.925 15.280 22.625 15.610 ;
        RECT 23.045 15.610 23.185 26.970 ;
        RECT 23.605 15.610 23.745 26.500 ;
        RECT 23.045 15.280 23.745 15.610 ;
        RECT 24.165 15.610 24.305 26.970 ;
        RECT 24.725 15.610 24.865 26.500 ;
        RECT 24.165 15.280 24.865 15.610 ;
        RECT 25.285 15.610 25.425 26.970 ;
        RECT 25.845 15.610 25.985 26.500 ;
        RECT 25.285 15.280 25.985 15.610 ;
        RECT 26.405 15.610 26.545 26.970 ;
        RECT 26.965 15.610 27.105 26.500 ;
        RECT 26.405 15.280 27.105 15.610 ;
        RECT 27.525 15.610 27.665 26.970 ;
        RECT 28.085 15.610 28.225 26.500 ;
        RECT 27.525 15.280 28.225 15.610 ;
        RECT 28.645 15.610 28.785 26.970 ;
        RECT 29.205 15.610 29.345 26.500 ;
        RECT 28.645 15.280 29.345 15.610 ;
        RECT 29.765 15.610 29.905 26.500 ;
        RECT 30.325 15.610 30.465 26.500 ;
        RECT 30.885 15.610 31.095 26.500 ;
        RECT 29.765 15.280 31.095 15.610 ;
        RECT 32.775 15.590 32.915 26.950 ;
        RECT 33.335 15.590 33.475 26.480 ;
        RECT 32.775 15.260 33.475 15.590 ;
        RECT 33.895 15.590 34.035 26.950 ;
        RECT 34.455 15.590 34.595 26.480 ;
        RECT 33.895 15.260 34.595 15.590 ;
        RECT 35.015 15.590 35.155 26.950 ;
        RECT 35.575 15.590 35.715 26.480 ;
        RECT 35.015 15.260 35.715 15.590 ;
        RECT 36.135 15.590 36.275 26.950 ;
        RECT 36.695 15.590 36.835 26.480 ;
        RECT 36.135 15.260 36.835 15.590 ;
        RECT 37.255 15.590 37.395 26.950 ;
        RECT 37.815 15.590 37.955 26.480 ;
        RECT 37.255 15.260 37.955 15.590 ;
        RECT 38.375 15.590 38.515 26.950 ;
        RECT 38.935 15.590 39.075 26.480 ;
        RECT 38.375 15.260 39.075 15.590 ;
        RECT 39.495 15.590 39.635 26.950 ;
        RECT 40.055 15.590 40.195 26.480 ;
        RECT 39.495 15.260 40.195 15.590 ;
        RECT 40.615 15.590 40.755 26.950 ;
        RECT 41.175 15.590 41.315 26.480 ;
        RECT 40.615 15.260 41.315 15.590 ;
        RECT 41.735 15.590 41.875 26.950 ;
        RECT 42.295 15.590 42.435 26.480 ;
        RECT 41.735 15.260 42.435 15.590 ;
        RECT 42.855 15.590 42.995 26.480 ;
        RECT 43.415 15.590 43.555 26.480 ;
        RECT 43.975 15.590 44.185 26.480 ;
        RECT 42.855 15.260 44.185 15.590 ;
        RECT 45.865 15.590 46.005 26.950 ;
        RECT 46.425 15.590 46.565 26.480 ;
        RECT 45.865 15.260 46.565 15.590 ;
        RECT 46.985 15.590 47.125 26.950 ;
        RECT 47.545 15.590 47.685 26.480 ;
        RECT 46.985 15.260 47.685 15.590 ;
        RECT 48.105 15.590 48.245 26.950 ;
        RECT 48.665 15.590 48.805 26.480 ;
        RECT 48.105 15.260 48.805 15.590 ;
        RECT 49.225 15.590 49.365 26.950 ;
        RECT 49.785 15.590 49.925 26.480 ;
        RECT 49.225 15.260 49.925 15.590 ;
        RECT 50.345 15.590 50.485 26.950 ;
        RECT 50.905 15.590 51.045 26.480 ;
        RECT 50.345 15.260 51.045 15.590 ;
        RECT 51.465 15.590 51.605 26.950 ;
        RECT 52.025 15.590 52.165 26.480 ;
        RECT 51.465 15.260 52.165 15.590 ;
        RECT 52.585 15.590 52.725 26.950 ;
        RECT 53.145 15.590 53.285 26.480 ;
        RECT 52.585 15.260 53.285 15.590 ;
        RECT 53.705 15.590 53.845 26.950 ;
        RECT 54.265 15.590 54.405 26.480 ;
        RECT 53.705 15.260 54.405 15.590 ;
        RECT 54.825 15.590 54.965 26.950 ;
        RECT 55.385 15.590 55.525 26.480 ;
        RECT 54.825 15.260 55.525 15.590 ;
        RECT 55.945 15.590 56.085 26.480 ;
        RECT 56.505 15.590 56.645 26.480 ;
        RECT 57.065 15.590 57.275 26.480 ;
        RECT 55.945 15.260 57.275 15.590 ;
        RECT 58.915 15.590 59.055 26.950 ;
        RECT 59.475 15.590 59.615 26.480 ;
        RECT 58.915 15.260 59.615 15.590 ;
        RECT 60.035 15.590 60.175 26.950 ;
        RECT 60.595 15.590 60.735 26.480 ;
        RECT 60.035 15.260 60.735 15.590 ;
        RECT 61.155 15.590 61.295 26.950 ;
        RECT 61.715 15.590 61.855 26.480 ;
        RECT 61.155 15.260 61.855 15.590 ;
        RECT 62.275 15.590 62.415 26.950 ;
        RECT 62.835 15.590 62.975 26.480 ;
        RECT 62.275 15.260 62.975 15.590 ;
        RECT 63.395 15.590 63.535 26.950 ;
        RECT 63.955 15.590 64.095 26.480 ;
        RECT 63.395 15.260 64.095 15.590 ;
        RECT 64.515 15.590 64.655 26.950 ;
        RECT 65.075 15.590 65.215 26.480 ;
        RECT 64.515 15.260 65.215 15.590 ;
        RECT 65.635 15.590 65.775 26.950 ;
        RECT 66.195 15.590 66.335 26.480 ;
        RECT 65.635 15.260 66.335 15.590 ;
        RECT 66.755 15.590 66.895 26.950 ;
        RECT 67.315 15.590 67.455 26.480 ;
        RECT 66.755 15.260 67.455 15.590 ;
        RECT 67.875 15.590 68.015 26.950 ;
        RECT 68.435 15.590 68.575 26.480 ;
        RECT 67.875 15.260 68.575 15.590 ;
        RECT 68.995 15.590 69.135 26.480 ;
        RECT 69.555 15.590 69.695 26.480 ;
        RECT 70.115 15.590 70.325 26.480 ;
        RECT 68.995 15.260 70.325 15.590 ;
        RECT 72.005 15.590 72.145 26.950 ;
        RECT 72.565 15.590 72.705 26.480 ;
        RECT 72.005 15.260 72.705 15.590 ;
        RECT 73.125 15.590 73.265 26.950 ;
        RECT 73.685 15.590 73.825 26.480 ;
        RECT 73.125 15.260 73.825 15.590 ;
        RECT 74.245 15.590 74.385 26.950 ;
        RECT 74.805 15.590 74.945 26.480 ;
        RECT 74.245 15.260 74.945 15.590 ;
        RECT 75.365 15.590 75.505 26.950 ;
        RECT 75.925 15.590 76.065 26.480 ;
        RECT 75.365 15.260 76.065 15.590 ;
        RECT 76.485 15.590 76.625 26.950 ;
        RECT 77.045 15.590 77.185 26.480 ;
        RECT 76.485 15.260 77.185 15.590 ;
        RECT 77.605 15.590 77.745 26.950 ;
        RECT 78.165 15.590 78.305 26.480 ;
        RECT 77.605 15.260 78.305 15.590 ;
        RECT 78.725 15.590 78.865 26.950 ;
        RECT 79.285 15.590 79.425 26.480 ;
        RECT 78.725 15.260 79.425 15.590 ;
        RECT 79.845 15.590 79.985 26.950 ;
        RECT 80.405 15.590 80.545 26.480 ;
        RECT 79.845 15.260 80.545 15.590 ;
        RECT 80.965 15.590 81.105 26.950 ;
        RECT 81.525 15.590 81.665 26.480 ;
        RECT 80.965 15.260 81.665 15.590 ;
        RECT 82.085 15.590 82.225 26.480 ;
        RECT 82.645 15.590 82.785 26.480 ;
        RECT 83.205 15.590 83.415 26.480 ;
        RECT 82.085 15.260 83.415 15.590 ;
        RECT 85.095 15.570 85.235 26.930 ;
        RECT 85.655 15.570 85.795 26.460 ;
        RECT 85.095 15.240 85.795 15.570 ;
        RECT 86.215 15.570 86.355 26.930 ;
        RECT 86.775 15.570 86.915 26.460 ;
        RECT 86.215 15.240 86.915 15.570 ;
        RECT 87.335 15.570 87.475 26.930 ;
        RECT 87.895 15.570 88.035 26.460 ;
        RECT 87.335 15.240 88.035 15.570 ;
        RECT 88.455 15.570 88.595 26.930 ;
        RECT 89.015 15.570 89.155 26.460 ;
        RECT 88.455 15.240 89.155 15.570 ;
        RECT 89.575 15.570 89.715 26.930 ;
        RECT 90.135 15.570 90.275 26.460 ;
        RECT 89.575 15.240 90.275 15.570 ;
        RECT 90.695 15.570 90.835 26.930 ;
        RECT 91.255 15.570 91.395 26.460 ;
        RECT 90.695 15.240 91.395 15.570 ;
        RECT 91.815 15.570 91.955 26.930 ;
        RECT 92.375 15.570 92.515 26.460 ;
        RECT 91.815 15.240 92.515 15.570 ;
        RECT 92.935 15.570 93.075 26.930 ;
        RECT 93.495 15.570 93.635 26.460 ;
        RECT 92.935 15.240 93.635 15.570 ;
        RECT 94.055 15.570 94.195 26.930 ;
        RECT 94.615 15.570 94.755 26.460 ;
        RECT 94.055 15.240 94.755 15.570 ;
        RECT 95.175 15.570 95.315 26.460 ;
        RECT 95.735 15.570 95.875 26.460 ;
        RECT 96.295 15.570 96.505 26.460 ;
        RECT 95.175 15.240 96.505 15.570 ;
        RECT 98.185 15.570 98.325 26.930 ;
        RECT 98.745 15.570 98.885 26.460 ;
        RECT 98.185 15.240 98.885 15.570 ;
        RECT 99.305 15.570 99.445 26.930 ;
        RECT 99.865 15.570 100.005 26.460 ;
        RECT 99.305 15.240 100.005 15.570 ;
        RECT 100.425 15.570 100.565 26.930 ;
        RECT 100.985 15.570 101.125 26.460 ;
        RECT 100.425 15.240 101.125 15.570 ;
        RECT 101.545 15.570 101.685 26.930 ;
        RECT 102.105 15.570 102.245 26.460 ;
        RECT 101.545 15.240 102.245 15.570 ;
        RECT 102.665 15.570 102.805 26.930 ;
        RECT 103.225 15.570 103.365 26.460 ;
        RECT 102.665 15.240 103.365 15.570 ;
        RECT 103.785 15.570 103.925 26.930 ;
        RECT 104.345 15.570 104.485 26.460 ;
        RECT 103.785 15.240 104.485 15.570 ;
        RECT 104.905 15.570 105.045 26.930 ;
        RECT 105.465 15.570 105.605 26.460 ;
        RECT 104.905 15.240 105.605 15.570 ;
        RECT 106.025 15.570 106.165 26.930 ;
        RECT 106.585 15.570 106.725 26.460 ;
        RECT 106.025 15.240 106.725 15.570 ;
        RECT 107.145 15.570 107.285 26.930 ;
        RECT 107.705 15.570 107.845 26.460 ;
        RECT 107.145 15.240 107.845 15.570 ;
        RECT 108.265 15.570 108.405 26.460 ;
        RECT 108.825 15.570 108.965 26.460 ;
        RECT 109.385 15.570 109.595 26.460 ;
        RECT 108.265 15.240 109.595 15.570 ;
        RECT 111.275 15.570 111.415 26.930 ;
        RECT 111.835 15.570 111.975 26.460 ;
        RECT 111.275 15.240 111.975 15.570 ;
        RECT 112.395 15.570 112.535 26.930 ;
        RECT 112.955 15.570 113.095 26.460 ;
        RECT 112.395 15.240 113.095 15.570 ;
        RECT 113.515 15.570 113.655 26.930 ;
        RECT 114.075 15.570 114.215 26.460 ;
        RECT 113.515 15.240 114.215 15.570 ;
        RECT 114.635 15.570 114.775 26.930 ;
        RECT 115.195 15.570 115.335 26.460 ;
        RECT 114.635 15.240 115.335 15.570 ;
        RECT 115.755 15.570 115.895 26.930 ;
        RECT 116.315 15.570 116.455 26.460 ;
        RECT 115.755 15.240 116.455 15.570 ;
        RECT 116.875 15.570 117.015 26.930 ;
        RECT 117.435 15.570 117.575 26.460 ;
        RECT 116.875 15.240 117.575 15.570 ;
        RECT 117.995 15.570 118.135 26.930 ;
        RECT 118.555 15.570 118.695 26.460 ;
        RECT 117.995 15.240 118.695 15.570 ;
        RECT 119.115 15.570 119.255 26.930 ;
        RECT 119.675 15.570 119.815 26.460 ;
        RECT 119.115 15.240 119.815 15.570 ;
        RECT 120.235 15.570 120.375 26.930 ;
        RECT 120.795 15.570 120.935 26.460 ;
        RECT 120.235 15.240 120.935 15.570 ;
        RECT 121.355 15.570 121.495 26.460 ;
        RECT 121.915 15.570 122.055 26.460 ;
        RECT 122.475 15.570 122.685 26.460 ;
        RECT 121.355 15.240 122.685 15.570 ;
        RECT 124.365 15.570 124.505 26.930 ;
        RECT 124.925 15.570 125.065 26.460 ;
        RECT 124.365 15.240 125.065 15.570 ;
        RECT 125.485 15.570 125.625 26.930 ;
        RECT 126.045 15.570 126.185 26.460 ;
        RECT 125.485 15.240 126.185 15.570 ;
        RECT 126.605 15.570 126.745 26.930 ;
        RECT 127.165 15.570 127.305 26.460 ;
        RECT 126.605 15.240 127.305 15.570 ;
        RECT 127.725 15.570 127.865 26.930 ;
        RECT 128.285 15.570 128.425 26.460 ;
        RECT 127.725 15.240 128.425 15.570 ;
        RECT 128.845 15.570 128.985 26.930 ;
        RECT 129.405 15.570 129.545 26.460 ;
        RECT 128.845 15.240 129.545 15.570 ;
        RECT 129.965 15.570 130.105 26.930 ;
        RECT 130.525 15.570 130.665 26.460 ;
        RECT 129.965 15.240 130.665 15.570 ;
        RECT 131.085 15.570 131.225 26.930 ;
        RECT 131.645 15.570 131.785 26.460 ;
        RECT 131.085 15.240 131.785 15.570 ;
        RECT 132.205 15.570 132.345 26.930 ;
        RECT 132.765 15.570 132.905 26.460 ;
        RECT 132.205 15.240 132.905 15.570 ;
        RECT 133.325 15.570 133.465 26.930 ;
        RECT 133.885 15.570 134.025 26.460 ;
        RECT 133.325 15.240 134.025 15.570 ;
        RECT 134.445 15.570 134.585 26.460 ;
        RECT 135.005 15.570 135.145 26.460 ;
        RECT 135.565 15.570 135.775 26.460 ;
        RECT 134.445 15.240 135.775 15.570 ;
        RECT 137.455 15.550 137.595 26.910 ;
        RECT 138.015 15.550 138.155 26.440 ;
        RECT 137.455 15.220 138.155 15.550 ;
        RECT 138.575 15.550 138.715 26.910 ;
        RECT 139.135 15.550 139.275 26.440 ;
        RECT 138.575 15.220 139.275 15.550 ;
        RECT 139.695 15.550 139.835 26.910 ;
        RECT 140.255 15.550 140.395 26.440 ;
        RECT 139.695 15.220 140.395 15.550 ;
        RECT 140.815 15.550 140.955 26.910 ;
        RECT 141.375 15.550 141.515 26.440 ;
        RECT 140.815 15.220 141.515 15.550 ;
        RECT 141.935 15.550 142.075 26.910 ;
        RECT 142.495 15.550 142.635 26.440 ;
        RECT 141.935 15.220 142.635 15.550 ;
        RECT 143.055 15.550 143.195 26.910 ;
        RECT 143.615 15.550 143.755 26.440 ;
        RECT 143.055 15.220 143.755 15.550 ;
        RECT 144.175 15.550 144.315 26.910 ;
        RECT 144.735 15.550 144.875 26.440 ;
        RECT 144.175 15.220 144.875 15.550 ;
        RECT 145.295 15.550 145.435 26.910 ;
        RECT 145.855 15.550 145.995 26.440 ;
        RECT 145.295 15.220 145.995 15.550 ;
        RECT 146.415 15.550 146.555 26.910 ;
        RECT 146.975 15.550 147.115 26.440 ;
        RECT 146.415 15.220 147.115 15.550 ;
        RECT 147.535 15.550 147.675 26.440 ;
        RECT 148.095 15.550 148.235 26.440 ;
        RECT 148.655 15.550 148.865 26.440 ;
        RECT 147.535 15.220 148.865 15.550 ;
        RECT 150.545 15.550 150.685 26.910 ;
        RECT 151.105 15.550 151.245 26.440 ;
        RECT 150.545 15.220 151.245 15.550 ;
        RECT 151.665 15.550 151.805 26.910 ;
        RECT 152.225 15.550 152.365 26.440 ;
        RECT 151.665 15.220 152.365 15.550 ;
        RECT 152.785 15.550 152.925 26.910 ;
        RECT 153.345 15.550 153.485 26.440 ;
        RECT 152.785 15.220 153.485 15.550 ;
        RECT 153.905 15.550 154.045 26.910 ;
        RECT 154.465 15.550 154.605 26.440 ;
        RECT 153.905 15.220 154.605 15.550 ;
        RECT 155.025 15.550 155.165 26.910 ;
        RECT 155.585 15.550 155.725 26.440 ;
        RECT 155.025 15.220 155.725 15.550 ;
        RECT 156.145 15.550 156.285 26.910 ;
        RECT 156.705 15.550 156.845 26.440 ;
        RECT 156.145 15.220 156.845 15.550 ;
        RECT 157.265 15.550 157.405 26.910 ;
        RECT 157.825 15.550 157.965 26.440 ;
        RECT 157.265 15.220 157.965 15.550 ;
        RECT 158.385 15.550 158.525 26.910 ;
        RECT 158.945 15.550 159.085 26.440 ;
        RECT 158.385 15.220 159.085 15.550 ;
        RECT 159.505 15.550 159.645 26.910 ;
        RECT 160.065 15.550 160.205 26.440 ;
        RECT 159.505 15.220 160.205 15.550 ;
        RECT 160.625 15.550 160.765 26.440 ;
        RECT 161.185 15.550 161.325 26.440 ;
        RECT 161.745 15.550 161.955 26.440 ;
        RECT 160.625 15.220 161.955 15.550 ;
        RECT 6.625 13.230 7.325 13.560 ;
        RECT 6.625 1.870 6.765 13.230 ;
        RECT 7.185 2.340 7.325 13.230 ;
        RECT 7.745 13.230 8.445 13.560 ;
        RECT 7.745 1.870 7.885 13.230 ;
        RECT 8.305 2.340 8.445 13.230 ;
        RECT 8.865 13.230 9.565 13.560 ;
        RECT 8.865 1.870 9.005 13.230 ;
        RECT 9.425 2.340 9.565 13.230 ;
        RECT 9.985 13.230 10.685 13.560 ;
        RECT 9.985 1.870 10.125 13.230 ;
        RECT 10.545 2.340 10.685 13.230 ;
        RECT 11.105 13.230 11.805 13.560 ;
        RECT 11.105 1.870 11.245 13.230 ;
        RECT 11.665 2.340 11.805 13.230 ;
        RECT 12.225 13.230 12.925 13.560 ;
        RECT 12.225 1.870 12.365 13.230 ;
        RECT 12.785 2.340 12.925 13.230 ;
        RECT 13.345 13.230 14.045 13.560 ;
        RECT 13.345 1.870 13.485 13.230 ;
        RECT 13.905 2.340 14.045 13.230 ;
        RECT 14.465 13.230 15.165 13.560 ;
        RECT 14.465 1.870 14.605 13.230 ;
        RECT 15.025 2.340 15.165 13.230 ;
        RECT 15.585 13.230 16.285 13.560 ;
        RECT 15.585 1.870 15.725 13.230 ;
        RECT 16.145 2.340 16.285 13.230 ;
        RECT 16.705 13.230 18.035 13.560 ;
        RECT 16.705 2.340 16.845 13.230 ;
        RECT 17.265 2.340 17.405 13.230 ;
        RECT 17.825 2.340 18.035 13.230 ;
        RECT 19.715 13.230 20.415 13.560 ;
        RECT 19.715 1.870 19.855 13.230 ;
        RECT 20.275 2.340 20.415 13.230 ;
        RECT 20.835 13.230 21.535 13.560 ;
        RECT 20.835 1.870 20.975 13.230 ;
        RECT 21.395 2.340 21.535 13.230 ;
        RECT 21.955 13.230 22.655 13.560 ;
        RECT 21.955 1.870 22.095 13.230 ;
        RECT 22.515 2.340 22.655 13.230 ;
        RECT 23.075 13.230 23.775 13.560 ;
        RECT 23.075 1.870 23.215 13.230 ;
        RECT 23.635 2.340 23.775 13.230 ;
        RECT 24.195 13.230 24.895 13.560 ;
        RECT 24.195 1.870 24.335 13.230 ;
        RECT 24.755 2.340 24.895 13.230 ;
        RECT 25.315 13.230 26.015 13.560 ;
        RECT 25.315 1.870 25.455 13.230 ;
        RECT 25.875 2.340 26.015 13.230 ;
        RECT 26.435 13.230 27.135 13.560 ;
        RECT 26.435 1.870 26.575 13.230 ;
        RECT 26.995 2.340 27.135 13.230 ;
        RECT 27.555 13.230 28.255 13.560 ;
        RECT 27.555 1.870 27.695 13.230 ;
        RECT 28.115 2.340 28.255 13.230 ;
        RECT 28.675 13.230 29.375 13.560 ;
        RECT 28.675 1.870 28.815 13.230 ;
        RECT 29.235 2.340 29.375 13.230 ;
        RECT 29.795 13.230 31.125 13.560 ;
        RECT 29.795 2.340 29.935 13.230 ;
        RECT 30.355 2.340 30.495 13.230 ;
        RECT 30.915 2.340 31.125 13.230 ;
        RECT 32.805 13.250 33.505 13.580 ;
        RECT 32.805 1.890 32.945 13.250 ;
        RECT 33.365 2.360 33.505 13.250 ;
        RECT 33.925 13.250 34.625 13.580 ;
        RECT 33.925 1.890 34.065 13.250 ;
        RECT 34.485 2.360 34.625 13.250 ;
        RECT 35.045 13.250 35.745 13.580 ;
        RECT 35.045 1.890 35.185 13.250 ;
        RECT 35.605 2.360 35.745 13.250 ;
        RECT 36.165 13.250 36.865 13.580 ;
        RECT 36.165 1.890 36.305 13.250 ;
        RECT 36.725 2.360 36.865 13.250 ;
        RECT 37.285 13.250 37.985 13.580 ;
        RECT 37.285 1.890 37.425 13.250 ;
        RECT 37.845 2.360 37.985 13.250 ;
        RECT 38.405 13.250 39.105 13.580 ;
        RECT 38.405 1.890 38.545 13.250 ;
        RECT 38.965 2.360 39.105 13.250 ;
        RECT 39.525 13.250 40.225 13.580 ;
        RECT 39.525 1.890 39.665 13.250 ;
        RECT 40.085 2.360 40.225 13.250 ;
        RECT 40.645 13.250 41.345 13.580 ;
        RECT 40.645 1.890 40.785 13.250 ;
        RECT 41.205 2.360 41.345 13.250 ;
        RECT 41.765 13.250 42.465 13.580 ;
        RECT 41.765 1.890 41.905 13.250 ;
        RECT 42.325 2.360 42.465 13.250 ;
        RECT 42.885 13.250 44.215 13.580 ;
        RECT 42.885 2.360 43.025 13.250 ;
        RECT 43.445 2.360 43.585 13.250 ;
        RECT 44.005 2.360 44.215 13.250 ;
        RECT 45.895 13.250 46.595 13.580 ;
        RECT 45.895 1.890 46.035 13.250 ;
        RECT 46.455 2.360 46.595 13.250 ;
        RECT 47.015 13.250 47.715 13.580 ;
        RECT 47.015 1.890 47.155 13.250 ;
        RECT 47.575 2.360 47.715 13.250 ;
        RECT 48.135 13.250 48.835 13.580 ;
        RECT 48.135 1.890 48.275 13.250 ;
        RECT 48.695 2.360 48.835 13.250 ;
        RECT 49.255 13.250 49.955 13.580 ;
        RECT 49.255 1.890 49.395 13.250 ;
        RECT 49.815 2.360 49.955 13.250 ;
        RECT 50.375 13.250 51.075 13.580 ;
        RECT 50.375 1.890 50.515 13.250 ;
        RECT 50.935 2.360 51.075 13.250 ;
        RECT 51.495 13.250 52.195 13.580 ;
        RECT 51.495 1.890 51.635 13.250 ;
        RECT 52.055 2.360 52.195 13.250 ;
        RECT 52.615 13.250 53.315 13.580 ;
        RECT 52.615 1.890 52.755 13.250 ;
        RECT 53.175 2.360 53.315 13.250 ;
        RECT 53.735 13.250 54.435 13.580 ;
        RECT 53.735 1.890 53.875 13.250 ;
        RECT 54.295 2.360 54.435 13.250 ;
        RECT 54.855 13.250 55.555 13.580 ;
        RECT 54.855 1.890 54.995 13.250 ;
        RECT 55.415 2.360 55.555 13.250 ;
        RECT 55.975 13.250 57.305 13.580 ;
        RECT 55.975 2.360 56.115 13.250 ;
        RECT 56.535 2.360 56.675 13.250 ;
        RECT 57.095 2.360 57.305 13.250 ;
        RECT 58.945 13.250 59.645 13.580 ;
        RECT 58.945 1.890 59.085 13.250 ;
        RECT 59.505 2.360 59.645 13.250 ;
        RECT 60.065 13.250 60.765 13.580 ;
        RECT 60.065 1.890 60.205 13.250 ;
        RECT 60.625 2.360 60.765 13.250 ;
        RECT 61.185 13.250 61.885 13.580 ;
        RECT 61.185 1.890 61.325 13.250 ;
        RECT 61.745 2.360 61.885 13.250 ;
        RECT 62.305 13.250 63.005 13.580 ;
        RECT 62.305 1.890 62.445 13.250 ;
        RECT 62.865 2.360 63.005 13.250 ;
        RECT 63.425 13.250 64.125 13.580 ;
        RECT 63.425 1.890 63.565 13.250 ;
        RECT 63.985 2.360 64.125 13.250 ;
        RECT 64.545 13.250 65.245 13.580 ;
        RECT 64.545 1.890 64.685 13.250 ;
        RECT 65.105 2.360 65.245 13.250 ;
        RECT 65.665 13.250 66.365 13.580 ;
        RECT 65.665 1.890 65.805 13.250 ;
        RECT 66.225 2.360 66.365 13.250 ;
        RECT 66.785 13.250 67.485 13.580 ;
        RECT 66.785 1.890 66.925 13.250 ;
        RECT 67.345 2.360 67.485 13.250 ;
        RECT 67.905 13.250 68.605 13.580 ;
        RECT 67.905 1.890 68.045 13.250 ;
        RECT 68.465 2.360 68.605 13.250 ;
        RECT 69.025 13.250 70.355 13.580 ;
        RECT 69.025 2.360 69.165 13.250 ;
        RECT 69.585 2.360 69.725 13.250 ;
        RECT 70.145 2.360 70.355 13.250 ;
        RECT 72.035 13.250 72.735 13.580 ;
        RECT 72.035 1.890 72.175 13.250 ;
        RECT 72.595 2.360 72.735 13.250 ;
        RECT 73.155 13.250 73.855 13.580 ;
        RECT 73.155 1.890 73.295 13.250 ;
        RECT 73.715 2.360 73.855 13.250 ;
        RECT 74.275 13.250 74.975 13.580 ;
        RECT 74.275 1.890 74.415 13.250 ;
        RECT 74.835 2.360 74.975 13.250 ;
        RECT 75.395 13.250 76.095 13.580 ;
        RECT 75.395 1.890 75.535 13.250 ;
        RECT 75.955 2.360 76.095 13.250 ;
        RECT 76.515 13.250 77.215 13.580 ;
        RECT 76.515 1.890 76.655 13.250 ;
        RECT 77.075 2.360 77.215 13.250 ;
        RECT 77.635 13.250 78.335 13.580 ;
        RECT 77.635 1.890 77.775 13.250 ;
        RECT 78.195 2.360 78.335 13.250 ;
        RECT 78.755 13.250 79.455 13.580 ;
        RECT 78.755 1.890 78.895 13.250 ;
        RECT 79.315 2.360 79.455 13.250 ;
        RECT 79.875 13.250 80.575 13.580 ;
        RECT 79.875 1.890 80.015 13.250 ;
        RECT 80.435 2.360 80.575 13.250 ;
        RECT 80.995 13.250 81.695 13.580 ;
        RECT 80.995 1.890 81.135 13.250 ;
        RECT 81.555 2.360 81.695 13.250 ;
        RECT 82.115 13.250 83.445 13.580 ;
        RECT 82.115 2.360 82.255 13.250 ;
        RECT 82.675 2.360 82.815 13.250 ;
        RECT 83.235 2.360 83.445 13.250 ;
        RECT 85.125 13.270 85.825 13.600 ;
        RECT 85.125 1.910 85.265 13.270 ;
        RECT 85.685 2.380 85.825 13.270 ;
        RECT 86.245 13.270 86.945 13.600 ;
        RECT 86.245 1.910 86.385 13.270 ;
        RECT 86.805 2.380 86.945 13.270 ;
        RECT 87.365 13.270 88.065 13.600 ;
        RECT 87.365 1.910 87.505 13.270 ;
        RECT 87.925 2.380 88.065 13.270 ;
        RECT 88.485 13.270 89.185 13.600 ;
        RECT 88.485 1.910 88.625 13.270 ;
        RECT 89.045 2.380 89.185 13.270 ;
        RECT 89.605 13.270 90.305 13.600 ;
        RECT 89.605 1.910 89.745 13.270 ;
        RECT 90.165 2.380 90.305 13.270 ;
        RECT 90.725 13.270 91.425 13.600 ;
        RECT 90.725 1.910 90.865 13.270 ;
        RECT 91.285 2.380 91.425 13.270 ;
        RECT 91.845 13.270 92.545 13.600 ;
        RECT 91.845 1.910 91.985 13.270 ;
        RECT 92.405 2.380 92.545 13.270 ;
        RECT 92.965 13.270 93.665 13.600 ;
        RECT 92.965 1.910 93.105 13.270 ;
        RECT 93.525 2.380 93.665 13.270 ;
        RECT 94.085 13.270 94.785 13.600 ;
        RECT 94.085 1.910 94.225 13.270 ;
        RECT 94.645 2.380 94.785 13.270 ;
        RECT 95.205 13.270 96.535 13.600 ;
        RECT 95.205 2.380 95.345 13.270 ;
        RECT 95.765 2.380 95.905 13.270 ;
        RECT 96.325 2.380 96.535 13.270 ;
        RECT 98.215 13.270 98.915 13.600 ;
        RECT 98.215 1.910 98.355 13.270 ;
        RECT 98.775 2.380 98.915 13.270 ;
        RECT 99.335 13.270 100.035 13.600 ;
        RECT 99.335 1.910 99.475 13.270 ;
        RECT 99.895 2.380 100.035 13.270 ;
        RECT 100.455 13.270 101.155 13.600 ;
        RECT 100.455 1.910 100.595 13.270 ;
        RECT 101.015 2.380 101.155 13.270 ;
        RECT 101.575 13.270 102.275 13.600 ;
        RECT 101.575 1.910 101.715 13.270 ;
        RECT 102.135 2.380 102.275 13.270 ;
        RECT 102.695 13.270 103.395 13.600 ;
        RECT 102.695 1.910 102.835 13.270 ;
        RECT 103.255 2.380 103.395 13.270 ;
        RECT 103.815 13.270 104.515 13.600 ;
        RECT 103.815 1.910 103.955 13.270 ;
        RECT 104.375 2.380 104.515 13.270 ;
        RECT 104.935 13.270 105.635 13.600 ;
        RECT 104.935 1.910 105.075 13.270 ;
        RECT 105.495 2.380 105.635 13.270 ;
        RECT 106.055 13.270 106.755 13.600 ;
        RECT 106.055 1.910 106.195 13.270 ;
        RECT 106.615 2.380 106.755 13.270 ;
        RECT 107.175 13.270 107.875 13.600 ;
        RECT 107.175 1.910 107.315 13.270 ;
        RECT 107.735 2.380 107.875 13.270 ;
        RECT 108.295 13.270 109.625 13.600 ;
        RECT 108.295 2.380 108.435 13.270 ;
        RECT 108.855 2.380 108.995 13.270 ;
        RECT 109.415 2.380 109.625 13.270 ;
        RECT 111.305 13.270 112.005 13.600 ;
        RECT 111.305 1.910 111.445 13.270 ;
        RECT 111.865 2.380 112.005 13.270 ;
        RECT 112.425 13.270 113.125 13.600 ;
        RECT 112.425 1.910 112.565 13.270 ;
        RECT 112.985 2.380 113.125 13.270 ;
        RECT 113.545 13.270 114.245 13.600 ;
        RECT 113.545 1.910 113.685 13.270 ;
        RECT 114.105 2.380 114.245 13.270 ;
        RECT 114.665 13.270 115.365 13.600 ;
        RECT 114.665 1.910 114.805 13.270 ;
        RECT 115.225 2.380 115.365 13.270 ;
        RECT 115.785 13.270 116.485 13.600 ;
        RECT 115.785 1.910 115.925 13.270 ;
        RECT 116.345 2.380 116.485 13.270 ;
        RECT 116.905 13.270 117.605 13.600 ;
        RECT 116.905 1.910 117.045 13.270 ;
        RECT 117.465 2.380 117.605 13.270 ;
        RECT 118.025 13.270 118.725 13.600 ;
        RECT 118.025 1.910 118.165 13.270 ;
        RECT 118.585 2.380 118.725 13.270 ;
        RECT 119.145 13.270 119.845 13.600 ;
        RECT 119.145 1.910 119.285 13.270 ;
        RECT 119.705 2.380 119.845 13.270 ;
        RECT 120.265 13.270 120.965 13.600 ;
        RECT 120.265 1.910 120.405 13.270 ;
        RECT 120.825 2.380 120.965 13.270 ;
        RECT 121.385 13.270 122.715 13.600 ;
        RECT 121.385 2.380 121.525 13.270 ;
        RECT 121.945 2.380 122.085 13.270 ;
        RECT 122.505 2.380 122.715 13.270 ;
        RECT 124.395 13.270 125.095 13.600 ;
        RECT 124.395 1.910 124.535 13.270 ;
        RECT 124.955 2.380 125.095 13.270 ;
        RECT 125.515 13.270 126.215 13.600 ;
        RECT 125.515 1.910 125.655 13.270 ;
        RECT 126.075 2.380 126.215 13.270 ;
        RECT 126.635 13.270 127.335 13.600 ;
        RECT 126.635 1.910 126.775 13.270 ;
        RECT 127.195 2.380 127.335 13.270 ;
        RECT 127.755 13.270 128.455 13.600 ;
        RECT 127.755 1.910 127.895 13.270 ;
        RECT 128.315 2.380 128.455 13.270 ;
        RECT 128.875 13.270 129.575 13.600 ;
        RECT 128.875 1.910 129.015 13.270 ;
        RECT 129.435 2.380 129.575 13.270 ;
        RECT 129.995 13.270 130.695 13.600 ;
        RECT 129.995 1.910 130.135 13.270 ;
        RECT 130.555 2.380 130.695 13.270 ;
        RECT 131.115 13.270 131.815 13.600 ;
        RECT 131.115 1.910 131.255 13.270 ;
        RECT 131.675 2.380 131.815 13.270 ;
        RECT 132.235 13.270 132.935 13.600 ;
        RECT 132.235 1.910 132.375 13.270 ;
        RECT 132.795 2.380 132.935 13.270 ;
        RECT 133.355 13.270 134.055 13.600 ;
        RECT 133.355 1.910 133.495 13.270 ;
        RECT 133.915 2.380 134.055 13.270 ;
        RECT 134.475 13.270 135.805 13.600 ;
        RECT 134.475 2.380 134.615 13.270 ;
        RECT 135.035 2.380 135.175 13.270 ;
        RECT 135.595 2.380 135.805 13.270 ;
        RECT 137.485 13.290 138.185 13.620 ;
        RECT 137.485 1.930 137.625 13.290 ;
        RECT 138.045 2.400 138.185 13.290 ;
        RECT 138.605 13.290 139.305 13.620 ;
        RECT 138.605 1.930 138.745 13.290 ;
        RECT 139.165 2.400 139.305 13.290 ;
        RECT 139.725 13.290 140.425 13.620 ;
        RECT 139.725 1.930 139.865 13.290 ;
        RECT 140.285 2.400 140.425 13.290 ;
        RECT 140.845 13.290 141.545 13.620 ;
        RECT 140.845 1.930 140.985 13.290 ;
        RECT 141.405 2.400 141.545 13.290 ;
        RECT 141.965 13.290 142.665 13.620 ;
        RECT 141.965 1.930 142.105 13.290 ;
        RECT 142.525 2.400 142.665 13.290 ;
        RECT 143.085 13.290 143.785 13.620 ;
        RECT 143.085 1.930 143.225 13.290 ;
        RECT 143.645 2.400 143.785 13.290 ;
        RECT 144.205 13.290 144.905 13.620 ;
        RECT 144.205 1.930 144.345 13.290 ;
        RECT 144.765 2.400 144.905 13.290 ;
        RECT 145.325 13.290 146.025 13.620 ;
        RECT 145.325 1.930 145.465 13.290 ;
        RECT 145.885 2.400 146.025 13.290 ;
        RECT 146.445 13.290 147.145 13.620 ;
        RECT 146.445 1.930 146.585 13.290 ;
        RECT 147.005 2.400 147.145 13.290 ;
        RECT 147.565 13.290 148.895 13.620 ;
        RECT 147.565 2.400 147.705 13.290 ;
        RECT 148.125 2.400 148.265 13.290 ;
        RECT 148.685 2.400 148.895 13.290 ;
        RECT 150.575 13.290 151.275 13.620 ;
        RECT 150.575 1.930 150.715 13.290 ;
        RECT 151.135 2.400 151.275 13.290 ;
        RECT 151.695 13.290 152.395 13.620 ;
        RECT 151.695 1.930 151.835 13.290 ;
        RECT 152.255 2.400 152.395 13.290 ;
        RECT 152.815 13.290 153.515 13.620 ;
        RECT 152.815 1.930 152.955 13.290 ;
        RECT 153.375 2.400 153.515 13.290 ;
        RECT 153.935 13.290 154.635 13.620 ;
        RECT 153.935 1.930 154.075 13.290 ;
        RECT 154.495 2.400 154.635 13.290 ;
        RECT 155.055 13.290 155.755 13.620 ;
        RECT 155.055 1.930 155.195 13.290 ;
        RECT 155.615 2.400 155.755 13.290 ;
        RECT 156.175 13.290 156.875 13.620 ;
        RECT 156.175 1.930 156.315 13.290 ;
        RECT 156.735 2.400 156.875 13.290 ;
        RECT 157.295 13.290 157.995 13.620 ;
        RECT 157.295 1.930 157.435 13.290 ;
        RECT 157.855 2.400 157.995 13.290 ;
        RECT 158.415 13.290 159.115 13.620 ;
        RECT 158.415 1.930 158.555 13.290 ;
        RECT 158.975 2.400 159.115 13.290 ;
        RECT 159.535 13.290 160.235 13.620 ;
        RECT 159.535 1.930 159.675 13.290 ;
        RECT 160.095 2.400 160.235 13.290 ;
        RECT 160.655 13.290 161.985 13.620 ;
        RECT 160.655 2.400 160.795 13.290 ;
        RECT 161.215 2.400 161.355 13.290 ;
        RECT 161.775 2.400 161.985 13.290 ;
      LAYER via2 ;
        RECT 6.365 106.945 6.645 107.225 ;
        RECT 7.485 106.945 7.765 107.225 ;
        RECT 8.605 106.945 8.885 107.225 ;
        RECT 9.725 106.945 10.005 107.225 ;
        RECT 10.845 106.945 11.125 107.225 ;
        RECT 11.965 106.945 12.245 107.225 ;
        RECT 13.085 106.945 13.365 107.225 ;
        RECT 14.205 106.945 14.485 107.225 ;
        RECT 15.325 106.945 15.605 107.225 ;
        RECT 16.445 106.945 16.725 107.225 ;
        RECT 19.455 106.945 19.735 107.225 ;
        RECT 20.575 106.945 20.855 107.225 ;
        RECT 21.695 106.945 21.975 107.225 ;
        RECT 22.815 106.945 23.095 107.225 ;
        RECT 23.935 106.945 24.215 107.225 ;
        RECT 25.055 106.945 25.335 107.225 ;
        RECT 26.175 106.945 26.455 107.225 ;
        RECT 27.295 106.945 27.575 107.225 ;
        RECT 28.415 106.945 28.695 107.225 ;
        RECT 29.535 106.945 29.815 107.225 ;
        RECT 32.545 106.925 32.825 107.205 ;
        RECT 33.665 106.925 33.945 107.205 ;
        RECT 34.785 106.925 35.065 107.205 ;
        RECT 35.905 106.925 36.185 107.205 ;
        RECT 37.025 106.925 37.305 107.205 ;
        RECT 38.145 106.925 38.425 107.205 ;
        RECT 39.265 106.925 39.545 107.205 ;
        RECT 40.385 106.925 40.665 107.205 ;
        RECT 41.505 106.925 41.785 107.205 ;
        RECT 42.625 106.925 42.905 107.205 ;
        RECT 45.635 106.925 45.915 107.205 ;
        RECT 46.755 106.925 47.035 107.205 ;
        RECT 47.875 106.925 48.155 107.205 ;
        RECT 48.995 106.925 49.275 107.205 ;
        RECT 50.115 106.925 50.395 107.205 ;
        RECT 51.235 106.925 51.515 107.205 ;
        RECT 52.355 106.925 52.635 107.205 ;
        RECT 53.475 106.925 53.755 107.205 ;
        RECT 54.595 106.925 54.875 107.205 ;
        RECT 55.715 106.925 55.995 107.205 ;
        RECT 58.685 106.925 58.965 107.205 ;
        RECT 59.805 106.925 60.085 107.205 ;
        RECT 60.925 106.925 61.205 107.205 ;
        RECT 62.045 106.925 62.325 107.205 ;
        RECT 63.165 106.925 63.445 107.205 ;
        RECT 64.285 106.925 64.565 107.205 ;
        RECT 65.405 106.925 65.685 107.205 ;
        RECT 66.525 106.925 66.805 107.205 ;
        RECT 67.645 106.925 67.925 107.205 ;
        RECT 68.765 106.925 69.045 107.205 ;
        RECT 71.775 106.925 72.055 107.205 ;
        RECT 72.895 106.925 73.175 107.205 ;
        RECT 74.015 106.925 74.295 107.205 ;
        RECT 75.135 106.925 75.415 107.205 ;
        RECT 76.255 106.925 76.535 107.205 ;
        RECT 77.375 106.925 77.655 107.205 ;
        RECT 78.495 106.925 78.775 107.205 ;
        RECT 79.615 106.925 79.895 107.205 ;
        RECT 80.735 106.925 81.015 107.205 ;
        RECT 81.855 106.925 82.135 107.205 ;
        RECT 84.865 106.905 85.145 107.185 ;
        RECT 85.985 106.905 86.265 107.185 ;
        RECT 87.105 106.905 87.385 107.185 ;
        RECT 88.225 106.905 88.505 107.185 ;
        RECT 89.345 106.905 89.625 107.185 ;
        RECT 90.465 106.905 90.745 107.185 ;
        RECT 91.585 106.905 91.865 107.185 ;
        RECT 92.705 106.905 92.985 107.185 ;
        RECT 93.825 106.905 94.105 107.185 ;
        RECT 94.945 106.905 95.225 107.185 ;
        RECT 97.955 106.905 98.235 107.185 ;
        RECT 99.075 106.905 99.355 107.185 ;
        RECT 100.195 106.905 100.475 107.185 ;
        RECT 101.315 106.905 101.595 107.185 ;
        RECT 102.435 106.905 102.715 107.185 ;
        RECT 103.555 106.905 103.835 107.185 ;
        RECT 104.675 106.905 104.955 107.185 ;
        RECT 105.795 106.905 106.075 107.185 ;
        RECT 106.915 106.905 107.195 107.185 ;
        RECT 108.035 106.905 108.315 107.185 ;
        RECT 111.045 106.905 111.325 107.185 ;
        RECT 112.165 106.905 112.445 107.185 ;
        RECT 113.285 106.905 113.565 107.185 ;
        RECT 114.405 106.905 114.685 107.185 ;
        RECT 115.525 106.905 115.805 107.185 ;
        RECT 116.645 106.905 116.925 107.185 ;
        RECT 117.765 106.905 118.045 107.185 ;
        RECT 118.885 106.905 119.165 107.185 ;
        RECT 120.005 106.905 120.285 107.185 ;
        RECT 121.125 106.905 121.405 107.185 ;
        RECT 124.135 106.905 124.415 107.185 ;
        RECT 125.255 106.905 125.535 107.185 ;
        RECT 126.375 106.905 126.655 107.185 ;
        RECT 127.495 106.905 127.775 107.185 ;
        RECT 128.615 106.905 128.895 107.185 ;
        RECT 129.735 106.905 130.015 107.185 ;
        RECT 130.855 106.905 131.135 107.185 ;
        RECT 131.975 106.905 132.255 107.185 ;
        RECT 133.095 106.905 133.375 107.185 ;
        RECT 134.215 106.905 134.495 107.185 ;
        RECT 137.225 106.885 137.505 107.165 ;
        RECT 138.345 106.885 138.625 107.165 ;
        RECT 139.465 106.885 139.745 107.165 ;
        RECT 140.585 106.885 140.865 107.165 ;
        RECT 141.705 106.885 141.985 107.165 ;
        RECT 142.825 106.885 143.105 107.165 ;
        RECT 143.945 106.885 144.225 107.165 ;
        RECT 145.065 106.885 145.345 107.165 ;
        RECT 146.185 106.885 146.465 107.165 ;
        RECT 147.305 106.885 147.585 107.165 ;
        RECT 150.315 106.885 150.595 107.165 ;
        RECT 151.435 106.885 151.715 107.165 ;
        RECT 152.555 106.885 152.835 107.165 ;
        RECT 153.675 106.885 153.955 107.165 ;
        RECT 154.795 106.885 155.075 107.165 ;
        RECT 155.915 106.885 156.195 107.165 ;
        RECT 157.035 106.885 157.315 107.165 ;
        RECT 158.155 106.885 158.435 107.165 ;
        RECT 159.275 106.885 159.555 107.165 ;
        RECT 160.395 106.885 160.675 107.165 ;
        RECT 6.395 104.895 6.675 105.175 ;
        RECT 7.515 104.895 7.795 105.175 ;
        RECT 8.635 104.895 8.915 105.175 ;
        RECT 9.755 104.895 10.035 105.175 ;
        RECT 10.875 104.895 11.155 105.175 ;
        RECT 11.995 104.895 12.275 105.175 ;
        RECT 13.115 104.895 13.395 105.175 ;
        RECT 14.235 104.895 14.515 105.175 ;
        RECT 15.355 104.895 15.635 105.175 ;
        RECT 16.475 104.895 16.755 105.175 ;
        RECT 19.485 104.895 19.765 105.175 ;
        RECT 20.605 104.895 20.885 105.175 ;
        RECT 21.725 104.895 22.005 105.175 ;
        RECT 22.845 104.895 23.125 105.175 ;
        RECT 23.965 104.895 24.245 105.175 ;
        RECT 25.085 104.895 25.365 105.175 ;
        RECT 26.205 104.895 26.485 105.175 ;
        RECT 27.325 104.895 27.605 105.175 ;
        RECT 28.445 104.895 28.725 105.175 ;
        RECT 29.565 104.895 29.845 105.175 ;
        RECT 32.575 104.915 32.855 105.195 ;
        RECT 33.695 104.915 33.975 105.195 ;
        RECT 34.815 104.915 35.095 105.195 ;
        RECT 35.935 104.915 36.215 105.195 ;
        RECT 37.055 104.915 37.335 105.195 ;
        RECT 38.175 104.915 38.455 105.195 ;
        RECT 39.295 104.915 39.575 105.195 ;
        RECT 40.415 104.915 40.695 105.195 ;
        RECT 41.535 104.915 41.815 105.195 ;
        RECT 42.655 104.915 42.935 105.195 ;
        RECT 45.665 104.915 45.945 105.195 ;
        RECT 46.785 104.915 47.065 105.195 ;
        RECT 47.905 104.915 48.185 105.195 ;
        RECT 49.025 104.915 49.305 105.195 ;
        RECT 50.145 104.915 50.425 105.195 ;
        RECT 51.265 104.915 51.545 105.195 ;
        RECT 52.385 104.915 52.665 105.195 ;
        RECT 53.505 104.915 53.785 105.195 ;
        RECT 54.625 104.915 54.905 105.195 ;
        RECT 55.745 104.915 56.025 105.195 ;
        RECT 58.715 104.915 58.995 105.195 ;
        RECT 59.835 104.915 60.115 105.195 ;
        RECT 60.955 104.915 61.235 105.195 ;
        RECT 62.075 104.915 62.355 105.195 ;
        RECT 63.195 104.915 63.475 105.195 ;
        RECT 64.315 104.915 64.595 105.195 ;
        RECT 65.435 104.915 65.715 105.195 ;
        RECT 66.555 104.915 66.835 105.195 ;
        RECT 67.675 104.915 67.955 105.195 ;
        RECT 68.795 104.915 69.075 105.195 ;
        RECT 71.805 104.915 72.085 105.195 ;
        RECT 72.925 104.915 73.205 105.195 ;
        RECT 74.045 104.915 74.325 105.195 ;
        RECT 75.165 104.915 75.445 105.195 ;
        RECT 76.285 104.915 76.565 105.195 ;
        RECT 77.405 104.915 77.685 105.195 ;
        RECT 78.525 104.915 78.805 105.195 ;
        RECT 79.645 104.915 79.925 105.195 ;
        RECT 80.765 104.915 81.045 105.195 ;
        RECT 81.885 104.915 82.165 105.195 ;
        RECT 84.895 104.935 85.175 105.215 ;
        RECT 86.015 104.935 86.295 105.215 ;
        RECT 87.135 104.935 87.415 105.215 ;
        RECT 88.255 104.935 88.535 105.215 ;
        RECT 89.375 104.935 89.655 105.215 ;
        RECT 90.495 104.935 90.775 105.215 ;
        RECT 91.615 104.935 91.895 105.215 ;
        RECT 92.735 104.935 93.015 105.215 ;
        RECT 93.855 104.935 94.135 105.215 ;
        RECT 94.975 104.935 95.255 105.215 ;
        RECT 97.985 104.935 98.265 105.215 ;
        RECT 99.105 104.935 99.385 105.215 ;
        RECT 100.225 104.935 100.505 105.215 ;
        RECT 101.345 104.935 101.625 105.215 ;
        RECT 102.465 104.935 102.745 105.215 ;
        RECT 103.585 104.935 103.865 105.215 ;
        RECT 104.705 104.935 104.985 105.215 ;
        RECT 105.825 104.935 106.105 105.215 ;
        RECT 106.945 104.935 107.225 105.215 ;
        RECT 108.065 104.935 108.345 105.215 ;
        RECT 111.075 104.935 111.355 105.215 ;
        RECT 112.195 104.935 112.475 105.215 ;
        RECT 113.315 104.935 113.595 105.215 ;
        RECT 114.435 104.935 114.715 105.215 ;
        RECT 115.555 104.935 115.835 105.215 ;
        RECT 116.675 104.935 116.955 105.215 ;
        RECT 117.795 104.935 118.075 105.215 ;
        RECT 118.915 104.935 119.195 105.215 ;
        RECT 120.035 104.935 120.315 105.215 ;
        RECT 121.155 104.935 121.435 105.215 ;
        RECT 124.165 104.935 124.445 105.215 ;
        RECT 125.285 104.935 125.565 105.215 ;
        RECT 126.405 104.935 126.685 105.215 ;
        RECT 127.525 104.935 127.805 105.215 ;
        RECT 128.645 104.935 128.925 105.215 ;
        RECT 129.765 104.935 130.045 105.215 ;
        RECT 130.885 104.935 131.165 105.215 ;
        RECT 132.005 104.935 132.285 105.215 ;
        RECT 133.125 104.935 133.405 105.215 ;
        RECT 134.245 104.935 134.525 105.215 ;
        RECT 137.255 104.955 137.535 105.235 ;
        RECT 138.375 104.955 138.655 105.235 ;
        RECT 139.495 104.955 139.775 105.235 ;
        RECT 140.615 104.955 140.895 105.235 ;
        RECT 141.735 104.955 142.015 105.235 ;
        RECT 142.855 104.955 143.135 105.235 ;
        RECT 143.975 104.955 144.255 105.235 ;
        RECT 145.095 104.955 145.375 105.235 ;
        RECT 146.215 104.955 146.495 105.235 ;
        RECT 147.335 104.955 147.615 105.235 ;
        RECT 150.345 104.955 150.625 105.235 ;
        RECT 151.465 104.955 151.745 105.235 ;
        RECT 152.585 104.955 152.865 105.235 ;
        RECT 153.705 104.955 153.985 105.235 ;
        RECT 154.825 104.955 155.105 105.235 ;
        RECT 155.945 104.955 156.225 105.235 ;
        RECT 157.065 104.955 157.345 105.235 ;
        RECT 158.185 104.955 158.465 105.235 ;
        RECT 159.305 104.955 159.585 105.235 ;
        RECT 160.425 104.955 160.705 105.235 ;
        RECT 162.875 90.270 163.350 90.745 ;
        RECT 4.760 88.675 5.230 89.145 ;
        RECT 4.750 33.215 5.220 33.685 ;
        RECT 163.275 29.215 163.750 29.690 ;
        RECT 6.805 15.305 7.085 15.585 ;
        RECT 7.925 15.305 8.205 15.585 ;
        RECT 9.045 15.305 9.325 15.585 ;
        RECT 10.165 15.305 10.445 15.585 ;
        RECT 11.285 15.305 11.565 15.585 ;
        RECT 12.405 15.305 12.685 15.585 ;
        RECT 13.525 15.305 13.805 15.585 ;
        RECT 14.645 15.305 14.925 15.585 ;
        RECT 15.765 15.305 16.045 15.585 ;
        RECT 16.885 15.305 17.165 15.585 ;
        RECT 19.895 15.305 20.175 15.585 ;
        RECT 21.015 15.305 21.295 15.585 ;
        RECT 22.135 15.305 22.415 15.585 ;
        RECT 23.255 15.305 23.535 15.585 ;
        RECT 24.375 15.305 24.655 15.585 ;
        RECT 25.495 15.305 25.775 15.585 ;
        RECT 26.615 15.305 26.895 15.585 ;
        RECT 27.735 15.305 28.015 15.585 ;
        RECT 28.855 15.305 29.135 15.585 ;
        RECT 29.975 15.305 30.255 15.585 ;
        RECT 32.985 15.285 33.265 15.565 ;
        RECT 34.105 15.285 34.385 15.565 ;
        RECT 35.225 15.285 35.505 15.565 ;
        RECT 36.345 15.285 36.625 15.565 ;
        RECT 37.465 15.285 37.745 15.565 ;
        RECT 38.585 15.285 38.865 15.565 ;
        RECT 39.705 15.285 39.985 15.565 ;
        RECT 40.825 15.285 41.105 15.565 ;
        RECT 41.945 15.285 42.225 15.565 ;
        RECT 43.065 15.285 43.345 15.565 ;
        RECT 46.075 15.285 46.355 15.565 ;
        RECT 47.195 15.285 47.475 15.565 ;
        RECT 48.315 15.285 48.595 15.565 ;
        RECT 49.435 15.285 49.715 15.565 ;
        RECT 50.555 15.285 50.835 15.565 ;
        RECT 51.675 15.285 51.955 15.565 ;
        RECT 52.795 15.285 53.075 15.565 ;
        RECT 53.915 15.285 54.195 15.565 ;
        RECT 55.035 15.285 55.315 15.565 ;
        RECT 56.155 15.285 56.435 15.565 ;
        RECT 59.125 15.285 59.405 15.565 ;
        RECT 60.245 15.285 60.525 15.565 ;
        RECT 61.365 15.285 61.645 15.565 ;
        RECT 62.485 15.285 62.765 15.565 ;
        RECT 63.605 15.285 63.885 15.565 ;
        RECT 64.725 15.285 65.005 15.565 ;
        RECT 65.845 15.285 66.125 15.565 ;
        RECT 66.965 15.285 67.245 15.565 ;
        RECT 68.085 15.285 68.365 15.565 ;
        RECT 69.205 15.285 69.485 15.565 ;
        RECT 72.215 15.285 72.495 15.565 ;
        RECT 73.335 15.285 73.615 15.565 ;
        RECT 74.455 15.285 74.735 15.565 ;
        RECT 75.575 15.285 75.855 15.565 ;
        RECT 76.695 15.285 76.975 15.565 ;
        RECT 77.815 15.285 78.095 15.565 ;
        RECT 78.935 15.285 79.215 15.565 ;
        RECT 80.055 15.285 80.335 15.565 ;
        RECT 81.175 15.285 81.455 15.565 ;
        RECT 82.295 15.285 82.575 15.565 ;
        RECT 85.305 15.265 85.585 15.545 ;
        RECT 86.425 15.265 86.705 15.545 ;
        RECT 87.545 15.265 87.825 15.545 ;
        RECT 88.665 15.265 88.945 15.545 ;
        RECT 89.785 15.265 90.065 15.545 ;
        RECT 90.905 15.265 91.185 15.545 ;
        RECT 92.025 15.265 92.305 15.545 ;
        RECT 93.145 15.265 93.425 15.545 ;
        RECT 94.265 15.265 94.545 15.545 ;
        RECT 95.385 15.265 95.665 15.545 ;
        RECT 98.395 15.265 98.675 15.545 ;
        RECT 99.515 15.265 99.795 15.545 ;
        RECT 100.635 15.265 100.915 15.545 ;
        RECT 101.755 15.265 102.035 15.545 ;
        RECT 102.875 15.265 103.155 15.545 ;
        RECT 103.995 15.265 104.275 15.545 ;
        RECT 105.115 15.265 105.395 15.545 ;
        RECT 106.235 15.265 106.515 15.545 ;
        RECT 107.355 15.265 107.635 15.545 ;
        RECT 108.475 15.265 108.755 15.545 ;
        RECT 111.485 15.265 111.765 15.545 ;
        RECT 112.605 15.265 112.885 15.545 ;
        RECT 113.725 15.265 114.005 15.545 ;
        RECT 114.845 15.265 115.125 15.545 ;
        RECT 115.965 15.265 116.245 15.545 ;
        RECT 117.085 15.265 117.365 15.545 ;
        RECT 118.205 15.265 118.485 15.545 ;
        RECT 119.325 15.265 119.605 15.545 ;
        RECT 120.445 15.265 120.725 15.545 ;
        RECT 121.565 15.265 121.845 15.545 ;
        RECT 124.575 15.265 124.855 15.545 ;
        RECT 125.695 15.265 125.975 15.545 ;
        RECT 126.815 15.265 127.095 15.545 ;
        RECT 127.935 15.265 128.215 15.545 ;
        RECT 129.055 15.265 129.335 15.545 ;
        RECT 130.175 15.265 130.455 15.545 ;
        RECT 131.295 15.265 131.575 15.545 ;
        RECT 132.415 15.265 132.695 15.545 ;
        RECT 133.535 15.265 133.815 15.545 ;
        RECT 134.655 15.265 134.935 15.545 ;
        RECT 137.665 15.245 137.945 15.525 ;
        RECT 138.785 15.245 139.065 15.525 ;
        RECT 139.905 15.245 140.185 15.525 ;
        RECT 141.025 15.245 141.305 15.525 ;
        RECT 142.145 15.245 142.425 15.525 ;
        RECT 143.265 15.245 143.545 15.525 ;
        RECT 144.385 15.245 144.665 15.525 ;
        RECT 145.505 15.245 145.785 15.525 ;
        RECT 146.625 15.245 146.905 15.525 ;
        RECT 147.745 15.245 148.025 15.525 ;
        RECT 150.755 15.245 151.035 15.525 ;
        RECT 151.875 15.245 152.155 15.525 ;
        RECT 152.995 15.245 153.275 15.525 ;
        RECT 154.115 15.245 154.395 15.525 ;
        RECT 155.235 15.245 155.515 15.525 ;
        RECT 156.355 15.245 156.635 15.525 ;
        RECT 157.475 15.245 157.755 15.525 ;
        RECT 158.595 15.245 158.875 15.525 ;
        RECT 159.715 15.245 159.995 15.525 ;
        RECT 160.835 15.245 161.115 15.525 ;
        RECT 6.835 13.255 7.115 13.535 ;
        RECT 7.955 13.255 8.235 13.535 ;
        RECT 9.075 13.255 9.355 13.535 ;
        RECT 10.195 13.255 10.475 13.535 ;
        RECT 11.315 13.255 11.595 13.535 ;
        RECT 12.435 13.255 12.715 13.535 ;
        RECT 13.555 13.255 13.835 13.535 ;
        RECT 14.675 13.255 14.955 13.535 ;
        RECT 15.795 13.255 16.075 13.535 ;
        RECT 16.915 13.255 17.195 13.535 ;
        RECT 19.925 13.255 20.205 13.535 ;
        RECT 21.045 13.255 21.325 13.535 ;
        RECT 22.165 13.255 22.445 13.535 ;
        RECT 23.285 13.255 23.565 13.535 ;
        RECT 24.405 13.255 24.685 13.535 ;
        RECT 25.525 13.255 25.805 13.535 ;
        RECT 26.645 13.255 26.925 13.535 ;
        RECT 27.765 13.255 28.045 13.535 ;
        RECT 28.885 13.255 29.165 13.535 ;
        RECT 30.005 13.255 30.285 13.535 ;
        RECT 33.015 13.275 33.295 13.555 ;
        RECT 34.135 13.275 34.415 13.555 ;
        RECT 35.255 13.275 35.535 13.555 ;
        RECT 36.375 13.275 36.655 13.555 ;
        RECT 37.495 13.275 37.775 13.555 ;
        RECT 38.615 13.275 38.895 13.555 ;
        RECT 39.735 13.275 40.015 13.555 ;
        RECT 40.855 13.275 41.135 13.555 ;
        RECT 41.975 13.275 42.255 13.555 ;
        RECT 43.095 13.275 43.375 13.555 ;
        RECT 46.105 13.275 46.385 13.555 ;
        RECT 47.225 13.275 47.505 13.555 ;
        RECT 48.345 13.275 48.625 13.555 ;
        RECT 49.465 13.275 49.745 13.555 ;
        RECT 50.585 13.275 50.865 13.555 ;
        RECT 51.705 13.275 51.985 13.555 ;
        RECT 52.825 13.275 53.105 13.555 ;
        RECT 53.945 13.275 54.225 13.555 ;
        RECT 55.065 13.275 55.345 13.555 ;
        RECT 56.185 13.275 56.465 13.555 ;
        RECT 59.155 13.275 59.435 13.555 ;
        RECT 60.275 13.275 60.555 13.555 ;
        RECT 61.395 13.275 61.675 13.555 ;
        RECT 62.515 13.275 62.795 13.555 ;
        RECT 63.635 13.275 63.915 13.555 ;
        RECT 64.755 13.275 65.035 13.555 ;
        RECT 65.875 13.275 66.155 13.555 ;
        RECT 66.995 13.275 67.275 13.555 ;
        RECT 68.115 13.275 68.395 13.555 ;
        RECT 69.235 13.275 69.515 13.555 ;
        RECT 72.245 13.275 72.525 13.555 ;
        RECT 73.365 13.275 73.645 13.555 ;
        RECT 74.485 13.275 74.765 13.555 ;
        RECT 75.605 13.275 75.885 13.555 ;
        RECT 76.725 13.275 77.005 13.555 ;
        RECT 77.845 13.275 78.125 13.555 ;
        RECT 78.965 13.275 79.245 13.555 ;
        RECT 80.085 13.275 80.365 13.555 ;
        RECT 81.205 13.275 81.485 13.555 ;
        RECT 82.325 13.275 82.605 13.555 ;
        RECT 85.335 13.295 85.615 13.575 ;
        RECT 86.455 13.295 86.735 13.575 ;
        RECT 87.575 13.295 87.855 13.575 ;
        RECT 88.695 13.295 88.975 13.575 ;
        RECT 89.815 13.295 90.095 13.575 ;
        RECT 90.935 13.295 91.215 13.575 ;
        RECT 92.055 13.295 92.335 13.575 ;
        RECT 93.175 13.295 93.455 13.575 ;
        RECT 94.295 13.295 94.575 13.575 ;
        RECT 95.415 13.295 95.695 13.575 ;
        RECT 98.425 13.295 98.705 13.575 ;
        RECT 99.545 13.295 99.825 13.575 ;
        RECT 100.665 13.295 100.945 13.575 ;
        RECT 101.785 13.295 102.065 13.575 ;
        RECT 102.905 13.295 103.185 13.575 ;
        RECT 104.025 13.295 104.305 13.575 ;
        RECT 105.145 13.295 105.425 13.575 ;
        RECT 106.265 13.295 106.545 13.575 ;
        RECT 107.385 13.295 107.665 13.575 ;
        RECT 108.505 13.295 108.785 13.575 ;
        RECT 111.515 13.295 111.795 13.575 ;
        RECT 112.635 13.295 112.915 13.575 ;
        RECT 113.755 13.295 114.035 13.575 ;
        RECT 114.875 13.295 115.155 13.575 ;
        RECT 115.995 13.295 116.275 13.575 ;
        RECT 117.115 13.295 117.395 13.575 ;
        RECT 118.235 13.295 118.515 13.575 ;
        RECT 119.355 13.295 119.635 13.575 ;
        RECT 120.475 13.295 120.755 13.575 ;
        RECT 121.595 13.295 121.875 13.575 ;
        RECT 124.605 13.295 124.885 13.575 ;
        RECT 125.725 13.295 126.005 13.575 ;
        RECT 126.845 13.295 127.125 13.575 ;
        RECT 127.965 13.295 128.245 13.575 ;
        RECT 129.085 13.295 129.365 13.575 ;
        RECT 130.205 13.295 130.485 13.575 ;
        RECT 131.325 13.295 131.605 13.575 ;
        RECT 132.445 13.295 132.725 13.575 ;
        RECT 133.565 13.295 133.845 13.575 ;
        RECT 134.685 13.295 134.965 13.575 ;
        RECT 137.695 13.315 137.975 13.595 ;
        RECT 138.815 13.315 139.095 13.595 ;
        RECT 139.935 13.315 140.215 13.595 ;
        RECT 141.055 13.315 141.335 13.595 ;
        RECT 142.175 13.315 142.455 13.595 ;
        RECT 143.295 13.315 143.575 13.595 ;
        RECT 144.415 13.315 144.695 13.595 ;
        RECT 145.535 13.315 145.815 13.595 ;
        RECT 146.655 13.315 146.935 13.595 ;
        RECT 147.775 13.315 148.055 13.595 ;
        RECT 150.785 13.315 151.065 13.595 ;
        RECT 151.905 13.315 152.185 13.595 ;
        RECT 153.025 13.315 153.305 13.595 ;
        RECT 154.145 13.315 154.425 13.595 ;
        RECT 155.265 13.315 155.545 13.595 ;
        RECT 156.385 13.315 156.665 13.595 ;
        RECT 157.505 13.315 157.785 13.595 ;
        RECT 158.625 13.315 158.905 13.595 ;
        RECT 159.745 13.315 160.025 13.595 ;
        RECT 160.865 13.315 161.145 13.595 ;
      LAYER met3 ;
        RECT 6.755 107.250 7.055 117.980 ;
        RECT 7.955 107.250 8.255 117.980 ;
        RECT 9.155 107.250 9.455 117.980 ;
        RECT 10.355 107.250 10.655 117.980 ;
        RECT 11.555 107.250 11.855 117.980 ;
        RECT 12.755 107.250 13.055 117.980 ;
        RECT 13.955 107.250 14.255 117.980 ;
        RECT 15.155 107.250 15.455 117.980 ;
        RECT 16.355 107.250 16.655 117.980 ;
        RECT 19.845 107.250 20.145 117.980 ;
        RECT 21.045 107.250 21.345 117.980 ;
        RECT 22.245 107.250 22.545 117.980 ;
        RECT 23.445 107.250 23.745 117.980 ;
        RECT 24.645 107.250 24.945 117.980 ;
        RECT 25.845 107.250 26.145 117.980 ;
        RECT 27.045 107.250 27.345 117.980 ;
        RECT 28.245 107.250 28.545 117.980 ;
        RECT 29.445 107.250 29.745 117.980 ;
        RECT 6.155 106.920 17.565 107.250 ;
        RECT 19.245 106.920 30.655 107.250 ;
        RECT 32.935 107.230 33.235 117.960 ;
        RECT 34.135 107.230 34.435 117.960 ;
        RECT 35.335 107.230 35.635 117.960 ;
        RECT 36.535 107.230 36.835 117.960 ;
        RECT 37.735 107.230 38.035 117.960 ;
        RECT 38.935 107.230 39.235 117.960 ;
        RECT 40.135 107.230 40.435 117.960 ;
        RECT 41.335 107.230 41.635 117.960 ;
        RECT 42.535 107.230 42.835 117.960 ;
        RECT 46.025 107.230 46.325 117.960 ;
        RECT 47.225 107.230 47.525 117.960 ;
        RECT 48.425 107.230 48.725 117.960 ;
        RECT 49.625 107.230 49.925 117.960 ;
        RECT 50.825 107.230 51.125 117.960 ;
        RECT 52.025 107.230 52.325 117.960 ;
        RECT 53.225 107.230 53.525 117.960 ;
        RECT 54.425 107.230 54.725 117.960 ;
        RECT 55.625 107.230 55.925 117.960 ;
        RECT 59.075 107.230 59.375 117.960 ;
        RECT 60.275 107.230 60.575 117.960 ;
        RECT 61.475 107.230 61.775 117.960 ;
        RECT 62.675 107.230 62.975 117.960 ;
        RECT 63.875 107.230 64.175 117.960 ;
        RECT 65.075 107.230 65.375 117.960 ;
        RECT 66.275 107.230 66.575 117.960 ;
        RECT 67.475 107.230 67.775 117.960 ;
        RECT 68.675 107.230 68.975 117.960 ;
        RECT 72.165 107.230 72.465 117.960 ;
        RECT 73.365 107.230 73.665 117.960 ;
        RECT 74.565 107.230 74.865 117.960 ;
        RECT 75.765 107.230 76.065 117.960 ;
        RECT 76.965 107.230 77.265 117.960 ;
        RECT 78.165 107.230 78.465 117.960 ;
        RECT 79.365 107.230 79.665 117.960 ;
        RECT 80.565 107.230 80.865 117.960 ;
        RECT 81.765 107.230 82.065 117.960 ;
        RECT 32.335 106.900 43.745 107.230 ;
        RECT 45.425 106.900 56.835 107.230 ;
        RECT 58.475 106.900 69.885 107.230 ;
        RECT 71.565 106.900 82.975 107.230 ;
        RECT 85.255 107.210 85.555 117.940 ;
        RECT 86.455 107.210 86.755 117.940 ;
        RECT 87.655 107.210 87.955 117.940 ;
        RECT 88.855 107.210 89.155 117.940 ;
        RECT 90.055 107.210 90.355 117.940 ;
        RECT 91.255 107.210 91.555 117.940 ;
        RECT 92.455 107.210 92.755 117.940 ;
        RECT 93.655 107.210 93.955 117.940 ;
        RECT 94.855 107.210 95.155 117.940 ;
        RECT 98.345 107.210 98.645 117.940 ;
        RECT 99.545 107.210 99.845 117.940 ;
        RECT 100.745 107.210 101.045 117.940 ;
        RECT 101.945 107.210 102.245 117.940 ;
        RECT 103.145 107.210 103.445 117.940 ;
        RECT 104.345 107.210 104.645 117.940 ;
        RECT 105.545 107.210 105.845 117.940 ;
        RECT 106.745 107.210 107.045 117.940 ;
        RECT 107.945 107.210 108.245 117.940 ;
        RECT 111.435 107.210 111.735 117.940 ;
        RECT 112.635 107.210 112.935 117.940 ;
        RECT 113.835 107.210 114.135 117.940 ;
        RECT 115.035 107.210 115.335 117.940 ;
        RECT 116.235 107.210 116.535 117.940 ;
        RECT 117.435 107.210 117.735 117.940 ;
        RECT 118.635 107.210 118.935 117.940 ;
        RECT 119.835 107.210 120.135 117.940 ;
        RECT 121.035 107.210 121.335 117.940 ;
        RECT 124.525 107.210 124.825 117.940 ;
        RECT 125.725 107.210 126.025 117.940 ;
        RECT 126.925 107.210 127.225 117.940 ;
        RECT 128.125 107.210 128.425 117.940 ;
        RECT 129.325 107.210 129.625 117.940 ;
        RECT 130.525 107.210 130.825 117.940 ;
        RECT 131.725 107.210 132.025 117.940 ;
        RECT 132.925 107.210 133.225 117.940 ;
        RECT 134.125 107.210 134.425 117.940 ;
        RECT 84.655 106.880 96.065 107.210 ;
        RECT 97.745 106.880 109.155 107.210 ;
        RECT 110.835 106.880 122.245 107.210 ;
        RECT 123.925 106.880 135.335 107.210 ;
        RECT 137.615 107.190 137.915 117.920 ;
        RECT 138.815 107.190 139.115 117.920 ;
        RECT 140.015 107.190 140.315 117.920 ;
        RECT 141.215 107.190 141.515 117.920 ;
        RECT 142.415 107.190 142.715 117.920 ;
        RECT 143.615 107.190 143.915 117.920 ;
        RECT 144.815 107.190 145.115 117.920 ;
        RECT 146.015 107.190 146.315 117.920 ;
        RECT 147.215 107.190 147.515 117.920 ;
        RECT 150.705 107.190 151.005 117.920 ;
        RECT 151.905 107.190 152.205 117.920 ;
        RECT 153.105 107.190 153.405 117.920 ;
        RECT 154.305 107.190 154.605 117.920 ;
        RECT 155.505 107.190 155.805 117.920 ;
        RECT 156.705 107.190 157.005 117.920 ;
        RECT 157.905 107.190 158.205 117.920 ;
        RECT 159.105 107.190 159.405 117.920 ;
        RECT 160.305 107.190 160.605 117.920 ;
        RECT 137.015 106.860 148.425 107.190 ;
        RECT 150.105 106.860 161.515 107.190 ;
        RECT 6.185 104.870 17.595 105.200 ;
        RECT 19.275 104.870 30.685 105.200 ;
        RECT 32.365 104.890 43.775 105.220 ;
        RECT 45.455 104.890 56.865 105.220 ;
        RECT 58.505 104.890 69.915 105.220 ;
        RECT 71.595 104.890 83.005 105.220 ;
        RECT 84.685 104.910 96.095 105.240 ;
        RECT 97.775 104.910 109.185 105.240 ;
        RECT 110.865 104.910 122.275 105.240 ;
        RECT 123.955 104.910 135.365 105.240 ;
        RECT 137.045 104.930 148.455 105.260 ;
        RECT 150.135 104.930 161.545 105.260 ;
        RECT 6.785 94.140 7.085 104.870 ;
        RECT 7.985 94.140 8.285 104.870 ;
        RECT 9.185 94.140 9.485 104.870 ;
        RECT 10.385 94.140 10.685 104.870 ;
        RECT 11.585 94.140 11.885 104.870 ;
        RECT 12.785 94.140 13.085 104.870 ;
        RECT 13.985 94.140 14.285 104.870 ;
        RECT 15.185 94.140 15.485 104.870 ;
        RECT 16.385 94.140 16.685 104.870 ;
        RECT 19.875 94.140 20.175 104.870 ;
        RECT 21.075 94.140 21.375 104.870 ;
        RECT 22.275 94.140 22.575 104.870 ;
        RECT 23.475 94.140 23.775 104.870 ;
        RECT 24.675 94.140 24.975 104.870 ;
        RECT 25.875 94.140 26.175 104.870 ;
        RECT 27.075 94.140 27.375 104.870 ;
        RECT 28.275 94.140 28.575 104.870 ;
        RECT 29.475 94.140 29.775 104.870 ;
        RECT 32.965 94.160 33.265 104.890 ;
        RECT 34.165 94.160 34.465 104.890 ;
        RECT 35.365 94.160 35.665 104.890 ;
        RECT 36.565 94.160 36.865 104.890 ;
        RECT 37.765 94.160 38.065 104.890 ;
        RECT 38.965 94.160 39.265 104.890 ;
        RECT 40.165 94.160 40.465 104.890 ;
        RECT 41.365 94.160 41.665 104.890 ;
        RECT 42.565 94.160 42.865 104.890 ;
        RECT 46.055 94.160 46.355 104.890 ;
        RECT 47.255 94.160 47.555 104.890 ;
        RECT 48.455 94.160 48.755 104.890 ;
        RECT 49.655 94.160 49.955 104.890 ;
        RECT 50.855 94.160 51.155 104.890 ;
        RECT 52.055 94.160 52.355 104.890 ;
        RECT 53.255 94.160 53.555 104.890 ;
        RECT 54.455 94.160 54.755 104.890 ;
        RECT 55.655 94.160 55.955 104.890 ;
        RECT 59.105 94.160 59.405 104.890 ;
        RECT 60.305 94.160 60.605 104.890 ;
        RECT 61.505 94.160 61.805 104.890 ;
        RECT 62.705 94.160 63.005 104.890 ;
        RECT 63.905 94.160 64.205 104.890 ;
        RECT 65.105 94.160 65.405 104.890 ;
        RECT 66.305 94.160 66.605 104.890 ;
        RECT 67.505 94.160 67.805 104.890 ;
        RECT 68.705 94.160 69.005 104.890 ;
        RECT 72.195 94.160 72.495 104.890 ;
        RECT 73.395 94.160 73.695 104.890 ;
        RECT 74.595 94.160 74.895 104.890 ;
        RECT 75.795 94.160 76.095 104.890 ;
        RECT 76.995 94.160 77.295 104.890 ;
        RECT 78.195 94.160 78.495 104.890 ;
        RECT 79.395 94.160 79.695 104.890 ;
        RECT 80.595 94.160 80.895 104.890 ;
        RECT 81.795 94.160 82.095 104.890 ;
        RECT 85.285 94.180 85.585 104.910 ;
        RECT 86.485 94.180 86.785 104.910 ;
        RECT 87.685 94.180 87.985 104.910 ;
        RECT 88.885 94.180 89.185 104.910 ;
        RECT 90.085 94.180 90.385 104.910 ;
        RECT 91.285 94.180 91.585 104.910 ;
        RECT 92.485 94.180 92.785 104.910 ;
        RECT 93.685 94.180 93.985 104.910 ;
        RECT 94.885 94.180 95.185 104.910 ;
        RECT 98.375 94.180 98.675 104.910 ;
        RECT 99.575 94.180 99.875 104.910 ;
        RECT 100.775 94.180 101.075 104.910 ;
        RECT 101.975 94.180 102.275 104.910 ;
        RECT 103.175 94.180 103.475 104.910 ;
        RECT 104.375 94.180 104.675 104.910 ;
        RECT 105.575 94.180 105.875 104.910 ;
        RECT 106.775 94.180 107.075 104.910 ;
        RECT 107.975 94.180 108.275 104.910 ;
        RECT 111.465 94.180 111.765 104.910 ;
        RECT 112.665 94.180 112.965 104.910 ;
        RECT 113.865 94.180 114.165 104.910 ;
        RECT 115.065 94.180 115.365 104.910 ;
        RECT 116.265 94.180 116.565 104.910 ;
        RECT 117.465 94.180 117.765 104.910 ;
        RECT 118.665 94.180 118.965 104.910 ;
        RECT 119.865 94.180 120.165 104.910 ;
        RECT 121.065 94.180 121.365 104.910 ;
        RECT 124.555 94.180 124.855 104.910 ;
        RECT 125.755 94.180 126.055 104.910 ;
        RECT 126.955 94.180 127.255 104.910 ;
        RECT 128.155 94.180 128.455 104.910 ;
        RECT 129.355 94.180 129.655 104.910 ;
        RECT 130.555 94.180 130.855 104.910 ;
        RECT 131.755 94.180 132.055 104.910 ;
        RECT 132.955 94.180 133.255 104.910 ;
        RECT 134.155 94.180 134.455 104.910 ;
        RECT 137.645 94.200 137.945 104.930 ;
        RECT 138.845 94.200 139.145 104.930 ;
        RECT 140.045 94.200 140.345 104.930 ;
        RECT 141.245 94.200 141.545 104.930 ;
        RECT 142.445 94.200 142.745 104.930 ;
        RECT 143.645 94.200 143.945 104.930 ;
        RECT 144.845 94.200 145.145 104.930 ;
        RECT 146.045 94.200 146.345 104.930 ;
        RECT 147.245 94.200 147.545 104.930 ;
        RECT 150.735 94.200 151.035 104.930 ;
        RECT 151.935 94.200 152.235 104.930 ;
        RECT 153.135 94.200 153.435 104.930 ;
        RECT 154.335 94.200 154.635 104.930 ;
        RECT 155.535 94.200 155.835 104.930 ;
        RECT 156.735 94.200 157.035 104.930 ;
        RECT 157.935 94.200 158.235 104.930 ;
        RECT 159.135 94.200 159.435 104.930 ;
        RECT 160.335 94.200 160.635 104.930 ;
        RECT 162.850 90.245 163.405 90.770 ;
        RECT 4.735 88.650 5.255 89.200 ;
        RECT 4.725 33.160 5.245 33.710 ;
        RECT 163.250 29.190 163.775 29.745 ;
        RECT 7.195 15.610 7.495 26.340 ;
        RECT 8.395 15.610 8.695 26.340 ;
        RECT 9.595 15.610 9.895 26.340 ;
        RECT 10.795 15.610 11.095 26.340 ;
        RECT 11.995 15.610 12.295 26.340 ;
        RECT 13.195 15.610 13.495 26.340 ;
        RECT 14.395 15.610 14.695 26.340 ;
        RECT 15.595 15.610 15.895 26.340 ;
        RECT 16.795 15.610 17.095 26.340 ;
        RECT 20.285 15.610 20.585 26.340 ;
        RECT 21.485 15.610 21.785 26.340 ;
        RECT 22.685 15.610 22.985 26.340 ;
        RECT 23.885 15.610 24.185 26.340 ;
        RECT 25.085 15.610 25.385 26.340 ;
        RECT 26.285 15.610 26.585 26.340 ;
        RECT 27.485 15.610 27.785 26.340 ;
        RECT 28.685 15.610 28.985 26.340 ;
        RECT 29.885 15.610 30.185 26.340 ;
        RECT 6.595 15.280 18.005 15.610 ;
        RECT 19.685 15.280 31.095 15.610 ;
        RECT 33.375 15.590 33.675 26.320 ;
        RECT 34.575 15.590 34.875 26.320 ;
        RECT 35.775 15.590 36.075 26.320 ;
        RECT 36.975 15.590 37.275 26.320 ;
        RECT 38.175 15.590 38.475 26.320 ;
        RECT 39.375 15.590 39.675 26.320 ;
        RECT 40.575 15.590 40.875 26.320 ;
        RECT 41.775 15.590 42.075 26.320 ;
        RECT 42.975 15.590 43.275 26.320 ;
        RECT 46.465 15.590 46.765 26.320 ;
        RECT 47.665 15.590 47.965 26.320 ;
        RECT 48.865 15.590 49.165 26.320 ;
        RECT 50.065 15.590 50.365 26.320 ;
        RECT 51.265 15.590 51.565 26.320 ;
        RECT 52.465 15.590 52.765 26.320 ;
        RECT 53.665 15.590 53.965 26.320 ;
        RECT 54.865 15.590 55.165 26.320 ;
        RECT 56.065 15.590 56.365 26.320 ;
        RECT 59.515 15.590 59.815 26.320 ;
        RECT 60.715 15.590 61.015 26.320 ;
        RECT 61.915 15.590 62.215 26.320 ;
        RECT 63.115 15.590 63.415 26.320 ;
        RECT 64.315 15.590 64.615 26.320 ;
        RECT 65.515 15.590 65.815 26.320 ;
        RECT 66.715 15.590 67.015 26.320 ;
        RECT 67.915 15.590 68.215 26.320 ;
        RECT 69.115 15.590 69.415 26.320 ;
        RECT 72.605 15.590 72.905 26.320 ;
        RECT 73.805 15.590 74.105 26.320 ;
        RECT 75.005 15.590 75.305 26.320 ;
        RECT 76.205 15.590 76.505 26.320 ;
        RECT 77.405 15.590 77.705 26.320 ;
        RECT 78.605 15.590 78.905 26.320 ;
        RECT 79.805 15.590 80.105 26.320 ;
        RECT 81.005 15.590 81.305 26.320 ;
        RECT 82.205 15.590 82.505 26.320 ;
        RECT 32.775 15.260 44.185 15.590 ;
        RECT 45.865 15.260 57.275 15.590 ;
        RECT 58.915 15.260 70.325 15.590 ;
        RECT 72.005 15.260 83.415 15.590 ;
        RECT 85.695 15.570 85.995 26.300 ;
        RECT 86.895 15.570 87.195 26.300 ;
        RECT 88.095 15.570 88.395 26.300 ;
        RECT 89.295 15.570 89.595 26.300 ;
        RECT 90.495 15.570 90.795 26.300 ;
        RECT 91.695 15.570 91.995 26.300 ;
        RECT 92.895 15.570 93.195 26.300 ;
        RECT 94.095 15.570 94.395 26.300 ;
        RECT 95.295 15.570 95.595 26.300 ;
        RECT 98.785 15.570 99.085 26.300 ;
        RECT 99.985 15.570 100.285 26.300 ;
        RECT 101.185 15.570 101.485 26.300 ;
        RECT 102.385 15.570 102.685 26.300 ;
        RECT 103.585 15.570 103.885 26.300 ;
        RECT 104.785 15.570 105.085 26.300 ;
        RECT 105.985 15.570 106.285 26.300 ;
        RECT 107.185 15.570 107.485 26.300 ;
        RECT 108.385 15.570 108.685 26.300 ;
        RECT 111.875 15.570 112.175 26.300 ;
        RECT 113.075 15.570 113.375 26.300 ;
        RECT 114.275 15.570 114.575 26.300 ;
        RECT 115.475 15.570 115.775 26.300 ;
        RECT 116.675 15.570 116.975 26.300 ;
        RECT 117.875 15.570 118.175 26.300 ;
        RECT 119.075 15.570 119.375 26.300 ;
        RECT 120.275 15.570 120.575 26.300 ;
        RECT 121.475 15.570 121.775 26.300 ;
        RECT 124.965 15.570 125.265 26.300 ;
        RECT 126.165 15.570 126.465 26.300 ;
        RECT 127.365 15.570 127.665 26.300 ;
        RECT 128.565 15.570 128.865 26.300 ;
        RECT 129.765 15.570 130.065 26.300 ;
        RECT 130.965 15.570 131.265 26.300 ;
        RECT 132.165 15.570 132.465 26.300 ;
        RECT 133.365 15.570 133.665 26.300 ;
        RECT 134.565 15.570 134.865 26.300 ;
        RECT 85.095 15.240 96.505 15.570 ;
        RECT 98.185 15.240 109.595 15.570 ;
        RECT 111.275 15.240 122.685 15.570 ;
        RECT 124.365 15.240 135.775 15.570 ;
        RECT 138.055 15.550 138.355 26.280 ;
        RECT 139.255 15.550 139.555 26.280 ;
        RECT 140.455 15.550 140.755 26.280 ;
        RECT 141.655 15.550 141.955 26.280 ;
        RECT 142.855 15.550 143.155 26.280 ;
        RECT 144.055 15.550 144.355 26.280 ;
        RECT 145.255 15.550 145.555 26.280 ;
        RECT 146.455 15.550 146.755 26.280 ;
        RECT 147.655 15.550 147.955 26.280 ;
        RECT 151.145 15.550 151.445 26.280 ;
        RECT 152.345 15.550 152.645 26.280 ;
        RECT 153.545 15.550 153.845 26.280 ;
        RECT 154.745 15.550 155.045 26.280 ;
        RECT 155.945 15.550 156.245 26.280 ;
        RECT 157.145 15.550 157.445 26.280 ;
        RECT 158.345 15.550 158.645 26.280 ;
        RECT 159.545 15.550 159.845 26.280 ;
        RECT 160.745 15.550 161.045 26.280 ;
        RECT 137.455 15.220 148.865 15.550 ;
        RECT 150.545 15.220 161.955 15.550 ;
        RECT 6.625 13.230 18.035 13.560 ;
        RECT 19.715 13.230 31.125 13.560 ;
        RECT 32.805 13.250 44.215 13.580 ;
        RECT 45.895 13.250 57.305 13.580 ;
        RECT 58.945 13.250 70.355 13.580 ;
        RECT 72.035 13.250 83.445 13.580 ;
        RECT 85.125 13.270 96.535 13.600 ;
        RECT 98.215 13.270 109.625 13.600 ;
        RECT 111.305 13.270 122.715 13.600 ;
        RECT 124.395 13.270 135.805 13.600 ;
        RECT 137.485 13.290 148.895 13.620 ;
        RECT 150.575 13.290 161.985 13.620 ;
        RECT 7.225 2.500 7.525 13.230 ;
        RECT 8.425 2.500 8.725 13.230 ;
        RECT 9.625 2.500 9.925 13.230 ;
        RECT 10.825 2.500 11.125 13.230 ;
        RECT 12.025 2.500 12.325 13.230 ;
        RECT 13.225 2.500 13.525 13.230 ;
        RECT 14.425 2.500 14.725 13.230 ;
        RECT 15.625 2.500 15.925 13.230 ;
        RECT 16.825 2.500 17.125 13.230 ;
        RECT 20.315 2.500 20.615 13.230 ;
        RECT 21.515 2.500 21.815 13.230 ;
        RECT 22.715 2.500 23.015 13.230 ;
        RECT 23.915 2.500 24.215 13.230 ;
        RECT 25.115 2.500 25.415 13.230 ;
        RECT 26.315 2.500 26.615 13.230 ;
        RECT 27.515 2.500 27.815 13.230 ;
        RECT 28.715 2.500 29.015 13.230 ;
        RECT 29.915 2.500 30.215 13.230 ;
        RECT 33.405 2.520 33.705 13.250 ;
        RECT 34.605 2.520 34.905 13.250 ;
        RECT 35.805 2.520 36.105 13.250 ;
        RECT 37.005 2.520 37.305 13.250 ;
        RECT 38.205 2.520 38.505 13.250 ;
        RECT 39.405 2.520 39.705 13.250 ;
        RECT 40.605 2.520 40.905 13.250 ;
        RECT 41.805 2.520 42.105 13.250 ;
        RECT 43.005 2.520 43.305 13.250 ;
        RECT 46.495 2.520 46.795 13.250 ;
        RECT 47.695 2.520 47.995 13.250 ;
        RECT 48.895 2.520 49.195 13.250 ;
        RECT 50.095 2.520 50.395 13.250 ;
        RECT 51.295 2.520 51.595 13.250 ;
        RECT 52.495 2.520 52.795 13.250 ;
        RECT 53.695 2.520 53.995 13.250 ;
        RECT 54.895 2.520 55.195 13.250 ;
        RECT 56.095 2.520 56.395 13.250 ;
        RECT 59.545 2.520 59.845 13.250 ;
        RECT 60.745 2.520 61.045 13.250 ;
        RECT 61.945 2.520 62.245 13.250 ;
        RECT 63.145 2.520 63.445 13.250 ;
        RECT 64.345 2.520 64.645 13.250 ;
        RECT 65.545 2.520 65.845 13.250 ;
        RECT 66.745 2.520 67.045 13.250 ;
        RECT 67.945 2.520 68.245 13.250 ;
        RECT 69.145 2.520 69.445 13.250 ;
        RECT 72.635 2.520 72.935 13.250 ;
        RECT 73.835 2.520 74.135 13.250 ;
        RECT 75.035 2.520 75.335 13.250 ;
        RECT 76.235 2.520 76.535 13.250 ;
        RECT 77.435 2.520 77.735 13.250 ;
        RECT 78.635 2.520 78.935 13.250 ;
        RECT 79.835 2.520 80.135 13.250 ;
        RECT 81.035 2.520 81.335 13.250 ;
        RECT 82.235 2.520 82.535 13.250 ;
        RECT 85.725 2.540 86.025 13.270 ;
        RECT 86.925 2.540 87.225 13.270 ;
        RECT 88.125 2.540 88.425 13.270 ;
        RECT 89.325 2.540 89.625 13.270 ;
        RECT 90.525 2.540 90.825 13.270 ;
        RECT 91.725 2.540 92.025 13.270 ;
        RECT 92.925 2.540 93.225 13.270 ;
        RECT 94.125 2.540 94.425 13.270 ;
        RECT 95.325 2.540 95.625 13.270 ;
        RECT 98.815 2.540 99.115 13.270 ;
        RECT 100.015 2.540 100.315 13.270 ;
        RECT 101.215 2.540 101.515 13.270 ;
        RECT 102.415 2.540 102.715 13.270 ;
        RECT 103.615 2.540 103.915 13.270 ;
        RECT 104.815 2.540 105.115 13.270 ;
        RECT 106.015 2.540 106.315 13.270 ;
        RECT 107.215 2.540 107.515 13.270 ;
        RECT 108.415 2.540 108.715 13.270 ;
        RECT 111.905 2.540 112.205 13.270 ;
        RECT 113.105 2.540 113.405 13.270 ;
        RECT 114.305 2.540 114.605 13.270 ;
        RECT 115.505 2.540 115.805 13.270 ;
        RECT 116.705 2.540 117.005 13.270 ;
        RECT 117.905 2.540 118.205 13.270 ;
        RECT 119.105 2.540 119.405 13.270 ;
        RECT 120.305 2.540 120.605 13.270 ;
        RECT 121.505 2.540 121.805 13.270 ;
        RECT 124.995 2.540 125.295 13.270 ;
        RECT 126.195 2.540 126.495 13.270 ;
        RECT 127.395 2.540 127.695 13.270 ;
        RECT 128.595 2.540 128.895 13.270 ;
        RECT 129.795 2.540 130.095 13.270 ;
        RECT 130.995 2.540 131.295 13.270 ;
        RECT 132.195 2.540 132.495 13.270 ;
        RECT 133.395 2.540 133.695 13.270 ;
        RECT 134.595 2.540 134.895 13.270 ;
        RECT 138.085 2.560 138.385 13.290 ;
        RECT 139.285 2.560 139.585 13.290 ;
        RECT 140.485 2.560 140.785 13.290 ;
        RECT 141.685 2.560 141.985 13.290 ;
        RECT 142.885 2.560 143.185 13.290 ;
        RECT 144.085 2.560 144.385 13.290 ;
        RECT 145.285 2.560 145.585 13.290 ;
        RECT 146.485 2.560 146.785 13.290 ;
        RECT 147.685 2.560 147.985 13.290 ;
        RECT 151.175 2.560 151.475 13.290 ;
        RECT 152.375 2.560 152.675 13.290 ;
        RECT 153.575 2.560 153.875 13.290 ;
        RECT 154.775 2.560 155.075 13.290 ;
        RECT 155.975 2.560 156.275 13.290 ;
        RECT 157.175 2.560 157.475 13.290 ;
        RECT 158.375 2.560 158.675 13.290 ;
        RECT 159.575 2.560 159.875 13.290 ;
        RECT 160.775 2.560 161.075 13.290 ;
      LAYER via3 ;
        RECT 6.295 106.925 6.615 107.245 ;
        RECT 6.695 106.925 7.015 107.245 ;
        RECT 7.095 106.925 7.415 107.245 ;
        RECT 7.495 106.925 7.815 107.245 ;
        RECT 7.895 106.925 8.215 107.245 ;
        RECT 8.295 106.925 8.615 107.245 ;
        RECT 8.695 106.925 9.015 107.245 ;
        RECT 9.095 106.925 9.415 107.245 ;
        RECT 9.495 106.925 9.815 107.245 ;
        RECT 9.895 106.925 10.215 107.245 ;
        RECT 10.295 106.925 10.615 107.245 ;
        RECT 10.695 106.925 11.015 107.245 ;
        RECT 11.095 106.925 11.415 107.245 ;
        RECT 11.495 106.925 11.815 107.245 ;
        RECT 11.895 106.925 12.215 107.245 ;
        RECT 12.295 106.925 12.615 107.245 ;
        RECT 12.695 106.925 13.015 107.245 ;
        RECT 13.095 106.925 13.415 107.245 ;
        RECT 13.495 106.925 13.815 107.245 ;
        RECT 13.895 106.925 14.215 107.245 ;
        RECT 14.295 106.925 14.615 107.245 ;
        RECT 14.695 106.925 15.015 107.245 ;
        RECT 15.095 106.925 15.415 107.245 ;
        RECT 15.495 106.925 15.815 107.245 ;
        RECT 15.895 106.925 16.215 107.245 ;
        RECT 16.295 106.925 16.615 107.245 ;
        RECT 16.695 106.925 17.015 107.245 ;
        RECT 17.095 106.925 17.415 107.245 ;
        RECT 19.385 106.925 19.705 107.245 ;
        RECT 19.785 106.925 20.105 107.245 ;
        RECT 20.185 106.925 20.505 107.245 ;
        RECT 20.585 106.925 20.905 107.245 ;
        RECT 20.985 106.925 21.305 107.245 ;
        RECT 21.385 106.925 21.705 107.245 ;
        RECT 21.785 106.925 22.105 107.245 ;
        RECT 22.185 106.925 22.505 107.245 ;
        RECT 22.585 106.925 22.905 107.245 ;
        RECT 22.985 106.925 23.305 107.245 ;
        RECT 23.385 106.925 23.705 107.245 ;
        RECT 23.785 106.925 24.105 107.245 ;
        RECT 24.185 106.925 24.505 107.245 ;
        RECT 24.585 106.925 24.905 107.245 ;
        RECT 24.985 106.925 25.305 107.245 ;
        RECT 25.385 106.925 25.705 107.245 ;
        RECT 25.785 106.925 26.105 107.245 ;
        RECT 26.185 106.925 26.505 107.245 ;
        RECT 26.585 106.925 26.905 107.245 ;
        RECT 26.985 106.925 27.305 107.245 ;
        RECT 27.385 106.925 27.705 107.245 ;
        RECT 27.785 106.925 28.105 107.245 ;
        RECT 28.185 106.925 28.505 107.245 ;
        RECT 28.585 106.925 28.905 107.245 ;
        RECT 28.985 106.925 29.305 107.245 ;
        RECT 29.385 106.925 29.705 107.245 ;
        RECT 29.785 106.925 30.105 107.245 ;
        RECT 30.185 106.925 30.505 107.245 ;
        RECT 32.475 106.905 32.795 107.225 ;
        RECT 32.875 106.905 33.195 107.225 ;
        RECT 33.275 106.905 33.595 107.225 ;
        RECT 33.675 106.905 33.995 107.225 ;
        RECT 34.075 106.905 34.395 107.225 ;
        RECT 34.475 106.905 34.795 107.225 ;
        RECT 34.875 106.905 35.195 107.225 ;
        RECT 35.275 106.905 35.595 107.225 ;
        RECT 35.675 106.905 35.995 107.225 ;
        RECT 36.075 106.905 36.395 107.225 ;
        RECT 36.475 106.905 36.795 107.225 ;
        RECT 36.875 106.905 37.195 107.225 ;
        RECT 37.275 106.905 37.595 107.225 ;
        RECT 37.675 106.905 37.995 107.225 ;
        RECT 38.075 106.905 38.395 107.225 ;
        RECT 38.475 106.905 38.795 107.225 ;
        RECT 38.875 106.905 39.195 107.225 ;
        RECT 39.275 106.905 39.595 107.225 ;
        RECT 39.675 106.905 39.995 107.225 ;
        RECT 40.075 106.905 40.395 107.225 ;
        RECT 40.475 106.905 40.795 107.225 ;
        RECT 40.875 106.905 41.195 107.225 ;
        RECT 41.275 106.905 41.595 107.225 ;
        RECT 41.675 106.905 41.995 107.225 ;
        RECT 42.075 106.905 42.395 107.225 ;
        RECT 42.475 106.905 42.795 107.225 ;
        RECT 42.875 106.905 43.195 107.225 ;
        RECT 43.275 106.905 43.595 107.225 ;
        RECT 45.565 106.905 45.885 107.225 ;
        RECT 45.965 106.905 46.285 107.225 ;
        RECT 46.365 106.905 46.685 107.225 ;
        RECT 46.765 106.905 47.085 107.225 ;
        RECT 47.165 106.905 47.485 107.225 ;
        RECT 47.565 106.905 47.885 107.225 ;
        RECT 47.965 106.905 48.285 107.225 ;
        RECT 48.365 106.905 48.685 107.225 ;
        RECT 48.765 106.905 49.085 107.225 ;
        RECT 49.165 106.905 49.485 107.225 ;
        RECT 49.565 106.905 49.885 107.225 ;
        RECT 49.965 106.905 50.285 107.225 ;
        RECT 50.365 106.905 50.685 107.225 ;
        RECT 50.765 106.905 51.085 107.225 ;
        RECT 51.165 106.905 51.485 107.225 ;
        RECT 51.565 106.905 51.885 107.225 ;
        RECT 51.965 106.905 52.285 107.225 ;
        RECT 52.365 106.905 52.685 107.225 ;
        RECT 52.765 106.905 53.085 107.225 ;
        RECT 53.165 106.905 53.485 107.225 ;
        RECT 53.565 106.905 53.885 107.225 ;
        RECT 53.965 106.905 54.285 107.225 ;
        RECT 54.365 106.905 54.685 107.225 ;
        RECT 54.765 106.905 55.085 107.225 ;
        RECT 55.165 106.905 55.485 107.225 ;
        RECT 55.565 106.905 55.885 107.225 ;
        RECT 55.965 106.905 56.285 107.225 ;
        RECT 56.365 106.905 56.685 107.225 ;
        RECT 58.615 106.905 58.935 107.225 ;
        RECT 59.015 106.905 59.335 107.225 ;
        RECT 59.415 106.905 59.735 107.225 ;
        RECT 59.815 106.905 60.135 107.225 ;
        RECT 60.215 106.905 60.535 107.225 ;
        RECT 60.615 106.905 60.935 107.225 ;
        RECT 61.015 106.905 61.335 107.225 ;
        RECT 61.415 106.905 61.735 107.225 ;
        RECT 61.815 106.905 62.135 107.225 ;
        RECT 62.215 106.905 62.535 107.225 ;
        RECT 62.615 106.905 62.935 107.225 ;
        RECT 63.015 106.905 63.335 107.225 ;
        RECT 63.415 106.905 63.735 107.225 ;
        RECT 63.815 106.905 64.135 107.225 ;
        RECT 64.215 106.905 64.535 107.225 ;
        RECT 64.615 106.905 64.935 107.225 ;
        RECT 65.015 106.905 65.335 107.225 ;
        RECT 65.415 106.905 65.735 107.225 ;
        RECT 65.815 106.905 66.135 107.225 ;
        RECT 66.215 106.905 66.535 107.225 ;
        RECT 66.615 106.905 66.935 107.225 ;
        RECT 67.015 106.905 67.335 107.225 ;
        RECT 67.415 106.905 67.735 107.225 ;
        RECT 67.815 106.905 68.135 107.225 ;
        RECT 68.215 106.905 68.535 107.225 ;
        RECT 68.615 106.905 68.935 107.225 ;
        RECT 69.015 106.905 69.335 107.225 ;
        RECT 69.415 106.905 69.735 107.225 ;
        RECT 71.705 106.905 72.025 107.225 ;
        RECT 72.105 106.905 72.425 107.225 ;
        RECT 72.505 106.905 72.825 107.225 ;
        RECT 72.905 106.905 73.225 107.225 ;
        RECT 73.305 106.905 73.625 107.225 ;
        RECT 73.705 106.905 74.025 107.225 ;
        RECT 74.105 106.905 74.425 107.225 ;
        RECT 74.505 106.905 74.825 107.225 ;
        RECT 74.905 106.905 75.225 107.225 ;
        RECT 75.305 106.905 75.625 107.225 ;
        RECT 75.705 106.905 76.025 107.225 ;
        RECT 76.105 106.905 76.425 107.225 ;
        RECT 76.505 106.905 76.825 107.225 ;
        RECT 76.905 106.905 77.225 107.225 ;
        RECT 77.305 106.905 77.625 107.225 ;
        RECT 77.705 106.905 78.025 107.225 ;
        RECT 78.105 106.905 78.425 107.225 ;
        RECT 78.505 106.905 78.825 107.225 ;
        RECT 78.905 106.905 79.225 107.225 ;
        RECT 79.305 106.905 79.625 107.225 ;
        RECT 79.705 106.905 80.025 107.225 ;
        RECT 80.105 106.905 80.425 107.225 ;
        RECT 80.505 106.905 80.825 107.225 ;
        RECT 80.905 106.905 81.225 107.225 ;
        RECT 81.305 106.905 81.625 107.225 ;
        RECT 81.705 106.905 82.025 107.225 ;
        RECT 82.105 106.905 82.425 107.225 ;
        RECT 82.505 106.905 82.825 107.225 ;
        RECT 84.795 106.885 85.115 107.205 ;
        RECT 85.195 106.885 85.515 107.205 ;
        RECT 85.595 106.885 85.915 107.205 ;
        RECT 85.995 106.885 86.315 107.205 ;
        RECT 86.395 106.885 86.715 107.205 ;
        RECT 86.795 106.885 87.115 107.205 ;
        RECT 87.195 106.885 87.515 107.205 ;
        RECT 87.595 106.885 87.915 107.205 ;
        RECT 87.995 106.885 88.315 107.205 ;
        RECT 88.395 106.885 88.715 107.205 ;
        RECT 88.795 106.885 89.115 107.205 ;
        RECT 89.195 106.885 89.515 107.205 ;
        RECT 89.595 106.885 89.915 107.205 ;
        RECT 89.995 106.885 90.315 107.205 ;
        RECT 90.395 106.885 90.715 107.205 ;
        RECT 90.795 106.885 91.115 107.205 ;
        RECT 91.195 106.885 91.515 107.205 ;
        RECT 91.595 106.885 91.915 107.205 ;
        RECT 91.995 106.885 92.315 107.205 ;
        RECT 92.395 106.885 92.715 107.205 ;
        RECT 92.795 106.885 93.115 107.205 ;
        RECT 93.195 106.885 93.515 107.205 ;
        RECT 93.595 106.885 93.915 107.205 ;
        RECT 93.995 106.885 94.315 107.205 ;
        RECT 94.395 106.885 94.715 107.205 ;
        RECT 94.795 106.885 95.115 107.205 ;
        RECT 95.195 106.885 95.515 107.205 ;
        RECT 95.595 106.885 95.915 107.205 ;
        RECT 97.885 106.885 98.205 107.205 ;
        RECT 98.285 106.885 98.605 107.205 ;
        RECT 98.685 106.885 99.005 107.205 ;
        RECT 99.085 106.885 99.405 107.205 ;
        RECT 99.485 106.885 99.805 107.205 ;
        RECT 99.885 106.885 100.205 107.205 ;
        RECT 100.285 106.885 100.605 107.205 ;
        RECT 100.685 106.885 101.005 107.205 ;
        RECT 101.085 106.885 101.405 107.205 ;
        RECT 101.485 106.885 101.805 107.205 ;
        RECT 101.885 106.885 102.205 107.205 ;
        RECT 102.285 106.885 102.605 107.205 ;
        RECT 102.685 106.885 103.005 107.205 ;
        RECT 103.085 106.885 103.405 107.205 ;
        RECT 103.485 106.885 103.805 107.205 ;
        RECT 103.885 106.885 104.205 107.205 ;
        RECT 104.285 106.885 104.605 107.205 ;
        RECT 104.685 106.885 105.005 107.205 ;
        RECT 105.085 106.885 105.405 107.205 ;
        RECT 105.485 106.885 105.805 107.205 ;
        RECT 105.885 106.885 106.205 107.205 ;
        RECT 106.285 106.885 106.605 107.205 ;
        RECT 106.685 106.885 107.005 107.205 ;
        RECT 107.085 106.885 107.405 107.205 ;
        RECT 107.485 106.885 107.805 107.205 ;
        RECT 107.885 106.885 108.205 107.205 ;
        RECT 108.285 106.885 108.605 107.205 ;
        RECT 108.685 106.885 109.005 107.205 ;
        RECT 110.975 106.885 111.295 107.205 ;
        RECT 111.375 106.885 111.695 107.205 ;
        RECT 111.775 106.885 112.095 107.205 ;
        RECT 112.175 106.885 112.495 107.205 ;
        RECT 112.575 106.885 112.895 107.205 ;
        RECT 112.975 106.885 113.295 107.205 ;
        RECT 113.375 106.885 113.695 107.205 ;
        RECT 113.775 106.885 114.095 107.205 ;
        RECT 114.175 106.885 114.495 107.205 ;
        RECT 114.575 106.885 114.895 107.205 ;
        RECT 114.975 106.885 115.295 107.205 ;
        RECT 115.375 106.885 115.695 107.205 ;
        RECT 115.775 106.885 116.095 107.205 ;
        RECT 116.175 106.885 116.495 107.205 ;
        RECT 116.575 106.885 116.895 107.205 ;
        RECT 116.975 106.885 117.295 107.205 ;
        RECT 117.375 106.885 117.695 107.205 ;
        RECT 117.775 106.885 118.095 107.205 ;
        RECT 118.175 106.885 118.495 107.205 ;
        RECT 118.575 106.885 118.895 107.205 ;
        RECT 118.975 106.885 119.295 107.205 ;
        RECT 119.375 106.885 119.695 107.205 ;
        RECT 119.775 106.885 120.095 107.205 ;
        RECT 120.175 106.885 120.495 107.205 ;
        RECT 120.575 106.885 120.895 107.205 ;
        RECT 120.975 106.885 121.295 107.205 ;
        RECT 121.375 106.885 121.695 107.205 ;
        RECT 121.775 106.885 122.095 107.205 ;
        RECT 124.065 106.885 124.385 107.205 ;
        RECT 124.465 106.885 124.785 107.205 ;
        RECT 124.865 106.885 125.185 107.205 ;
        RECT 125.265 106.885 125.585 107.205 ;
        RECT 125.665 106.885 125.985 107.205 ;
        RECT 126.065 106.885 126.385 107.205 ;
        RECT 126.465 106.885 126.785 107.205 ;
        RECT 126.865 106.885 127.185 107.205 ;
        RECT 127.265 106.885 127.585 107.205 ;
        RECT 127.665 106.885 127.985 107.205 ;
        RECT 128.065 106.885 128.385 107.205 ;
        RECT 128.465 106.885 128.785 107.205 ;
        RECT 128.865 106.885 129.185 107.205 ;
        RECT 129.265 106.885 129.585 107.205 ;
        RECT 129.665 106.885 129.985 107.205 ;
        RECT 130.065 106.885 130.385 107.205 ;
        RECT 130.465 106.885 130.785 107.205 ;
        RECT 130.865 106.885 131.185 107.205 ;
        RECT 131.265 106.885 131.585 107.205 ;
        RECT 131.665 106.885 131.985 107.205 ;
        RECT 132.065 106.885 132.385 107.205 ;
        RECT 132.465 106.885 132.785 107.205 ;
        RECT 132.865 106.885 133.185 107.205 ;
        RECT 133.265 106.885 133.585 107.205 ;
        RECT 133.665 106.885 133.985 107.205 ;
        RECT 134.065 106.885 134.385 107.205 ;
        RECT 134.465 106.885 134.785 107.205 ;
        RECT 134.865 106.885 135.185 107.205 ;
        RECT 137.155 106.865 137.475 107.185 ;
        RECT 137.555 106.865 137.875 107.185 ;
        RECT 137.955 106.865 138.275 107.185 ;
        RECT 138.355 106.865 138.675 107.185 ;
        RECT 138.755 106.865 139.075 107.185 ;
        RECT 139.155 106.865 139.475 107.185 ;
        RECT 139.555 106.865 139.875 107.185 ;
        RECT 139.955 106.865 140.275 107.185 ;
        RECT 140.355 106.865 140.675 107.185 ;
        RECT 140.755 106.865 141.075 107.185 ;
        RECT 141.155 106.865 141.475 107.185 ;
        RECT 141.555 106.865 141.875 107.185 ;
        RECT 141.955 106.865 142.275 107.185 ;
        RECT 142.355 106.865 142.675 107.185 ;
        RECT 142.755 106.865 143.075 107.185 ;
        RECT 143.155 106.865 143.475 107.185 ;
        RECT 143.555 106.865 143.875 107.185 ;
        RECT 143.955 106.865 144.275 107.185 ;
        RECT 144.355 106.865 144.675 107.185 ;
        RECT 144.755 106.865 145.075 107.185 ;
        RECT 145.155 106.865 145.475 107.185 ;
        RECT 145.555 106.865 145.875 107.185 ;
        RECT 145.955 106.865 146.275 107.185 ;
        RECT 146.355 106.865 146.675 107.185 ;
        RECT 146.755 106.865 147.075 107.185 ;
        RECT 147.155 106.865 147.475 107.185 ;
        RECT 147.555 106.865 147.875 107.185 ;
        RECT 147.955 106.865 148.275 107.185 ;
        RECT 150.245 106.865 150.565 107.185 ;
        RECT 150.645 106.865 150.965 107.185 ;
        RECT 151.045 106.865 151.365 107.185 ;
        RECT 151.445 106.865 151.765 107.185 ;
        RECT 151.845 106.865 152.165 107.185 ;
        RECT 152.245 106.865 152.565 107.185 ;
        RECT 152.645 106.865 152.965 107.185 ;
        RECT 153.045 106.865 153.365 107.185 ;
        RECT 153.445 106.865 153.765 107.185 ;
        RECT 153.845 106.865 154.165 107.185 ;
        RECT 154.245 106.865 154.565 107.185 ;
        RECT 154.645 106.865 154.965 107.185 ;
        RECT 155.045 106.865 155.365 107.185 ;
        RECT 155.445 106.865 155.765 107.185 ;
        RECT 155.845 106.865 156.165 107.185 ;
        RECT 156.245 106.865 156.565 107.185 ;
        RECT 156.645 106.865 156.965 107.185 ;
        RECT 157.045 106.865 157.365 107.185 ;
        RECT 157.445 106.865 157.765 107.185 ;
        RECT 157.845 106.865 158.165 107.185 ;
        RECT 158.245 106.865 158.565 107.185 ;
        RECT 158.645 106.865 158.965 107.185 ;
        RECT 159.045 106.865 159.365 107.185 ;
        RECT 159.445 106.865 159.765 107.185 ;
        RECT 159.845 106.865 160.165 107.185 ;
        RECT 160.245 106.865 160.565 107.185 ;
        RECT 160.645 106.865 160.965 107.185 ;
        RECT 161.045 106.865 161.365 107.185 ;
        RECT 6.325 104.875 6.645 105.195 ;
        RECT 6.725 104.875 7.045 105.195 ;
        RECT 7.125 104.875 7.445 105.195 ;
        RECT 7.525 104.875 7.845 105.195 ;
        RECT 7.925 104.875 8.245 105.195 ;
        RECT 8.325 104.875 8.645 105.195 ;
        RECT 8.725 104.875 9.045 105.195 ;
        RECT 9.125 104.875 9.445 105.195 ;
        RECT 9.525 104.875 9.845 105.195 ;
        RECT 9.925 104.875 10.245 105.195 ;
        RECT 10.325 104.875 10.645 105.195 ;
        RECT 10.725 104.875 11.045 105.195 ;
        RECT 11.125 104.875 11.445 105.195 ;
        RECT 11.525 104.875 11.845 105.195 ;
        RECT 11.925 104.875 12.245 105.195 ;
        RECT 12.325 104.875 12.645 105.195 ;
        RECT 12.725 104.875 13.045 105.195 ;
        RECT 13.125 104.875 13.445 105.195 ;
        RECT 13.525 104.875 13.845 105.195 ;
        RECT 13.925 104.875 14.245 105.195 ;
        RECT 14.325 104.875 14.645 105.195 ;
        RECT 14.725 104.875 15.045 105.195 ;
        RECT 15.125 104.875 15.445 105.195 ;
        RECT 15.525 104.875 15.845 105.195 ;
        RECT 15.925 104.875 16.245 105.195 ;
        RECT 16.325 104.875 16.645 105.195 ;
        RECT 16.725 104.875 17.045 105.195 ;
        RECT 17.125 104.875 17.445 105.195 ;
        RECT 19.415 104.875 19.735 105.195 ;
        RECT 19.815 104.875 20.135 105.195 ;
        RECT 20.215 104.875 20.535 105.195 ;
        RECT 20.615 104.875 20.935 105.195 ;
        RECT 21.015 104.875 21.335 105.195 ;
        RECT 21.415 104.875 21.735 105.195 ;
        RECT 21.815 104.875 22.135 105.195 ;
        RECT 22.215 104.875 22.535 105.195 ;
        RECT 22.615 104.875 22.935 105.195 ;
        RECT 23.015 104.875 23.335 105.195 ;
        RECT 23.415 104.875 23.735 105.195 ;
        RECT 23.815 104.875 24.135 105.195 ;
        RECT 24.215 104.875 24.535 105.195 ;
        RECT 24.615 104.875 24.935 105.195 ;
        RECT 25.015 104.875 25.335 105.195 ;
        RECT 25.415 104.875 25.735 105.195 ;
        RECT 25.815 104.875 26.135 105.195 ;
        RECT 26.215 104.875 26.535 105.195 ;
        RECT 26.615 104.875 26.935 105.195 ;
        RECT 27.015 104.875 27.335 105.195 ;
        RECT 27.415 104.875 27.735 105.195 ;
        RECT 27.815 104.875 28.135 105.195 ;
        RECT 28.215 104.875 28.535 105.195 ;
        RECT 28.615 104.875 28.935 105.195 ;
        RECT 29.015 104.875 29.335 105.195 ;
        RECT 29.415 104.875 29.735 105.195 ;
        RECT 29.815 104.875 30.135 105.195 ;
        RECT 30.215 104.875 30.535 105.195 ;
        RECT 32.505 104.895 32.825 105.215 ;
        RECT 32.905 104.895 33.225 105.215 ;
        RECT 33.305 104.895 33.625 105.215 ;
        RECT 33.705 104.895 34.025 105.215 ;
        RECT 34.105 104.895 34.425 105.215 ;
        RECT 34.505 104.895 34.825 105.215 ;
        RECT 34.905 104.895 35.225 105.215 ;
        RECT 35.305 104.895 35.625 105.215 ;
        RECT 35.705 104.895 36.025 105.215 ;
        RECT 36.105 104.895 36.425 105.215 ;
        RECT 36.505 104.895 36.825 105.215 ;
        RECT 36.905 104.895 37.225 105.215 ;
        RECT 37.305 104.895 37.625 105.215 ;
        RECT 37.705 104.895 38.025 105.215 ;
        RECT 38.105 104.895 38.425 105.215 ;
        RECT 38.505 104.895 38.825 105.215 ;
        RECT 38.905 104.895 39.225 105.215 ;
        RECT 39.305 104.895 39.625 105.215 ;
        RECT 39.705 104.895 40.025 105.215 ;
        RECT 40.105 104.895 40.425 105.215 ;
        RECT 40.505 104.895 40.825 105.215 ;
        RECT 40.905 104.895 41.225 105.215 ;
        RECT 41.305 104.895 41.625 105.215 ;
        RECT 41.705 104.895 42.025 105.215 ;
        RECT 42.105 104.895 42.425 105.215 ;
        RECT 42.505 104.895 42.825 105.215 ;
        RECT 42.905 104.895 43.225 105.215 ;
        RECT 43.305 104.895 43.625 105.215 ;
        RECT 45.595 104.895 45.915 105.215 ;
        RECT 45.995 104.895 46.315 105.215 ;
        RECT 46.395 104.895 46.715 105.215 ;
        RECT 46.795 104.895 47.115 105.215 ;
        RECT 47.195 104.895 47.515 105.215 ;
        RECT 47.595 104.895 47.915 105.215 ;
        RECT 47.995 104.895 48.315 105.215 ;
        RECT 48.395 104.895 48.715 105.215 ;
        RECT 48.795 104.895 49.115 105.215 ;
        RECT 49.195 104.895 49.515 105.215 ;
        RECT 49.595 104.895 49.915 105.215 ;
        RECT 49.995 104.895 50.315 105.215 ;
        RECT 50.395 104.895 50.715 105.215 ;
        RECT 50.795 104.895 51.115 105.215 ;
        RECT 51.195 104.895 51.515 105.215 ;
        RECT 51.595 104.895 51.915 105.215 ;
        RECT 51.995 104.895 52.315 105.215 ;
        RECT 52.395 104.895 52.715 105.215 ;
        RECT 52.795 104.895 53.115 105.215 ;
        RECT 53.195 104.895 53.515 105.215 ;
        RECT 53.595 104.895 53.915 105.215 ;
        RECT 53.995 104.895 54.315 105.215 ;
        RECT 54.395 104.895 54.715 105.215 ;
        RECT 54.795 104.895 55.115 105.215 ;
        RECT 55.195 104.895 55.515 105.215 ;
        RECT 55.595 104.895 55.915 105.215 ;
        RECT 55.995 104.895 56.315 105.215 ;
        RECT 56.395 104.895 56.715 105.215 ;
        RECT 58.645 104.895 58.965 105.215 ;
        RECT 59.045 104.895 59.365 105.215 ;
        RECT 59.445 104.895 59.765 105.215 ;
        RECT 59.845 104.895 60.165 105.215 ;
        RECT 60.245 104.895 60.565 105.215 ;
        RECT 60.645 104.895 60.965 105.215 ;
        RECT 61.045 104.895 61.365 105.215 ;
        RECT 61.445 104.895 61.765 105.215 ;
        RECT 61.845 104.895 62.165 105.215 ;
        RECT 62.245 104.895 62.565 105.215 ;
        RECT 62.645 104.895 62.965 105.215 ;
        RECT 63.045 104.895 63.365 105.215 ;
        RECT 63.445 104.895 63.765 105.215 ;
        RECT 63.845 104.895 64.165 105.215 ;
        RECT 64.245 104.895 64.565 105.215 ;
        RECT 64.645 104.895 64.965 105.215 ;
        RECT 65.045 104.895 65.365 105.215 ;
        RECT 65.445 104.895 65.765 105.215 ;
        RECT 65.845 104.895 66.165 105.215 ;
        RECT 66.245 104.895 66.565 105.215 ;
        RECT 66.645 104.895 66.965 105.215 ;
        RECT 67.045 104.895 67.365 105.215 ;
        RECT 67.445 104.895 67.765 105.215 ;
        RECT 67.845 104.895 68.165 105.215 ;
        RECT 68.245 104.895 68.565 105.215 ;
        RECT 68.645 104.895 68.965 105.215 ;
        RECT 69.045 104.895 69.365 105.215 ;
        RECT 69.445 104.895 69.765 105.215 ;
        RECT 71.735 104.895 72.055 105.215 ;
        RECT 72.135 104.895 72.455 105.215 ;
        RECT 72.535 104.895 72.855 105.215 ;
        RECT 72.935 104.895 73.255 105.215 ;
        RECT 73.335 104.895 73.655 105.215 ;
        RECT 73.735 104.895 74.055 105.215 ;
        RECT 74.135 104.895 74.455 105.215 ;
        RECT 74.535 104.895 74.855 105.215 ;
        RECT 74.935 104.895 75.255 105.215 ;
        RECT 75.335 104.895 75.655 105.215 ;
        RECT 75.735 104.895 76.055 105.215 ;
        RECT 76.135 104.895 76.455 105.215 ;
        RECT 76.535 104.895 76.855 105.215 ;
        RECT 76.935 104.895 77.255 105.215 ;
        RECT 77.335 104.895 77.655 105.215 ;
        RECT 77.735 104.895 78.055 105.215 ;
        RECT 78.135 104.895 78.455 105.215 ;
        RECT 78.535 104.895 78.855 105.215 ;
        RECT 78.935 104.895 79.255 105.215 ;
        RECT 79.335 104.895 79.655 105.215 ;
        RECT 79.735 104.895 80.055 105.215 ;
        RECT 80.135 104.895 80.455 105.215 ;
        RECT 80.535 104.895 80.855 105.215 ;
        RECT 80.935 104.895 81.255 105.215 ;
        RECT 81.335 104.895 81.655 105.215 ;
        RECT 81.735 104.895 82.055 105.215 ;
        RECT 82.135 104.895 82.455 105.215 ;
        RECT 82.535 104.895 82.855 105.215 ;
        RECT 84.825 104.915 85.145 105.235 ;
        RECT 85.225 104.915 85.545 105.235 ;
        RECT 85.625 104.915 85.945 105.235 ;
        RECT 86.025 104.915 86.345 105.235 ;
        RECT 86.425 104.915 86.745 105.235 ;
        RECT 86.825 104.915 87.145 105.235 ;
        RECT 87.225 104.915 87.545 105.235 ;
        RECT 87.625 104.915 87.945 105.235 ;
        RECT 88.025 104.915 88.345 105.235 ;
        RECT 88.425 104.915 88.745 105.235 ;
        RECT 88.825 104.915 89.145 105.235 ;
        RECT 89.225 104.915 89.545 105.235 ;
        RECT 89.625 104.915 89.945 105.235 ;
        RECT 90.025 104.915 90.345 105.235 ;
        RECT 90.425 104.915 90.745 105.235 ;
        RECT 90.825 104.915 91.145 105.235 ;
        RECT 91.225 104.915 91.545 105.235 ;
        RECT 91.625 104.915 91.945 105.235 ;
        RECT 92.025 104.915 92.345 105.235 ;
        RECT 92.425 104.915 92.745 105.235 ;
        RECT 92.825 104.915 93.145 105.235 ;
        RECT 93.225 104.915 93.545 105.235 ;
        RECT 93.625 104.915 93.945 105.235 ;
        RECT 94.025 104.915 94.345 105.235 ;
        RECT 94.425 104.915 94.745 105.235 ;
        RECT 94.825 104.915 95.145 105.235 ;
        RECT 95.225 104.915 95.545 105.235 ;
        RECT 95.625 104.915 95.945 105.235 ;
        RECT 97.915 104.915 98.235 105.235 ;
        RECT 98.315 104.915 98.635 105.235 ;
        RECT 98.715 104.915 99.035 105.235 ;
        RECT 99.115 104.915 99.435 105.235 ;
        RECT 99.515 104.915 99.835 105.235 ;
        RECT 99.915 104.915 100.235 105.235 ;
        RECT 100.315 104.915 100.635 105.235 ;
        RECT 100.715 104.915 101.035 105.235 ;
        RECT 101.115 104.915 101.435 105.235 ;
        RECT 101.515 104.915 101.835 105.235 ;
        RECT 101.915 104.915 102.235 105.235 ;
        RECT 102.315 104.915 102.635 105.235 ;
        RECT 102.715 104.915 103.035 105.235 ;
        RECT 103.115 104.915 103.435 105.235 ;
        RECT 103.515 104.915 103.835 105.235 ;
        RECT 103.915 104.915 104.235 105.235 ;
        RECT 104.315 104.915 104.635 105.235 ;
        RECT 104.715 104.915 105.035 105.235 ;
        RECT 105.115 104.915 105.435 105.235 ;
        RECT 105.515 104.915 105.835 105.235 ;
        RECT 105.915 104.915 106.235 105.235 ;
        RECT 106.315 104.915 106.635 105.235 ;
        RECT 106.715 104.915 107.035 105.235 ;
        RECT 107.115 104.915 107.435 105.235 ;
        RECT 107.515 104.915 107.835 105.235 ;
        RECT 107.915 104.915 108.235 105.235 ;
        RECT 108.315 104.915 108.635 105.235 ;
        RECT 108.715 104.915 109.035 105.235 ;
        RECT 111.005 104.915 111.325 105.235 ;
        RECT 111.405 104.915 111.725 105.235 ;
        RECT 111.805 104.915 112.125 105.235 ;
        RECT 112.205 104.915 112.525 105.235 ;
        RECT 112.605 104.915 112.925 105.235 ;
        RECT 113.005 104.915 113.325 105.235 ;
        RECT 113.405 104.915 113.725 105.235 ;
        RECT 113.805 104.915 114.125 105.235 ;
        RECT 114.205 104.915 114.525 105.235 ;
        RECT 114.605 104.915 114.925 105.235 ;
        RECT 115.005 104.915 115.325 105.235 ;
        RECT 115.405 104.915 115.725 105.235 ;
        RECT 115.805 104.915 116.125 105.235 ;
        RECT 116.205 104.915 116.525 105.235 ;
        RECT 116.605 104.915 116.925 105.235 ;
        RECT 117.005 104.915 117.325 105.235 ;
        RECT 117.405 104.915 117.725 105.235 ;
        RECT 117.805 104.915 118.125 105.235 ;
        RECT 118.205 104.915 118.525 105.235 ;
        RECT 118.605 104.915 118.925 105.235 ;
        RECT 119.005 104.915 119.325 105.235 ;
        RECT 119.405 104.915 119.725 105.235 ;
        RECT 119.805 104.915 120.125 105.235 ;
        RECT 120.205 104.915 120.525 105.235 ;
        RECT 120.605 104.915 120.925 105.235 ;
        RECT 121.005 104.915 121.325 105.235 ;
        RECT 121.405 104.915 121.725 105.235 ;
        RECT 121.805 104.915 122.125 105.235 ;
        RECT 124.095 104.915 124.415 105.235 ;
        RECT 124.495 104.915 124.815 105.235 ;
        RECT 124.895 104.915 125.215 105.235 ;
        RECT 125.295 104.915 125.615 105.235 ;
        RECT 125.695 104.915 126.015 105.235 ;
        RECT 126.095 104.915 126.415 105.235 ;
        RECT 126.495 104.915 126.815 105.235 ;
        RECT 126.895 104.915 127.215 105.235 ;
        RECT 127.295 104.915 127.615 105.235 ;
        RECT 127.695 104.915 128.015 105.235 ;
        RECT 128.095 104.915 128.415 105.235 ;
        RECT 128.495 104.915 128.815 105.235 ;
        RECT 128.895 104.915 129.215 105.235 ;
        RECT 129.295 104.915 129.615 105.235 ;
        RECT 129.695 104.915 130.015 105.235 ;
        RECT 130.095 104.915 130.415 105.235 ;
        RECT 130.495 104.915 130.815 105.235 ;
        RECT 130.895 104.915 131.215 105.235 ;
        RECT 131.295 104.915 131.615 105.235 ;
        RECT 131.695 104.915 132.015 105.235 ;
        RECT 132.095 104.915 132.415 105.235 ;
        RECT 132.495 104.915 132.815 105.235 ;
        RECT 132.895 104.915 133.215 105.235 ;
        RECT 133.295 104.915 133.615 105.235 ;
        RECT 133.695 104.915 134.015 105.235 ;
        RECT 134.095 104.915 134.415 105.235 ;
        RECT 134.495 104.915 134.815 105.235 ;
        RECT 134.895 104.915 135.215 105.235 ;
        RECT 137.185 104.935 137.505 105.255 ;
        RECT 137.585 104.935 137.905 105.255 ;
        RECT 137.985 104.935 138.305 105.255 ;
        RECT 138.385 104.935 138.705 105.255 ;
        RECT 138.785 104.935 139.105 105.255 ;
        RECT 139.185 104.935 139.505 105.255 ;
        RECT 139.585 104.935 139.905 105.255 ;
        RECT 139.985 104.935 140.305 105.255 ;
        RECT 140.385 104.935 140.705 105.255 ;
        RECT 140.785 104.935 141.105 105.255 ;
        RECT 141.185 104.935 141.505 105.255 ;
        RECT 141.585 104.935 141.905 105.255 ;
        RECT 141.985 104.935 142.305 105.255 ;
        RECT 142.385 104.935 142.705 105.255 ;
        RECT 142.785 104.935 143.105 105.255 ;
        RECT 143.185 104.935 143.505 105.255 ;
        RECT 143.585 104.935 143.905 105.255 ;
        RECT 143.985 104.935 144.305 105.255 ;
        RECT 144.385 104.935 144.705 105.255 ;
        RECT 144.785 104.935 145.105 105.255 ;
        RECT 145.185 104.935 145.505 105.255 ;
        RECT 145.585 104.935 145.905 105.255 ;
        RECT 145.985 104.935 146.305 105.255 ;
        RECT 146.385 104.935 146.705 105.255 ;
        RECT 146.785 104.935 147.105 105.255 ;
        RECT 147.185 104.935 147.505 105.255 ;
        RECT 147.585 104.935 147.905 105.255 ;
        RECT 147.985 104.935 148.305 105.255 ;
        RECT 150.275 104.935 150.595 105.255 ;
        RECT 150.675 104.935 150.995 105.255 ;
        RECT 151.075 104.935 151.395 105.255 ;
        RECT 151.475 104.935 151.795 105.255 ;
        RECT 151.875 104.935 152.195 105.255 ;
        RECT 152.275 104.935 152.595 105.255 ;
        RECT 152.675 104.935 152.995 105.255 ;
        RECT 153.075 104.935 153.395 105.255 ;
        RECT 153.475 104.935 153.795 105.255 ;
        RECT 153.875 104.935 154.195 105.255 ;
        RECT 154.275 104.935 154.595 105.255 ;
        RECT 154.675 104.935 154.995 105.255 ;
        RECT 155.075 104.935 155.395 105.255 ;
        RECT 155.475 104.935 155.795 105.255 ;
        RECT 155.875 104.935 156.195 105.255 ;
        RECT 156.275 104.935 156.595 105.255 ;
        RECT 156.675 104.935 156.995 105.255 ;
        RECT 157.075 104.935 157.395 105.255 ;
        RECT 157.475 104.935 157.795 105.255 ;
        RECT 157.875 104.935 158.195 105.255 ;
        RECT 158.275 104.935 158.595 105.255 ;
        RECT 158.675 104.935 158.995 105.255 ;
        RECT 159.075 104.935 159.395 105.255 ;
        RECT 159.475 104.935 159.795 105.255 ;
        RECT 159.875 104.935 160.195 105.255 ;
        RECT 160.275 104.935 160.595 105.255 ;
        RECT 160.675 104.935 160.995 105.255 ;
        RECT 161.075 104.935 161.395 105.255 ;
        RECT 162.900 90.245 163.375 90.770 ;
        RECT 4.735 88.700 5.255 89.170 ;
        RECT 4.725 33.190 5.245 33.660 ;
        RECT 163.250 29.240 163.775 29.715 ;
        RECT 6.735 15.285 7.055 15.605 ;
        RECT 7.135 15.285 7.455 15.605 ;
        RECT 7.535 15.285 7.855 15.605 ;
        RECT 7.935 15.285 8.255 15.605 ;
        RECT 8.335 15.285 8.655 15.605 ;
        RECT 8.735 15.285 9.055 15.605 ;
        RECT 9.135 15.285 9.455 15.605 ;
        RECT 9.535 15.285 9.855 15.605 ;
        RECT 9.935 15.285 10.255 15.605 ;
        RECT 10.335 15.285 10.655 15.605 ;
        RECT 10.735 15.285 11.055 15.605 ;
        RECT 11.135 15.285 11.455 15.605 ;
        RECT 11.535 15.285 11.855 15.605 ;
        RECT 11.935 15.285 12.255 15.605 ;
        RECT 12.335 15.285 12.655 15.605 ;
        RECT 12.735 15.285 13.055 15.605 ;
        RECT 13.135 15.285 13.455 15.605 ;
        RECT 13.535 15.285 13.855 15.605 ;
        RECT 13.935 15.285 14.255 15.605 ;
        RECT 14.335 15.285 14.655 15.605 ;
        RECT 14.735 15.285 15.055 15.605 ;
        RECT 15.135 15.285 15.455 15.605 ;
        RECT 15.535 15.285 15.855 15.605 ;
        RECT 15.935 15.285 16.255 15.605 ;
        RECT 16.335 15.285 16.655 15.605 ;
        RECT 16.735 15.285 17.055 15.605 ;
        RECT 17.135 15.285 17.455 15.605 ;
        RECT 17.535 15.285 17.855 15.605 ;
        RECT 19.825 15.285 20.145 15.605 ;
        RECT 20.225 15.285 20.545 15.605 ;
        RECT 20.625 15.285 20.945 15.605 ;
        RECT 21.025 15.285 21.345 15.605 ;
        RECT 21.425 15.285 21.745 15.605 ;
        RECT 21.825 15.285 22.145 15.605 ;
        RECT 22.225 15.285 22.545 15.605 ;
        RECT 22.625 15.285 22.945 15.605 ;
        RECT 23.025 15.285 23.345 15.605 ;
        RECT 23.425 15.285 23.745 15.605 ;
        RECT 23.825 15.285 24.145 15.605 ;
        RECT 24.225 15.285 24.545 15.605 ;
        RECT 24.625 15.285 24.945 15.605 ;
        RECT 25.025 15.285 25.345 15.605 ;
        RECT 25.425 15.285 25.745 15.605 ;
        RECT 25.825 15.285 26.145 15.605 ;
        RECT 26.225 15.285 26.545 15.605 ;
        RECT 26.625 15.285 26.945 15.605 ;
        RECT 27.025 15.285 27.345 15.605 ;
        RECT 27.425 15.285 27.745 15.605 ;
        RECT 27.825 15.285 28.145 15.605 ;
        RECT 28.225 15.285 28.545 15.605 ;
        RECT 28.625 15.285 28.945 15.605 ;
        RECT 29.025 15.285 29.345 15.605 ;
        RECT 29.425 15.285 29.745 15.605 ;
        RECT 29.825 15.285 30.145 15.605 ;
        RECT 30.225 15.285 30.545 15.605 ;
        RECT 30.625 15.285 30.945 15.605 ;
        RECT 32.915 15.265 33.235 15.585 ;
        RECT 33.315 15.265 33.635 15.585 ;
        RECT 33.715 15.265 34.035 15.585 ;
        RECT 34.115 15.265 34.435 15.585 ;
        RECT 34.515 15.265 34.835 15.585 ;
        RECT 34.915 15.265 35.235 15.585 ;
        RECT 35.315 15.265 35.635 15.585 ;
        RECT 35.715 15.265 36.035 15.585 ;
        RECT 36.115 15.265 36.435 15.585 ;
        RECT 36.515 15.265 36.835 15.585 ;
        RECT 36.915 15.265 37.235 15.585 ;
        RECT 37.315 15.265 37.635 15.585 ;
        RECT 37.715 15.265 38.035 15.585 ;
        RECT 38.115 15.265 38.435 15.585 ;
        RECT 38.515 15.265 38.835 15.585 ;
        RECT 38.915 15.265 39.235 15.585 ;
        RECT 39.315 15.265 39.635 15.585 ;
        RECT 39.715 15.265 40.035 15.585 ;
        RECT 40.115 15.265 40.435 15.585 ;
        RECT 40.515 15.265 40.835 15.585 ;
        RECT 40.915 15.265 41.235 15.585 ;
        RECT 41.315 15.265 41.635 15.585 ;
        RECT 41.715 15.265 42.035 15.585 ;
        RECT 42.115 15.265 42.435 15.585 ;
        RECT 42.515 15.265 42.835 15.585 ;
        RECT 42.915 15.265 43.235 15.585 ;
        RECT 43.315 15.265 43.635 15.585 ;
        RECT 43.715 15.265 44.035 15.585 ;
        RECT 46.005 15.265 46.325 15.585 ;
        RECT 46.405 15.265 46.725 15.585 ;
        RECT 46.805 15.265 47.125 15.585 ;
        RECT 47.205 15.265 47.525 15.585 ;
        RECT 47.605 15.265 47.925 15.585 ;
        RECT 48.005 15.265 48.325 15.585 ;
        RECT 48.405 15.265 48.725 15.585 ;
        RECT 48.805 15.265 49.125 15.585 ;
        RECT 49.205 15.265 49.525 15.585 ;
        RECT 49.605 15.265 49.925 15.585 ;
        RECT 50.005 15.265 50.325 15.585 ;
        RECT 50.405 15.265 50.725 15.585 ;
        RECT 50.805 15.265 51.125 15.585 ;
        RECT 51.205 15.265 51.525 15.585 ;
        RECT 51.605 15.265 51.925 15.585 ;
        RECT 52.005 15.265 52.325 15.585 ;
        RECT 52.405 15.265 52.725 15.585 ;
        RECT 52.805 15.265 53.125 15.585 ;
        RECT 53.205 15.265 53.525 15.585 ;
        RECT 53.605 15.265 53.925 15.585 ;
        RECT 54.005 15.265 54.325 15.585 ;
        RECT 54.405 15.265 54.725 15.585 ;
        RECT 54.805 15.265 55.125 15.585 ;
        RECT 55.205 15.265 55.525 15.585 ;
        RECT 55.605 15.265 55.925 15.585 ;
        RECT 56.005 15.265 56.325 15.585 ;
        RECT 56.405 15.265 56.725 15.585 ;
        RECT 56.805 15.265 57.125 15.585 ;
        RECT 59.055 15.265 59.375 15.585 ;
        RECT 59.455 15.265 59.775 15.585 ;
        RECT 59.855 15.265 60.175 15.585 ;
        RECT 60.255 15.265 60.575 15.585 ;
        RECT 60.655 15.265 60.975 15.585 ;
        RECT 61.055 15.265 61.375 15.585 ;
        RECT 61.455 15.265 61.775 15.585 ;
        RECT 61.855 15.265 62.175 15.585 ;
        RECT 62.255 15.265 62.575 15.585 ;
        RECT 62.655 15.265 62.975 15.585 ;
        RECT 63.055 15.265 63.375 15.585 ;
        RECT 63.455 15.265 63.775 15.585 ;
        RECT 63.855 15.265 64.175 15.585 ;
        RECT 64.255 15.265 64.575 15.585 ;
        RECT 64.655 15.265 64.975 15.585 ;
        RECT 65.055 15.265 65.375 15.585 ;
        RECT 65.455 15.265 65.775 15.585 ;
        RECT 65.855 15.265 66.175 15.585 ;
        RECT 66.255 15.265 66.575 15.585 ;
        RECT 66.655 15.265 66.975 15.585 ;
        RECT 67.055 15.265 67.375 15.585 ;
        RECT 67.455 15.265 67.775 15.585 ;
        RECT 67.855 15.265 68.175 15.585 ;
        RECT 68.255 15.265 68.575 15.585 ;
        RECT 68.655 15.265 68.975 15.585 ;
        RECT 69.055 15.265 69.375 15.585 ;
        RECT 69.455 15.265 69.775 15.585 ;
        RECT 69.855 15.265 70.175 15.585 ;
        RECT 72.145 15.265 72.465 15.585 ;
        RECT 72.545 15.265 72.865 15.585 ;
        RECT 72.945 15.265 73.265 15.585 ;
        RECT 73.345 15.265 73.665 15.585 ;
        RECT 73.745 15.265 74.065 15.585 ;
        RECT 74.145 15.265 74.465 15.585 ;
        RECT 74.545 15.265 74.865 15.585 ;
        RECT 74.945 15.265 75.265 15.585 ;
        RECT 75.345 15.265 75.665 15.585 ;
        RECT 75.745 15.265 76.065 15.585 ;
        RECT 76.145 15.265 76.465 15.585 ;
        RECT 76.545 15.265 76.865 15.585 ;
        RECT 76.945 15.265 77.265 15.585 ;
        RECT 77.345 15.265 77.665 15.585 ;
        RECT 77.745 15.265 78.065 15.585 ;
        RECT 78.145 15.265 78.465 15.585 ;
        RECT 78.545 15.265 78.865 15.585 ;
        RECT 78.945 15.265 79.265 15.585 ;
        RECT 79.345 15.265 79.665 15.585 ;
        RECT 79.745 15.265 80.065 15.585 ;
        RECT 80.145 15.265 80.465 15.585 ;
        RECT 80.545 15.265 80.865 15.585 ;
        RECT 80.945 15.265 81.265 15.585 ;
        RECT 81.345 15.265 81.665 15.585 ;
        RECT 81.745 15.265 82.065 15.585 ;
        RECT 82.145 15.265 82.465 15.585 ;
        RECT 82.545 15.265 82.865 15.585 ;
        RECT 82.945 15.265 83.265 15.585 ;
        RECT 85.235 15.245 85.555 15.565 ;
        RECT 85.635 15.245 85.955 15.565 ;
        RECT 86.035 15.245 86.355 15.565 ;
        RECT 86.435 15.245 86.755 15.565 ;
        RECT 86.835 15.245 87.155 15.565 ;
        RECT 87.235 15.245 87.555 15.565 ;
        RECT 87.635 15.245 87.955 15.565 ;
        RECT 88.035 15.245 88.355 15.565 ;
        RECT 88.435 15.245 88.755 15.565 ;
        RECT 88.835 15.245 89.155 15.565 ;
        RECT 89.235 15.245 89.555 15.565 ;
        RECT 89.635 15.245 89.955 15.565 ;
        RECT 90.035 15.245 90.355 15.565 ;
        RECT 90.435 15.245 90.755 15.565 ;
        RECT 90.835 15.245 91.155 15.565 ;
        RECT 91.235 15.245 91.555 15.565 ;
        RECT 91.635 15.245 91.955 15.565 ;
        RECT 92.035 15.245 92.355 15.565 ;
        RECT 92.435 15.245 92.755 15.565 ;
        RECT 92.835 15.245 93.155 15.565 ;
        RECT 93.235 15.245 93.555 15.565 ;
        RECT 93.635 15.245 93.955 15.565 ;
        RECT 94.035 15.245 94.355 15.565 ;
        RECT 94.435 15.245 94.755 15.565 ;
        RECT 94.835 15.245 95.155 15.565 ;
        RECT 95.235 15.245 95.555 15.565 ;
        RECT 95.635 15.245 95.955 15.565 ;
        RECT 96.035 15.245 96.355 15.565 ;
        RECT 98.325 15.245 98.645 15.565 ;
        RECT 98.725 15.245 99.045 15.565 ;
        RECT 99.125 15.245 99.445 15.565 ;
        RECT 99.525 15.245 99.845 15.565 ;
        RECT 99.925 15.245 100.245 15.565 ;
        RECT 100.325 15.245 100.645 15.565 ;
        RECT 100.725 15.245 101.045 15.565 ;
        RECT 101.125 15.245 101.445 15.565 ;
        RECT 101.525 15.245 101.845 15.565 ;
        RECT 101.925 15.245 102.245 15.565 ;
        RECT 102.325 15.245 102.645 15.565 ;
        RECT 102.725 15.245 103.045 15.565 ;
        RECT 103.125 15.245 103.445 15.565 ;
        RECT 103.525 15.245 103.845 15.565 ;
        RECT 103.925 15.245 104.245 15.565 ;
        RECT 104.325 15.245 104.645 15.565 ;
        RECT 104.725 15.245 105.045 15.565 ;
        RECT 105.125 15.245 105.445 15.565 ;
        RECT 105.525 15.245 105.845 15.565 ;
        RECT 105.925 15.245 106.245 15.565 ;
        RECT 106.325 15.245 106.645 15.565 ;
        RECT 106.725 15.245 107.045 15.565 ;
        RECT 107.125 15.245 107.445 15.565 ;
        RECT 107.525 15.245 107.845 15.565 ;
        RECT 107.925 15.245 108.245 15.565 ;
        RECT 108.325 15.245 108.645 15.565 ;
        RECT 108.725 15.245 109.045 15.565 ;
        RECT 109.125 15.245 109.445 15.565 ;
        RECT 111.415 15.245 111.735 15.565 ;
        RECT 111.815 15.245 112.135 15.565 ;
        RECT 112.215 15.245 112.535 15.565 ;
        RECT 112.615 15.245 112.935 15.565 ;
        RECT 113.015 15.245 113.335 15.565 ;
        RECT 113.415 15.245 113.735 15.565 ;
        RECT 113.815 15.245 114.135 15.565 ;
        RECT 114.215 15.245 114.535 15.565 ;
        RECT 114.615 15.245 114.935 15.565 ;
        RECT 115.015 15.245 115.335 15.565 ;
        RECT 115.415 15.245 115.735 15.565 ;
        RECT 115.815 15.245 116.135 15.565 ;
        RECT 116.215 15.245 116.535 15.565 ;
        RECT 116.615 15.245 116.935 15.565 ;
        RECT 117.015 15.245 117.335 15.565 ;
        RECT 117.415 15.245 117.735 15.565 ;
        RECT 117.815 15.245 118.135 15.565 ;
        RECT 118.215 15.245 118.535 15.565 ;
        RECT 118.615 15.245 118.935 15.565 ;
        RECT 119.015 15.245 119.335 15.565 ;
        RECT 119.415 15.245 119.735 15.565 ;
        RECT 119.815 15.245 120.135 15.565 ;
        RECT 120.215 15.245 120.535 15.565 ;
        RECT 120.615 15.245 120.935 15.565 ;
        RECT 121.015 15.245 121.335 15.565 ;
        RECT 121.415 15.245 121.735 15.565 ;
        RECT 121.815 15.245 122.135 15.565 ;
        RECT 122.215 15.245 122.535 15.565 ;
        RECT 124.505 15.245 124.825 15.565 ;
        RECT 124.905 15.245 125.225 15.565 ;
        RECT 125.305 15.245 125.625 15.565 ;
        RECT 125.705 15.245 126.025 15.565 ;
        RECT 126.105 15.245 126.425 15.565 ;
        RECT 126.505 15.245 126.825 15.565 ;
        RECT 126.905 15.245 127.225 15.565 ;
        RECT 127.305 15.245 127.625 15.565 ;
        RECT 127.705 15.245 128.025 15.565 ;
        RECT 128.105 15.245 128.425 15.565 ;
        RECT 128.505 15.245 128.825 15.565 ;
        RECT 128.905 15.245 129.225 15.565 ;
        RECT 129.305 15.245 129.625 15.565 ;
        RECT 129.705 15.245 130.025 15.565 ;
        RECT 130.105 15.245 130.425 15.565 ;
        RECT 130.505 15.245 130.825 15.565 ;
        RECT 130.905 15.245 131.225 15.565 ;
        RECT 131.305 15.245 131.625 15.565 ;
        RECT 131.705 15.245 132.025 15.565 ;
        RECT 132.105 15.245 132.425 15.565 ;
        RECT 132.505 15.245 132.825 15.565 ;
        RECT 132.905 15.245 133.225 15.565 ;
        RECT 133.305 15.245 133.625 15.565 ;
        RECT 133.705 15.245 134.025 15.565 ;
        RECT 134.105 15.245 134.425 15.565 ;
        RECT 134.505 15.245 134.825 15.565 ;
        RECT 134.905 15.245 135.225 15.565 ;
        RECT 135.305 15.245 135.625 15.565 ;
        RECT 137.595 15.225 137.915 15.545 ;
        RECT 137.995 15.225 138.315 15.545 ;
        RECT 138.395 15.225 138.715 15.545 ;
        RECT 138.795 15.225 139.115 15.545 ;
        RECT 139.195 15.225 139.515 15.545 ;
        RECT 139.595 15.225 139.915 15.545 ;
        RECT 139.995 15.225 140.315 15.545 ;
        RECT 140.395 15.225 140.715 15.545 ;
        RECT 140.795 15.225 141.115 15.545 ;
        RECT 141.195 15.225 141.515 15.545 ;
        RECT 141.595 15.225 141.915 15.545 ;
        RECT 141.995 15.225 142.315 15.545 ;
        RECT 142.395 15.225 142.715 15.545 ;
        RECT 142.795 15.225 143.115 15.545 ;
        RECT 143.195 15.225 143.515 15.545 ;
        RECT 143.595 15.225 143.915 15.545 ;
        RECT 143.995 15.225 144.315 15.545 ;
        RECT 144.395 15.225 144.715 15.545 ;
        RECT 144.795 15.225 145.115 15.545 ;
        RECT 145.195 15.225 145.515 15.545 ;
        RECT 145.595 15.225 145.915 15.545 ;
        RECT 145.995 15.225 146.315 15.545 ;
        RECT 146.395 15.225 146.715 15.545 ;
        RECT 146.795 15.225 147.115 15.545 ;
        RECT 147.195 15.225 147.515 15.545 ;
        RECT 147.595 15.225 147.915 15.545 ;
        RECT 147.995 15.225 148.315 15.545 ;
        RECT 148.395 15.225 148.715 15.545 ;
        RECT 150.685 15.225 151.005 15.545 ;
        RECT 151.085 15.225 151.405 15.545 ;
        RECT 151.485 15.225 151.805 15.545 ;
        RECT 151.885 15.225 152.205 15.545 ;
        RECT 152.285 15.225 152.605 15.545 ;
        RECT 152.685 15.225 153.005 15.545 ;
        RECT 153.085 15.225 153.405 15.545 ;
        RECT 153.485 15.225 153.805 15.545 ;
        RECT 153.885 15.225 154.205 15.545 ;
        RECT 154.285 15.225 154.605 15.545 ;
        RECT 154.685 15.225 155.005 15.545 ;
        RECT 155.085 15.225 155.405 15.545 ;
        RECT 155.485 15.225 155.805 15.545 ;
        RECT 155.885 15.225 156.205 15.545 ;
        RECT 156.285 15.225 156.605 15.545 ;
        RECT 156.685 15.225 157.005 15.545 ;
        RECT 157.085 15.225 157.405 15.545 ;
        RECT 157.485 15.225 157.805 15.545 ;
        RECT 157.885 15.225 158.205 15.545 ;
        RECT 158.285 15.225 158.605 15.545 ;
        RECT 158.685 15.225 159.005 15.545 ;
        RECT 159.085 15.225 159.405 15.545 ;
        RECT 159.485 15.225 159.805 15.545 ;
        RECT 159.885 15.225 160.205 15.545 ;
        RECT 160.285 15.225 160.605 15.545 ;
        RECT 160.685 15.225 161.005 15.545 ;
        RECT 161.085 15.225 161.405 15.545 ;
        RECT 161.485 15.225 161.805 15.545 ;
        RECT 6.765 13.235 7.085 13.555 ;
        RECT 7.165 13.235 7.485 13.555 ;
        RECT 7.565 13.235 7.885 13.555 ;
        RECT 7.965 13.235 8.285 13.555 ;
        RECT 8.365 13.235 8.685 13.555 ;
        RECT 8.765 13.235 9.085 13.555 ;
        RECT 9.165 13.235 9.485 13.555 ;
        RECT 9.565 13.235 9.885 13.555 ;
        RECT 9.965 13.235 10.285 13.555 ;
        RECT 10.365 13.235 10.685 13.555 ;
        RECT 10.765 13.235 11.085 13.555 ;
        RECT 11.165 13.235 11.485 13.555 ;
        RECT 11.565 13.235 11.885 13.555 ;
        RECT 11.965 13.235 12.285 13.555 ;
        RECT 12.365 13.235 12.685 13.555 ;
        RECT 12.765 13.235 13.085 13.555 ;
        RECT 13.165 13.235 13.485 13.555 ;
        RECT 13.565 13.235 13.885 13.555 ;
        RECT 13.965 13.235 14.285 13.555 ;
        RECT 14.365 13.235 14.685 13.555 ;
        RECT 14.765 13.235 15.085 13.555 ;
        RECT 15.165 13.235 15.485 13.555 ;
        RECT 15.565 13.235 15.885 13.555 ;
        RECT 15.965 13.235 16.285 13.555 ;
        RECT 16.365 13.235 16.685 13.555 ;
        RECT 16.765 13.235 17.085 13.555 ;
        RECT 17.165 13.235 17.485 13.555 ;
        RECT 17.565 13.235 17.885 13.555 ;
        RECT 19.855 13.235 20.175 13.555 ;
        RECT 20.255 13.235 20.575 13.555 ;
        RECT 20.655 13.235 20.975 13.555 ;
        RECT 21.055 13.235 21.375 13.555 ;
        RECT 21.455 13.235 21.775 13.555 ;
        RECT 21.855 13.235 22.175 13.555 ;
        RECT 22.255 13.235 22.575 13.555 ;
        RECT 22.655 13.235 22.975 13.555 ;
        RECT 23.055 13.235 23.375 13.555 ;
        RECT 23.455 13.235 23.775 13.555 ;
        RECT 23.855 13.235 24.175 13.555 ;
        RECT 24.255 13.235 24.575 13.555 ;
        RECT 24.655 13.235 24.975 13.555 ;
        RECT 25.055 13.235 25.375 13.555 ;
        RECT 25.455 13.235 25.775 13.555 ;
        RECT 25.855 13.235 26.175 13.555 ;
        RECT 26.255 13.235 26.575 13.555 ;
        RECT 26.655 13.235 26.975 13.555 ;
        RECT 27.055 13.235 27.375 13.555 ;
        RECT 27.455 13.235 27.775 13.555 ;
        RECT 27.855 13.235 28.175 13.555 ;
        RECT 28.255 13.235 28.575 13.555 ;
        RECT 28.655 13.235 28.975 13.555 ;
        RECT 29.055 13.235 29.375 13.555 ;
        RECT 29.455 13.235 29.775 13.555 ;
        RECT 29.855 13.235 30.175 13.555 ;
        RECT 30.255 13.235 30.575 13.555 ;
        RECT 30.655 13.235 30.975 13.555 ;
        RECT 32.945 13.255 33.265 13.575 ;
        RECT 33.345 13.255 33.665 13.575 ;
        RECT 33.745 13.255 34.065 13.575 ;
        RECT 34.145 13.255 34.465 13.575 ;
        RECT 34.545 13.255 34.865 13.575 ;
        RECT 34.945 13.255 35.265 13.575 ;
        RECT 35.345 13.255 35.665 13.575 ;
        RECT 35.745 13.255 36.065 13.575 ;
        RECT 36.145 13.255 36.465 13.575 ;
        RECT 36.545 13.255 36.865 13.575 ;
        RECT 36.945 13.255 37.265 13.575 ;
        RECT 37.345 13.255 37.665 13.575 ;
        RECT 37.745 13.255 38.065 13.575 ;
        RECT 38.145 13.255 38.465 13.575 ;
        RECT 38.545 13.255 38.865 13.575 ;
        RECT 38.945 13.255 39.265 13.575 ;
        RECT 39.345 13.255 39.665 13.575 ;
        RECT 39.745 13.255 40.065 13.575 ;
        RECT 40.145 13.255 40.465 13.575 ;
        RECT 40.545 13.255 40.865 13.575 ;
        RECT 40.945 13.255 41.265 13.575 ;
        RECT 41.345 13.255 41.665 13.575 ;
        RECT 41.745 13.255 42.065 13.575 ;
        RECT 42.145 13.255 42.465 13.575 ;
        RECT 42.545 13.255 42.865 13.575 ;
        RECT 42.945 13.255 43.265 13.575 ;
        RECT 43.345 13.255 43.665 13.575 ;
        RECT 43.745 13.255 44.065 13.575 ;
        RECT 46.035 13.255 46.355 13.575 ;
        RECT 46.435 13.255 46.755 13.575 ;
        RECT 46.835 13.255 47.155 13.575 ;
        RECT 47.235 13.255 47.555 13.575 ;
        RECT 47.635 13.255 47.955 13.575 ;
        RECT 48.035 13.255 48.355 13.575 ;
        RECT 48.435 13.255 48.755 13.575 ;
        RECT 48.835 13.255 49.155 13.575 ;
        RECT 49.235 13.255 49.555 13.575 ;
        RECT 49.635 13.255 49.955 13.575 ;
        RECT 50.035 13.255 50.355 13.575 ;
        RECT 50.435 13.255 50.755 13.575 ;
        RECT 50.835 13.255 51.155 13.575 ;
        RECT 51.235 13.255 51.555 13.575 ;
        RECT 51.635 13.255 51.955 13.575 ;
        RECT 52.035 13.255 52.355 13.575 ;
        RECT 52.435 13.255 52.755 13.575 ;
        RECT 52.835 13.255 53.155 13.575 ;
        RECT 53.235 13.255 53.555 13.575 ;
        RECT 53.635 13.255 53.955 13.575 ;
        RECT 54.035 13.255 54.355 13.575 ;
        RECT 54.435 13.255 54.755 13.575 ;
        RECT 54.835 13.255 55.155 13.575 ;
        RECT 55.235 13.255 55.555 13.575 ;
        RECT 55.635 13.255 55.955 13.575 ;
        RECT 56.035 13.255 56.355 13.575 ;
        RECT 56.435 13.255 56.755 13.575 ;
        RECT 56.835 13.255 57.155 13.575 ;
        RECT 59.085 13.255 59.405 13.575 ;
        RECT 59.485 13.255 59.805 13.575 ;
        RECT 59.885 13.255 60.205 13.575 ;
        RECT 60.285 13.255 60.605 13.575 ;
        RECT 60.685 13.255 61.005 13.575 ;
        RECT 61.085 13.255 61.405 13.575 ;
        RECT 61.485 13.255 61.805 13.575 ;
        RECT 61.885 13.255 62.205 13.575 ;
        RECT 62.285 13.255 62.605 13.575 ;
        RECT 62.685 13.255 63.005 13.575 ;
        RECT 63.085 13.255 63.405 13.575 ;
        RECT 63.485 13.255 63.805 13.575 ;
        RECT 63.885 13.255 64.205 13.575 ;
        RECT 64.285 13.255 64.605 13.575 ;
        RECT 64.685 13.255 65.005 13.575 ;
        RECT 65.085 13.255 65.405 13.575 ;
        RECT 65.485 13.255 65.805 13.575 ;
        RECT 65.885 13.255 66.205 13.575 ;
        RECT 66.285 13.255 66.605 13.575 ;
        RECT 66.685 13.255 67.005 13.575 ;
        RECT 67.085 13.255 67.405 13.575 ;
        RECT 67.485 13.255 67.805 13.575 ;
        RECT 67.885 13.255 68.205 13.575 ;
        RECT 68.285 13.255 68.605 13.575 ;
        RECT 68.685 13.255 69.005 13.575 ;
        RECT 69.085 13.255 69.405 13.575 ;
        RECT 69.485 13.255 69.805 13.575 ;
        RECT 69.885 13.255 70.205 13.575 ;
        RECT 72.175 13.255 72.495 13.575 ;
        RECT 72.575 13.255 72.895 13.575 ;
        RECT 72.975 13.255 73.295 13.575 ;
        RECT 73.375 13.255 73.695 13.575 ;
        RECT 73.775 13.255 74.095 13.575 ;
        RECT 74.175 13.255 74.495 13.575 ;
        RECT 74.575 13.255 74.895 13.575 ;
        RECT 74.975 13.255 75.295 13.575 ;
        RECT 75.375 13.255 75.695 13.575 ;
        RECT 75.775 13.255 76.095 13.575 ;
        RECT 76.175 13.255 76.495 13.575 ;
        RECT 76.575 13.255 76.895 13.575 ;
        RECT 76.975 13.255 77.295 13.575 ;
        RECT 77.375 13.255 77.695 13.575 ;
        RECT 77.775 13.255 78.095 13.575 ;
        RECT 78.175 13.255 78.495 13.575 ;
        RECT 78.575 13.255 78.895 13.575 ;
        RECT 78.975 13.255 79.295 13.575 ;
        RECT 79.375 13.255 79.695 13.575 ;
        RECT 79.775 13.255 80.095 13.575 ;
        RECT 80.175 13.255 80.495 13.575 ;
        RECT 80.575 13.255 80.895 13.575 ;
        RECT 80.975 13.255 81.295 13.575 ;
        RECT 81.375 13.255 81.695 13.575 ;
        RECT 81.775 13.255 82.095 13.575 ;
        RECT 82.175 13.255 82.495 13.575 ;
        RECT 82.575 13.255 82.895 13.575 ;
        RECT 82.975 13.255 83.295 13.575 ;
        RECT 85.265 13.275 85.585 13.595 ;
        RECT 85.665 13.275 85.985 13.595 ;
        RECT 86.065 13.275 86.385 13.595 ;
        RECT 86.465 13.275 86.785 13.595 ;
        RECT 86.865 13.275 87.185 13.595 ;
        RECT 87.265 13.275 87.585 13.595 ;
        RECT 87.665 13.275 87.985 13.595 ;
        RECT 88.065 13.275 88.385 13.595 ;
        RECT 88.465 13.275 88.785 13.595 ;
        RECT 88.865 13.275 89.185 13.595 ;
        RECT 89.265 13.275 89.585 13.595 ;
        RECT 89.665 13.275 89.985 13.595 ;
        RECT 90.065 13.275 90.385 13.595 ;
        RECT 90.465 13.275 90.785 13.595 ;
        RECT 90.865 13.275 91.185 13.595 ;
        RECT 91.265 13.275 91.585 13.595 ;
        RECT 91.665 13.275 91.985 13.595 ;
        RECT 92.065 13.275 92.385 13.595 ;
        RECT 92.465 13.275 92.785 13.595 ;
        RECT 92.865 13.275 93.185 13.595 ;
        RECT 93.265 13.275 93.585 13.595 ;
        RECT 93.665 13.275 93.985 13.595 ;
        RECT 94.065 13.275 94.385 13.595 ;
        RECT 94.465 13.275 94.785 13.595 ;
        RECT 94.865 13.275 95.185 13.595 ;
        RECT 95.265 13.275 95.585 13.595 ;
        RECT 95.665 13.275 95.985 13.595 ;
        RECT 96.065 13.275 96.385 13.595 ;
        RECT 98.355 13.275 98.675 13.595 ;
        RECT 98.755 13.275 99.075 13.595 ;
        RECT 99.155 13.275 99.475 13.595 ;
        RECT 99.555 13.275 99.875 13.595 ;
        RECT 99.955 13.275 100.275 13.595 ;
        RECT 100.355 13.275 100.675 13.595 ;
        RECT 100.755 13.275 101.075 13.595 ;
        RECT 101.155 13.275 101.475 13.595 ;
        RECT 101.555 13.275 101.875 13.595 ;
        RECT 101.955 13.275 102.275 13.595 ;
        RECT 102.355 13.275 102.675 13.595 ;
        RECT 102.755 13.275 103.075 13.595 ;
        RECT 103.155 13.275 103.475 13.595 ;
        RECT 103.555 13.275 103.875 13.595 ;
        RECT 103.955 13.275 104.275 13.595 ;
        RECT 104.355 13.275 104.675 13.595 ;
        RECT 104.755 13.275 105.075 13.595 ;
        RECT 105.155 13.275 105.475 13.595 ;
        RECT 105.555 13.275 105.875 13.595 ;
        RECT 105.955 13.275 106.275 13.595 ;
        RECT 106.355 13.275 106.675 13.595 ;
        RECT 106.755 13.275 107.075 13.595 ;
        RECT 107.155 13.275 107.475 13.595 ;
        RECT 107.555 13.275 107.875 13.595 ;
        RECT 107.955 13.275 108.275 13.595 ;
        RECT 108.355 13.275 108.675 13.595 ;
        RECT 108.755 13.275 109.075 13.595 ;
        RECT 109.155 13.275 109.475 13.595 ;
        RECT 111.445 13.275 111.765 13.595 ;
        RECT 111.845 13.275 112.165 13.595 ;
        RECT 112.245 13.275 112.565 13.595 ;
        RECT 112.645 13.275 112.965 13.595 ;
        RECT 113.045 13.275 113.365 13.595 ;
        RECT 113.445 13.275 113.765 13.595 ;
        RECT 113.845 13.275 114.165 13.595 ;
        RECT 114.245 13.275 114.565 13.595 ;
        RECT 114.645 13.275 114.965 13.595 ;
        RECT 115.045 13.275 115.365 13.595 ;
        RECT 115.445 13.275 115.765 13.595 ;
        RECT 115.845 13.275 116.165 13.595 ;
        RECT 116.245 13.275 116.565 13.595 ;
        RECT 116.645 13.275 116.965 13.595 ;
        RECT 117.045 13.275 117.365 13.595 ;
        RECT 117.445 13.275 117.765 13.595 ;
        RECT 117.845 13.275 118.165 13.595 ;
        RECT 118.245 13.275 118.565 13.595 ;
        RECT 118.645 13.275 118.965 13.595 ;
        RECT 119.045 13.275 119.365 13.595 ;
        RECT 119.445 13.275 119.765 13.595 ;
        RECT 119.845 13.275 120.165 13.595 ;
        RECT 120.245 13.275 120.565 13.595 ;
        RECT 120.645 13.275 120.965 13.595 ;
        RECT 121.045 13.275 121.365 13.595 ;
        RECT 121.445 13.275 121.765 13.595 ;
        RECT 121.845 13.275 122.165 13.595 ;
        RECT 122.245 13.275 122.565 13.595 ;
        RECT 124.535 13.275 124.855 13.595 ;
        RECT 124.935 13.275 125.255 13.595 ;
        RECT 125.335 13.275 125.655 13.595 ;
        RECT 125.735 13.275 126.055 13.595 ;
        RECT 126.135 13.275 126.455 13.595 ;
        RECT 126.535 13.275 126.855 13.595 ;
        RECT 126.935 13.275 127.255 13.595 ;
        RECT 127.335 13.275 127.655 13.595 ;
        RECT 127.735 13.275 128.055 13.595 ;
        RECT 128.135 13.275 128.455 13.595 ;
        RECT 128.535 13.275 128.855 13.595 ;
        RECT 128.935 13.275 129.255 13.595 ;
        RECT 129.335 13.275 129.655 13.595 ;
        RECT 129.735 13.275 130.055 13.595 ;
        RECT 130.135 13.275 130.455 13.595 ;
        RECT 130.535 13.275 130.855 13.595 ;
        RECT 130.935 13.275 131.255 13.595 ;
        RECT 131.335 13.275 131.655 13.595 ;
        RECT 131.735 13.275 132.055 13.595 ;
        RECT 132.135 13.275 132.455 13.595 ;
        RECT 132.535 13.275 132.855 13.595 ;
        RECT 132.935 13.275 133.255 13.595 ;
        RECT 133.335 13.275 133.655 13.595 ;
        RECT 133.735 13.275 134.055 13.595 ;
        RECT 134.135 13.275 134.455 13.595 ;
        RECT 134.535 13.275 134.855 13.595 ;
        RECT 134.935 13.275 135.255 13.595 ;
        RECT 135.335 13.275 135.655 13.595 ;
        RECT 137.625 13.295 137.945 13.615 ;
        RECT 138.025 13.295 138.345 13.615 ;
        RECT 138.425 13.295 138.745 13.615 ;
        RECT 138.825 13.295 139.145 13.615 ;
        RECT 139.225 13.295 139.545 13.615 ;
        RECT 139.625 13.295 139.945 13.615 ;
        RECT 140.025 13.295 140.345 13.615 ;
        RECT 140.425 13.295 140.745 13.615 ;
        RECT 140.825 13.295 141.145 13.615 ;
        RECT 141.225 13.295 141.545 13.615 ;
        RECT 141.625 13.295 141.945 13.615 ;
        RECT 142.025 13.295 142.345 13.615 ;
        RECT 142.425 13.295 142.745 13.615 ;
        RECT 142.825 13.295 143.145 13.615 ;
        RECT 143.225 13.295 143.545 13.615 ;
        RECT 143.625 13.295 143.945 13.615 ;
        RECT 144.025 13.295 144.345 13.615 ;
        RECT 144.425 13.295 144.745 13.615 ;
        RECT 144.825 13.295 145.145 13.615 ;
        RECT 145.225 13.295 145.545 13.615 ;
        RECT 145.625 13.295 145.945 13.615 ;
        RECT 146.025 13.295 146.345 13.615 ;
        RECT 146.425 13.295 146.745 13.615 ;
        RECT 146.825 13.295 147.145 13.615 ;
        RECT 147.225 13.295 147.545 13.615 ;
        RECT 147.625 13.295 147.945 13.615 ;
        RECT 148.025 13.295 148.345 13.615 ;
        RECT 148.425 13.295 148.745 13.615 ;
        RECT 150.715 13.295 151.035 13.615 ;
        RECT 151.115 13.295 151.435 13.615 ;
        RECT 151.515 13.295 151.835 13.615 ;
        RECT 151.915 13.295 152.235 13.615 ;
        RECT 152.315 13.295 152.635 13.615 ;
        RECT 152.715 13.295 153.035 13.615 ;
        RECT 153.115 13.295 153.435 13.615 ;
        RECT 153.515 13.295 153.835 13.615 ;
        RECT 153.915 13.295 154.235 13.615 ;
        RECT 154.315 13.295 154.635 13.615 ;
        RECT 154.715 13.295 155.035 13.615 ;
        RECT 155.115 13.295 155.435 13.615 ;
        RECT 155.515 13.295 155.835 13.615 ;
        RECT 155.915 13.295 156.235 13.615 ;
        RECT 156.315 13.295 156.635 13.615 ;
        RECT 156.715 13.295 157.035 13.615 ;
        RECT 157.115 13.295 157.435 13.615 ;
        RECT 157.515 13.295 157.835 13.615 ;
        RECT 157.915 13.295 158.235 13.615 ;
        RECT 158.315 13.295 158.635 13.615 ;
        RECT 158.715 13.295 159.035 13.615 ;
        RECT 159.115 13.295 159.435 13.615 ;
        RECT 159.515 13.295 159.835 13.615 ;
        RECT 159.915 13.295 160.235 13.615 ;
        RECT 160.315 13.295 160.635 13.615 ;
        RECT 160.715 13.295 161.035 13.615 ;
        RECT 161.115 13.295 161.435 13.615 ;
        RECT 161.515 13.295 161.835 13.615 ;
      LAYER met4 ;
        RECT 6.155 107.250 6.455 117.980 ;
        RECT 7.355 108.475 7.655 116.755 ;
        RECT 8.555 108.475 8.855 117.980 ;
        RECT 7.355 107.250 8.855 108.475 ;
        RECT 9.755 107.250 10.055 117.980 ;
        RECT 10.955 107.250 11.255 117.980 ;
        RECT 12.155 107.250 12.455 117.980 ;
        RECT 13.355 107.250 13.655 117.980 ;
        RECT 14.555 108.475 14.855 116.755 ;
        RECT 15.755 108.475 16.055 117.980 ;
        RECT 14.555 107.250 16.055 108.475 ;
        RECT 16.955 107.250 17.565 117.980 ;
        RECT 6.155 106.920 17.565 107.250 ;
        RECT 19.245 107.250 19.545 117.980 ;
        RECT 20.445 108.475 20.745 116.755 ;
        RECT 21.645 108.475 21.945 117.980 ;
        RECT 20.445 107.250 21.945 108.475 ;
        RECT 22.845 107.250 23.145 117.980 ;
        RECT 24.045 107.250 24.345 117.980 ;
        RECT 25.245 107.250 25.545 117.980 ;
        RECT 26.445 107.250 26.745 117.980 ;
        RECT 27.645 108.475 27.945 116.755 ;
        RECT 28.845 108.475 29.145 117.980 ;
        RECT 27.645 107.250 29.145 108.475 ;
        RECT 30.045 107.250 30.655 117.980 ;
        RECT 19.245 106.920 30.655 107.250 ;
        RECT 32.335 107.230 32.635 117.960 ;
        RECT 33.535 108.455 33.835 116.735 ;
        RECT 34.735 108.455 35.035 117.960 ;
        RECT 33.535 107.230 35.035 108.455 ;
        RECT 35.935 107.230 36.235 117.960 ;
        RECT 37.135 107.230 37.435 117.960 ;
        RECT 38.335 107.230 38.635 117.960 ;
        RECT 39.535 107.230 39.835 117.960 ;
        RECT 40.735 108.455 41.035 116.735 ;
        RECT 41.935 108.455 42.235 117.960 ;
        RECT 40.735 107.230 42.235 108.455 ;
        RECT 43.135 107.230 43.745 117.960 ;
        RECT 32.335 106.900 43.745 107.230 ;
        RECT 45.425 107.230 45.725 117.960 ;
        RECT 46.625 108.455 46.925 116.735 ;
        RECT 47.825 108.455 48.125 117.960 ;
        RECT 46.625 107.230 48.125 108.455 ;
        RECT 49.025 107.230 49.325 117.960 ;
        RECT 50.225 107.230 50.525 117.960 ;
        RECT 51.425 107.230 51.725 117.960 ;
        RECT 52.625 107.230 52.925 117.960 ;
        RECT 53.825 108.455 54.125 116.735 ;
        RECT 55.025 108.455 55.325 117.960 ;
        RECT 53.825 107.230 55.325 108.455 ;
        RECT 56.225 107.230 56.835 117.960 ;
        RECT 45.425 106.900 56.835 107.230 ;
        RECT 58.475 107.230 58.775 117.960 ;
        RECT 59.675 108.455 59.975 116.735 ;
        RECT 60.875 108.455 61.175 117.960 ;
        RECT 59.675 107.230 61.175 108.455 ;
        RECT 62.075 107.230 62.375 117.960 ;
        RECT 63.275 107.230 63.575 117.960 ;
        RECT 64.475 107.230 64.775 117.960 ;
        RECT 65.675 107.230 65.975 117.960 ;
        RECT 66.875 108.455 67.175 116.735 ;
        RECT 68.075 108.455 68.375 117.960 ;
        RECT 66.875 107.230 68.375 108.455 ;
        RECT 69.275 107.230 69.885 117.960 ;
        RECT 58.475 106.900 69.885 107.230 ;
        RECT 71.565 107.230 71.865 117.960 ;
        RECT 72.765 108.455 73.065 116.735 ;
        RECT 73.965 108.455 74.265 117.960 ;
        RECT 72.765 107.230 74.265 108.455 ;
        RECT 75.165 107.230 75.465 117.960 ;
        RECT 76.365 107.230 76.665 117.960 ;
        RECT 77.565 107.230 77.865 117.960 ;
        RECT 78.765 107.230 79.065 117.960 ;
        RECT 79.965 108.455 80.265 116.735 ;
        RECT 81.165 108.455 81.465 117.960 ;
        RECT 79.965 107.230 81.465 108.455 ;
        RECT 82.365 107.230 82.975 117.960 ;
        RECT 71.565 106.900 82.975 107.230 ;
        RECT 84.655 107.210 84.955 117.940 ;
        RECT 85.855 108.435 86.155 116.715 ;
        RECT 87.055 108.435 87.355 117.940 ;
        RECT 85.855 107.210 87.355 108.435 ;
        RECT 88.255 107.210 88.555 117.940 ;
        RECT 89.455 107.210 89.755 117.940 ;
        RECT 90.655 107.210 90.955 117.940 ;
        RECT 91.855 107.210 92.155 117.940 ;
        RECT 93.055 108.435 93.355 116.715 ;
        RECT 94.255 108.435 94.555 117.940 ;
        RECT 93.055 107.210 94.555 108.435 ;
        RECT 95.455 107.210 96.065 117.940 ;
        RECT 84.655 106.880 96.065 107.210 ;
        RECT 97.745 107.210 98.045 117.940 ;
        RECT 98.945 108.435 99.245 116.715 ;
        RECT 100.145 108.435 100.445 117.940 ;
        RECT 98.945 107.210 100.445 108.435 ;
        RECT 101.345 107.210 101.645 117.940 ;
        RECT 102.545 107.210 102.845 117.940 ;
        RECT 103.745 107.210 104.045 117.940 ;
        RECT 104.945 107.210 105.245 117.940 ;
        RECT 106.145 108.435 106.445 116.715 ;
        RECT 107.345 108.435 107.645 117.940 ;
        RECT 106.145 107.210 107.645 108.435 ;
        RECT 108.545 107.210 109.155 117.940 ;
        RECT 97.745 106.880 109.155 107.210 ;
        RECT 110.835 107.210 111.135 117.940 ;
        RECT 112.035 108.435 112.335 116.715 ;
        RECT 113.235 108.435 113.535 117.940 ;
        RECT 112.035 107.210 113.535 108.435 ;
        RECT 114.435 107.210 114.735 117.940 ;
        RECT 115.635 107.210 115.935 117.940 ;
        RECT 116.835 107.210 117.135 117.940 ;
        RECT 118.035 107.210 118.335 117.940 ;
        RECT 119.235 108.435 119.535 116.715 ;
        RECT 120.435 108.435 120.735 117.940 ;
        RECT 119.235 107.210 120.735 108.435 ;
        RECT 121.635 107.210 122.245 117.940 ;
        RECT 110.835 106.880 122.245 107.210 ;
        RECT 123.925 107.210 124.225 117.940 ;
        RECT 125.125 108.435 125.425 116.715 ;
        RECT 126.325 108.435 126.625 117.940 ;
        RECT 125.125 107.210 126.625 108.435 ;
        RECT 127.525 107.210 127.825 117.940 ;
        RECT 128.725 107.210 129.025 117.940 ;
        RECT 129.925 107.210 130.225 117.940 ;
        RECT 131.125 107.210 131.425 117.940 ;
        RECT 132.325 108.435 132.625 116.715 ;
        RECT 133.525 108.435 133.825 117.940 ;
        RECT 132.325 107.210 133.825 108.435 ;
        RECT 134.725 107.210 135.335 117.940 ;
        RECT 123.925 106.880 135.335 107.210 ;
        RECT 137.015 107.190 137.315 117.920 ;
        RECT 138.215 108.415 138.515 116.695 ;
        RECT 139.415 108.415 139.715 117.920 ;
        RECT 138.215 107.190 139.715 108.415 ;
        RECT 140.615 107.190 140.915 117.920 ;
        RECT 141.815 107.190 142.115 117.920 ;
        RECT 143.015 107.190 143.315 117.920 ;
        RECT 144.215 107.190 144.515 117.920 ;
        RECT 145.415 108.415 145.715 116.695 ;
        RECT 146.615 108.415 146.915 117.920 ;
        RECT 145.415 107.190 146.915 108.415 ;
        RECT 147.815 107.190 148.425 117.920 ;
        RECT 137.015 106.860 148.425 107.190 ;
        RECT 150.105 107.190 150.405 117.920 ;
        RECT 151.305 108.415 151.605 116.695 ;
        RECT 152.505 108.415 152.805 117.920 ;
        RECT 151.305 107.190 152.805 108.415 ;
        RECT 153.705 107.190 154.005 117.920 ;
        RECT 154.905 107.190 155.205 117.920 ;
        RECT 156.105 107.190 156.405 117.920 ;
        RECT 157.305 107.190 157.605 117.920 ;
        RECT 158.505 108.415 158.805 116.695 ;
        RECT 159.705 108.415 160.005 117.920 ;
        RECT 158.505 107.190 160.005 108.415 ;
        RECT 160.905 107.190 161.515 117.920 ;
        RECT 150.105 106.860 161.515 107.190 ;
        RECT 4.235 105.180 5.835 106.780 ;
        RECT 162.345 105.380 163.945 106.980 ;
        RECT 4.435 15.390 5.635 105.180 ;
        RECT 6.185 104.870 17.595 105.200 ;
        RECT 6.185 94.140 6.485 104.870 ;
        RECT 7.385 103.645 8.885 104.870 ;
        RECT 7.385 95.365 7.685 103.645 ;
        RECT 8.585 94.140 8.885 103.645 ;
        RECT 9.785 94.140 10.085 104.870 ;
        RECT 10.985 94.140 11.285 104.870 ;
        RECT 12.185 94.140 12.485 104.870 ;
        RECT 13.385 94.140 13.685 104.870 ;
        RECT 14.585 103.645 16.085 104.870 ;
        RECT 14.585 95.365 14.885 103.645 ;
        RECT 15.785 94.140 16.085 103.645 ;
        RECT 16.985 94.140 17.595 104.870 ;
        RECT 19.275 104.870 30.685 105.200 ;
        RECT 19.275 94.140 19.575 104.870 ;
        RECT 20.475 103.645 21.975 104.870 ;
        RECT 20.475 95.365 20.775 103.645 ;
        RECT 21.675 94.140 21.975 103.645 ;
        RECT 22.875 94.140 23.175 104.870 ;
        RECT 24.075 94.140 24.375 104.870 ;
        RECT 25.275 94.140 25.575 104.870 ;
        RECT 26.475 94.140 26.775 104.870 ;
        RECT 27.675 103.645 29.175 104.870 ;
        RECT 27.675 95.365 27.975 103.645 ;
        RECT 28.875 94.140 29.175 103.645 ;
        RECT 30.075 94.140 30.685 104.870 ;
        RECT 32.365 104.890 43.775 105.220 ;
        RECT 32.365 94.160 32.665 104.890 ;
        RECT 33.565 103.665 35.065 104.890 ;
        RECT 33.565 95.385 33.865 103.665 ;
        RECT 34.765 94.160 35.065 103.665 ;
        RECT 35.965 94.160 36.265 104.890 ;
        RECT 37.165 94.160 37.465 104.890 ;
        RECT 38.365 94.160 38.665 104.890 ;
        RECT 39.565 94.160 39.865 104.890 ;
        RECT 40.765 103.665 42.265 104.890 ;
        RECT 40.765 95.385 41.065 103.665 ;
        RECT 41.965 94.160 42.265 103.665 ;
        RECT 43.165 94.160 43.775 104.890 ;
        RECT 45.455 104.890 56.865 105.220 ;
        RECT 45.455 94.160 45.755 104.890 ;
        RECT 46.655 103.665 48.155 104.890 ;
        RECT 46.655 95.385 46.955 103.665 ;
        RECT 47.855 94.160 48.155 103.665 ;
        RECT 49.055 94.160 49.355 104.890 ;
        RECT 50.255 94.160 50.555 104.890 ;
        RECT 51.455 94.160 51.755 104.890 ;
        RECT 52.655 94.160 52.955 104.890 ;
        RECT 53.855 103.665 55.355 104.890 ;
        RECT 53.855 95.385 54.155 103.665 ;
        RECT 55.055 94.160 55.355 103.665 ;
        RECT 56.255 94.160 56.865 104.890 ;
        RECT 58.505 104.890 69.915 105.220 ;
        RECT 58.505 94.160 58.805 104.890 ;
        RECT 59.705 103.665 61.205 104.890 ;
        RECT 59.705 95.385 60.005 103.665 ;
        RECT 60.905 94.160 61.205 103.665 ;
        RECT 62.105 94.160 62.405 104.890 ;
        RECT 63.305 94.160 63.605 104.890 ;
        RECT 64.505 94.160 64.805 104.890 ;
        RECT 65.705 94.160 66.005 104.890 ;
        RECT 66.905 103.665 68.405 104.890 ;
        RECT 66.905 95.385 67.205 103.665 ;
        RECT 68.105 94.160 68.405 103.665 ;
        RECT 69.305 94.160 69.915 104.890 ;
        RECT 71.595 104.890 83.005 105.220 ;
        RECT 71.595 94.160 71.895 104.890 ;
        RECT 72.795 103.665 74.295 104.890 ;
        RECT 72.795 95.385 73.095 103.665 ;
        RECT 73.995 94.160 74.295 103.665 ;
        RECT 75.195 94.160 75.495 104.890 ;
        RECT 76.395 94.160 76.695 104.890 ;
        RECT 77.595 94.160 77.895 104.890 ;
        RECT 78.795 94.160 79.095 104.890 ;
        RECT 79.995 103.665 81.495 104.890 ;
        RECT 79.995 95.385 80.295 103.665 ;
        RECT 81.195 94.160 81.495 103.665 ;
        RECT 82.395 94.160 83.005 104.890 ;
        RECT 84.685 104.910 96.095 105.240 ;
        RECT 84.685 94.180 84.985 104.910 ;
        RECT 85.885 103.685 87.385 104.910 ;
        RECT 85.885 95.405 86.185 103.685 ;
        RECT 87.085 94.180 87.385 103.685 ;
        RECT 88.285 94.180 88.585 104.910 ;
        RECT 89.485 94.180 89.785 104.910 ;
        RECT 90.685 94.180 90.985 104.910 ;
        RECT 91.885 94.180 92.185 104.910 ;
        RECT 93.085 103.685 94.585 104.910 ;
        RECT 93.085 95.405 93.385 103.685 ;
        RECT 94.285 94.180 94.585 103.685 ;
        RECT 95.485 94.180 96.095 104.910 ;
        RECT 97.775 104.910 109.185 105.240 ;
        RECT 97.775 94.180 98.075 104.910 ;
        RECT 98.975 103.685 100.475 104.910 ;
        RECT 98.975 95.405 99.275 103.685 ;
        RECT 100.175 94.180 100.475 103.685 ;
        RECT 101.375 94.180 101.675 104.910 ;
        RECT 102.575 94.180 102.875 104.910 ;
        RECT 103.775 94.180 104.075 104.910 ;
        RECT 104.975 94.180 105.275 104.910 ;
        RECT 106.175 103.685 107.675 104.910 ;
        RECT 106.175 95.405 106.475 103.685 ;
        RECT 107.375 94.180 107.675 103.685 ;
        RECT 108.575 94.180 109.185 104.910 ;
        RECT 110.865 104.910 122.275 105.240 ;
        RECT 110.865 94.180 111.165 104.910 ;
        RECT 112.065 103.685 113.565 104.910 ;
        RECT 112.065 95.405 112.365 103.685 ;
        RECT 113.265 94.180 113.565 103.685 ;
        RECT 114.465 94.180 114.765 104.910 ;
        RECT 115.665 94.180 115.965 104.910 ;
        RECT 116.865 94.180 117.165 104.910 ;
        RECT 118.065 94.180 118.365 104.910 ;
        RECT 119.265 103.685 120.765 104.910 ;
        RECT 119.265 95.405 119.565 103.685 ;
        RECT 120.465 94.180 120.765 103.685 ;
        RECT 121.665 94.180 122.275 104.910 ;
        RECT 123.955 104.910 135.365 105.240 ;
        RECT 123.955 94.180 124.255 104.910 ;
        RECT 125.155 103.685 126.655 104.910 ;
        RECT 125.155 95.405 125.455 103.685 ;
        RECT 126.355 94.180 126.655 103.685 ;
        RECT 127.555 94.180 127.855 104.910 ;
        RECT 128.755 94.180 129.055 104.910 ;
        RECT 129.955 94.180 130.255 104.910 ;
        RECT 131.155 94.180 131.455 104.910 ;
        RECT 132.355 103.685 133.855 104.910 ;
        RECT 132.355 95.405 132.655 103.685 ;
        RECT 133.555 94.180 133.855 103.685 ;
        RECT 134.755 94.180 135.365 104.910 ;
        RECT 137.045 104.930 148.455 105.260 ;
        RECT 137.045 94.200 137.345 104.930 ;
        RECT 138.245 103.705 139.745 104.930 ;
        RECT 138.245 95.425 138.545 103.705 ;
        RECT 139.445 94.200 139.745 103.705 ;
        RECT 140.645 94.200 140.945 104.930 ;
        RECT 141.845 94.200 142.145 104.930 ;
        RECT 143.045 94.200 143.345 104.930 ;
        RECT 144.245 94.200 144.545 104.930 ;
        RECT 145.445 103.705 146.945 104.930 ;
        RECT 145.445 95.425 145.745 103.705 ;
        RECT 146.645 94.200 146.945 103.705 ;
        RECT 147.845 94.200 148.455 104.930 ;
        RECT 150.135 104.930 161.545 105.260 ;
        RECT 150.135 94.200 150.435 104.930 ;
        RECT 151.335 103.705 152.835 104.930 ;
        RECT 151.335 95.425 151.635 103.705 ;
        RECT 152.535 94.200 152.835 103.705 ;
        RECT 153.735 94.200 154.035 104.930 ;
        RECT 154.935 94.200 155.235 104.930 ;
        RECT 156.135 94.200 156.435 104.930 ;
        RECT 157.335 94.200 157.635 104.930 ;
        RECT 158.535 103.705 160.035 104.930 ;
        RECT 158.535 95.425 158.835 103.705 ;
        RECT 159.735 94.200 160.035 103.705 ;
        RECT 160.935 94.200 161.545 104.930 ;
        RECT 162.545 90.140 163.745 105.380 ;
        RECT 6.595 15.610 6.895 26.340 ;
        RECT 7.795 16.835 8.095 25.115 ;
        RECT 8.995 16.835 9.295 26.340 ;
        RECT 7.795 15.610 9.295 16.835 ;
        RECT 10.195 15.610 10.495 26.340 ;
        RECT 11.395 15.610 11.695 26.340 ;
        RECT 12.595 15.610 12.895 26.340 ;
        RECT 13.795 15.610 14.095 26.340 ;
        RECT 14.995 16.835 15.295 25.115 ;
        RECT 16.195 16.835 16.495 26.340 ;
        RECT 14.995 15.610 16.495 16.835 ;
        RECT 17.395 15.610 18.005 26.340 ;
        RECT 4.235 13.790 5.835 15.390 ;
        RECT 6.595 15.280 18.005 15.610 ;
        RECT 19.685 15.610 19.985 26.340 ;
        RECT 20.885 16.835 21.185 25.115 ;
        RECT 22.085 16.835 22.385 26.340 ;
        RECT 20.885 15.610 22.385 16.835 ;
        RECT 23.285 15.610 23.585 26.340 ;
        RECT 24.485 15.610 24.785 26.340 ;
        RECT 25.685 15.610 25.985 26.340 ;
        RECT 26.885 15.610 27.185 26.340 ;
        RECT 28.085 16.835 28.385 25.115 ;
        RECT 29.285 16.835 29.585 26.340 ;
        RECT 28.085 15.610 29.585 16.835 ;
        RECT 30.485 15.610 31.095 26.340 ;
        RECT 19.685 15.280 31.095 15.610 ;
        RECT 32.775 15.590 33.075 26.320 ;
        RECT 33.975 16.815 34.275 25.095 ;
        RECT 35.175 16.815 35.475 26.320 ;
        RECT 33.975 15.590 35.475 16.815 ;
        RECT 36.375 15.590 36.675 26.320 ;
        RECT 37.575 15.590 37.875 26.320 ;
        RECT 38.775 15.590 39.075 26.320 ;
        RECT 39.975 15.590 40.275 26.320 ;
        RECT 41.175 16.815 41.475 25.095 ;
        RECT 42.375 16.815 42.675 26.320 ;
        RECT 41.175 15.590 42.675 16.815 ;
        RECT 43.575 15.590 44.185 26.320 ;
        RECT 32.775 15.260 44.185 15.590 ;
        RECT 45.865 15.590 46.165 26.320 ;
        RECT 47.065 16.815 47.365 25.095 ;
        RECT 48.265 16.815 48.565 26.320 ;
        RECT 47.065 15.590 48.565 16.815 ;
        RECT 49.465 15.590 49.765 26.320 ;
        RECT 50.665 15.590 50.965 26.320 ;
        RECT 51.865 15.590 52.165 26.320 ;
        RECT 53.065 15.590 53.365 26.320 ;
        RECT 54.265 16.815 54.565 25.095 ;
        RECT 55.465 16.815 55.765 26.320 ;
        RECT 54.265 15.590 55.765 16.815 ;
        RECT 56.665 15.590 57.275 26.320 ;
        RECT 45.865 15.260 57.275 15.590 ;
        RECT 58.915 15.590 59.215 26.320 ;
        RECT 60.115 16.815 60.415 25.095 ;
        RECT 61.315 16.815 61.615 26.320 ;
        RECT 60.115 15.590 61.615 16.815 ;
        RECT 62.515 15.590 62.815 26.320 ;
        RECT 63.715 15.590 64.015 26.320 ;
        RECT 64.915 15.590 65.215 26.320 ;
        RECT 66.115 15.590 66.415 26.320 ;
        RECT 67.315 16.815 67.615 25.095 ;
        RECT 68.515 16.815 68.815 26.320 ;
        RECT 67.315 15.590 68.815 16.815 ;
        RECT 69.715 15.590 70.325 26.320 ;
        RECT 58.915 15.260 70.325 15.590 ;
        RECT 72.005 15.590 72.305 26.320 ;
        RECT 73.205 16.815 73.505 25.095 ;
        RECT 74.405 16.815 74.705 26.320 ;
        RECT 73.205 15.590 74.705 16.815 ;
        RECT 75.605 15.590 75.905 26.320 ;
        RECT 76.805 15.590 77.105 26.320 ;
        RECT 78.005 15.590 78.305 26.320 ;
        RECT 79.205 15.590 79.505 26.320 ;
        RECT 80.405 16.815 80.705 25.095 ;
        RECT 81.605 16.815 81.905 26.320 ;
        RECT 80.405 15.590 81.905 16.815 ;
        RECT 82.805 15.590 83.415 26.320 ;
        RECT 72.005 15.260 83.415 15.590 ;
        RECT 85.095 15.570 85.395 26.300 ;
        RECT 86.295 16.795 86.595 25.075 ;
        RECT 87.495 16.795 87.795 26.300 ;
        RECT 86.295 15.570 87.795 16.795 ;
        RECT 88.695 15.570 88.995 26.300 ;
        RECT 89.895 15.570 90.195 26.300 ;
        RECT 91.095 15.570 91.395 26.300 ;
        RECT 92.295 15.570 92.595 26.300 ;
        RECT 93.495 16.795 93.795 25.075 ;
        RECT 94.695 16.795 94.995 26.300 ;
        RECT 93.495 15.570 94.995 16.795 ;
        RECT 95.895 15.570 96.505 26.300 ;
        RECT 85.095 15.240 96.505 15.570 ;
        RECT 98.185 15.570 98.485 26.300 ;
        RECT 99.385 16.795 99.685 25.075 ;
        RECT 100.585 16.795 100.885 26.300 ;
        RECT 99.385 15.570 100.885 16.795 ;
        RECT 101.785 15.570 102.085 26.300 ;
        RECT 102.985 15.570 103.285 26.300 ;
        RECT 104.185 15.570 104.485 26.300 ;
        RECT 105.385 15.570 105.685 26.300 ;
        RECT 106.585 16.795 106.885 25.075 ;
        RECT 107.785 16.795 108.085 26.300 ;
        RECT 106.585 15.570 108.085 16.795 ;
        RECT 108.985 15.570 109.595 26.300 ;
        RECT 98.185 15.240 109.595 15.570 ;
        RECT 111.275 15.570 111.575 26.300 ;
        RECT 112.475 16.795 112.775 25.075 ;
        RECT 113.675 16.795 113.975 26.300 ;
        RECT 112.475 15.570 113.975 16.795 ;
        RECT 114.875 15.570 115.175 26.300 ;
        RECT 116.075 15.570 116.375 26.300 ;
        RECT 117.275 15.570 117.575 26.300 ;
        RECT 118.475 15.570 118.775 26.300 ;
        RECT 119.675 16.795 119.975 25.075 ;
        RECT 120.875 16.795 121.175 26.300 ;
        RECT 119.675 15.570 121.175 16.795 ;
        RECT 122.075 15.570 122.685 26.300 ;
        RECT 111.275 15.240 122.685 15.570 ;
        RECT 124.365 15.570 124.665 26.300 ;
        RECT 125.565 16.795 125.865 25.075 ;
        RECT 126.765 16.795 127.065 26.300 ;
        RECT 125.565 15.570 127.065 16.795 ;
        RECT 127.965 15.570 128.265 26.300 ;
        RECT 129.165 15.570 129.465 26.300 ;
        RECT 130.365 15.570 130.665 26.300 ;
        RECT 131.565 15.570 131.865 26.300 ;
        RECT 132.765 16.795 133.065 25.075 ;
        RECT 133.965 16.795 134.265 26.300 ;
        RECT 132.765 15.570 134.265 16.795 ;
        RECT 135.165 15.570 135.775 26.300 ;
        RECT 124.365 15.240 135.775 15.570 ;
        RECT 137.455 15.550 137.755 26.280 ;
        RECT 138.655 16.775 138.955 25.055 ;
        RECT 139.855 16.775 140.155 26.280 ;
        RECT 138.655 15.550 140.155 16.775 ;
        RECT 141.055 15.550 141.355 26.280 ;
        RECT 142.255 15.550 142.555 26.280 ;
        RECT 143.455 15.550 143.755 26.280 ;
        RECT 144.655 15.550 144.955 26.280 ;
        RECT 145.855 16.775 146.155 25.055 ;
        RECT 147.055 16.775 147.355 26.280 ;
        RECT 145.855 15.550 147.355 16.775 ;
        RECT 148.255 15.550 148.865 26.280 ;
        RECT 137.455 15.220 148.865 15.550 ;
        RECT 150.545 15.550 150.845 26.280 ;
        RECT 151.745 16.775 152.045 25.055 ;
        RECT 152.945 16.775 153.245 26.280 ;
        RECT 151.745 15.550 153.245 16.775 ;
        RECT 154.145 15.550 154.445 26.280 ;
        RECT 155.345 15.550 155.645 26.280 ;
        RECT 156.545 15.550 156.845 26.280 ;
        RECT 157.745 15.550 158.045 26.280 ;
        RECT 158.945 16.775 159.245 25.055 ;
        RECT 160.145 16.775 160.445 26.280 ;
        RECT 158.945 15.550 160.445 16.775 ;
        RECT 161.345 15.550 161.955 26.280 ;
        RECT 150.545 15.220 161.955 15.550 ;
        RECT 162.975 15.110 164.175 29.920 ;
        RECT 6.625 13.230 18.035 13.560 ;
        RECT 6.625 2.500 6.925 13.230 ;
        RECT 7.825 12.005 9.325 13.230 ;
        RECT 7.825 3.725 8.125 12.005 ;
        RECT 9.025 2.500 9.325 12.005 ;
        RECT 10.225 2.500 10.525 13.230 ;
        RECT 11.425 2.500 11.725 13.230 ;
        RECT 12.625 2.500 12.925 13.230 ;
        RECT 13.825 2.500 14.125 13.230 ;
        RECT 15.025 12.005 16.525 13.230 ;
        RECT 15.025 3.725 15.325 12.005 ;
        RECT 16.225 2.500 16.525 12.005 ;
        RECT 17.425 2.500 18.035 13.230 ;
        RECT 19.715 13.230 31.125 13.560 ;
        RECT 19.715 2.500 20.015 13.230 ;
        RECT 20.915 12.005 22.415 13.230 ;
        RECT 20.915 3.725 21.215 12.005 ;
        RECT 22.115 2.500 22.415 12.005 ;
        RECT 23.315 2.500 23.615 13.230 ;
        RECT 24.515 2.500 24.815 13.230 ;
        RECT 25.715 2.500 26.015 13.230 ;
        RECT 26.915 2.500 27.215 13.230 ;
        RECT 28.115 12.005 29.615 13.230 ;
        RECT 28.115 3.725 28.415 12.005 ;
        RECT 29.315 2.500 29.615 12.005 ;
        RECT 30.515 2.500 31.125 13.230 ;
        RECT 32.805 13.250 44.215 13.580 ;
        RECT 32.805 2.520 33.105 13.250 ;
        RECT 34.005 12.025 35.505 13.250 ;
        RECT 34.005 3.745 34.305 12.025 ;
        RECT 35.205 2.520 35.505 12.025 ;
        RECT 36.405 2.520 36.705 13.250 ;
        RECT 37.605 2.520 37.905 13.250 ;
        RECT 38.805 2.520 39.105 13.250 ;
        RECT 40.005 2.520 40.305 13.250 ;
        RECT 41.205 12.025 42.705 13.250 ;
        RECT 41.205 3.745 41.505 12.025 ;
        RECT 42.405 2.520 42.705 12.025 ;
        RECT 43.605 2.520 44.215 13.250 ;
        RECT 45.895 13.250 57.305 13.580 ;
        RECT 45.895 2.520 46.195 13.250 ;
        RECT 47.095 12.025 48.595 13.250 ;
        RECT 47.095 3.745 47.395 12.025 ;
        RECT 48.295 2.520 48.595 12.025 ;
        RECT 49.495 2.520 49.795 13.250 ;
        RECT 50.695 2.520 50.995 13.250 ;
        RECT 51.895 2.520 52.195 13.250 ;
        RECT 53.095 2.520 53.395 13.250 ;
        RECT 54.295 12.025 55.795 13.250 ;
        RECT 54.295 3.745 54.595 12.025 ;
        RECT 55.495 2.520 55.795 12.025 ;
        RECT 56.695 2.520 57.305 13.250 ;
        RECT 58.945 13.250 70.355 13.580 ;
        RECT 58.945 2.520 59.245 13.250 ;
        RECT 60.145 12.025 61.645 13.250 ;
        RECT 60.145 3.745 60.445 12.025 ;
        RECT 61.345 2.520 61.645 12.025 ;
        RECT 62.545 2.520 62.845 13.250 ;
        RECT 63.745 2.520 64.045 13.250 ;
        RECT 64.945 2.520 65.245 13.250 ;
        RECT 66.145 2.520 66.445 13.250 ;
        RECT 67.345 12.025 68.845 13.250 ;
        RECT 67.345 3.745 67.645 12.025 ;
        RECT 68.545 2.520 68.845 12.025 ;
        RECT 69.745 2.520 70.355 13.250 ;
        RECT 72.035 13.250 83.445 13.580 ;
        RECT 72.035 2.520 72.335 13.250 ;
        RECT 73.235 12.025 74.735 13.250 ;
        RECT 73.235 3.745 73.535 12.025 ;
        RECT 74.435 2.520 74.735 12.025 ;
        RECT 75.635 2.520 75.935 13.250 ;
        RECT 76.835 2.520 77.135 13.250 ;
        RECT 78.035 2.520 78.335 13.250 ;
        RECT 79.235 2.520 79.535 13.250 ;
        RECT 80.435 12.025 81.935 13.250 ;
        RECT 80.435 3.745 80.735 12.025 ;
        RECT 81.635 2.520 81.935 12.025 ;
        RECT 82.835 2.520 83.445 13.250 ;
        RECT 85.125 13.270 96.535 13.600 ;
        RECT 85.125 2.540 85.425 13.270 ;
        RECT 86.325 12.045 87.825 13.270 ;
        RECT 86.325 3.765 86.625 12.045 ;
        RECT 87.525 2.540 87.825 12.045 ;
        RECT 88.725 2.540 89.025 13.270 ;
        RECT 89.925 2.540 90.225 13.270 ;
        RECT 91.125 2.540 91.425 13.270 ;
        RECT 92.325 2.540 92.625 13.270 ;
        RECT 93.525 12.045 95.025 13.270 ;
        RECT 93.525 3.765 93.825 12.045 ;
        RECT 94.725 2.540 95.025 12.045 ;
        RECT 95.925 2.540 96.535 13.270 ;
        RECT 98.215 13.270 109.625 13.600 ;
        RECT 98.215 2.540 98.515 13.270 ;
        RECT 99.415 12.045 100.915 13.270 ;
        RECT 99.415 3.765 99.715 12.045 ;
        RECT 100.615 2.540 100.915 12.045 ;
        RECT 101.815 2.540 102.115 13.270 ;
        RECT 103.015 2.540 103.315 13.270 ;
        RECT 104.215 2.540 104.515 13.270 ;
        RECT 105.415 2.540 105.715 13.270 ;
        RECT 106.615 12.045 108.115 13.270 ;
        RECT 106.615 3.765 106.915 12.045 ;
        RECT 107.815 2.540 108.115 12.045 ;
        RECT 109.015 2.540 109.625 13.270 ;
        RECT 111.305 13.270 122.715 13.600 ;
        RECT 111.305 2.540 111.605 13.270 ;
        RECT 112.505 12.045 114.005 13.270 ;
        RECT 112.505 3.765 112.805 12.045 ;
        RECT 113.705 2.540 114.005 12.045 ;
        RECT 114.905 2.540 115.205 13.270 ;
        RECT 116.105 2.540 116.405 13.270 ;
        RECT 117.305 2.540 117.605 13.270 ;
        RECT 118.505 2.540 118.805 13.270 ;
        RECT 119.705 12.045 121.205 13.270 ;
        RECT 119.705 3.765 120.005 12.045 ;
        RECT 120.905 2.540 121.205 12.045 ;
        RECT 122.105 2.540 122.715 13.270 ;
        RECT 124.395 13.270 135.805 13.600 ;
        RECT 124.395 2.540 124.695 13.270 ;
        RECT 125.595 12.045 127.095 13.270 ;
        RECT 125.595 3.765 125.895 12.045 ;
        RECT 126.795 2.540 127.095 12.045 ;
        RECT 127.995 2.540 128.295 13.270 ;
        RECT 129.195 2.540 129.495 13.270 ;
        RECT 130.395 2.540 130.695 13.270 ;
        RECT 131.595 2.540 131.895 13.270 ;
        RECT 132.795 12.045 134.295 13.270 ;
        RECT 132.795 3.765 133.095 12.045 ;
        RECT 133.995 2.540 134.295 12.045 ;
        RECT 135.195 2.540 135.805 13.270 ;
        RECT 137.485 13.290 148.895 13.620 ;
        RECT 137.485 2.560 137.785 13.290 ;
        RECT 138.685 12.065 140.185 13.290 ;
        RECT 138.685 3.785 138.985 12.065 ;
        RECT 139.885 2.560 140.185 12.065 ;
        RECT 141.085 2.560 141.385 13.290 ;
        RECT 142.285 2.560 142.585 13.290 ;
        RECT 143.485 2.560 143.785 13.290 ;
        RECT 144.685 2.560 144.985 13.290 ;
        RECT 145.885 12.065 147.385 13.290 ;
        RECT 145.885 3.785 146.185 12.065 ;
        RECT 147.085 2.560 147.385 12.065 ;
        RECT 148.285 2.560 148.895 13.290 ;
        RECT 150.575 13.290 161.985 13.620 ;
        RECT 162.775 13.510 164.375 15.110 ;
        RECT 150.575 2.560 150.875 13.290 ;
        RECT 151.775 12.065 153.275 13.290 ;
        RECT 151.775 3.785 152.075 12.065 ;
        RECT 152.975 2.560 153.275 12.065 ;
        RECT 154.175 2.560 154.475 13.290 ;
        RECT 155.375 2.560 155.675 13.290 ;
        RECT 156.575 2.560 156.875 13.290 ;
        RECT 157.775 2.560 158.075 13.290 ;
        RECT 158.975 12.065 160.475 13.290 ;
        RECT 158.975 3.785 159.275 12.065 ;
        RECT 160.175 2.560 160.475 12.065 ;
        RECT 161.375 2.560 161.985 13.290 ;
      LAYER via4 ;
        RECT 7.515 107.295 8.695 108.475 ;
        RECT 14.715 107.295 15.895 108.475 ;
        RECT 20.605 107.295 21.785 108.475 ;
        RECT 27.805 107.295 28.985 108.475 ;
        RECT 33.695 107.275 34.875 108.455 ;
        RECT 40.895 107.275 42.075 108.455 ;
        RECT 46.785 107.275 47.965 108.455 ;
        RECT 53.985 107.275 55.165 108.455 ;
        RECT 59.835 107.275 61.015 108.455 ;
        RECT 67.035 107.275 68.215 108.455 ;
        RECT 72.925 107.275 74.105 108.455 ;
        RECT 80.125 107.275 81.305 108.455 ;
        RECT 86.015 107.255 87.195 108.435 ;
        RECT 93.215 107.255 94.395 108.435 ;
        RECT 99.105 107.255 100.285 108.435 ;
        RECT 106.305 107.255 107.485 108.435 ;
        RECT 112.195 107.255 113.375 108.435 ;
        RECT 119.395 107.255 120.575 108.435 ;
        RECT 125.285 107.255 126.465 108.435 ;
        RECT 132.485 107.255 133.665 108.435 ;
        RECT 138.375 107.235 139.555 108.415 ;
        RECT 145.575 107.235 146.755 108.415 ;
        RECT 151.465 107.235 152.645 108.415 ;
        RECT 158.665 107.235 159.845 108.415 ;
        RECT 7.545 103.645 8.725 104.825 ;
        RECT 14.745 103.645 15.925 104.825 ;
        RECT 20.635 103.645 21.815 104.825 ;
        RECT 27.835 103.645 29.015 104.825 ;
        RECT 33.725 103.665 34.905 104.845 ;
        RECT 40.925 103.665 42.105 104.845 ;
        RECT 46.815 103.665 47.995 104.845 ;
        RECT 54.015 103.665 55.195 104.845 ;
        RECT 59.865 103.665 61.045 104.845 ;
        RECT 67.065 103.665 68.245 104.845 ;
        RECT 72.955 103.665 74.135 104.845 ;
        RECT 80.155 103.665 81.335 104.845 ;
        RECT 86.045 103.685 87.225 104.865 ;
        RECT 93.245 103.685 94.425 104.865 ;
        RECT 99.135 103.685 100.315 104.865 ;
        RECT 106.335 103.685 107.515 104.865 ;
        RECT 112.225 103.685 113.405 104.865 ;
        RECT 119.425 103.685 120.605 104.865 ;
        RECT 125.315 103.685 126.495 104.865 ;
        RECT 132.515 103.685 133.695 104.865 ;
        RECT 138.405 103.705 139.585 104.885 ;
        RECT 145.605 103.705 146.785 104.885 ;
        RECT 151.495 103.705 152.675 104.885 ;
        RECT 158.695 103.705 159.875 104.885 ;
        RECT 7.955 15.655 9.135 16.835 ;
        RECT 15.155 15.655 16.335 16.835 ;
        RECT 21.045 15.655 22.225 16.835 ;
        RECT 28.245 15.655 29.425 16.835 ;
        RECT 34.135 15.635 35.315 16.815 ;
        RECT 41.335 15.635 42.515 16.815 ;
        RECT 47.225 15.635 48.405 16.815 ;
        RECT 54.425 15.635 55.605 16.815 ;
        RECT 60.275 15.635 61.455 16.815 ;
        RECT 67.475 15.635 68.655 16.815 ;
        RECT 73.365 15.635 74.545 16.815 ;
        RECT 80.565 15.635 81.745 16.815 ;
        RECT 86.455 15.615 87.635 16.795 ;
        RECT 93.655 15.615 94.835 16.795 ;
        RECT 99.545 15.615 100.725 16.795 ;
        RECT 106.745 15.615 107.925 16.795 ;
        RECT 112.635 15.615 113.815 16.795 ;
        RECT 119.835 15.615 121.015 16.795 ;
        RECT 125.725 15.615 126.905 16.795 ;
        RECT 132.925 15.615 134.105 16.795 ;
        RECT 138.815 15.595 139.995 16.775 ;
        RECT 146.015 15.595 147.195 16.775 ;
        RECT 151.905 15.595 153.085 16.775 ;
        RECT 159.105 15.595 160.285 16.775 ;
        RECT 7.985 12.005 9.165 13.185 ;
        RECT 15.185 12.005 16.365 13.185 ;
        RECT 21.075 12.005 22.255 13.185 ;
        RECT 28.275 12.005 29.455 13.185 ;
        RECT 34.165 12.025 35.345 13.205 ;
        RECT 41.365 12.025 42.545 13.205 ;
        RECT 47.255 12.025 48.435 13.205 ;
        RECT 54.455 12.025 55.635 13.205 ;
        RECT 60.305 12.025 61.485 13.205 ;
        RECT 67.505 12.025 68.685 13.205 ;
        RECT 73.395 12.025 74.575 13.205 ;
        RECT 80.595 12.025 81.775 13.205 ;
        RECT 86.485 12.045 87.665 13.225 ;
        RECT 93.685 12.045 94.865 13.225 ;
        RECT 99.575 12.045 100.755 13.225 ;
        RECT 106.775 12.045 107.955 13.225 ;
        RECT 112.665 12.045 113.845 13.225 ;
        RECT 119.865 12.045 121.045 13.225 ;
        RECT 125.755 12.045 126.935 13.225 ;
        RECT 132.955 12.045 134.135 13.225 ;
        RECT 138.845 12.065 140.025 13.245 ;
        RECT 146.045 12.065 147.225 13.245 ;
        RECT 151.935 12.065 153.115 13.245 ;
        RECT 159.135 12.065 160.315 13.245 ;
      LAYER met5 ;
        RECT 9.355 108.595 10.955 115.335 ;
        RECT 15.755 108.595 17.565 115.335 ;
        RECT 22.445 108.595 24.045 115.335 ;
        RECT 28.845 108.595 30.655 115.335 ;
        RECT 6.155 107.700 17.565 108.595 ;
        RECT 19.245 107.700 30.655 108.595 ;
        RECT 35.535 108.575 37.135 115.315 ;
        RECT 41.935 108.575 43.745 115.315 ;
        RECT 48.625 108.575 50.225 115.315 ;
        RECT 55.025 108.575 56.835 115.315 ;
        RECT 61.675 108.575 63.275 115.315 ;
        RECT 68.075 108.575 69.885 115.315 ;
        RECT 74.765 108.575 76.365 115.315 ;
        RECT 81.165 108.575 82.975 115.315 ;
        RECT 32.335 107.700 43.745 108.575 ;
        RECT 45.425 107.700 56.835 108.575 ;
        RECT 58.475 107.700 69.885 108.575 ;
        RECT 71.565 107.700 82.975 108.575 ;
        RECT 87.855 108.555 89.455 115.295 ;
        RECT 94.255 108.555 96.065 115.295 ;
        RECT 100.945 108.555 102.545 115.295 ;
        RECT 107.345 108.555 109.155 115.295 ;
        RECT 114.035 108.555 115.635 115.295 ;
        RECT 120.435 108.555 122.245 115.295 ;
        RECT 127.125 108.555 128.725 115.295 ;
        RECT 133.525 108.555 135.335 115.295 ;
        RECT 84.655 107.700 96.065 108.555 ;
        RECT 97.745 107.700 109.155 108.555 ;
        RECT 110.835 107.700 122.245 108.555 ;
        RECT 123.925 107.700 135.335 108.555 ;
        RECT 140.215 108.535 141.815 115.275 ;
        RECT 146.615 108.535 148.425 115.275 ;
        RECT 153.305 108.535 154.905 115.275 ;
        RECT 159.705 108.535 161.515 115.275 ;
        RECT 137.015 107.700 148.425 108.535 ;
        RECT 150.105 107.700 161.515 108.535 ;
        RECT 3.330 104.390 164.710 107.700 ;
        RECT 6.185 103.525 17.595 104.390 ;
        RECT 19.275 103.525 30.685 104.390 ;
        RECT 32.365 103.545 43.775 104.390 ;
        RECT 45.455 103.545 56.865 104.390 ;
        RECT 58.505 103.545 69.915 104.390 ;
        RECT 71.595 103.545 83.005 104.390 ;
        RECT 84.685 103.565 96.095 104.390 ;
        RECT 97.775 103.565 109.185 104.390 ;
        RECT 110.865 103.565 122.275 104.390 ;
        RECT 123.955 103.565 135.365 104.390 ;
        RECT 137.045 103.585 148.455 104.390 ;
        RECT 150.135 103.585 161.545 104.390 ;
        RECT 9.385 96.785 10.985 103.525 ;
        RECT 15.785 96.785 17.595 103.525 ;
        RECT 22.475 96.785 24.075 103.525 ;
        RECT 28.875 96.785 30.685 103.525 ;
        RECT 35.565 96.805 37.165 103.545 ;
        RECT 41.965 96.805 43.775 103.545 ;
        RECT 48.655 96.805 50.255 103.545 ;
        RECT 55.055 96.805 56.865 103.545 ;
        RECT 61.705 96.805 63.305 103.545 ;
        RECT 68.105 96.805 69.915 103.545 ;
        RECT 74.795 96.805 76.395 103.545 ;
        RECT 81.195 96.805 83.005 103.545 ;
        RECT 87.885 96.825 89.485 103.565 ;
        RECT 94.285 96.825 96.095 103.565 ;
        RECT 100.975 96.825 102.575 103.565 ;
        RECT 107.375 96.825 109.185 103.565 ;
        RECT 114.065 96.825 115.665 103.565 ;
        RECT 120.465 96.825 122.275 103.565 ;
        RECT 127.155 96.825 128.755 103.565 ;
        RECT 133.555 96.825 135.365 103.565 ;
        RECT 140.245 96.845 141.845 103.585 ;
        RECT 146.645 96.845 148.455 103.585 ;
        RECT 153.335 96.845 154.935 103.585 ;
        RECT 159.735 96.845 161.545 103.585 ;
        RECT 9.795 16.955 11.395 23.695 ;
        RECT 16.195 16.955 18.005 23.695 ;
        RECT 22.885 16.955 24.485 23.695 ;
        RECT 29.285 16.955 31.095 23.695 ;
        RECT 6.595 16.120 18.005 16.955 ;
        RECT 19.685 16.120 31.095 16.955 ;
        RECT 35.975 16.935 37.575 23.675 ;
        RECT 42.375 16.935 44.185 23.675 ;
        RECT 49.065 16.935 50.665 23.675 ;
        RECT 55.465 16.935 57.275 23.675 ;
        RECT 62.115 16.935 63.715 23.675 ;
        RECT 68.515 16.935 70.325 23.675 ;
        RECT 75.205 16.935 76.805 23.675 ;
        RECT 81.605 16.935 83.415 23.675 ;
        RECT 32.775 16.120 44.185 16.935 ;
        RECT 45.865 16.120 57.275 16.935 ;
        RECT 58.915 16.120 70.325 16.935 ;
        RECT 72.005 16.120 83.415 16.935 ;
        RECT 88.295 16.915 89.895 23.655 ;
        RECT 94.695 16.915 96.505 23.655 ;
        RECT 101.385 16.915 102.985 23.655 ;
        RECT 107.785 16.915 109.595 23.655 ;
        RECT 114.475 16.915 116.075 23.655 ;
        RECT 120.875 16.915 122.685 23.655 ;
        RECT 127.565 16.915 129.165 23.655 ;
        RECT 133.965 16.915 135.775 23.655 ;
        RECT 85.095 16.120 96.505 16.915 ;
        RECT 98.185 16.120 109.595 16.915 ;
        RECT 111.275 16.120 122.685 16.915 ;
        RECT 124.365 16.120 135.775 16.915 ;
        RECT 140.655 16.895 142.255 23.635 ;
        RECT 147.055 16.895 148.865 23.635 ;
        RECT 153.745 16.895 155.345 23.635 ;
        RECT 160.145 16.895 161.955 23.635 ;
        RECT 137.455 16.120 148.865 16.895 ;
        RECT 150.545 16.120 161.955 16.895 ;
        RECT 3.655 12.810 164.540 16.120 ;
        RECT 6.625 11.885 18.035 12.810 ;
        RECT 19.715 11.885 31.125 12.810 ;
        RECT 32.805 11.905 44.215 12.810 ;
        RECT 45.895 11.905 57.305 12.810 ;
        RECT 58.945 11.905 70.355 12.810 ;
        RECT 72.035 11.905 83.445 12.810 ;
        RECT 85.125 11.925 96.535 12.810 ;
        RECT 98.215 11.925 109.625 12.810 ;
        RECT 111.305 11.925 122.715 12.810 ;
        RECT 124.395 11.925 135.805 12.810 ;
        RECT 137.485 11.945 148.895 12.810 ;
        RECT 150.575 11.945 161.985 12.810 ;
        RECT 9.825 5.145 11.425 11.885 ;
        RECT 16.225 5.145 18.035 11.885 ;
        RECT 22.915 5.145 24.515 11.885 ;
        RECT 29.315 5.145 31.125 11.885 ;
        RECT 36.005 5.165 37.605 11.905 ;
        RECT 42.405 5.165 44.215 11.905 ;
        RECT 49.095 5.165 50.695 11.905 ;
        RECT 55.495 5.165 57.305 11.905 ;
        RECT 62.145 5.165 63.745 11.905 ;
        RECT 68.545 5.165 70.355 11.905 ;
        RECT 75.235 5.165 76.835 11.905 ;
        RECT 81.635 5.165 83.445 11.905 ;
        RECT 88.325 5.185 89.925 11.925 ;
        RECT 94.725 5.185 96.535 11.925 ;
        RECT 101.415 5.185 103.015 11.925 ;
        RECT 107.815 5.185 109.625 11.925 ;
        RECT 114.505 5.185 116.105 11.925 ;
        RECT 120.905 5.185 122.715 11.925 ;
        RECT 127.595 5.185 129.195 11.925 ;
        RECT 133.995 5.185 135.805 11.925 ;
        RECT 140.685 5.205 142.285 11.945 ;
        RECT 147.085 5.205 148.895 11.945 ;
        RECT 153.775 5.205 155.375 11.945 ;
        RECT 160.175 5.205 161.985 11.945 ;
    END
  END avss
  OBS
      LAYER pwell ;
        RECT 147.900 88.585 148.685 89.475 ;
        RECT 147.815 88.440 148.725 88.570 ;
        RECT 147.625 88.270 148.725 88.440 ;
        RECT 147.815 87.220 148.725 88.270 ;
        RECT 147.815 87.065 148.725 87.195 ;
        RECT 147.625 86.895 148.725 87.065 ;
        RECT 147.815 85.845 148.725 86.895 ;
        RECT 147.815 85.695 148.725 85.825 ;
        RECT 147.625 85.525 148.725 85.695 ;
        RECT 147.815 84.475 148.725 85.525 ;
        RECT 147.815 84.320 148.725 84.450 ;
        RECT 147.625 84.150 148.725 84.320 ;
        RECT 147.815 83.100 148.725 84.150 ;
        RECT 147.815 82.940 148.725 83.070 ;
        RECT 147.625 82.770 148.725 82.940 ;
        RECT 10.890 81.645 11.060 81.835 ;
        RECT 14.560 81.645 14.730 81.835 ;
        RECT 16.825 81.645 16.995 81.835 ;
        RECT 19.125 81.645 19.295 81.835 ;
        RECT 20.505 81.645 20.675 81.835 ;
        RECT 24.175 81.645 24.345 81.835 ;
        RECT 26.440 81.645 26.610 81.835 ;
        RECT 28.740 81.645 28.910 81.835 ;
        RECT 30.120 81.645 30.290 81.835 ;
        RECT 33.790 81.645 33.960 81.835 ;
        RECT 36.055 81.645 36.225 81.835 ;
        RECT 38.355 81.645 38.525 81.835 ;
        RECT 39.735 81.645 39.905 81.835 ;
        RECT 43.405 81.645 43.575 81.835 ;
        RECT 45.670 81.645 45.840 81.835 ;
        RECT 47.970 81.645 48.140 81.835 ;
        RECT 147.815 81.720 148.725 82.770 ;
        RECT 9.840 80.775 10.730 81.560 ;
        RECT 10.750 80.835 14.420 81.645 ;
        RECT 14.470 80.735 16.660 81.645 ;
        RECT 16.735 80.735 18.925 81.645 ;
        RECT 18.985 80.835 20.355 81.645 ;
        RECT 20.365 80.835 24.035 81.645 ;
        RECT 24.085 80.735 26.275 81.645 ;
        RECT 26.350 80.735 28.540 81.645 ;
        RECT 28.600 80.835 29.970 81.645 ;
        RECT 29.980 80.835 33.650 81.645 ;
        RECT 33.700 80.735 35.890 81.645 ;
        RECT 35.965 80.735 38.155 81.645 ;
        RECT 38.215 80.835 39.585 81.645 ;
        RECT 39.595 80.835 43.265 81.645 ;
        RECT 43.315 80.735 45.505 81.645 ;
        RECT 45.580 80.735 47.770 81.645 ;
        RECT 47.830 80.835 49.200 81.645 ;
        RECT 147.815 81.565 148.725 81.695 ;
        RECT 49.220 80.775 50.110 81.560 ;
        RECT 147.625 81.395 148.725 81.565 ;
        RECT 147.815 80.345 148.725 81.395 ;
        RECT 147.815 80.190 148.725 80.320 ;
        RECT 147.625 80.020 148.725 80.190 ;
        RECT 147.815 78.970 148.725 80.020 ;
        RECT 147.815 78.820 148.725 78.950 ;
        RECT 147.625 78.650 148.725 78.820 ;
        RECT 147.815 77.600 148.725 78.650 ;
        RECT 147.815 77.445 148.725 77.575 ;
        RECT 147.625 77.275 148.725 77.445 ;
        RECT 147.815 76.225 148.725 77.275 ;
        RECT 147.900 75.320 148.685 76.210 ;
      LAYER nwell ;
        RECT 149.015 75.115 150.620 89.680 ;
      LAYER pwell ;
        RECT 172.785 64.455 174.045 65.695 ;
        RECT 172.785 62.885 174.045 64.125 ;
        RECT 172.785 61.315 174.045 62.555 ;
        RECT 172.785 58.955 174.045 60.195 ;
        RECT 172.785 57.385 174.045 58.625 ;
        RECT 172.785 55.815 174.045 57.055 ;
        RECT 147.900 43.640 148.685 44.530 ;
        RECT 147.815 42.575 148.725 43.625 ;
        RECT 147.625 42.405 148.725 42.575 ;
        RECT 147.815 42.275 148.725 42.405 ;
        RECT 147.815 41.200 148.725 42.250 ;
        RECT 147.625 41.030 148.725 41.200 ;
        RECT 147.815 40.900 148.725 41.030 ;
        RECT 147.815 39.830 148.725 40.880 ;
        RECT 147.625 39.660 148.725 39.830 ;
        RECT 147.815 39.530 148.725 39.660 ;
        RECT 9.840 38.290 10.730 39.075 ;
        RECT 10.750 38.205 14.420 39.015 ;
        RECT 14.470 38.205 16.660 39.115 ;
        RECT 16.735 38.205 18.925 39.115 ;
        RECT 18.985 38.205 20.355 39.015 ;
        RECT 20.365 38.205 24.035 39.015 ;
        RECT 24.085 38.205 26.275 39.115 ;
        RECT 26.350 38.205 28.540 39.115 ;
        RECT 28.600 38.205 29.970 39.015 ;
        RECT 29.980 38.205 33.650 39.015 ;
        RECT 33.700 38.205 35.890 39.115 ;
        RECT 35.965 38.205 38.155 39.115 ;
        RECT 38.215 38.205 39.585 39.015 ;
        RECT 39.595 38.205 43.265 39.015 ;
        RECT 43.315 38.205 45.505 39.115 ;
        RECT 45.580 38.205 47.770 39.115 ;
        RECT 47.830 38.205 49.200 39.015 ;
        RECT 49.220 38.290 50.110 39.075 ;
        RECT 147.815 38.455 148.725 39.505 ;
        RECT 147.625 38.285 148.725 38.455 ;
        RECT 10.890 38.015 11.060 38.205 ;
        RECT 14.560 38.015 14.730 38.205 ;
        RECT 16.825 38.015 16.995 38.205 ;
        RECT 19.125 38.015 19.295 38.205 ;
        RECT 20.505 38.015 20.675 38.205 ;
        RECT 24.175 38.015 24.345 38.205 ;
        RECT 26.440 38.015 26.610 38.205 ;
        RECT 28.740 38.015 28.910 38.205 ;
        RECT 30.120 38.015 30.290 38.205 ;
        RECT 33.790 38.015 33.960 38.205 ;
        RECT 36.055 38.015 36.225 38.205 ;
        RECT 38.355 38.015 38.525 38.205 ;
        RECT 39.735 38.015 39.905 38.205 ;
        RECT 43.405 38.015 43.575 38.205 ;
        RECT 45.670 38.015 45.840 38.205 ;
        RECT 47.970 38.015 48.140 38.205 ;
        RECT 147.815 38.155 148.725 38.285 ;
        RECT 147.815 37.080 148.725 38.130 ;
        RECT 147.625 36.910 148.725 37.080 ;
        RECT 147.815 36.780 148.725 36.910 ;
        RECT 147.815 35.700 148.725 36.750 ;
        RECT 147.625 35.530 148.725 35.700 ;
        RECT 147.815 35.400 148.725 35.530 ;
        RECT 147.815 34.325 148.725 35.375 ;
        RECT 147.625 34.155 148.725 34.325 ;
        RECT 147.815 34.025 148.725 34.155 ;
        RECT 147.815 32.955 148.725 34.005 ;
        RECT 147.625 32.785 148.725 32.955 ;
        RECT 147.815 32.655 148.725 32.785 ;
        RECT 147.815 31.580 148.725 32.630 ;
        RECT 147.625 31.410 148.725 31.580 ;
        RECT 147.815 31.280 148.725 31.410 ;
        RECT 147.900 30.375 148.685 31.265 ;
      LAYER nwell ;
        RECT 149.015 30.170 150.620 44.735 ;
      LAYER li1 ;
        RECT 147.975 88.655 148.520 89.405 ;
        RECT 149.180 88.655 150.165 89.405 ;
        RECT 147.965 87.980 148.595 88.060 ;
        RECT 149.195 87.980 150.175 88.060 ;
        RECT 147.965 87.730 150.175 87.980 ;
        RECT 147.965 86.605 148.595 86.685 ;
        RECT 149.195 86.605 150.175 86.685 ;
        RECT 147.965 86.355 150.175 86.605 ;
        RECT 147.965 85.235 148.595 85.315 ;
        RECT 149.195 85.235 150.175 85.315 ;
        RECT 147.965 84.985 150.175 85.235 ;
        RECT 147.965 83.860 148.595 83.940 ;
        RECT 149.195 83.860 150.175 83.940 ;
        RECT 147.965 83.610 150.175 83.860 ;
        RECT 147.965 82.480 148.595 82.560 ;
        RECT 149.195 82.480 150.175 82.560 ;
        RECT 147.965 82.230 150.175 82.480 ;
        RECT 9.910 80.940 10.660 81.485 ;
        RECT 14.980 81.025 15.310 81.495 ;
        RECT 15.820 81.025 16.150 81.495 ;
        RECT 17.245 81.025 17.575 81.495 ;
        RECT 18.085 81.025 18.415 81.495 ;
        RECT 24.595 81.025 24.925 81.495 ;
        RECT 25.435 81.025 25.765 81.495 ;
        RECT 26.860 81.025 27.190 81.495 ;
        RECT 27.700 81.025 28.030 81.495 ;
        RECT 34.210 81.025 34.540 81.495 ;
        RECT 35.050 81.025 35.380 81.495 ;
        RECT 36.475 81.025 36.805 81.495 ;
        RECT 37.315 81.025 37.645 81.495 ;
        RECT 43.825 81.025 44.155 81.495 ;
        RECT 44.665 81.025 44.995 81.495 ;
        RECT 46.090 81.025 46.420 81.495 ;
        RECT 46.930 81.025 47.260 81.495 ;
        RECT 14.980 80.930 16.585 81.025 ;
        RECT 14.980 80.845 16.595 80.930 ;
        RECT 17.245 80.845 18.850 81.025 ;
        RECT 24.595 80.930 26.200 81.025 ;
        RECT 24.595 80.845 26.210 80.930 ;
        RECT 26.860 80.845 28.465 81.025 ;
        RECT 34.210 80.930 35.815 81.025 ;
        RECT 34.210 80.845 35.825 80.930 ;
        RECT 36.475 80.845 38.080 81.025 ;
        RECT 43.825 80.930 45.430 81.025 ;
        RECT 43.825 80.845 45.440 80.930 ;
        RECT 46.090 80.845 47.695 81.025 ;
        RECT 49.290 80.940 50.040 81.485 ;
        RECT 147.965 81.105 148.595 81.185 ;
        RECT 149.195 81.105 150.175 81.185 ;
        RECT 147.965 80.855 150.175 81.105 ;
        RECT 16.320 80.255 16.595 80.845 ;
        RECT 16.785 80.425 18.415 80.675 ;
        RECT 18.585 80.255 18.850 80.845 ;
        RECT 25.935 80.255 26.210 80.845 ;
        RECT 26.400 80.425 28.030 80.675 ;
        RECT 28.200 80.255 28.465 80.845 ;
        RECT 35.550 80.255 35.825 80.845 ;
        RECT 36.015 80.425 37.645 80.675 ;
        RECT 37.815 80.255 38.080 80.845 ;
        RECT 45.165 80.255 45.440 80.845 ;
        RECT 45.630 80.425 47.260 80.675 ;
        RECT 47.430 80.255 47.695 80.845 ;
        RECT 14.980 80.130 16.595 80.255 ;
        RECT 14.980 80.085 16.585 80.130 ;
        RECT 14.980 79.285 15.310 80.085 ;
        RECT 15.820 80.065 16.585 80.085 ;
        RECT 17.245 80.085 18.850 80.255 ;
        RECT 15.820 79.285 16.150 80.065 ;
        RECT 17.245 79.285 17.575 80.085 ;
        RECT 18.085 80.065 18.850 80.085 ;
        RECT 24.595 80.130 26.210 80.255 ;
        RECT 24.595 80.085 26.200 80.130 ;
        RECT 18.085 79.285 18.415 80.065 ;
        RECT 24.595 79.285 24.925 80.085 ;
        RECT 25.435 80.065 26.200 80.085 ;
        RECT 26.860 80.085 28.465 80.255 ;
        RECT 25.435 79.285 25.765 80.065 ;
        RECT 26.860 79.285 27.190 80.085 ;
        RECT 27.700 80.065 28.465 80.085 ;
        RECT 34.210 80.130 35.825 80.255 ;
        RECT 34.210 80.085 35.815 80.130 ;
        RECT 27.700 79.285 28.030 80.065 ;
        RECT 34.210 79.285 34.540 80.085 ;
        RECT 35.050 80.065 35.815 80.085 ;
        RECT 36.475 80.085 38.080 80.255 ;
        RECT 35.050 79.285 35.380 80.065 ;
        RECT 36.475 79.285 36.805 80.085 ;
        RECT 37.315 80.065 38.080 80.085 ;
        RECT 43.825 80.130 45.440 80.255 ;
        RECT 43.825 80.085 45.430 80.130 ;
        RECT 37.315 79.285 37.645 80.065 ;
        RECT 43.825 79.285 44.155 80.085 ;
        RECT 44.665 80.065 45.430 80.085 ;
        RECT 46.090 80.085 47.695 80.255 ;
        RECT 44.665 79.285 44.995 80.065 ;
        RECT 46.090 79.285 46.420 80.085 ;
        RECT 46.930 80.065 47.695 80.085 ;
        RECT 46.930 79.285 47.260 80.065 ;
        RECT 147.965 79.730 148.595 79.810 ;
        RECT 149.195 79.730 150.175 79.810 ;
        RECT 147.965 79.480 150.175 79.730 ;
        RECT 147.965 78.360 148.595 78.440 ;
        RECT 149.195 78.360 150.175 78.440 ;
        RECT 147.965 78.110 150.175 78.360 ;
        RECT 12.400 77.490 12.730 77.660 ;
        RECT 12.990 77.490 13.320 77.660 ;
        RECT 13.580 77.490 13.910 77.660 ;
        RECT 14.170 77.490 14.500 77.660 ;
        RECT 14.760 77.490 15.090 77.660 ;
        RECT 15.350 77.490 15.680 77.660 ;
        RECT 15.940 77.490 16.270 77.660 ;
        RECT 16.530 77.490 16.860 77.660 ;
        RECT 17.120 77.490 17.450 77.660 ;
        RECT 17.710 77.490 18.040 77.660 ;
        RECT 22.015 77.490 22.345 77.660 ;
        RECT 22.605 77.490 22.935 77.660 ;
        RECT 23.195 77.490 23.525 77.660 ;
        RECT 23.785 77.490 24.115 77.660 ;
        RECT 24.375 77.490 24.705 77.660 ;
        RECT 24.965 77.490 25.295 77.660 ;
        RECT 25.555 77.490 25.885 77.660 ;
        RECT 26.145 77.490 26.475 77.660 ;
        RECT 26.735 77.490 27.065 77.660 ;
        RECT 27.325 77.490 27.655 77.660 ;
        RECT 31.630 77.490 31.960 77.660 ;
        RECT 32.220 77.490 32.550 77.660 ;
        RECT 32.810 77.490 33.140 77.660 ;
        RECT 33.400 77.490 33.730 77.660 ;
        RECT 33.990 77.490 34.320 77.660 ;
        RECT 34.580 77.490 34.910 77.660 ;
        RECT 35.170 77.490 35.500 77.660 ;
        RECT 35.760 77.490 36.090 77.660 ;
        RECT 36.350 77.490 36.680 77.660 ;
        RECT 36.940 77.490 37.270 77.660 ;
        RECT 41.245 77.490 41.575 77.660 ;
        RECT 41.835 77.490 42.165 77.660 ;
        RECT 42.425 77.490 42.755 77.660 ;
        RECT 43.015 77.490 43.345 77.660 ;
        RECT 43.605 77.490 43.935 77.660 ;
        RECT 44.195 77.490 44.525 77.660 ;
        RECT 44.785 77.490 45.115 77.660 ;
        RECT 45.375 77.490 45.705 77.660 ;
        RECT 45.965 77.490 46.295 77.660 ;
        RECT 46.555 77.490 46.885 77.660 ;
        RECT 12.775 76.370 12.945 77.230 ;
        RECT 13.955 76.370 14.125 77.230 ;
        RECT 15.135 76.370 15.305 77.230 ;
        RECT 16.315 76.370 16.485 77.230 ;
        RECT 17.495 76.370 17.665 77.230 ;
        RECT 22.390 76.370 22.560 77.230 ;
        RECT 23.570 76.370 23.740 77.230 ;
        RECT 24.750 76.370 24.920 77.230 ;
        RECT 25.930 76.370 26.100 77.230 ;
        RECT 27.110 76.370 27.280 77.230 ;
        RECT 32.005 76.370 32.175 77.230 ;
        RECT 33.185 76.370 33.355 77.230 ;
        RECT 34.365 76.370 34.535 77.230 ;
        RECT 35.545 76.370 35.715 77.230 ;
        RECT 36.725 76.370 36.895 77.230 ;
        RECT 41.620 76.370 41.790 77.230 ;
        RECT 42.800 76.370 42.970 77.230 ;
        RECT 43.980 76.370 44.150 77.230 ;
        RECT 45.160 76.370 45.330 77.230 ;
        RECT 46.340 76.370 46.510 77.230 ;
        RECT 147.965 76.985 148.595 77.065 ;
        RECT 149.195 76.985 150.175 77.065 ;
        RECT 147.965 76.735 150.175 76.985 ;
        RECT 147.975 75.390 148.520 76.140 ;
        RECT 149.180 75.390 150.165 76.140 ;
        RECT 12.785 73.885 12.955 74.745 ;
        RECT 13.965 73.885 14.135 74.745 ;
        RECT 15.145 73.885 15.315 74.745 ;
        RECT 16.325 73.885 16.495 74.745 ;
        RECT 17.505 73.885 17.675 74.745 ;
        RECT 22.400 73.885 22.570 74.745 ;
        RECT 23.580 73.885 23.750 74.745 ;
        RECT 24.760 73.885 24.930 74.745 ;
        RECT 25.940 73.885 26.110 74.745 ;
        RECT 27.120 73.885 27.290 74.745 ;
        RECT 32.015 73.885 32.185 74.745 ;
        RECT 33.195 73.885 33.365 74.745 ;
        RECT 34.375 73.885 34.545 74.745 ;
        RECT 35.555 73.885 35.725 74.745 ;
        RECT 36.735 73.885 36.905 74.745 ;
        RECT 41.630 73.885 41.800 74.745 ;
        RECT 42.810 73.885 42.980 74.745 ;
        RECT 43.990 73.885 44.160 74.745 ;
        RECT 45.170 73.885 45.340 74.745 ;
        RECT 46.350 73.885 46.520 74.745 ;
        RECT 12.410 73.410 12.740 73.580 ;
        RECT 13.000 73.410 13.330 73.580 ;
        RECT 13.590 73.410 13.920 73.580 ;
        RECT 14.180 73.410 14.510 73.580 ;
        RECT 14.770 73.410 15.100 73.580 ;
        RECT 15.360 73.410 15.690 73.580 ;
        RECT 15.950 73.410 16.280 73.580 ;
        RECT 16.540 73.410 16.870 73.580 ;
        RECT 17.130 73.410 17.460 73.580 ;
        RECT 17.720 73.410 18.050 73.580 ;
        RECT 22.025 73.410 22.355 73.580 ;
        RECT 22.615 73.410 22.945 73.580 ;
        RECT 23.205 73.410 23.535 73.580 ;
        RECT 23.795 73.410 24.125 73.580 ;
        RECT 24.385 73.410 24.715 73.580 ;
        RECT 24.975 73.410 25.305 73.580 ;
        RECT 25.565 73.410 25.895 73.580 ;
        RECT 26.155 73.410 26.485 73.580 ;
        RECT 26.745 73.410 27.075 73.580 ;
        RECT 27.335 73.410 27.665 73.580 ;
        RECT 31.640 73.410 31.970 73.580 ;
        RECT 32.230 73.410 32.560 73.580 ;
        RECT 32.820 73.410 33.150 73.580 ;
        RECT 33.410 73.410 33.740 73.580 ;
        RECT 34.000 73.410 34.330 73.580 ;
        RECT 34.590 73.410 34.920 73.580 ;
        RECT 35.180 73.410 35.510 73.580 ;
        RECT 35.770 73.410 36.100 73.580 ;
        RECT 36.360 73.410 36.690 73.580 ;
        RECT 36.950 73.410 37.280 73.580 ;
        RECT 41.255 73.410 41.585 73.580 ;
        RECT 41.845 73.410 42.175 73.580 ;
        RECT 42.435 73.410 42.765 73.580 ;
        RECT 43.025 73.410 43.355 73.580 ;
        RECT 43.615 73.410 43.945 73.580 ;
        RECT 44.205 73.410 44.535 73.580 ;
        RECT 44.795 73.410 45.125 73.580 ;
        RECT 45.385 73.410 45.715 73.580 ;
        RECT 45.975 73.410 46.305 73.580 ;
        RECT 46.565 73.410 46.895 73.580 ;
        RECT 166.665 68.885 167.525 69.055 ;
        RECT 169.460 68.950 170.320 69.120 ;
        RECT 150.590 68.025 150.760 68.885 ;
        RECT 151.770 68.025 151.940 68.885 ;
        RECT 152.950 68.025 153.120 68.885 ;
        RECT 154.130 68.025 154.300 68.885 ;
        RECT 155.310 68.025 155.480 68.885 ;
        RECT 158.580 68.025 158.750 68.885 ;
        RECT 159.760 68.025 159.930 68.885 ;
        RECT 160.940 68.025 161.110 68.885 ;
        RECT 163.485 68.025 163.655 68.885 ;
        RECT 164.665 68.025 164.835 68.885 ;
        RECT 174.105 64.875 174.275 65.275 ;
        RECT 175.935 64.875 176.105 65.275 ;
        RECT 172.895 64.645 173.935 64.815 ;
        RECT 176.320 64.645 177.360 64.815 ;
        RECT 174.105 63.305 174.275 63.705 ;
        RECT 172.895 63.075 173.935 63.245 ;
        RECT 174.105 61.735 174.275 62.135 ;
        RECT 175.935 61.735 176.105 62.135 ;
        RECT 154.295 60.755 154.465 61.615 ;
        RECT 155.995 60.780 156.165 61.640 ;
        RECT 156.585 60.780 156.755 61.640 ;
        RECT 158.295 60.795 158.465 61.655 ;
        RECT 158.885 60.795 159.055 61.655 ;
        RECT 160.985 61.265 161.845 61.435 ;
        RECT 162.490 61.265 163.350 61.435 ;
        RECT 164.315 61.265 165.175 61.435 ;
        RECT 160.510 60.890 160.680 61.220 ;
        RECT 156.200 60.355 156.540 60.530 ;
        RECT 158.510 60.365 158.840 60.535 ;
        RECT 156.210 60.350 156.540 60.355 ;
        RECT 156.210 59.770 156.550 59.940 ;
        RECT 158.510 59.785 158.840 59.955 ;
        RECT 172.895 59.835 173.935 60.005 ;
        RECT 176.320 59.835 177.360 60.005 ;
        RECT 154.295 58.625 154.465 59.485 ;
        RECT 155.995 58.650 156.165 59.510 ;
        RECT 156.585 58.650 156.755 59.510 ;
        RECT 158.295 58.665 158.465 59.525 ;
        RECT 158.885 58.665 159.055 59.525 ;
        RECT 160.510 59.095 160.680 59.425 ;
        RECT 160.985 58.880 161.845 59.050 ;
        RECT 162.490 58.880 163.350 59.050 ;
        RECT 164.315 58.880 165.175 59.050 ;
        RECT 174.105 57.805 174.275 58.205 ;
        RECT 172.895 56.695 173.935 56.865 ;
        RECT 176.320 56.695 177.360 56.865 ;
        RECT 174.105 56.235 174.275 56.635 ;
        RECT 175.935 56.235 176.105 56.635 ;
        RECT 150.705 51.095 150.875 51.955 ;
        RECT 151.885 51.095 152.055 51.955 ;
        RECT 153.065 51.095 153.235 51.955 ;
        RECT 154.245 51.095 154.415 51.955 ;
        RECT 155.425 51.095 155.595 51.955 ;
        RECT 158.695 51.095 158.865 51.955 ;
        RECT 159.875 51.095 160.045 51.955 ;
        RECT 161.055 51.095 161.225 51.955 ;
        RECT 163.600 51.095 163.770 51.955 ;
        RECT 164.780 51.095 164.950 51.955 ;
        RECT 166.780 50.925 167.640 51.095 ;
        RECT 169.575 50.860 170.435 51.030 ;
        RECT 12.410 46.270 12.740 46.440 ;
        RECT 13.000 46.270 13.330 46.440 ;
        RECT 13.590 46.270 13.920 46.440 ;
        RECT 14.180 46.270 14.510 46.440 ;
        RECT 14.770 46.270 15.100 46.440 ;
        RECT 15.360 46.270 15.690 46.440 ;
        RECT 15.950 46.270 16.280 46.440 ;
        RECT 16.540 46.270 16.870 46.440 ;
        RECT 17.130 46.270 17.460 46.440 ;
        RECT 17.720 46.270 18.050 46.440 ;
        RECT 22.025 46.270 22.355 46.440 ;
        RECT 22.615 46.270 22.945 46.440 ;
        RECT 23.205 46.270 23.535 46.440 ;
        RECT 23.795 46.270 24.125 46.440 ;
        RECT 24.385 46.270 24.715 46.440 ;
        RECT 24.975 46.270 25.305 46.440 ;
        RECT 25.565 46.270 25.895 46.440 ;
        RECT 26.155 46.270 26.485 46.440 ;
        RECT 26.745 46.270 27.075 46.440 ;
        RECT 27.335 46.270 27.665 46.440 ;
        RECT 31.640 46.270 31.970 46.440 ;
        RECT 32.230 46.270 32.560 46.440 ;
        RECT 32.820 46.270 33.150 46.440 ;
        RECT 33.410 46.270 33.740 46.440 ;
        RECT 34.000 46.270 34.330 46.440 ;
        RECT 34.590 46.270 34.920 46.440 ;
        RECT 35.180 46.270 35.510 46.440 ;
        RECT 35.770 46.270 36.100 46.440 ;
        RECT 36.360 46.270 36.690 46.440 ;
        RECT 36.950 46.270 37.280 46.440 ;
        RECT 41.255 46.270 41.585 46.440 ;
        RECT 41.845 46.270 42.175 46.440 ;
        RECT 42.435 46.270 42.765 46.440 ;
        RECT 43.025 46.270 43.355 46.440 ;
        RECT 43.615 46.270 43.945 46.440 ;
        RECT 44.205 46.270 44.535 46.440 ;
        RECT 44.795 46.270 45.125 46.440 ;
        RECT 45.385 46.270 45.715 46.440 ;
        RECT 45.975 46.270 46.305 46.440 ;
        RECT 46.565 46.270 46.895 46.440 ;
        RECT 12.785 45.105 12.955 45.965 ;
        RECT 13.965 45.105 14.135 45.965 ;
        RECT 15.145 45.105 15.315 45.965 ;
        RECT 16.325 45.105 16.495 45.965 ;
        RECT 17.505 45.105 17.675 45.965 ;
        RECT 22.400 45.105 22.570 45.965 ;
        RECT 23.580 45.105 23.750 45.965 ;
        RECT 24.760 45.105 24.930 45.965 ;
        RECT 25.940 45.105 26.110 45.965 ;
        RECT 27.120 45.105 27.290 45.965 ;
        RECT 32.015 45.105 32.185 45.965 ;
        RECT 33.195 45.105 33.365 45.965 ;
        RECT 34.375 45.105 34.545 45.965 ;
        RECT 35.555 45.105 35.725 45.965 ;
        RECT 36.735 45.105 36.905 45.965 ;
        RECT 41.630 45.105 41.800 45.965 ;
        RECT 42.810 45.105 42.980 45.965 ;
        RECT 43.990 45.105 44.160 45.965 ;
        RECT 45.170 45.105 45.340 45.965 ;
        RECT 46.350 45.105 46.520 45.965 ;
        RECT 147.975 43.710 148.520 44.460 ;
        RECT 149.180 43.710 150.165 44.460 ;
        RECT 12.775 42.620 12.945 43.480 ;
        RECT 13.955 42.620 14.125 43.480 ;
        RECT 15.135 42.620 15.305 43.480 ;
        RECT 16.315 42.620 16.485 43.480 ;
        RECT 17.495 42.620 17.665 43.480 ;
        RECT 22.390 42.620 22.560 43.480 ;
        RECT 23.570 42.620 23.740 43.480 ;
        RECT 24.750 42.620 24.920 43.480 ;
        RECT 25.930 42.620 26.100 43.480 ;
        RECT 27.110 42.620 27.280 43.480 ;
        RECT 32.005 42.620 32.175 43.480 ;
        RECT 33.185 42.620 33.355 43.480 ;
        RECT 34.365 42.620 34.535 43.480 ;
        RECT 35.545 42.620 35.715 43.480 ;
        RECT 36.725 42.620 36.895 43.480 ;
        RECT 41.620 42.620 41.790 43.480 ;
        RECT 42.800 42.620 42.970 43.480 ;
        RECT 43.980 42.620 44.150 43.480 ;
        RECT 45.160 42.620 45.330 43.480 ;
        RECT 46.340 42.620 46.510 43.480 ;
        RECT 147.965 42.865 150.175 43.115 ;
        RECT 147.965 42.785 148.595 42.865 ;
        RECT 149.195 42.785 150.175 42.865 ;
        RECT 12.400 42.190 12.730 42.360 ;
        RECT 12.990 42.190 13.320 42.360 ;
        RECT 13.580 42.190 13.910 42.360 ;
        RECT 14.170 42.190 14.500 42.360 ;
        RECT 14.760 42.190 15.090 42.360 ;
        RECT 15.350 42.190 15.680 42.360 ;
        RECT 15.940 42.190 16.270 42.360 ;
        RECT 16.530 42.190 16.860 42.360 ;
        RECT 17.120 42.190 17.450 42.360 ;
        RECT 17.710 42.190 18.040 42.360 ;
        RECT 22.015 42.190 22.345 42.360 ;
        RECT 22.605 42.190 22.935 42.360 ;
        RECT 23.195 42.190 23.525 42.360 ;
        RECT 23.785 42.190 24.115 42.360 ;
        RECT 24.375 42.190 24.705 42.360 ;
        RECT 24.965 42.190 25.295 42.360 ;
        RECT 25.555 42.190 25.885 42.360 ;
        RECT 26.145 42.190 26.475 42.360 ;
        RECT 26.735 42.190 27.065 42.360 ;
        RECT 27.325 42.190 27.655 42.360 ;
        RECT 31.630 42.190 31.960 42.360 ;
        RECT 32.220 42.190 32.550 42.360 ;
        RECT 32.810 42.190 33.140 42.360 ;
        RECT 33.400 42.190 33.730 42.360 ;
        RECT 33.990 42.190 34.320 42.360 ;
        RECT 34.580 42.190 34.910 42.360 ;
        RECT 35.170 42.190 35.500 42.360 ;
        RECT 35.760 42.190 36.090 42.360 ;
        RECT 36.350 42.190 36.680 42.360 ;
        RECT 36.940 42.190 37.270 42.360 ;
        RECT 41.245 42.190 41.575 42.360 ;
        RECT 41.835 42.190 42.165 42.360 ;
        RECT 42.425 42.190 42.755 42.360 ;
        RECT 43.015 42.190 43.345 42.360 ;
        RECT 43.605 42.190 43.935 42.360 ;
        RECT 44.195 42.190 44.525 42.360 ;
        RECT 44.785 42.190 45.115 42.360 ;
        RECT 45.375 42.190 45.705 42.360 ;
        RECT 45.965 42.190 46.295 42.360 ;
        RECT 46.555 42.190 46.885 42.360 ;
        RECT 147.965 41.490 150.175 41.740 ;
        RECT 147.965 41.410 148.595 41.490 ;
        RECT 149.195 41.410 150.175 41.490 ;
        RECT 14.980 39.765 15.310 40.565 ;
        RECT 15.820 39.785 16.150 40.565 ;
        RECT 15.820 39.765 16.585 39.785 ;
        RECT 14.980 39.720 16.585 39.765 ;
        RECT 17.245 39.765 17.575 40.565 ;
        RECT 18.085 39.785 18.415 40.565 ;
        RECT 18.085 39.765 18.850 39.785 ;
        RECT 14.980 39.595 16.595 39.720 ;
        RECT 17.245 39.595 18.850 39.765 ;
        RECT 24.595 39.765 24.925 40.565 ;
        RECT 25.435 39.785 25.765 40.565 ;
        RECT 25.435 39.765 26.200 39.785 ;
        RECT 24.595 39.720 26.200 39.765 ;
        RECT 26.860 39.765 27.190 40.565 ;
        RECT 27.700 39.785 28.030 40.565 ;
        RECT 27.700 39.765 28.465 39.785 ;
        RECT 24.595 39.595 26.210 39.720 ;
        RECT 26.860 39.595 28.465 39.765 ;
        RECT 34.210 39.765 34.540 40.565 ;
        RECT 35.050 39.785 35.380 40.565 ;
        RECT 35.050 39.765 35.815 39.785 ;
        RECT 34.210 39.720 35.815 39.765 ;
        RECT 36.475 39.765 36.805 40.565 ;
        RECT 37.315 39.785 37.645 40.565 ;
        RECT 37.315 39.765 38.080 39.785 ;
        RECT 34.210 39.595 35.825 39.720 ;
        RECT 36.475 39.595 38.080 39.765 ;
        RECT 43.825 39.765 44.155 40.565 ;
        RECT 44.665 39.785 44.995 40.565 ;
        RECT 44.665 39.765 45.430 39.785 ;
        RECT 43.825 39.720 45.430 39.765 ;
        RECT 46.090 39.765 46.420 40.565 ;
        RECT 46.930 39.785 47.260 40.565 ;
        RECT 147.965 40.120 150.175 40.370 ;
        RECT 147.965 40.040 148.595 40.120 ;
        RECT 149.195 40.040 150.175 40.120 ;
        RECT 46.930 39.765 47.695 39.785 ;
        RECT 43.825 39.595 45.440 39.720 ;
        RECT 46.090 39.595 47.695 39.765 ;
        RECT 16.320 39.005 16.595 39.595 ;
        RECT 16.785 39.175 18.415 39.425 ;
        RECT 18.585 39.005 18.850 39.595 ;
        RECT 25.935 39.005 26.210 39.595 ;
        RECT 26.400 39.175 28.030 39.425 ;
        RECT 28.200 39.005 28.465 39.595 ;
        RECT 35.550 39.005 35.825 39.595 ;
        RECT 36.015 39.175 37.645 39.425 ;
        RECT 37.815 39.005 38.080 39.595 ;
        RECT 45.165 39.005 45.440 39.595 ;
        RECT 45.630 39.175 47.260 39.425 ;
        RECT 47.430 39.005 47.695 39.595 ;
        RECT 14.980 38.920 16.595 39.005 ;
        RECT 9.910 38.365 10.660 38.910 ;
        RECT 14.980 38.825 16.585 38.920 ;
        RECT 17.245 38.825 18.850 39.005 ;
        RECT 24.595 38.920 26.210 39.005 ;
        RECT 24.595 38.825 26.200 38.920 ;
        RECT 26.860 38.825 28.465 39.005 ;
        RECT 34.210 38.920 35.825 39.005 ;
        RECT 34.210 38.825 35.815 38.920 ;
        RECT 36.475 38.825 38.080 39.005 ;
        RECT 43.825 38.920 45.440 39.005 ;
        RECT 43.825 38.825 45.430 38.920 ;
        RECT 46.090 38.825 47.695 39.005 ;
        RECT 14.980 38.355 15.310 38.825 ;
        RECT 15.820 38.355 16.150 38.825 ;
        RECT 17.245 38.355 17.575 38.825 ;
        RECT 18.085 38.355 18.415 38.825 ;
        RECT 24.595 38.355 24.925 38.825 ;
        RECT 25.435 38.355 25.765 38.825 ;
        RECT 26.860 38.355 27.190 38.825 ;
        RECT 27.700 38.355 28.030 38.825 ;
        RECT 34.210 38.355 34.540 38.825 ;
        RECT 35.050 38.355 35.380 38.825 ;
        RECT 36.475 38.355 36.805 38.825 ;
        RECT 37.315 38.355 37.645 38.825 ;
        RECT 43.825 38.355 44.155 38.825 ;
        RECT 44.665 38.355 44.995 38.825 ;
        RECT 46.090 38.355 46.420 38.825 ;
        RECT 46.930 38.355 47.260 38.825 ;
        RECT 49.290 38.365 50.040 38.910 ;
        RECT 147.965 38.745 150.175 38.995 ;
        RECT 147.965 38.665 148.595 38.745 ;
        RECT 149.195 38.665 150.175 38.745 ;
        RECT 147.965 37.370 150.175 37.620 ;
        RECT 147.965 37.290 148.595 37.370 ;
        RECT 149.195 37.290 150.175 37.370 ;
        RECT 147.965 35.990 150.175 36.240 ;
        RECT 147.965 35.910 148.595 35.990 ;
        RECT 149.195 35.910 150.175 35.990 ;
        RECT 147.965 34.615 150.175 34.865 ;
        RECT 147.965 34.535 148.595 34.615 ;
        RECT 149.195 34.535 150.175 34.615 ;
        RECT 147.965 33.245 150.175 33.495 ;
        RECT 147.965 33.165 148.595 33.245 ;
        RECT 149.195 33.165 150.175 33.245 ;
        RECT 147.965 31.870 150.175 32.120 ;
        RECT 147.965 31.790 148.595 31.870 ;
        RECT 149.195 31.790 150.175 31.870 ;
        RECT 147.975 30.445 148.520 31.195 ;
        RECT 149.180 30.445 150.165 31.195 ;
      LAYER mcon ;
        RECT 148.820 87.770 149.020 87.970 ;
        RECT 148.810 86.385 149.010 86.585 ;
        RECT 148.825 85.035 149.025 85.235 ;
        RECT 148.790 83.645 148.990 83.845 ;
        RECT 148.795 82.275 148.995 82.475 ;
        RECT 148.820 80.885 149.020 81.085 ;
        RECT 17.295 80.475 17.495 80.675 ;
        RECT 18.635 80.485 18.835 80.685 ;
        RECT 16.410 80.130 16.580 80.330 ;
        RECT 26.910 80.475 27.110 80.675 ;
        RECT 28.250 80.485 28.450 80.685 ;
        RECT 26.025 80.130 26.195 80.330 ;
        RECT 36.525 80.475 36.725 80.675 ;
        RECT 37.865 80.485 38.065 80.685 ;
        RECT 35.640 80.130 35.810 80.330 ;
        RECT 46.140 80.475 46.340 80.675 ;
        RECT 47.480 80.485 47.680 80.685 ;
        RECT 45.255 80.130 45.425 80.330 ;
        RECT 148.820 79.530 149.020 79.730 ;
        RECT 148.800 78.135 149.000 78.335 ;
        RECT 12.480 77.490 12.650 77.660 ;
        RECT 13.070 77.490 13.240 77.660 ;
        RECT 13.660 77.490 13.830 77.660 ;
        RECT 14.250 77.490 14.420 77.660 ;
        RECT 14.840 77.490 15.010 77.660 ;
        RECT 15.430 77.490 15.600 77.660 ;
        RECT 16.020 77.490 16.190 77.660 ;
        RECT 16.610 77.490 16.780 77.660 ;
        RECT 17.200 77.490 17.370 77.660 ;
        RECT 17.790 77.490 17.960 77.660 ;
        RECT 22.095 77.490 22.265 77.660 ;
        RECT 22.685 77.490 22.855 77.660 ;
        RECT 23.275 77.490 23.445 77.660 ;
        RECT 23.865 77.490 24.035 77.660 ;
        RECT 24.455 77.490 24.625 77.660 ;
        RECT 25.045 77.490 25.215 77.660 ;
        RECT 25.635 77.490 25.805 77.660 ;
        RECT 26.225 77.490 26.395 77.660 ;
        RECT 26.815 77.490 26.985 77.660 ;
        RECT 27.405 77.490 27.575 77.660 ;
        RECT 31.710 77.490 31.880 77.660 ;
        RECT 32.300 77.490 32.470 77.660 ;
        RECT 32.890 77.490 33.060 77.660 ;
        RECT 33.480 77.490 33.650 77.660 ;
        RECT 34.070 77.490 34.240 77.660 ;
        RECT 34.660 77.490 34.830 77.660 ;
        RECT 35.250 77.490 35.420 77.660 ;
        RECT 35.840 77.490 36.010 77.660 ;
        RECT 36.430 77.490 36.600 77.660 ;
        RECT 37.020 77.490 37.190 77.660 ;
        RECT 41.325 77.490 41.495 77.660 ;
        RECT 41.915 77.490 42.085 77.660 ;
        RECT 42.505 77.490 42.675 77.660 ;
        RECT 43.095 77.490 43.265 77.660 ;
        RECT 43.685 77.490 43.855 77.660 ;
        RECT 44.275 77.490 44.445 77.660 ;
        RECT 44.865 77.490 45.035 77.660 ;
        RECT 45.455 77.490 45.625 77.660 ;
        RECT 46.045 77.490 46.215 77.660 ;
        RECT 46.635 77.490 46.805 77.660 ;
        RECT 12.775 76.535 12.945 77.065 ;
        RECT 13.955 76.535 14.125 77.065 ;
        RECT 15.135 76.535 15.305 77.065 ;
        RECT 16.315 76.535 16.485 77.065 ;
        RECT 17.495 76.535 17.665 77.065 ;
        RECT 22.390 76.535 22.560 77.065 ;
        RECT 23.570 76.535 23.740 77.065 ;
        RECT 24.750 76.535 24.920 77.065 ;
        RECT 25.930 76.535 26.100 77.065 ;
        RECT 27.110 76.535 27.280 77.065 ;
        RECT 32.005 76.535 32.175 77.065 ;
        RECT 33.185 76.535 33.355 77.065 ;
        RECT 34.365 76.535 34.535 77.065 ;
        RECT 35.545 76.535 35.715 77.065 ;
        RECT 36.725 76.535 36.895 77.065 ;
        RECT 41.620 76.535 41.790 77.065 ;
        RECT 42.800 76.535 42.970 77.065 ;
        RECT 43.980 76.535 44.150 77.065 ;
        RECT 45.160 76.535 45.330 77.065 ;
        RECT 46.340 76.535 46.510 77.065 ;
        RECT 148.790 76.765 148.990 76.965 ;
        RECT 12.785 74.050 12.955 74.580 ;
        RECT 13.965 74.050 14.135 74.580 ;
        RECT 15.145 74.050 15.315 74.580 ;
        RECT 16.325 74.050 16.495 74.580 ;
        RECT 17.505 74.050 17.675 74.580 ;
        RECT 22.400 74.050 22.570 74.580 ;
        RECT 23.580 74.050 23.750 74.580 ;
        RECT 24.760 74.050 24.930 74.580 ;
        RECT 25.940 74.050 26.110 74.580 ;
        RECT 27.120 74.050 27.290 74.580 ;
        RECT 32.015 74.050 32.185 74.580 ;
        RECT 33.195 74.050 33.365 74.580 ;
        RECT 34.375 74.050 34.545 74.580 ;
        RECT 35.555 74.050 35.725 74.580 ;
        RECT 36.735 74.050 36.905 74.580 ;
        RECT 41.630 74.050 41.800 74.580 ;
        RECT 42.810 74.050 42.980 74.580 ;
        RECT 43.990 74.050 44.160 74.580 ;
        RECT 45.170 74.050 45.340 74.580 ;
        RECT 46.350 74.050 46.520 74.580 ;
        RECT 12.490 73.410 12.660 73.580 ;
        RECT 13.080 73.410 13.250 73.580 ;
        RECT 13.670 73.410 13.840 73.580 ;
        RECT 14.260 73.410 14.430 73.580 ;
        RECT 14.850 73.410 15.020 73.580 ;
        RECT 15.440 73.410 15.610 73.580 ;
        RECT 16.030 73.410 16.200 73.580 ;
        RECT 16.620 73.410 16.790 73.580 ;
        RECT 17.210 73.410 17.380 73.580 ;
        RECT 17.800 73.410 17.970 73.580 ;
        RECT 22.105 73.410 22.275 73.580 ;
        RECT 22.695 73.410 22.865 73.580 ;
        RECT 23.285 73.410 23.455 73.580 ;
        RECT 23.875 73.410 24.045 73.580 ;
        RECT 24.465 73.410 24.635 73.580 ;
        RECT 25.055 73.410 25.225 73.580 ;
        RECT 25.645 73.410 25.815 73.580 ;
        RECT 26.235 73.410 26.405 73.580 ;
        RECT 26.825 73.410 26.995 73.580 ;
        RECT 27.415 73.410 27.585 73.580 ;
        RECT 31.720 73.410 31.890 73.580 ;
        RECT 32.310 73.410 32.480 73.580 ;
        RECT 32.900 73.410 33.070 73.580 ;
        RECT 33.490 73.410 33.660 73.580 ;
        RECT 34.080 73.410 34.250 73.580 ;
        RECT 34.670 73.410 34.840 73.580 ;
        RECT 35.260 73.410 35.430 73.580 ;
        RECT 35.850 73.410 36.020 73.580 ;
        RECT 36.440 73.410 36.610 73.580 ;
        RECT 37.030 73.410 37.200 73.580 ;
        RECT 41.335 73.410 41.505 73.580 ;
        RECT 41.925 73.410 42.095 73.580 ;
        RECT 42.515 73.410 42.685 73.580 ;
        RECT 43.105 73.410 43.275 73.580 ;
        RECT 43.695 73.410 43.865 73.580 ;
        RECT 44.285 73.410 44.455 73.580 ;
        RECT 44.875 73.410 45.045 73.580 ;
        RECT 45.465 73.410 45.635 73.580 ;
        RECT 46.055 73.410 46.225 73.580 ;
        RECT 46.645 73.410 46.815 73.580 ;
        RECT 166.745 68.885 167.445 69.055 ;
        RECT 169.540 68.950 170.240 69.120 ;
        RECT 150.590 68.105 150.760 68.805 ;
        RECT 151.770 68.105 151.940 68.805 ;
        RECT 152.950 68.105 153.120 68.805 ;
        RECT 154.130 68.105 154.300 68.805 ;
        RECT 155.310 68.105 155.480 68.805 ;
        RECT 158.580 68.060 158.750 68.850 ;
        RECT 159.760 68.060 159.930 68.850 ;
        RECT 160.940 68.060 161.110 68.850 ;
        RECT 163.485 68.105 163.655 68.805 ;
        RECT 164.665 68.105 164.835 68.805 ;
        RECT 174.105 64.990 174.275 65.160 ;
        RECT 175.935 64.990 176.105 65.160 ;
        RECT 173.150 64.645 173.320 64.815 ;
        RECT 173.510 64.645 173.680 64.815 ;
        RECT 176.575 64.645 176.745 64.815 ;
        RECT 176.935 64.645 177.105 64.815 ;
        RECT 174.105 63.420 174.275 63.590 ;
        RECT 173.150 63.075 173.320 63.245 ;
        RECT 173.510 63.075 173.680 63.245 ;
        RECT 174.105 61.850 174.275 62.020 ;
        RECT 175.935 61.850 176.105 62.020 ;
        RECT 154.295 60.835 154.465 61.535 ;
        RECT 155.995 60.945 156.165 61.475 ;
        RECT 156.585 60.860 156.755 61.560 ;
        RECT 158.295 60.960 158.465 61.490 ;
        RECT 158.885 60.875 159.055 61.575 ;
        RECT 161.065 61.265 161.765 61.435 ;
        RECT 162.570 61.265 163.270 61.435 ;
        RECT 164.395 61.265 165.095 61.435 ;
        RECT 160.510 60.970 160.680 61.140 ;
        RECT 156.290 60.350 156.460 60.520 ;
        RECT 158.590 60.365 158.760 60.535 ;
        RECT 156.290 59.770 156.460 59.940 ;
        RECT 158.590 59.785 158.760 59.955 ;
        RECT 173.150 59.835 173.320 60.005 ;
        RECT 173.510 59.835 173.680 60.005 ;
        RECT 176.575 59.835 176.745 60.005 ;
        RECT 176.935 59.835 177.105 60.005 ;
        RECT 154.295 58.705 154.465 59.405 ;
        RECT 155.995 58.815 156.165 59.345 ;
        RECT 156.585 58.730 156.755 59.430 ;
        RECT 158.295 58.830 158.465 59.360 ;
        RECT 158.885 58.745 159.055 59.445 ;
        RECT 160.510 59.175 160.680 59.345 ;
        RECT 161.065 58.880 161.765 59.050 ;
        RECT 162.570 58.880 163.270 59.050 ;
        RECT 164.395 58.880 165.095 59.050 ;
        RECT 174.105 57.920 174.275 58.090 ;
        RECT 173.150 56.695 173.320 56.865 ;
        RECT 173.510 56.695 173.680 56.865 ;
        RECT 176.575 56.695 176.745 56.865 ;
        RECT 176.935 56.695 177.105 56.865 ;
        RECT 174.105 56.350 174.275 56.520 ;
        RECT 175.935 56.350 176.105 56.520 ;
        RECT 150.705 51.175 150.875 51.875 ;
        RECT 151.885 51.175 152.055 51.875 ;
        RECT 153.065 51.175 153.235 51.875 ;
        RECT 154.245 51.175 154.415 51.875 ;
        RECT 155.425 51.175 155.595 51.875 ;
        RECT 158.695 51.130 158.865 51.920 ;
        RECT 159.875 51.130 160.045 51.920 ;
        RECT 161.055 51.130 161.225 51.920 ;
        RECT 163.600 51.175 163.770 51.875 ;
        RECT 164.780 51.175 164.950 51.875 ;
        RECT 166.860 50.925 167.560 51.095 ;
        RECT 169.655 50.860 170.355 51.030 ;
        RECT 12.490 46.270 12.660 46.440 ;
        RECT 13.080 46.270 13.250 46.440 ;
        RECT 13.670 46.270 13.840 46.440 ;
        RECT 14.260 46.270 14.430 46.440 ;
        RECT 14.850 46.270 15.020 46.440 ;
        RECT 15.440 46.270 15.610 46.440 ;
        RECT 16.030 46.270 16.200 46.440 ;
        RECT 16.620 46.270 16.790 46.440 ;
        RECT 17.210 46.270 17.380 46.440 ;
        RECT 17.800 46.270 17.970 46.440 ;
        RECT 22.105 46.270 22.275 46.440 ;
        RECT 22.695 46.270 22.865 46.440 ;
        RECT 23.285 46.270 23.455 46.440 ;
        RECT 23.875 46.270 24.045 46.440 ;
        RECT 24.465 46.270 24.635 46.440 ;
        RECT 25.055 46.270 25.225 46.440 ;
        RECT 25.645 46.270 25.815 46.440 ;
        RECT 26.235 46.270 26.405 46.440 ;
        RECT 26.825 46.270 26.995 46.440 ;
        RECT 27.415 46.270 27.585 46.440 ;
        RECT 31.720 46.270 31.890 46.440 ;
        RECT 32.310 46.270 32.480 46.440 ;
        RECT 32.900 46.270 33.070 46.440 ;
        RECT 33.490 46.270 33.660 46.440 ;
        RECT 34.080 46.270 34.250 46.440 ;
        RECT 34.670 46.270 34.840 46.440 ;
        RECT 35.260 46.270 35.430 46.440 ;
        RECT 35.850 46.270 36.020 46.440 ;
        RECT 36.440 46.270 36.610 46.440 ;
        RECT 37.030 46.270 37.200 46.440 ;
        RECT 41.335 46.270 41.505 46.440 ;
        RECT 41.925 46.270 42.095 46.440 ;
        RECT 42.515 46.270 42.685 46.440 ;
        RECT 43.105 46.270 43.275 46.440 ;
        RECT 43.695 46.270 43.865 46.440 ;
        RECT 44.285 46.270 44.455 46.440 ;
        RECT 44.875 46.270 45.045 46.440 ;
        RECT 45.465 46.270 45.635 46.440 ;
        RECT 46.055 46.270 46.225 46.440 ;
        RECT 46.645 46.270 46.815 46.440 ;
        RECT 12.785 45.270 12.955 45.800 ;
        RECT 13.965 45.270 14.135 45.800 ;
        RECT 15.145 45.270 15.315 45.800 ;
        RECT 16.325 45.270 16.495 45.800 ;
        RECT 17.505 45.270 17.675 45.800 ;
        RECT 22.400 45.270 22.570 45.800 ;
        RECT 23.580 45.270 23.750 45.800 ;
        RECT 24.760 45.270 24.930 45.800 ;
        RECT 25.940 45.270 26.110 45.800 ;
        RECT 27.120 45.270 27.290 45.800 ;
        RECT 32.015 45.270 32.185 45.800 ;
        RECT 33.195 45.270 33.365 45.800 ;
        RECT 34.375 45.270 34.545 45.800 ;
        RECT 35.555 45.270 35.725 45.800 ;
        RECT 36.735 45.270 36.905 45.800 ;
        RECT 41.630 45.270 41.800 45.800 ;
        RECT 42.810 45.270 42.980 45.800 ;
        RECT 43.990 45.270 44.160 45.800 ;
        RECT 45.170 45.270 45.340 45.800 ;
        RECT 46.350 45.270 46.520 45.800 ;
        RECT 12.775 42.785 12.945 43.315 ;
        RECT 13.955 42.785 14.125 43.315 ;
        RECT 15.135 42.785 15.305 43.315 ;
        RECT 16.315 42.785 16.485 43.315 ;
        RECT 17.495 42.785 17.665 43.315 ;
        RECT 22.390 42.785 22.560 43.315 ;
        RECT 23.570 42.785 23.740 43.315 ;
        RECT 24.750 42.785 24.920 43.315 ;
        RECT 25.930 42.785 26.100 43.315 ;
        RECT 27.110 42.785 27.280 43.315 ;
        RECT 32.005 42.785 32.175 43.315 ;
        RECT 33.185 42.785 33.355 43.315 ;
        RECT 34.365 42.785 34.535 43.315 ;
        RECT 35.545 42.785 35.715 43.315 ;
        RECT 36.725 42.785 36.895 43.315 ;
        RECT 41.620 42.785 41.790 43.315 ;
        RECT 42.800 42.785 42.970 43.315 ;
        RECT 43.980 42.785 44.150 43.315 ;
        RECT 45.160 42.785 45.330 43.315 ;
        RECT 46.340 42.785 46.510 43.315 ;
        RECT 148.790 42.885 148.990 43.085 ;
        RECT 12.480 42.190 12.650 42.360 ;
        RECT 13.070 42.190 13.240 42.360 ;
        RECT 13.660 42.190 13.830 42.360 ;
        RECT 14.250 42.190 14.420 42.360 ;
        RECT 14.840 42.190 15.010 42.360 ;
        RECT 15.430 42.190 15.600 42.360 ;
        RECT 16.020 42.190 16.190 42.360 ;
        RECT 16.610 42.190 16.780 42.360 ;
        RECT 17.200 42.190 17.370 42.360 ;
        RECT 17.790 42.190 17.960 42.360 ;
        RECT 22.095 42.190 22.265 42.360 ;
        RECT 22.685 42.190 22.855 42.360 ;
        RECT 23.275 42.190 23.445 42.360 ;
        RECT 23.865 42.190 24.035 42.360 ;
        RECT 24.455 42.190 24.625 42.360 ;
        RECT 25.045 42.190 25.215 42.360 ;
        RECT 25.635 42.190 25.805 42.360 ;
        RECT 26.225 42.190 26.395 42.360 ;
        RECT 26.815 42.190 26.985 42.360 ;
        RECT 27.405 42.190 27.575 42.360 ;
        RECT 31.710 42.190 31.880 42.360 ;
        RECT 32.300 42.190 32.470 42.360 ;
        RECT 32.890 42.190 33.060 42.360 ;
        RECT 33.480 42.190 33.650 42.360 ;
        RECT 34.070 42.190 34.240 42.360 ;
        RECT 34.660 42.190 34.830 42.360 ;
        RECT 35.250 42.190 35.420 42.360 ;
        RECT 35.840 42.190 36.010 42.360 ;
        RECT 36.430 42.190 36.600 42.360 ;
        RECT 37.020 42.190 37.190 42.360 ;
        RECT 41.325 42.190 41.495 42.360 ;
        RECT 41.915 42.190 42.085 42.360 ;
        RECT 42.505 42.190 42.675 42.360 ;
        RECT 43.095 42.190 43.265 42.360 ;
        RECT 43.685 42.190 43.855 42.360 ;
        RECT 44.275 42.190 44.445 42.360 ;
        RECT 44.865 42.190 45.035 42.360 ;
        RECT 45.455 42.190 45.625 42.360 ;
        RECT 46.045 42.190 46.215 42.360 ;
        RECT 46.635 42.190 46.805 42.360 ;
        RECT 148.800 41.515 149.000 41.715 ;
        RECT 16.410 39.520 16.580 39.720 ;
        RECT 17.295 39.175 17.495 39.375 ;
        RECT 18.635 39.165 18.835 39.365 ;
        RECT 26.025 39.520 26.195 39.720 ;
        RECT 26.910 39.175 27.110 39.375 ;
        RECT 28.250 39.165 28.450 39.365 ;
        RECT 35.640 39.520 35.810 39.720 ;
        RECT 148.820 40.120 149.020 40.320 ;
        RECT 36.525 39.175 36.725 39.375 ;
        RECT 37.865 39.165 38.065 39.365 ;
        RECT 45.255 39.520 45.425 39.720 ;
        RECT 46.140 39.175 46.340 39.375 ;
        RECT 47.480 39.165 47.680 39.365 ;
        RECT 148.820 38.765 149.020 38.965 ;
        RECT 148.795 37.375 148.995 37.575 ;
        RECT 148.790 36.005 148.990 36.205 ;
        RECT 148.825 34.615 149.025 34.815 ;
        RECT 148.810 33.265 149.010 33.465 ;
        RECT 148.820 31.880 149.020 32.080 ;
      LAYER met1 ;
        RECT 148.790 87.710 149.050 88.030 ;
        RECT 148.780 86.325 149.040 86.645 ;
        RECT 148.795 84.975 149.055 85.295 ;
        RECT 148.760 83.585 149.020 83.905 ;
        RECT 148.765 82.215 149.025 82.535 ;
        RECT 148.790 80.825 149.050 81.145 ;
        RECT 17.265 80.415 17.525 80.735 ;
        RECT 18.575 80.455 18.895 80.715 ;
        RECT 26.880 80.415 27.140 80.735 ;
        RECT 28.190 80.455 28.510 80.715 ;
        RECT 36.495 80.415 36.755 80.735 ;
        RECT 37.805 80.455 38.125 80.715 ;
        RECT 46.110 80.415 46.370 80.735 ;
        RECT 47.420 80.455 47.740 80.715 ;
        RECT 16.320 80.100 16.640 80.360 ;
        RECT 25.935 80.100 26.255 80.360 ;
        RECT 35.550 80.100 35.870 80.360 ;
        RECT 45.165 80.100 45.485 80.360 ;
        RECT 148.790 79.470 149.050 79.790 ;
        RECT 148.770 78.075 149.030 78.395 ;
        RECT 17.990 77.690 18.310 77.710 ;
        RECT 27.605 77.690 27.925 77.710 ;
        RECT 37.220 77.690 37.540 77.710 ;
        RECT 46.835 77.690 47.155 77.710 ;
        RECT 12.420 77.680 12.710 77.690 ;
        RECT 13.010 77.680 13.300 77.690 ;
        RECT 13.600 77.680 13.890 77.690 ;
        RECT 14.190 77.680 14.480 77.690 ;
        RECT 14.780 77.680 15.070 77.690 ;
        RECT 15.370 77.680 15.660 77.690 ;
        RECT 15.960 77.680 16.250 77.690 ;
        RECT 16.550 77.680 16.840 77.690 ;
        RECT 17.140 77.680 17.430 77.690 ;
        RECT 17.730 77.680 18.310 77.690 ;
        RECT 12.420 77.485 18.310 77.680 ;
        RECT 12.420 77.460 12.710 77.485 ;
        RECT 13.010 77.460 13.300 77.485 ;
        RECT 13.600 77.460 13.890 77.485 ;
        RECT 14.190 77.460 14.480 77.485 ;
        RECT 14.780 77.460 15.070 77.485 ;
        RECT 15.370 77.460 15.660 77.485 ;
        RECT 15.960 77.460 16.250 77.485 ;
        RECT 16.550 77.460 16.840 77.485 ;
        RECT 17.140 77.460 17.430 77.485 ;
        RECT 17.730 77.460 18.310 77.485 ;
        RECT 22.035 77.680 22.325 77.690 ;
        RECT 22.625 77.680 22.915 77.690 ;
        RECT 23.215 77.680 23.505 77.690 ;
        RECT 23.805 77.680 24.095 77.690 ;
        RECT 24.395 77.680 24.685 77.690 ;
        RECT 24.985 77.680 25.275 77.690 ;
        RECT 25.575 77.680 25.865 77.690 ;
        RECT 26.165 77.680 26.455 77.690 ;
        RECT 26.755 77.680 27.045 77.690 ;
        RECT 27.345 77.680 27.925 77.690 ;
        RECT 22.035 77.485 27.925 77.680 ;
        RECT 22.035 77.460 22.325 77.485 ;
        RECT 22.625 77.460 22.915 77.485 ;
        RECT 23.215 77.460 23.505 77.485 ;
        RECT 23.805 77.460 24.095 77.485 ;
        RECT 24.395 77.460 24.685 77.485 ;
        RECT 24.985 77.460 25.275 77.485 ;
        RECT 25.575 77.460 25.865 77.485 ;
        RECT 26.165 77.460 26.455 77.485 ;
        RECT 26.755 77.460 27.045 77.485 ;
        RECT 27.345 77.460 27.925 77.485 ;
        RECT 31.650 77.680 31.940 77.690 ;
        RECT 32.240 77.680 32.530 77.690 ;
        RECT 32.830 77.680 33.120 77.690 ;
        RECT 33.420 77.680 33.710 77.690 ;
        RECT 34.010 77.680 34.300 77.690 ;
        RECT 34.600 77.680 34.890 77.690 ;
        RECT 35.190 77.680 35.480 77.690 ;
        RECT 35.780 77.680 36.070 77.690 ;
        RECT 36.370 77.680 36.660 77.690 ;
        RECT 36.960 77.680 37.540 77.690 ;
        RECT 31.650 77.485 37.540 77.680 ;
        RECT 31.650 77.460 31.940 77.485 ;
        RECT 32.240 77.460 32.530 77.485 ;
        RECT 32.830 77.460 33.120 77.485 ;
        RECT 33.420 77.460 33.710 77.485 ;
        RECT 34.010 77.460 34.300 77.485 ;
        RECT 34.600 77.460 34.890 77.485 ;
        RECT 35.190 77.460 35.480 77.485 ;
        RECT 35.780 77.460 36.070 77.485 ;
        RECT 36.370 77.460 36.660 77.485 ;
        RECT 36.960 77.460 37.540 77.485 ;
        RECT 41.265 77.680 41.555 77.690 ;
        RECT 41.855 77.680 42.145 77.690 ;
        RECT 42.445 77.680 42.735 77.690 ;
        RECT 43.035 77.680 43.325 77.690 ;
        RECT 43.625 77.680 43.915 77.690 ;
        RECT 44.215 77.680 44.505 77.690 ;
        RECT 44.805 77.680 45.095 77.690 ;
        RECT 45.395 77.680 45.685 77.690 ;
        RECT 45.985 77.680 46.275 77.690 ;
        RECT 46.575 77.680 47.155 77.690 ;
        RECT 41.265 77.485 47.155 77.680 ;
        RECT 41.265 77.460 41.555 77.485 ;
        RECT 41.855 77.460 42.145 77.485 ;
        RECT 42.445 77.460 42.735 77.485 ;
        RECT 43.035 77.460 43.325 77.485 ;
        RECT 43.625 77.460 43.915 77.485 ;
        RECT 44.215 77.460 44.505 77.485 ;
        RECT 44.805 77.460 45.095 77.485 ;
        RECT 45.395 77.460 45.685 77.485 ;
        RECT 45.985 77.460 46.275 77.485 ;
        RECT 46.575 77.460 47.155 77.485 ;
        RECT 17.990 77.450 18.310 77.460 ;
        RECT 27.605 77.450 27.925 77.460 ;
        RECT 37.220 77.450 37.540 77.460 ;
        RECT 46.835 77.450 47.155 77.460 ;
        RECT 12.745 76.760 12.975 77.125 ;
        RECT 13.925 76.840 14.155 77.125 ;
        RECT 15.105 76.890 15.335 77.125 ;
        RECT 16.285 76.920 16.515 77.125 ;
        RECT 15.095 76.860 15.355 76.890 ;
        RECT 12.720 76.500 13.040 76.760 ;
        RECT 13.885 76.580 14.205 76.840 ;
        RECT 15.065 76.600 15.385 76.860 ;
        RECT 16.255 76.660 16.575 76.920 ;
        RECT 17.465 76.900 17.695 77.125 ;
        RECT 12.745 76.475 12.975 76.500 ;
        RECT 13.925 76.475 14.155 76.580 ;
        RECT 15.095 76.570 15.355 76.600 ;
        RECT 15.105 76.475 15.335 76.570 ;
        RECT 16.285 76.475 16.515 76.660 ;
        RECT 17.425 76.640 17.745 76.900 ;
        RECT 22.360 76.760 22.590 77.125 ;
        RECT 23.540 76.840 23.770 77.125 ;
        RECT 24.720 76.890 24.950 77.125 ;
        RECT 25.900 76.920 26.130 77.125 ;
        RECT 24.710 76.860 24.970 76.890 ;
        RECT 17.465 76.475 17.695 76.640 ;
        RECT 22.335 76.500 22.655 76.760 ;
        RECT 23.500 76.580 23.820 76.840 ;
        RECT 24.680 76.600 25.000 76.860 ;
        RECT 25.870 76.660 26.190 76.920 ;
        RECT 27.080 76.900 27.310 77.125 ;
        RECT 22.360 76.475 22.590 76.500 ;
        RECT 23.540 76.475 23.770 76.580 ;
        RECT 24.710 76.570 24.970 76.600 ;
        RECT 24.720 76.475 24.950 76.570 ;
        RECT 25.900 76.475 26.130 76.660 ;
        RECT 27.040 76.640 27.360 76.900 ;
        RECT 31.975 76.760 32.205 77.125 ;
        RECT 33.155 76.840 33.385 77.125 ;
        RECT 34.335 76.890 34.565 77.125 ;
        RECT 35.515 76.920 35.745 77.125 ;
        RECT 34.325 76.860 34.585 76.890 ;
        RECT 27.080 76.475 27.310 76.640 ;
        RECT 31.950 76.500 32.270 76.760 ;
        RECT 33.115 76.580 33.435 76.840 ;
        RECT 34.295 76.600 34.615 76.860 ;
        RECT 35.485 76.660 35.805 76.920 ;
        RECT 36.695 76.900 36.925 77.125 ;
        RECT 31.975 76.475 32.205 76.500 ;
        RECT 33.155 76.475 33.385 76.580 ;
        RECT 34.325 76.570 34.585 76.600 ;
        RECT 34.335 76.475 34.565 76.570 ;
        RECT 35.515 76.475 35.745 76.660 ;
        RECT 36.655 76.640 36.975 76.900 ;
        RECT 41.590 76.760 41.820 77.125 ;
        RECT 42.770 76.840 43.000 77.125 ;
        RECT 43.950 76.890 44.180 77.125 ;
        RECT 45.130 76.920 45.360 77.125 ;
        RECT 43.940 76.860 44.200 76.890 ;
        RECT 36.695 76.475 36.925 76.640 ;
        RECT 41.565 76.500 41.885 76.760 ;
        RECT 42.730 76.580 43.050 76.840 ;
        RECT 43.910 76.600 44.230 76.860 ;
        RECT 45.100 76.660 45.420 76.920 ;
        RECT 46.310 76.900 46.540 77.125 ;
        RECT 41.590 76.475 41.820 76.500 ;
        RECT 42.770 76.475 43.000 76.580 ;
        RECT 43.940 76.570 44.200 76.600 ;
        RECT 43.950 76.475 44.180 76.570 ;
        RECT 45.130 76.475 45.360 76.660 ;
        RECT 46.270 76.640 46.590 76.900 ;
        RECT 148.760 76.705 149.020 77.025 ;
        RECT 46.310 76.475 46.540 76.640 ;
        RECT 132.675 75.370 133.095 75.400 ;
        RECT 132.675 74.950 143.490 75.370 ;
        RECT 132.675 74.920 133.095 74.950 ;
        RECT 12.720 74.480 13.040 74.740 ;
        RECT 13.915 74.730 14.175 74.760 ;
        RECT 12.755 73.990 12.985 74.480 ;
        RECT 13.885 74.470 14.205 74.730 ;
        RECT 15.065 74.470 15.385 74.730 ;
        RECT 16.255 74.470 16.575 74.730 ;
        RECT 17.425 74.470 17.745 74.730 ;
        RECT 22.335 74.480 22.655 74.740 ;
        RECT 23.530 74.730 23.790 74.760 ;
        RECT 13.915 74.440 14.175 74.470 ;
        RECT 13.935 73.990 14.165 74.440 ;
        RECT 15.115 73.990 15.345 74.470 ;
        RECT 16.295 73.990 16.525 74.470 ;
        RECT 17.475 73.990 17.705 74.470 ;
        RECT 22.370 73.990 22.600 74.480 ;
        RECT 23.500 74.470 23.820 74.730 ;
        RECT 24.680 74.470 25.000 74.730 ;
        RECT 25.870 74.470 26.190 74.730 ;
        RECT 27.040 74.470 27.360 74.730 ;
        RECT 31.950 74.480 32.270 74.740 ;
        RECT 33.145 74.730 33.405 74.760 ;
        RECT 23.530 74.440 23.790 74.470 ;
        RECT 23.550 73.990 23.780 74.440 ;
        RECT 24.730 73.990 24.960 74.470 ;
        RECT 25.910 73.990 26.140 74.470 ;
        RECT 27.090 73.990 27.320 74.470 ;
        RECT 31.985 73.990 32.215 74.480 ;
        RECT 33.115 74.470 33.435 74.730 ;
        RECT 34.295 74.470 34.615 74.730 ;
        RECT 35.485 74.470 35.805 74.730 ;
        RECT 36.655 74.470 36.975 74.730 ;
        RECT 41.565 74.480 41.885 74.740 ;
        RECT 42.760 74.730 43.020 74.760 ;
        RECT 33.145 74.440 33.405 74.470 ;
        RECT 33.165 73.990 33.395 74.440 ;
        RECT 34.345 73.990 34.575 74.470 ;
        RECT 35.525 73.990 35.755 74.470 ;
        RECT 36.705 73.990 36.935 74.470 ;
        RECT 41.600 73.990 41.830 74.480 ;
        RECT 42.730 74.470 43.050 74.730 ;
        RECT 43.910 74.470 44.230 74.730 ;
        RECT 45.100 74.470 45.420 74.730 ;
        RECT 46.270 74.470 46.590 74.730 ;
        RECT 148.615 74.500 149.225 74.735 ;
        RECT 151.645 74.500 152.255 74.715 ;
        RECT 154.655 74.500 155.265 74.745 ;
        RECT 157.685 74.500 158.295 74.725 ;
        RECT 160.655 74.500 161.265 74.745 ;
        RECT 163.695 74.500 164.305 74.750 ;
        RECT 166.695 74.500 167.305 74.755 ;
        RECT 169.725 74.500 170.335 74.735 ;
        RECT 42.760 74.440 43.020 74.470 ;
        RECT 42.780 73.990 43.010 74.440 ;
        RECT 43.960 73.990 44.190 74.470 ;
        RECT 45.140 73.990 45.370 74.470 ;
        RECT 46.320 73.990 46.550 74.470 ;
        RECT 147.975 74.355 170.335 74.500 ;
        RECT 12.445 73.610 12.705 73.630 ;
        RECT 17.095 73.610 17.355 73.650 ;
        RECT 22.060 73.610 22.320 73.630 ;
        RECT 26.710 73.610 26.970 73.650 ;
        RECT 31.675 73.610 31.935 73.630 ;
        RECT 36.325 73.610 36.585 73.650 ;
        RECT 41.290 73.610 41.550 73.630 ;
        RECT 45.940 73.610 46.200 73.650 ;
        RECT 12.430 73.590 12.720 73.610 ;
        RECT 13.020 73.590 13.310 73.610 ;
        RECT 13.610 73.590 13.900 73.610 ;
        RECT 14.200 73.590 14.490 73.610 ;
        RECT 14.790 73.590 15.080 73.610 ;
        RECT 15.380 73.590 15.670 73.610 ;
        RECT 15.970 73.590 16.260 73.610 ;
        RECT 16.560 73.590 16.850 73.610 ;
        RECT 17.095 73.590 17.440 73.610 ;
        RECT 17.740 73.590 18.030 73.610 ;
        RECT 12.430 73.395 18.030 73.590 ;
        RECT 12.430 73.380 13.360 73.395 ;
        RECT 13.610 73.380 13.900 73.395 ;
        RECT 14.200 73.380 14.490 73.395 ;
        RECT 14.790 73.380 15.080 73.395 ;
        RECT 15.380 73.380 15.670 73.395 ;
        RECT 15.970 73.380 16.260 73.395 ;
        RECT 16.560 73.380 16.850 73.395 ;
        RECT 17.095 73.380 17.440 73.395 ;
        RECT 17.740 73.380 18.030 73.395 ;
        RECT 22.045 73.590 22.335 73.610 ;
        RECT 22.635 73.590 22.925 73.610 ;
        RECT 23.225 73.590 23.515 73.610 ;
        RECT 23.815 73.590 24.105 73.610 ;
        RECT 24.405 73.590 24.695 73.610 ;
        RECT 24.995 73.590 25.285 73.610 ;
        RECT 25.585 73.590 25.875 73.610 ;
        RECT 26.175 73.590 26.465 73.610 ;
        RECT 26.710 73.590 27.055 73.610 ;
        RECT 27.355 73.590 27.645 73.610 ;
        RECT 22.045 73.395 27.645 73.590 ;
        RECT 22.045 73.380 22.975 73.395 ;
        RECT 23.225 73.380 23.515 73.395 ;
        RECT 23.815 73.380 24.105 73.395 ;
        RECT 24.405 73.380 24.695 73.395 ;
        RECT 24.995 73.380 25.285 73.395 ;
        RECT 25.585 73.380 25.875 73.395 ;
        RECT 26.175 73.380 26.465 73.395 ;
        RECT 26.710 73.380 27.055 73.395 ;
        RECT 27.355 73.380 27.645 73.395 ;
        RECT 31.660 73.590 31.950 73.610 ;
        RECT 32.250 73.590 32.540 73.610 ;
        RECT 32.840 73.590 33.130 73.610 ;
        RECT 33.430 73.590 33.720 73.610 ;
        RECT 34.020 73.590 34.310 73.610 ;
        RECT 34.610 73.590 34.900 73.610 ;
        RECT 35.200 73.590 35.490 73.610 ;
        RECT 35.790 73.590 36.080 73.610 ;
        RECT 36.325 73.590 36.670 73.610 ;
        RECT 36.970 73.590 37.260 73.610 ;
        RECT 31.660 73.395 37.260 73.590 ;
        RECT 31.660 73.380 32.590 73.395 ;
        RECT 32.840 73.380 33.130 73.395 ;
        RECT 33.430 73.380 33.720 73.395 ;
        RECT 34.020 73.380 34.310 73.395 ;
        RECT 34.610 73.380 34.900 73.395 ;
        RECT 35.200 73.380 35.490 73.395 ;
        RECT 35.790 73.380 36.080 73.395 ;
        RECT 36.325 73.380 36.670 73.395 ;
        RECT 36.970 73.380 37.260 73.395 ;
        RECT 41.275 73.590 41.565 73.610 ;
        RECT 41.865 73.590 42.155 73.610 ;
        RECT 42.455 73.590 42.745 73.610 ;
        RECT 43.045 73.590 43.335 73.610 ;
        RECT 43.635 73.590 43.925 73.610 ;
        RECT 44.225 73.590 44.515 73.610 ;
        RECT 44.815 73.590 45.105 73.610 ;
        RECT 45.405 73.590 45.695 73.610 ;
        RECT 45.940 73.590 46.285 73.610 ;
        RECT 46.585 73.590 46.875 73.610 ;
        RECT 41.275 73.395 46.875 73.590 ;
        RECT 41.275 73.380 42.205 73.395 ;
        RECT 42.455 73.380 42.745 73.395 ;
        RECT 43.045 73.380 43.335 73.395 ;
        RECT 43.635 73.380 43.925 73.395 ;
        RECT 44.225 73.380 44.515 73.395 ;
        RECT 44.815 73.380 45.105 73.395 ;
        RECT 45.405 73.380 45.695 73.395 ;
        RECT 45.940 73.380 46.285 73.395 ;
        RECT 46.585 73.380 46.875 73.395 ;
        RECT 12.445 73.370 13.360 73.380 ;
        RECT 12.445 73.310 12.705 73.370 ;
        RECT 17.095 73.330 17.355 73.380 ;
        RECT 22.060 73.370 22.975 73.380 ;
        RECT 22.060 73.310 22.320 73.370 ;
        RECT 26.710 73.330 26.970 73.380 ;
        RECT 31.675 73.370 32.590 73.380 ;
        RECT 31.675 73.310 31.935 73.370 ;
        RECT 36.325 73.330 36.585 73.380 ;
        RECT 41.290 73.370 42.205 73.380 ;
        RECT 41.290 73.310 41.550 73.370 ;
        RECT 45.940 73.330 46.200 73.380 ;
        RECT 128.580 72.275 129.000 72.305 ;
        RECT 128.580 71.855 143.560 72.275 ;
        RECT 128.580 71.825 129.000 71.855 ;
        RECT 143.105 69.270 143.365 69.280 ;
        RECT 120.725 68.955 143.430 69.270 ;
        RECT 74.455 64.130 74.960 64.575 ;
        RECT 78.610 64.145 79.050 64.525 ;
        RECT 74.460 64.050 74.905 64.130 ;
        RECT 147.975 62.865 148.120 74.355 ;
        RECT 148.615 74.185 149.225 74.355 ;
        RECT 151.645 74.165 152.255 74.355 ;
        RECT 154.655 74.195 155.265 74.355 ;
        RECT 157.685 74.175 158.295 74.355 ;
        RECT 160.655 74.195 161.265 74.355 ;
        RECT 163.695 74.200 164.305 74.355 ;
        RECT 166.695 74.205 167.305 74.355 ;
        RECT 169.725 74.185 170.335 74.355 ;
        RECT 148.630 70.535 149.225 70.820 ;
        RECT 151.660 70.535 152.255 70.800 ;
        RECT 154.670 70.535 155.265 70.830 ;
        RECT 157.700 70.535 158.295 70.810 ;
        RECT 148.630 70.390 158.295 70.535 ;
        RECT 148.630 70.285 149.225 70.390 ;
        RECT 151.660 70.265 152.255 70.390 ;
        RECT 154.670 70.295 155.265 70.390 ;
        RECT 150.560 68.045 150.790 68.865 ;
        RECT 151.740 68.045 151.970 68.865 ;
        RECT 152.920 68.045 153.150 68.865 ;
        RECT 154.100 68.045 154.330 68.865 ;
        RECT 155.280 68.045 155.510 68.865 ;
        RECT 150.605 67.805 150.750 68.045 ;
        RECT 151.780 67.805 151.925 68.045 ;
        RECT 152.950 67.805 153.095 68.045 ;
        RECT 154.150 67.805 154.295 68.045 ;
        RECT 150.605 67.800 154.295 67.805 ;
        RECT 155.315 67.800 155.460 68.045 ;
        RECT 150.605 67.660 155.460 67.800 ;
        RECT 157.255 67.830 157.400 70.390 ;
        RECT 157.700 70.275 158.295 70.390 ;
        RECT 160.670 70.515 161.265 70.830 ;
        RECT 163.710 70.515 164.305 70.835 ;
        RECT 160.670 70.360 164.305 70.515 ;
        RECT 160.670 70.295 161.265 70.360 ;
        RECT 158.550 68.000 158.780 68.910 ;
        RECT 159.730 68.000 159.960 68.910 ;
        RECT 160.910 68.000 161.140 68.910 ;
        RECT 163.215 68.880 163.370 70.360 ;
        RECT 163.710 70.300 164.305 70.360 ;
        RECT 166.710 70.305 167.305 70.840 ;
        RECT 166.930 69.085 167.085 70.305 ;
        RECT 169.740 70.285 170.335 70.820 ;
        RECT 169.955 69.150 170.110 70.285 ;
        RECT 163.215 68.865 163.665 68.880 ;
        RECT 163.215 68.725 163.685 68.865 ;
        RECT 163.455 68.045 163.685 68.725 ;
        RECT 164.635 68.045 164.865 68.865 ;
        RECT 166.685 68.855 167.505 69.085 ;
        RECT 169.480 68.920 170.300 69.150 ;
        RECT 158.580 67.830 158.725 68.000 ;
        RECT 159.770 67.830 159.915 68.000 ;
        RECT 157.255 67.820 159.915 67.830 ;
        RECT 160.960 67.820 161.105 68.000 ;
        RECT 157.255 67.685 161.105 67.820 ;
        RECT 163.510 67.840 163.665 68.045 ;
        RECT 164.675 67.840 164.830 68.045 ;
        RECT 163.510 67.685 164.830 67.840 ;
        RECT 159.770 67.675 161.105 67.685 ;
        RECT 148.665 66.845 149.260 67.040 ;
        RECT 150.605 66.845 150.750 67.660 ;
        RECT 154.150 67.655 155.460 67.660 ;
        RECT 170.095 67.590 170.355 67.670 ;
        RECT 170.095 67.430 175.165 67.590 ;
        RECT 170.095 67.350 170.355 67.430 ;
        RECT 151.695 66.845 152.290 67.060 ;
        RECT 154.705 66.845 155.300 67.030 ;
        RECT 157.735 66.845 158.330 67.050 ;
        RECT 160.705 66.845 161.300 67.030 ;
        RECT 163.735 66.845 164.330 67.050 ;
        RECT 166.745 66.845 167.340 67.020 ;
        RECT 169.775 66.845 170.370 67.040 ;
        RECT 148.665 66.700 170.380 66.845 ;
        RECT 148.665 66.505 149.260 66.700 ;
        RECT 151.695 66.525 152.290 66.700 ;
        RECT 154.705 66.495 155.300 66.700 ;
        RECT 157.735 66.515 158.330 66.700 ;
        RECT 160.705 66.495 161.300 66.700 ;
        RECT 163.735 66.515 164.330 66.700 ;
        RECT 166.745 66.485 167.340 66.700 ;
        RECT 169.775 66.505 170.370 66.700 ;
        RECT 175.005 66.255 175.165 67.430 ;
        RECT 174.955 65.255 175.255 66.255 ;
        RECT 174.075 64.895 176.135 65.255 ;
        RECT 172.915 64.615 173.915 64.845 ;
        RECT 176.340 64.615 177.340 64.845 ;
        RECT 173.065 64.545 173.765 64.615 ;
        RECT 176.490 64.545 177.190 64.615 ;
        RECT 174.755 64.230 175.455 64.530 ;
        RECT 174.075 63.655 174.305 63.685 ;
        RECT 174.955 63.655 175.255 64.230 ;
        RECT 174.075 63.355 175.255 63.655 ;
        RECT 174.075 63.325 174.305 63.355 ;
        RECT 148.650 62.865 149.260 63.140 ;
        RECT 147.975 62.835 150.375 62.865 ;
        RECT 151.680 62.835 152.290 63.160 ;
        RECT 154.690 62.835 155.300 63.130 ;
        RECT 157.720 62.835 158.330 63.150 ;
        RECT 160.690 62.835 161.300 63.130 ;
        RECT 163.720 62.835 164.330 63.150 ;
        RECT 166.730 62.835 167.340 63.120 ;
        RECT 169.760 62.835 170.370 63.140 ;
        RECT 172.915 63.045 173.915 63.275 ;
        RECT 147.975 62.720 170.370 62.835 ;
        RECT 148.650 62.690 170.370 62.720 ;
        RECT 148.650 62.590 149.260 62.690 ;
        RECT 151.680 62.610 152.290 62.690 ;
        RECT 154.690 62.580 155.300 62.690 ;
        RECT 154.265 61.235 154.495 61.595 ;
        RECT 154.700 61.235 154.870 61.245 ;
        RECT 155.965 61.235 156.195 61.535 ;
        RECT 154.265 61.055 156.195 61.235 ;
        RECT 154.265 60.775 154.495 61.055 ;
        RECT 154.265 59.125 154.495 59.465 ;
        RECT 154.700 59.125 154.870 61.055 ;
        RECT 155.965 60.885 156.195 61.055 ;
        RECT 156.555 61.325 156.785 61.620 ;
        RECT 157.350 61.325 157.495 62.690 ;
        RECT 157.720 62.600 158.330 62.690 ;
        RECT 160.690 62.580 161.300 62.690 ;
        RECT 163.720 62.600 164.330 62.690 ;
        RECT 162.235 62.170 162.495 62.490 ;
        RECT 158.265 61.325 158.495 61.550 ;
        RECT 156.555 61.135 158.495 61.325 ;
        RECT 156.555 60.800 156.785 61.135 ;
        RECT 157.350 61.065 157.495 61.135 ;
        RECT 158.265 60.900 158.495 61.135 ;
        RECT 158.855 61.545 159.085 61.635 ;
        RECT 159.965 61.545 160.225 61.625 ;
        RECT 162.285 61.545 162.445 62.170 ;
        RECT 158.855 61.465 162.815 61.545 ;
        RECT 164.800 61.465 164.945 62.690 ;
        RECT 166.730 62.570 167.340 62.690 ;
        RECT 169.760 62.590 170.370 62.690 ;
        RECT 173.615 62.895 173.915 63.045 ;
        RECT 173.615 62.595 175.255 62.895 ;
        RECT 174.955 62.115 175.255 62.595 ;
        RECT 174.075 61.755 176.135 62.115 ;
        RECT 158.855 61.385 163.330 61.465 ;
        RECT 158.855 60.815 159.085 61.385 ;
        RECT 159.965 61.305 160.225 61.385 ;
        RECT 161.005 61.235 161.825 61.385 ;
        RECT 162.510 61.235 163.330 61.385 ;
        RECT 164.335 61.235 165.155 61.465 ;
        RECT 160.460 60.905 160.740 61.205 ;
        RECT 156.225 60.565 156.525 60.585 ;
        RECT 156.225 60.305 156.565 60.565 ;
        RECT 158.525 60.545 158.825 60.600 ;
        RECT 159.345 60.545 159.665 60.615 ;
        RECT 160.525 60.545 160.675 60.905 ;
        RECT 158.515 60.385 160.685 60.545 ;
        RECT 174.075 60.390 174.305 61.755 ;
        RECT 174.755 60.390 175.455 60.420 ;
        RECT 156.225 60.285 156.525 60.305 ;
        RECT 158.525 60.300 158.825 60.385 ;
        RECT 159.345 60.355 159.665 60.385 ;
        RECT 160.525 60.375 160.675 60.385 ;
        RECT 174.075 60.160 175.455 60.390 ;
        RECT 174.755 60.120 175.455 60.160 ;
        RECT 173.065 60.035 173.765 60.105 ;
        RECT 176.490 60.035 177.190 60.105 ;
        RECT 156.225 60.000 156.525 60.005 ;
        RECT 156.205 59.700 156.565 60.000 ;
        RECT 158.525 59.935 158.825 60.020 ;
        RECT 159.935 59.935 160.255 59.985 ;
        RECT 158.525 59.775 160.685 59.935 ;
        RECT 172.915 59.805 173.915 60.035 ;
        RECT 176.340 59.805 177.340 60.035 ;
        RECT 158.525 59.720 158.825 59.775 ;
        RECT 159.935 59.725 160.255 59.775 ;
        RECT 155.965 59.125 156.195 59.405 ;
        RECT 154.265 58.945 156.195 59.125 ;
        RECT 154.265 58.645 154.495 58.945 ;
        RECT 155.965 58.755 156.195 58.945 ;
        RECT 156.555 59.130 156.785 59.490 ;
        RECT 158.265 59.130 158.495 59.420 ;
        RECT 156.555 58.940 158.495 59.130 ;
        RECT 156.555 58.670 156.785 58.940 ;
        RECT 148.765 57.290 149.375 57.390 ;
        RECT 151.795 57.290 152.405 57.370 ;
        RECT 154.805 57.290 155.415 57.400 ;
        RECT 157.480 57.290 157.625 58.940 ;
        RECT 158.265 58.770 158.495 58.940 ;
        RECT 158.855 58.885 159.085 59.505 ;
        RECT 160.515 59.410 160.685 59.775 ;
        RECT 160.460 59.110 160.740 59.410 ;
        RECT 160.515 59.095 160.685 59.110 ;
        RECT 159.345 58.885 159.665 58.935 ;
        RECT 161.005 58.885 161.825 59.080 ;
        RECT 162.510 58.885 163.330 59.080 ;
        RECT 158.855 58.850 163.330 58.885 ;
        RECT 164.335 58.850 165.155 59.080 ;
        RECT 158.855 58.725 162.745 58.850 ;
        RECT 158.855 58.685 159.085 58.725 ;
        RECT 159.345 58.675 159.665 58.725 ;
        RECT 162.195 57.850 162.355 58.725 ;
        RECT 162.145 57.530 162.405 57.850 ;
        RECT 157.835 57.290 158.445 57.380 ;
        RECT 160.805 57.290 161.415 57.400 ;
        RECT 163.835 57.290 164.445 57.380 ;
        RECT 164.825 57.290 164.970 58.850 ;
        RECT 174.075 58.155 174.305 58.185 ;
        RECT 174.075 57.855 175.255 58.155 ;
        RECT 174.075 57.825 174.305 57.855 ;
        RECT 166.845 57.290 167.455 57.410 ;
        RECT 169.875 57.290 170.485 57.390 ;
        RECT 148.765 57.260 170.485 57.290 ;
        RECT 174.955 57.280 175.255 57.855 ;
        RECT 148.090 57.145 170.485 57.260 ;
        RECT 148.090 57.115 150.490 57.145 ;
        RECT 74.460 55.720 74.905 55.800 ;
        RECT 74.455 55.275 74.960 55.720 ;
        RECT 78.610 55.325 79.050 55.705 ;
        RECT 120.725 50.580 143.430 50.895 ;
        RECT 143.105 50.570 143.365 50.580 ;
        RECT 128.580 47.995 129.000 48.025 ;
        RECT 128.580 47.575 143.560 47.995 ;
        RECT 128.580 47.545 129.000 47.575 ;
        RECT 12.445 46.480 12.705 46.540 ;
        RECT 12.445 46.470 13.360 46.480 ;
        RECT 17.095 46.470 17.355 46.520 ;
        RECT 22.060 46.480 22.320 46.540 ;
        RECT 22.060 46.470 22.975 46.480 ;
        RECT 26.710 46.470 26.970 46.520 ;
        RECT 31.675 46.480 31.935 46.540 ;
        RECT 31.675 46.470 32.590 46.480 ;
        RECT 36.325 46.470 36.585 46.520 ;
        RECT 41.290 46.480 41.550 46.540 ;
        RECT 41.290 46.470 42.205 46.480 ;
        RECT 45.940 46.470 46.200 46.520 ;
        RECT 12.430 46.455 13.360 46.470 ;
        RECT 13.610 46.455 13.900 46.470 ;
        RECT 14.200 46.455 14.490 46.470 ;
        RECT 14.790 46.455 15.080 46.470 ;
        RECT 15.380 46.455 15.670 46.470 ;
        RECT 15.970 46.455 16.260 46.470 ;
        RECT 16.560 46.455 16.850 46.470 ;
        RECT 17.095 46.455 17.440 46.470 ;
        RECT 17.740 46.455 18.030 46.470 ;
        RECT 12.430 46.260 18.030 46.455 ;
        RECT 12.430 46.240 12.720 46.260 ;
        RECT 13.020 46.240 13.310 46.260 ;
        RECT 13.610 46.240 13.900 46.260 ;
        RECT 14.200 46.240 14.490 46.260 ;
        RECT 14.790 46.240 15.080 46.260 ;
        RECT 15.380 46.240 15.670 46.260 ;
        RECT 15.970 46.240 16.260 46.260 ;
        RECT 16.560 46.240 16.850 46.260 ;
        RECT 17.095 46.240 17.440 46.260 ;
        RECT 17.740 46.240 18.030 46.260 ;
        RECT 22.045 46.455 22.975 46.470 ;
        RECT 23.225 46.455 23.515 46.470 ;
        RECT 23.815 46.455 24.105 46.470 ;
        RECT 24.405 46.455 24.695 46.470 ;
        RECT 24.995 46.455 25.285 46.470 ;
        RECT 25.585 46.455 25.875 46.470 ;
        RECT 26.175 46.455 26.465 46.470 ;
        RECT 26.710 46.455 27.055 46.470 ;
        RECT 27.355 46.455 27.645 46.470 ;
        RECT 22.045 46.260 27.645 46.455 ;
        RECT 22.045 46.240 22.335 46.260 ;
        RECT 22.635 46.240 22.925 46.260 ;
        RECT 23.225 46.240 23.515 46.260 ;
        RECT 23.815 46.240 24.105 46.260 ;
        RECT 24.405 46.240 24.695 46.260 ;
        RECT 24.995 46.240 25.285 46.260 ;
        RECT 25.585 46.240 25.875 46.260 ;
        RECT 26.175 46.240 26.465 46.260 ;
        RECT 26.710 46.240 27.055 46.260 ;
        RECT 27.355 46.240 27.645 46.260 ;
        RECT 31.660 46.455 32.590 46.470 ;
        RECT 32.840 46.455 33.130 46.470 ;
        RECT 33.430 46.455 33.720 46.470 ;
        RECT 34.020 46.455 34.310 46.470 ;
        RECT 34.610 46.455 34.900 46.470 ;
        RECT 35.200 46.455 35.490 46.470 ;
        RECT 35.790 46.455 36.080 46.470 ;
        RECT 36.325 46.455 36.670 46.470 ;
        RECT 36.970 46.455 37.260 46.470 ;
        RECT 31.660 46.260 37.260 46.455 ;
        RECT 31.660 46.240 31.950 46.260 ;
        RECT 32.250 46.240 32.540 46.260 ;
        RECT 32.840 46.240 33.130 46.260 ;
        RECT 33.430 46.240 33.720 46.260 ;
        RECT 34.020 46.240 34.310 46.260 ;
        RECT 34.610 46.240 34.900 46.260 ;
        RECT 35.200 46.240 35.490 46.260 ;
        RECT 35.790 46.240 36.080 46.260 ;
        RECT 36.325 46.240 36.670 46.260 ;
        RECT 36.970 46.240 37.260 46.260 ;
        RECT 41.275 46.455 42.205 46.470 ;
        RECT 42.455 46.455 42.745 46.470 ;
        RECT 43.045 46.455 43.335 46.470 ;
        RECT 43.635 46.455 43.925 46.470 ;
        RECT 44.225 46.455 44.515 46.470 ;
        RECT 44.815 46.455 45.105 46.470 ;
        RECT 45.405 46.455 45.695 46.470 ;
        RECT 45.940 46.455 46.285 46.470 ;
        RECT 46.585 46.455 46.875 46.470 ;
        RECT 41.275 46.260 46.875 46.455 ;
        RECT 41.275 46.240 41.565 46.260 ;
        RECT 41.865 46.240 42.155 46.260 ;
        RECT 42.455 46.240 42.745 46.260 ;
        RECT 43.045 46.240 43.335 46.260 ;
        RECT 43.635 46.240 43.925 46.260 ;
        RECT 44.225 46.240 44.515 46.260 ;
        RECT 44.815 46.240 45.105 46.260 ;
        RECT 45.405 46.240 45.695 46.260 ;
        RECT 45.940 46.240 46.285 46.260 ;
        RECT 46.585 46.240 46.875 46.260 ;
        RECT 12.445 46.220 12.705 46.240 ;
        RECT 17.095 46.200 17.355 46.240 ;
        RECT 22.060 46.220 22.320 46.240 ;
        RECT 26.710 46.200 26.970 46.240 ;
        RECT 31.675 46.220 31.935 46.240 ;
        RECT 36.325 46.200 36.585 46.240 ;
        RECT 41.290 46.220 41.550 46.240 ;
        RECT 45.940 46.200 46.200 46.240 ;
        RECT 12.755 45.370 12.985 45.860 ;
        RECT 13.935 45.410 14.165 45.860 ;
        RECT 13.915 45.380 14.175 45.410 ;
        RECT 15.115 45.380 15.345 45.860 ;
        RECT 16.295 45.380 16.525 45.860 ;
        RECT 17.475 45.380 17.705 45.860 ;
        RECT 12.720 45.110 13.040 45.370 ;
        RECT 13.885 45.120 14.205 45.380 ;
        RECT 15.065 45.120 15.385 45.380 ;
        RECT 16.255 45.120 16.575 45.380 ;
        RECT 17.425 45.120 17.745 45.380 ;
        RECT 22.370 45.370 22.600 45.860 ;
        RECT 23.550 45.410 23.780 45.860 ;
        RECT 23.530 45.380 23.790 45.410 ;
        RECT 24.730 45.380 24.960 45.860 ;
        RECT 25.910 45.380 26.140 45.860 ;
        RECT 27.090 45.380 27.320 45.860 ;
        RECT 13.915 45.090 14.175 45.120 ;
        RECT 22.335 45.110 22.655 45.370 ;
        RECT 23.500 45.120 23.820 45.380 ;
        RECT 24.680 45.120 25.000 45.380 ;
        RECT 25.870 45.120 26.190 45.380 ;
        RECT 27.040 45.120 27.360 45.380 ;
        RECT 31.985 45.370 32.215 45.860 ;
        RECT 33.165 45.410 33.395 45.860 ;
        RECT 33.145 45.380 33.405 45.410 ;
        RECT 34.345 45.380 34.575 45.860 ;
        RECT 35.525 45.380 35.755 45.860 ;
        RECT 36.705 45.380 36.935 45.860 ;
        RECT 23.530 45.090 23.790 45.120 ;
        RECT 31.950 45.110 32.270 45.370 ;
        RECT 33.115 45.120 33.435 45.380 ;
        RECT 34.295 45.120 34.615 45.380 ;
        RECT 35.485 45.120 35.805 45.380 ;
        RECT 36.655 45.120 36.975 45.380 ;
        RECT 41.600 45.370 41.830 45.860 ;
        RECT 42.780 45.410 43.010 45.860 ;
        RECT 42.760 45.380 43.020 45.410 ;
        RECT 43.960 45.380 44.190 45.860 ;
        RECT 45.140 45.380 45.370 45.860 ;
        RECT 46.320 45.380 46.550 45.860 ;
        RECT 148.090 45.625 148.235 57.115 ;
        RECT 148.765 56.840 149.375 57.115 ;
        RECT 151.795 56.820 152.405 57.145 ;
        RECT 154.805 56.850 155.415 57.145 ;
        RECT 157.835 56.830 158.445 57.145 ;
        RECT 160.805 56.850 161.415 57.145 ;
        RECT 163.835 56.830 164.445 57.145 ;
        RECT 166.845 56.860 167.455 57.145 ;
        RECT 169.875 56.840 170.485 57.145 ;
        RECT 174.755 56.980 175.455 57.280 ;
        RECT 173.065 56.895 173.765 56.965 ;
        RECT 176.490 56.895 177.190 56.965 ;
        RECT 172.915 56.665 173.915 56.895 ;
        RECT 176.340 56.665 177.340 56.895 ;
        RECT 174.075 56.255 176.135 56.615 ;
        RECT 174.955 55.490 175.255 56.255 ;
        RECT 174.945 55.230 175.265 55.490 ;
        RECT 148.780 53.280 149.375 53.475 ;
        RECT 151.810 53.280 152.405 53.455 ;
        RECT 154.820 53.280 155.415 53.485 ;
        RECT 157.850 53.280 158.445 53.465 ;
        RECT 160.820 53.280 161.415 53.485 ;
        RECT 163.850 53.280 164.445 53.465 ;
        RECT 166.860 53.280 167.455 53.495 ;
        RECT 169.890 53.280 170.485 53.475 ;
        RECT 148.780 53.135 170.495 53.280 ;
        RECT 148.780 52.940 149.375 53.135 ;
        RECT 150.720 52.320 150.865 53.135 ;
        RECT 151.810 52.920 152.405 53.135 ;
        RECT 154.820 52.950 155.415 53.135 ;
        RECT 157.850 52.930 158.445 53.135 ;
        RECT 160.820 52.950 161.415 53.135 ;
        RECT 163.850 52.930 164.445 53.135 ;
        RECT 166.860 52.960 167.455 53.135 ;
        RECT 169.890 52.940 170.485 53.135 ;
        RECT 154.265 52.320 155.575 52.325 ;
        RECT 150.720 52.180 155.575 52.320 ;
        RECT 159.885 52.295 161.220 52.305 ;
        RECT 150.720 52.175 154.410 52.180 ;
        RECT 150.720 51.935 150.865 52.175 ;
        RECT 151.895 51.935 152.040 52.175 ;
        RECT 153.065 51.935 153.210 52.175 ;
        RECT 154.265 51.935 154.410 52.175 ;
        RECT 155.430 51.935 155.575 52.180 ;
        RECT 157.370 52.160 161.220 52.295 ;
        RECT 157.370 52.150 160.030 52.160 ;
        RECT 150.675 51.115 150.905 51.935 ;
        RECT 151.855 51.115 152.085 51.935 ;
        RECT 153.035 51.115 153.265 51.935 ;
        RECT 154.215 51.115 154.445 51.935 ;
        RECT 155.395 51.115 155.625 51.935 ;
        RECT 148.745 49.590 149.340 49.695 ;
        RECT 151.775 49.590 152.370 49.715 ;
        RECT 154.785 49.590 155.380 49.685 ;
        RECT 157.370 49.590 157.515 52.150 ;
        RECT 158.695 51.980 158.840 52.150 ;
        RECT 159.885 51.980 160.030 52.150 ;
        RECT 161.075 51.980 161.220 52.160 ;
        RECT 163.625 52.140 164.945 52.295 ;
        RECT 158.665 51.070 158.895 51.980 ;
        RECT 159.845 51.070 160.075 51.980 ;
        RECT 161.025 51.070 161.255 51.980 ;
        RECT 163.625 51.935 163.780 52.140 ;
        RECT 164.790 51.935 164.945 52.140 ;
        RECT 163.570 51.255 163.800 51.935 ;
        RECT 163.330 51.115 163.800 51.255 ;
        RECT 164.750 51.115 164.980 51.935 ;
        RECT 163.330 51.100 163.780 51.115 ;
        RECT 157.815 49.590 158.410 49.705 ;
        RECT 148.745 49.445 158.410 49.590 ;
        RECT 148.745 49.160 149.340 49.445 ;
        RECT 151.775 49.180 152.370 49.445 ;
        RECT 154.785 49.150 155.380 49.445 ;
        RECT 157.815 49.170 158.410 49.445 ;
        RECT 160.785 49.620 161.380 49.685 ;
        RECT 163.330 49.620 163.485 51.100 ;
        RECT 166.800 50.895 167.620 51.125 ;
        RECT 163.825 49.620 164.420 49.680 ;
        RECT 167.045 49.675 167.200 50.895 ;
        RECT 169.595 50.830 170.415 51.060 ;
        RECT 170.070 49.695 170.225 50.830 ;
        RECT 160.785 49.465 164.420 49.620 ;
        RECT 160.785 49.150 161.380 49.465 ;
        RECT 163.825 49.145 164.420 49.465 ;
        RECT 166.825 49.140 167.420 49.675 ;
        RECT 169.855 49.160 170.450 49.695 ;
        RECT 148.730 45.625 149.340 45.795 ;
        RECT 151.760 45.625 152.370 45.815 ;
        RECT 154.770 45.625 155.380 45.785 ;
        RECT 157.800 45.625 158.410 45.805 ;
        RECT 160.770 45.625 161.380 45.785 ;
        RECT 163.810 45.625 164.420 45.780 ;
        RECT 166.810 45.625 167.420 45.775 ;
        RECT 169.840 45.625 170.450 45.795 ;
        RECT 148.090 45.480 170.450 45.625 ;
        RECT 33.145 45.090 33.405 45.120 ;
        RECT 41.565 45.110 41.885 45.370 ;
        RECT 42.730 45.120 43.050 45.380 ;
        RECT 43.910 45.120 44.230 45.380 ;
        RECT 45.100 45.120 45.420 45.380 ;
        RECT 46.270 45.120 46.590 45.380 ;
        RECT 148.730 45.245 149.340 45.480 ;
        RECT 151.760 45.265 152.370 45.480 ;
        RECT 154.770 45.235 155.380 45.480 ;
        RECT 157.800 45.255 158.410 45.480 ;
        RECT 160.770 45.235 161.380 45.480 ;
        RECT 163.810 45.230 164.420 45.480 ;
        RECT 166.810 45.225 167.420 45.480 ;
        RECT 169.840 45.245 170.450 45.480 ;
        RECT 42.760 45.090 43.020 45.120 ;
        RECT 132.675 44.900 133.095 44.930 ;
        RECT 132.675 44.480 143.490 44.900 ;
        RECT 132.675 44.450 133.095 44.480 ;
        RECT 12.745 43.350 12.975 43.375 ;
        RECT 12.720 43.090 13.040 43.350 ;
        RECT 13.925 43.270 14.155 43.375 ;
        RECT 15.105 43.280 15.335 43.375 ;
        RECT 12.745 42.725 12.975 43.090 ;
        RECT 13.885 43.010 14.205 43.270 ;
        RECT 15.095 43.250 15.355 43.280 ;
        RECT 13.925 42.725 14.155 43.010 ;
        RECT 15.065 42.990 15.385 43.250 ;
        RECT 16.285 43.190 16.515 43.375 ;
        RECT 17.465 43.210 17.695 43.375 ;
        RECT 22.360 43.350 22.590 43.375 ;
        RECT 15.095 42.960 15.355 42.990 ;
        RECT 15.105 42.725 15.335 42.960 ;
        RECT 16.255 42.930 16.575 43.190 ;
        RECT 17.425 42.950 17.745 43.210 ;
        RECT 22.335 43.090 22.655 43.350 ;
        RECT 23.540 43.270 23.770 43.375 ;
        RECT 24.720 43.280 24.950 43.375 ;
        RECT 16.285 42.725 16.515 42.930 ;
        RECT 17.465 42.725 17.695 42.950 ;
        RECT 22.360 42.725 22.590 43.090 ;
        RECT 23.500 43.010 23.820 43.270 ;
        RECT 24.710 43.250 24.970 43.280 ;
        RECT 23.540 42.725 23.770 43.010 ;
        RECT 24.680 42.990 25.000 43.250 ;
        RECT 25.900 43.190 26.130 43.375 ;
        RECT 27.080 43.210 27.310 43.375 ;
        RECT 31.975 43.350 32.205 43.375 ;
        RECT 24.710 42.960 24.970 42.990 ;
        RECT 24.720 42.725 24.950 42.960 ;
        RECT 25.870 42.930 26.190 43.190 ;
        RECT 27.040 42.950 27.360 43.210 ;
        RECT 31.950 43.090 32.270 43.350 ;
        RECT 33.155 43.270 33.385 43.375 ;
        RECT 34.335 43.280 34.565 43.375 ;
        RECT 25.900 42.725 26.130 42.930 ;
        RECT 27.080 42.725 27.310 42.950 ;
        RECT 31.975 42.725 32.205 43.090 ;
        RECT 33.115 43.010 33.435 43.270 ;
        RECT 34.325 43.250 34.585 43.280 ;
        RECT 33.155 42.725 33.385 43.010 ;
        RECT 34.295 42.990 34.615 43.250 ;
        RECT 35.515 43.190 35.745 43.375 ;
        RECT 36.695 43.210 36.925 43.375 ;
        RECT 41.590 43.350 41.820 43.375 ;
        RECT 34.325 42.960 34.585 42.990 ;
        RECT 34.335 42.725 34.565 42.960 ;
        RECT 35.485 42.930 35.805 43.190 ;
        RECT 36.655 42.950 36.975 43.210 ;
        RECT 41.565 43.090 41.885 43.350 ;
        RECT 42.770 43.270 43.000 43.375 ;
        RECT 43.950 43.280 44.180 43.375 ;
        RECT 35.515 42.725 35.745 42.930 ;
        RECT 36.695 42.725 36.925 42.950 ;
        RECT 41.590 42.725 41.820 43.090 ;
        RECT 42.730 43.010 43.050 43.270 ;
        RECT 43.940 43.250 44.200 43.280 ;
        RECT 42.770 42.725 43.000 43.010 ;
        RECT 43.910 42.990 44.230 43.250 ;
        RECT 45.130 43.190 45.360 43.375 ;
        RECT 46.310 43.210 46.540 43.375 ;
        RECT 43.940 42.960 44.200 42.990 ;
        RECT 43.950 42.725 44.180 42.960 ;
        RECT 45.100 42.930 45.420 43.190 ;
        RECT 46.270 42.950 46.590 43.210 ;
        RECT 45.130 42.725 45.360 42.930 ;
        RECT 46.310 42.725 46.540 42.950 ;
        RECT 148.760 42.825 149.020 43.145 ;
        RECT 17.990 42.390 18.310 42.400 ;
        RECT 27.605 42.390 27.925 42.400 ;
        RECT 37.220 42.390 37.540 42.400 ;
        RECT 46.835 42.390 47.155 42.400 ;
        RECT 12.420 42.365 12.710 42.390 ;
        RECT 13.010 42.365 13.300 42.390 ;
        RECT 13.600 42.365 13.890 42.390 ;
        RECT 14.190 42.365 14.480 42.390 ;
        RECT 14.780 42.365 15.070 42.390 ;
        RECT 15.370 42.365 15.660 42.390 ;
        RECT 15.960 42.365 16.250 42.390 ;
        RECT 16.550 42.365 16.840 42.390 ;
        RECT 17.140 42.365 17.430 42.390 ;
        RECT 17.730 42.365 18.310 42.390 ;
        RECT 12.420 42.170 18.310 42.365 ;
        RECT 12.420 42.160 12.710 42.170 ;
        RECT 13.010 42.160 13.300 42.170 ;
        RECT 13.600 42.160 13.890 42.170 ;
        RECT 14.190 42.160 14.480 42.170 ;
        RECT 14.780 42.160 15.070 42.170 ;
        RECT 15.370 42.160 15.660 42.170 ;
        RECT 15.960 42.160 16.250 42.170 ;
        RECT 16.550 42.160 16.840 42.170 ;
        RECT 17.140 42.160 17.430 42.170 ;
        RECT 17.730 42.160 18.310 42.170 ;
        RECT 22.035 42.365 22.325 42.390 ;
        RECT 22.625 42.365 22.915 42.390 ;
        RECT 23.215 42.365 23.505 42.390 ;
        RECT 23.805 42.365 24.095 42.390 ;
        RECT 24.395 42.365 24.685 42.390 ;
        RECT 24.985 42.365 25.275 42.390 ;
        RECT 25.575 42.365 25.865 42.390 ;
        RECT 26.165 42.365 26.455 42.390 ;
        RECT 26.755 42.365 27.045 42.390 ;
        RECT 27.345 42.365 27.925 42.390 ;
        RECT 22.035 42.170 27.925 42.365 ;
        RECT 22.035 42.160 22.325 42.170 ;
        RECT 22.625 42.160 22.915 42.170 ;
        RECT 23.215 42.160 23.505 42.170 ;
        RECT 23.805 42.160 24.095 42.170 ;
        RECT 24.395 42.160 24.685 42.170 ;
        RECT 24.985 42.160 25.275 42.170 ;
        RECT 25.575 42.160 25.865 42.170 ;
        RECT 26.165 42.160 26.455 42.170 ;
        RECT 26.755 42.160 27.045 42.170 ;
        RECT 27.345 42.160 27.925 42.170 ;
        RECT 31.650 42.365 31.940 42.390 ;
        RECT 32.240 42.365 32.530 42.390 ;
        RECT 32.830 42.365 33.120 42.390 ;
        RECT 33.420 42.365 33.710 42.390 ;
        RECT 34.010 42.365 34.300 42.390 ;
        RECT 34.600 42.365 34.890 42.390 ;
        RECT 35.190 42.365 35.480 42.390 ;
        RECT 35.780 42.365 36.070 42.390 ;
        RECT 36.370 42.365 36.660 42.390 ;
        RECT 36.960 42.365 37.540 42.390 ;
        RECT 31.650 42.170 37.540 42.365 ;
        RECT 31.650 42.160 31.940 42.170 ;
        RECT 32.240 42.160 32.530 42.170 ;
        RECT 32.830 42.160 33.120 42.170 ;
        RECT 33.420 42.160 33.710 42.170 ;
        RECT 34.010 42.160 34.300 42.170 ;
        RECT 34.600 42.160 34.890 42.170 ;
        RECT 35.190 42.160 35.480 42.170 ;
        RECT 35.780 42.160 36.070 42.170 ;
        RECT 36.370 42.160 36.660 42.170 ;
        RECT 36.960 42.160 37.540 42.170 ;
        RECT 41.265 42.365 41.555 42.390 ;
        RECT 41.855 42.365 42.145 42.390 ;
        RECT 42.445 42.365 42.735 42.390 ;
        RECT 43.035 42.365 43.325 42.390 ;
        RECT 43.625 42.365 43.915 42.390 ;
        RECT 44.215 42.365 44.505 42.390 ;
        RECT 44.805 42.365 45.095 42.390 ;
        RECT 45.395 42.365 45.685 42.390 ;
        RECT 45.985 42.365 46.275 42.390 ;
        RECT 46.575 42.365 47.155 42.390 ;
        RECT 41.265 42.170 47.155 42.365 ;
        RECT 41.265 42.160 41.555 42.170 ;
        RECT 41.855 42.160 42.145 42.170 ;
        RECT 42.445 42.160 42.735 42.170 ;
        RECT 43.035 42.160 43.325 42.170 ;
        RECT 43.625 42.160 43.915 42.170 ;
        RECT 44.215 42.160 44.505 42.170 ;
        RECT 44.805 42.160 45.095 42.170 ;
        RECT 45.395 42.160 45.685 42.170 ;
        RECT 45.985 42.160 46.275 42.170 ;
        RECT 46.575 42.160 47.155 42.170 ;
        RECT 17.990 42.140 18.310 42.160 ;
        RECT 27.605 42.140 27.925 42.160 ;
        RECT 37.220 42.140 37.540 42.160 ;
        RECT 46.835 42.140 47.155 42.160 ;
        RECT 148.770 41.455 149.030 41.775 ;
        RECT 148.790 40.060 149.050 40.380 ;
        RECT 16.320 39.490 16.640 39.750 ;
        RECT 25.935 39.490 26.255 39.750 ;
        RECT 35.550 39.490 35.870 39.750 ;
        RECT 45.165 39.490 45.485 39.750 ;
        RECT 17.265 39.115 17.525 39.435 ;
        RECT 18.575 39.135 18.895 39.395 ;
        RECT 26.880 39.115 27.140 39.435 ;
        RECT 28.190 39.135 28.510 39.395 ;
        RECT 36.495 39.115 36.755 39.435 ;
        RECT 37.805 39.135 38.125 39.395 ;
        RECT 46.110 39.115 46.370 39.435 ;
        RECT 47.420 39.135 47.740 39.395 ;
        RECT 148.790 38.705 149.050 39.025 ;
        RECT 148.765 37.315 149.025 37.635 ;
        RECT 148.760 35.945 149.020 36.265 ;
        RECT 148.795 34.555 149.055 34.875 ;
        RECT 148.780 33.205 149.040 33.525 ;
        RECT 148.790 31.820 149.050 32.140 ;
      LAYER via ;
        RECT 148.790 87.740 149.050 88.000 ;
        RECT 148.780 86.355 149.040 86.615 ;
        RECT 148.795 85.005 149.055 85.265 ;
        RECT 148.760 83.615 149.020 83.875 ;
        RECT 148.765 82.245 149.025 82.505 ;
        RECT 148.790 80.855 149.050 81.115 ;
        RECT 17.265 80.445 17.525 80.705 ;
        RECT 18.605 80.455 18.865 80.715 ;
        RECT 26.880 80.445 27.140 80.705 ;
        RECT 28.220 80.455 28.480 80.715 ;
        RECT 36.495 80.445 36.755 80.705 ;
        RECT 37.835 80.455 38.095 80.715 ;
        RECT 46.110 80.445 46.370 80.705 ;
        RECT 47.450 80.455 47.710 80.715 ;
        RECT 16.350 80.100 16.610 80.360 ;
        RECT 25.965 80.100 26.225 80.360 ;
        RECT 35.580 80.100 35.840 80.360 ;
        RECT 45.195 80.100 45.455 80.360 ;
        RECT 148.790 79.500 149.050 79.760 ;
        RECT 148.770 78.105 149.030 78.365 ;
        RECT 18.020 77.450 18.280 77.710 ;
        RECT 27.635 77.450 27.895 77.710 ;
        RECT 37.250 77.450 37.510 77.710 ;
        RECT 46.865 77.450 47.125 77.710 ;
        RECT 12.750 76.500 13.010 76.760 ;
        RECT 13.915 76.580 14.175 76.840 ;
        RECT 15.095 76.600 15.355 76.860 ;
        RECT 16.285 76.660 16.545 76.920 ;
        RECT 17.455 76.640 17.715 76.900 ;
        RECT 22.365 76.500 22.625 76.760 ;
        RECT 23.530 76.580 23.790 76.840 ;
        RECT 24.710 76.600 24.970 76.860 ;
        RECT 25.900 76.660 26.160 76.920 ;
        RECT 27.070 76.640 27.330 76.900 ;
        RECT 31.980 76.500 32.240 76.760 ;
        RECT 33.145 76.580 33.405 76.840 ;
        RECT 34.325 76.600 34.585 76.860 ;
        RECT 35.515 76.660 35.775 76.920 ;
        RECT 36.685 76.640 36.945 76.900 ;
        RECT 41.595 76.500 41.855 76.760 ;
        RECT 42.760 76.580 43.020 76.840 ;
        RECT 43.940 76.600 44.200 76.860 ;
        RECT 45.130 76.660 45.390 76.920 ;
        RECT 46.300 76.640 46.560 76.900 ;
        RECT 148.760 76.735 149.020 76.995 ;
        RECT 143.065 75.040 143.325 75.300 ;
        RECT 12.750 74.480 13.010 74.740 ;
        RECT 13.915 74.470 14.175 74.730 ;
        RECT 15.095 74.470 15.355 74.730 ;
        RECT 16.285 74.470 16.545 74.730 ;
        RECT 17.455 74.470 17.715 74.730 ;
        RECT 22.365 74.480 22.625 74.740 ;
        RECT 23.530 74.470 23.790 74.730 ;
        RECT 24.710 74.470 24.970 74.730 ;
        RECT 25.900 74.470 26.160 74.730 ;
        RECT 27.070 74.470 27.330 74.730 ;
        RECT 31.980 74.480 32.240 74.740 ;
        RECT 33.145 74.470 33.405 74.730 ;
        RECT 34.325 74.470 34.585 74.730 ;
        RECT 35.515 74.470 35.775 74.730 ;
        RECT 36.685 74.470 36.945 74.730 ;
        RECT 41.595 74.480 41.855 74.740 ;
        RECT 42.760 74.470 43.020 74.730 ;
        RECT 43.940 74.470 44.200 74.730 ;
        RECT 45.130 74.470 45.390 74.730 ;
        RECT 46.300 74.470 46.560 74.730 ;
        RECT 12.445 73.340 12.705 73.600 ;
        RECT 17.095 73.360 17.355 73.620 ;
        RECT 22.060 73.340 22.320 73.600 ;
        RECT 26.710 73.360 26.970 73.620 ;
        RECT 31.675 73.340 31.935 73.600 ;
        RECT 36.325 73.360 36.585 73.620 ;
        RECT 41.290 73.340 41.550 73.600 ;
        RECT 45.940 73.360 46.200 73.620 ;
        RECT 143.150 71.970 143.410 72.230 ;
        RECT 122.535 68.955 122.850 69.270 ;
        RECT 143.105 68.990 143.365 69.250 ;
        RECT 74.485 64.130 74.930 64.575 ;
        RECT 78.640 64.145 79.020 64.525 ;
        RECT 148.645 74.185 149.195 74.735 ;
        RECT 151.675 74.165 152.225 74.715 ;
        RECT 154.685 74.195 155.235 74.745 ;
        RECT 157.715 74.175 158.265 74.725 ;
        RECT 160.685 74.195 161.235 74.745 ;
        RECT 163.725 74.200 164.275 74.750 ;
        RECT 166.725 74.205 167.275 74.755 ;
        RECT 169.755 74.185 170.305 74.735 ;
        RECT 148.660 70.285 149.195 70.820 ;
        RECT 151.690 70.265 152.225 70.800 ;
        RECT 154.700 70.295 155.235 70.830 ;
        RECT 157.730 70.275 158.265 70.810 ;
        RECT 160.700 70.295 161.235 70.830 ;
        RECT 163.740 70.300 164.275 70.835 ;
        RECT 166.740 70.305 167.275 70.840 ;
        RECT 169.770 70.285 170.305 70.820 ;
        RECT 148.695 66.505 149.230 67.040 ;
        RECT 170.095 67.380 170.355 67.640 ;
        RECT 151.725 66.525 152.260 67.060 ;
        RECT 154.735 66.495 155.270 67.030 ;
        RECT 157.765 66.515 158.300 67.050 ;
        RECT 160.735 66.495 161.270 67.030 ;
        RECT 163.765 66.515 164.300 67.050 ;
        RECT 166.775 66.485 167.310 67.020 ;
        RECT 169.805 66.505 170.340 67.040 ;
        RECT 173.125 64.565 173.385 64.825 ;
        RECT 173.445 64.565 173.705 64.825 ;
        RECT 176.550 64.565 176.810 64.825 ;
        RECT 176.870 64.565 177.130 64.825 ;
        RECT 174.815 64.250 175.075 64.510 ;
        RECT 175.135 64.250 175.395 64.510 ;
        RECT 148.680 62.590 149.230 63.140 ;
        RECT 151.710 62.610 152.260 63.160 ;
        RECT 154.720 62.580 155.270 63.130 ;
        RECT 157.750 62.600 158.300 63.150 ;
        RECT 160.720 62.580 161.270 63.130 ;
        RECT 163.750 62.600 164.300 63.150 ;
        RECT 162.235 62.200 162.495 62.460 ;
        RECT 159.965 61.335 160.225 61.595 ;
        RECT 166.760 62.570 167.310 63.120 ;
        RECT 169.790 62.590 170.340 63.140 ;
        RECT 156.275 60.305 156.535 60.565 ;
        RECT 159.375 60.355 159.635 60.615 ;
        RECT 174.815 60.140 175.075 60.400 ;
        RECT 175.135 60.140 175.395 60.400 ;
        RECT 156.235 59.700 156.535 60.000 ;
        RECT 159.965 59.725 160.225 59.985 ;
        RECT 173.125 59.825 173.385 60.085 ;
        RECT 173.445 59.825 173.705 60.085 ;
        RECT 176.550 59.825 176.810 60.085 ;
        RECT 176.870 59.825 177.130 60.085 ;
        RECT 74.485 55.275 74.930 55.720 ;
        RECT 78.640 55.325 79.020 55.705 ;
        RECT 122.535 50.580 122.850 50.895 ;
        RECT 143.105 50.600 143.365 50.860 ;
        RECT 143.150 47.620 143.410 47.880 ;
        RECT 12.445 46.250 12.705 46.510 ;
        RECT 17.095 46.230 17.355 46.490 ;
        RECT 22.060 46.250 22.320 46.510 ;
        RECT 26.710 46.230 26.970 46.490 ;
        RECT 31.675 46.250 31.935 46.510 ;
        RECT 36.325 46.230 36.585 46.490 ;
        RECT 41.290 46.250 41.550 46.510 ;
        RECT 45.940 46.230 46.200 46.490 ;
        RECT 12.750 45.110 13.010 45.370 ;
        RECT 13.915 45.120 14.175 45.380 ;
        RECT 15.095 45.120 15.355 45.380 ;
        RECT 16.285 45.120 16.545 45.380 ;
        RECT 17.455 45.120 17.715 45.380 ;
        RECT 22.365 45.110 22.625 45.370 ;
        RECT 23.530 45.120 23.790 45.380 ;
        RECT 24.710 45.120 24.970 45.380 ;
        RECT 25.900 45.120 26.160 45.380 ;
        RECT 27.070 45.120 27.330 45.380 ;
        RECT 31.980 45.110 32.240 45.370 ;
        RECT 33.145 45.120 33.405 45.380 ;
        RECT 34.325 45.120 34.585 45.380 ;
        RECT 35.515 45.120 35.775 45.380 ;
        RECT 36.685 45.120 36.945 45.380 ;
        RECT 148.795 56.840 149.345 57.390 ;
        RECT 151.825 56.820 152.375 57.370 ;
        RECT 154.835 56.850 155.385 57.400 ;
        RECT 159.375 58.675 159.635 58.935 ;
        RECT 162.145 57.560 162.405 57.820 ;
        RECT 157.865 56.830 158.415 57.380 ;
        RECT 160.835 56.850 161.385 57.400 ;
        RECT 163.865 56.830 164.415 57.380 ;
        RECT 166.875 56.860 167.425 57.410 ;
        RECT 169.905 56.840 170.455 57.390 ;
        RECT 174.815 57.000 175.075 57.260 ;
        RECT 175.135 57.000 175.395 57.260 ;
        RECT 173.125 56.685 173.385 56.945 ;
        RECT 173.445 56.685 173.705 56.945 ;
        RECT 176.550 56.685 176.810 56.945 ;
        RECT 176.870 56.685 177.130 56.945 ;
        RECT 174.975 55.230 175.235 55.490 ;
        RECT 148.810 52.940 149.345 53.475 ;
        RECT 151.840 52.920 152.375 53.455 ;
        RECT 154.850 52.950 155.385 53.485 ;
        RECT 157.880 52.930 158.415 53.465 ;
        RECT 160.850 52.950 161.385 53.485 ;
        RECT 163.880 52.930 164.415 53.465 ;
        RECT 166.890 52.960 167.425 53.495 ;
        RECT 169.920 52.940 170.455 53.475 ;
        RECT 148.775 49.160 149.310 49.695 ;
        RECT 151.805 49.180 152.340 49.715 ;
        RECT 154.815 49.150 155.350 49.685 ;
        RECT 157.845 49.170 158.380 49.705 ;
        RECT 160.815 49.150 161.350 49.685 ;
        RECT 163.855 49.145 164.390 49.680 ;
        RECT 166.855 49.140 167.390 49.675 ;
        RECT 169.885 49.160 170.420 49.695 ;
        RECT 41.595 45.110 41.855 45.370 ;
        RECT 42.760 45.120 43.020 45.380 ;
        RECT 43.940 45.120 44.200 45.380 ;
        RECT 45.130 45.120 45.390 45.380 ;
        RECT 46.300 45.120 46.560 45.380 ;
        RECT 148.760 45.245 149.310 45.795 ;
        RECT 151.790 45.265 152.340 45.815 ;
        RECT 154.800 45.235 155.350 45.785 ;
        RECT 157.830 45.255 158.380 45.805 ;
        RECT 160.800 45.235 161.350 45.785 ;
        RECT 163.840 45.230 164.390 45.780 ;
        RECT 166.840 45.225 167.390 45.775 ;
        RECT 169.870 45.245 170.420 45.795 ;
        RECT 143.065 44.550 143.325 44.810 ;
        RECT 12.750 43.090 13.010 43.350 ;
        RECT 13.915 43.010 14.175 43.270 ;
        RECT 15.095 42.990 15.355 43.250 ;
        RECT 16.285 42.930 16.545 43.190 ;
        RECT 17.455 42.950 17.715 43.210 ;
        RECT 22.365 43.090 22.625 43.350 ;
        RECT 23.530 43.010 23.790 43.270 ;
        RECT 24.710 42.990 24.970 43.250 ;
        RECT 25.900 42.930 26.160 43.190 ;
        RECT 27.070 42.950 27.330 43.210 ;
        RECT 31.980 43.090 32.240 43.350 ;
        RECT 33.145 43.010 33.405 43.270 ;
        RECT 34.325 42.990 34.585 43.250 ;
        RECT 35.515 42.930 35.775 43.190 ;
        RECT 36.685 42.950 36.945 43.210 ;
        RECT 41.595 43.090 41.855 43.350 ;
        RECT 42.760 43.010 43.020 43.270 ;
        RECT 43.940 42.990 44.200 43.250 ;
        RECT 45.130 42.930 45.390 43.190 ;
        RECT 46.300 42.950 46.560 43.210 ;
        RECT 148.760 42.855 149.020 43.115 ;
        RECT 18.020 42.140 18.280 42.400 ;
        RECT 27.635 42.140 27.895 42.400 ;
        RECT 37.250 42.140 37.510 42.400 ;
        RECT 46.865 42.140 47.125 42.400 ;
        RECT 148.770 41.485 149.030 41.745 ;
        RECT 148.790 40.090 149.050 40.350 ;
        RECT 16.350 39.490 16.610 39.750 ;
        RECT 25.965 39.490 26.225 39.750 ;
        RECT 35.580 39.490 35.840 39.750 ;
        RECT 45.195 39.490 45.455 39.750 ;
        RECT 17.265 39.145 17.525 39.405 ;
        RECT 18.605 39.135 18.865 39.395 ;
        RECT 26.880 39.145 27.140 39.405 ;
        RECT 28.220 39.135 28.480 39.395 ;
        RECT 36.495 39.145 36.755 39.405 ;
        RECT 37.835 39.135 38.095 39.395 ;
        RECT 46.110 39.145 46.370 39.405 ;
        RECT 47.450 39.135 47.710 39.395 ;
        RECT 148.790 38.735 149.050 38.995 ;
        RECT 148.765 37.345 149.025 37.605 ;
        RECT 148.760 35.975 149.020 36.235 ;
        RECT 148.795 34.585 149.055 34.845 ;
        RECT 148.780 33.235 149.040 33.495 ;
        RECT 148.790 31.850 149.050 32.110 ;
      LAYER met2 ;
        RECT 148.760 87.975 149.080 88.000 ;
        RECT 143.170 87.765 149.080 87.975 ;
        RECT 143.170 87.205 143.380 87.765 ;
        RECT 148.760 87.740 149.080 87.765 ;
        RECT 138.775 86.890 143.435 87.205 ;
        RECT 138.775 85.390 139.090 86.890 ;
        RECT 148.750 86.595 149.070 86.615 ;
        RECT 143.150 86.380 149.070 86.595 ;
        RECT 138.725 84.910 139.145 85.390 ;
        RECT 143.150 84.360 143.365 86.380 ;
        RECT 148.750 86.355 149.070 86.380 ;
        RECT 148.765 85.255 149.085 85.265 ;
        RECT 143.885 85.015 149.085 85.255 ;
        RECT 138.680 83.995 143.520 84.360 ;
        RECT 138.680 82.380 139.045 83.995 ;
        RECT 138.680 82.360 139.080 82.380 ;
        RECT 138.655 81.940 139.135 82.360 ;
        RECT 138.710 81.920 139.080 81.940 ;
        RECT 138.715 81.160 143.565 81.230 ;
        RECT 143.885 81.160 144.125 85.015 ;
        RECT 148.765 85.005 149.085 85.015 ;
        RECT 148.730 83.865 149.050 83.875 ;
        RECT 138.715 80.920 144.125 81.160 ;
        RECT 144.425 83.625 149.050 83.865 ;
        RECT 138.715 80.825 143.565 80.920 ;
        RECT 17.235 80.675 17.555 80.705 ;
        RECT 17.100 80.445 17.555 80.675 ;
        RECT 16.350 80.070 16.610 80.390 ;
        RECT 16.380 79.780 16.575 80.070 ;
        RECT 17.100 79.780 17.295 80.445 ;
        RECT 18.605 80.425 18.865 80.745 ;
        RECT 26.850 80.675 27.170 80.705 ;
        RECT 26.715 80.445 27.170 80.675 ;
        RECT 11.870 79.585 17.295 79.780 ;
        RECT 11.870 73.570 12.065 79.585 ;
        RECT 17.100 79.580 17.295 79.585 ;
        RECT 18.020 77.675 18.280 77.740 ;
        RECT 18.635 77.675 18.830 80.425 ;
        RECT 25.965 80.070 26.225 80.390 ;
        RECT 25.995 79.780 26.190 80.070 ;
        RECT 26.715 79.780 26.910 80.445 ;
        RECT 28.220 80.425 28.480 80.745 ;
        RECT 36.465 80.675 36.785 80.705 ;
        RECT 36.330 80.445 36.785 80.675 ;
        RECT 18.020 77.480 18.830 77.675 ;
        RECT 21.485 79.585 26.910 79.780 ;
        RECT 18.020 77.420 18.280 77.480 ;
        RECT 12.750 76.470 13.010 76.790 ;
        RECT 13.915 76.550 14.175 76.870 ;
        RECT 15.095 76.860 15.355 76.890 ;
        RECT 15.065 76.600 15.385 76.860 ;
        RECT 16.285 76.630 16.545 76.950 ;
        RECT 15.095 76.570 15.355 76.600 ;
        RECT 12.785 75.655 12.975 76.470 ;
        RECT 13.950 75.665 14.140 76.550 ;
        RECT 15.130 75.665 15.320 76.570 ;
        RECT 16.320 75.665 16.510 76.630 ;
        RECT 17.455 76.610 17.715 76.930 ;
        RECT 13.950 75.655 16.510 75.665 ;
        RECT 17.490 75.655 17.680 76.610 ;
        RECT 12.785 75.645 17.680 75.655 ;
        RECT 12.785 75.475 20.130 75.645 ;
        RECT 12.785 75.465 14.140 75.475 ;
        RECT 12.785 74.770 12.975 75.465 ;
        RECT 12.750 74.450 13.010 74.770 ;
        RECT 13.950 74.760 14.140 75.465 ;
        RECT 15.130 74.760 15.320 75.475 ;
        RECT 16.320 75.465 20.130 75.475 ;
        RECT 16.320 74.760 16.510 75.465 ;
        RECT 17.490 75.455 20.130 75.465 ;
        RECT 17.490 74.760 17.680 75.455 ;
        RECT 13.915 74.730 14.175 74.760 ;
        RECT 13.885 74.470 14.205 74.730 ;
        RECT 13.915 74.440 14.175 74.470 ;
        RECT 15.095 74.440 15.355 74.760 ;
        RECT 16.285 74.440 16.545 74.760 ;
        RECT 17.455 74.440 17.715 74.760 ;
        RECT 12.415 73.570 12.735 73.600 ;
        RECT 11.870 73.375 12.735 73.570 ;
        RECT 12.415 73.340 12.735 73.375 ;
        RECT 17.065 73.360 17.385 73.620 ;
        RECT 19.940 72.445 20.130 75.455 ;
        RECT 21.485 73.570 21.680 79.585 ;
        RECT 26.715 79.580 26.910 79.585 ;
        RECT 27.635 77.675 27.895 77.740 ;
        RECT 28.250 77.675 28.445 80.425 ;
        RECT 35.580 80.070 35.840 80.390 ;
        RECT 35.610 79.780 35.805 80.070 ;
        RECT 36.330 79.780 36.525 80.445 ;
        RECT 37.835 80.425 38.095 80.745 ;
        RECT 46.080 80.675 46.400 80.705 ;
        RECT 45.945 80.445 46.400 80.675 ;
        RECT 27.635 77.480 28.445 77.675 ;
        RECT 31.100 79.585 36.525 79.780 ;
        RECT 27.635 77.420 27.895 77.480 ;
        RECT 22.365 76.470 22.625 76.790 ;
        RECT 23.530 76.550 23.790 76.870 ;
        RECT 24.710 76.860 24.970 76.890 ;
        RECT 24.680 76.600 25.000 76.860 ;
        RECT 25.900 76.630 26.160 76.950 ;
        RECT 24.710 76.570 24.970 76.600 ;
        RECT 22.400 75.655 22.590 76.470 ;
        RECT 23.565 75.665 23.755 76.550 ;
        RECT 24.745 75.665 24.935 76.570 ;
        RECT 25.935 75.665 26.125 76.630 ;
        RECT 27.070 76.610 27.330 76.930 ;
        RECT 23.565 75.655 26.125 75.665 ;
        RECT 27.105 75.655 27.295 76.610 ;
        RECT 22.400 75.645 27.295 75.655 ;
        RECT 28.900 75.645 29.680 75.655 ;
        RECT 22.400 75.475 29.680 75.645 ;
        RECT 22.400 75.465 23.755 75.475 ;
        RECT 22.400 74.770 22.590 75.465 ;
        RECT 22.365 74.450 22.625 74.770 ;
        RECT 23.565 74.760 23.755 75.465 ;
        RECT 24.745 74.760 24.935 75.475 ;
        RECT 25.935 75.465 29.680 75.475 ;
        RECT 25.935 74.760 26.125 75.465 ;
        RECT 27.105 75.455 29.095 75.465 ;
        RECT 27.105 74.760 27.295 75.455 ;
        RECT 23.530 74.730 23.790 74.760 ;
        RECT 23.500 74.470 23.820 74.730 ;
        RECT 23.530 74.440 23.790 74.470 ;
        RECT 24.710 74.440 24.970 74.760 ;
        RECT 25.900 74.440 26.160 74.760 ;
        RECT 27.070 74.440 27.330 74.760 ;
        RECT 22.030 73.570 22.350 73.600 ;
        RECT 21.485 73.375 22.350 73.570 ;
        RECT 22.030 73.340 22.350 73.375 ;
        RECT 26.680 73.360 27.000 73.620 ;
        RECT 29.490 72.445 29.680 75.465 ;
        RECT 31.100 73.570 31.295 79.585 ;
        RECT 36.330 79.580 36.525 79.585 ;
        RECT 37.250 77.675 37.510 77.740 ;
        RECT 37.865 77.675 38.060 80.425 ;
        RECT 45.195 80.070 45.455 80.390 ;
        RECT 45.225 79.780 45.420 80.070 ;
        RECT 45.945 79.780 46.140 80.445 ;
        RECT 47.450 80.425 47.710 80.745 ;
        RECT 37.250 77.480 38.060 77.675 ;
        RECT 40.715 79.585 46.140 79.780 ;
        RECT 37.250 77.420 37.510 77.480 ;
        RECT 31.980 76.470 32.240 76.790 ;
        RECT 33.145 76.550 33.405 76.870 ;
        RECT 34.325 76.860 34.585 76.890 ;
        RECT 34.295 76.600 34.615 76.860 ;
        RECT 35.515 76.630 35.775 76.950 ;
        RECT 34.325 76.570 34.585 76.600 ;
        RECT 32.015 75.655 32.205 76.470 ;
        RECT 33.180 75.665 33.370 76.550 ;
        RECT 34.360 75.665 34.550 76.570 ;
        RECT 35.550 75.665 35.740 76.630 ;
        RECT 36.685 76.610 36.945 76.930 ;
        RECT 33.180 75.655 35.740 75.665 ;
        RECT 36.720 75.655 36.910 76.610 ;
        RECT 32.015 75.645 36.910 75.655 ;
        RECT 32.015 75.475 39.100 75.645 ;
        RECT 32.015 75.465 33.370 75.475 ;
        RECT 32.015 74.770 32.205 75.465 ;
        RECT 31.980 74.450 32.240 74.770 ;
        RECT 33.180 74.760 33.370 75.465 ;
        RECT 34.360 74.760 34.550 75.475 ;
        RECT 35.550 75.465 39.100 75.475 ;
        RECT 35.550 74.760 35.740 75.465 ;
        RECT 36.720 75.455 39.100 75.465 ;
        RECT 36.720 74.760 36.910 75.455 ;
        RECT 33.145 74.730 33.405 74.760 ;
        RECT 33.115 74.470 33.435 74.730 ;
        RECT 33.145 74.440 33.405 74.470 ;
        RECT 34.325 74.440 34.585 74.760 ;
        RECT 35.515 74.440 35.775 74.760 ;
        RECT 36.685 74.440 36.945 74.760 ;
        RECT 31.645 73.570 31.965 73.600 ;
        RECT 31.100 73.375 31.965 73.570 ;
        RECT 31.645 73.340 31.965 73.375 ;
        RECT 36.295 73.360 36.615 73.620 ;
        RECT 38.910 72.445 39.100 75.455 ;
        RECT 40.715 73.570 40.910 79.585 ;
        RECT 45.945 79.580 46.140 79.585 ;
        RECT 46.865 77.675 47.125 77.740 ;
        RECT 47.480 77.675 47.675 80.425 ;
        RECT 138.715 78.380 139.120 80.825 ;
        RECT 136.610 78.360 139.120 78.380 ;
        RECT 136.590 78.005 139.120 78.360 ;
        RECT 136.610 77.975 139.120 78.005 ;
        RECT 140.020 78.265 140.490 78.295 ;
        RECT 140.020 78.220 143.560 78.265 ;
        RECT 144.425 78.220 144.665 83.625 ;
        RECT 148.730 83.615 149.050 83.625 ;
        RECT 148.735 82.495 149.055 82.505 ;
        RECT 140.020 77.980 144.665 78.220 ;
        RECT 144.905 82.255 149.055 82.495 ;
        RECT 140.020 77.855 143.560 77.980 ;
        RECT 140.020 77.825 140.490 77.855 ;
        RECT 46.865 77.480 47.675 77.675 ;
        RECT 46.865 77.420 47.125 77.480 ;
        RECT 41.595 76.470 41.855 76.790 ;
        RECT 42.760 76.550 43.020 76.870 ;
        RECT 43.940 76.860 44.200 76.890 ;
        RECT 43.910 76.600 44.230 76.860 ;
        RECT 45.130 76.630 45.390 76.950 ;
        RECT 43.940 76.570 44.200 76.600 ;
        RECT 41.630 75.655 41.820 76.470 ;
        RECT 42.795 75.665 42.985 76.550 ;
        RECT 43.975 75.665 44.165 76.570 ;
        RECT 45.165 75.665 45.355 76.630 ;
        RECT 46.300 76.610 46.560 76.930 ;
        RECT 42.795 75.655 45.355 75.665 ;
        RECT 46.335 75.655 46.525 76.610 ;
        RECT 41.630 75.645 46.525 75.655 ;
        RECT 48.160 75.645 48.740 75.655 ;
        RECT 41.630 75.475 48.740 75.645 ;
        RECT 41.630 75.465 42.985 75.475 ;
        RECT 41.630 74.770 41.820 75.465 ;
        RECT 41.595 74.450 41.855 74.770 ;
        RECT 42.795 74.760 42.985 75.465 ;
        RECT 43.975 74.760 44.165 75.475 ;
        RECT 45.165 75.465 48.740 75.475 ;
        RECT 45.165 74.760 45.355 75.465 ;
        RECT 46.335 75.455 48.325 75.465 ;
        RECT 46.335 74.760 46.525 75.455 ;
        RECT 42.760 74.730 43.020 74.760 ;
        RECT 42.730 74.470 43.050 74.730 ;
        RECT 42.760 74.440 43.020 74.470 ;
        RECT 43.940 74.440 44.200 74.760 ;
        RECT 45.130 74.440 45.390 74.760 ;
        RECT 46.300 74.440 46.560 74.760 ;
        RECT 41.260 73.570 41.580 73.600 ;
        RECT 40.715 73.375 41.580 73.570 ;
        RECT 41.260 73.340 41.580 73.375 ;
        RECT 45.910 73.360 46.230 73.620 ;
        RECT 48.550 72.445 48.740 75.465 ;
        RECT 132.700 75.370 133.070 75.390 ;
        RECT 132.645 74.950 133.125 75.370 ;
        RECT 132.700 74.930 133.070 74.950 ;
        RECT 19.940 72.255 48.740 72.445 ;
        RECT 136.635 72.365 136.990 72.400 ;
        RECT 140.050 72.365 140.455 77.825 ;
        RECT 143.035 75.290 143.355 75.300 ;
        RECT 144.905 75.290 145.145 82.255 ;
        RECT 148.735 82.245 149.055 82.255 ;
        RECT 143.035 75.050 145.145 75.290 ;
        RECT 145.310 80.860 149.080 81.115 ;
        RECT 143.035 75.040 143.355 75.050 ;
        RECT 128.605 72.275 128.975 72.295 ;
        RECT 22.840 71.845 23.030 72.255 ;
        RECT 128.550 71.855 129.030 72.275 ;
        RECT 136.610 71.960 140.455 72.365 ;
        RECT 145.310 72.230 145.565 80.860 ;
        RECT 148.760 80.855 149.080 80.860 ;
        RECT 148.760 79.740 149.080 79.760 ;
        RECT 143.120 71.975 145.565 72.230 ;
        RECT 145.705 79.520 149.080 79.740 ;
        RECT 143.120 71.970 143.440 71.975 ;
        RECT 136.635 71.935 136.990 71.960 ;
        RECT 22.785 71.455 23.085 71.845 ;
        RECT 128.605 71.835 128.975 71.855 ;
        RECT 122.535 69.270 122.850 69.300 ;
        RECT 120.725 68.955 122.850 69.270 ;
        RECT 143.075 69.230 143.395 69.250 ;
        RECT 145.705 69.230 145.925 79.520 ;
        RECT 148.760 79.500 149.080 79.520 ;
        RECT 148.740 78.355 149.060 78.365 ;
        RECT 143.075 69.010 145.925 69.230 ;
        RECT 146.090 78.120 149.060 78.355 ;
        RECT 143.075 68.990 143.395 69.010 ;
        RECT 122.535 68.925 122.850 68.955 ;
        RECT 78.640 66.290 143.460 66.350 ;
        RECT 146.090 66.290 146.325 78.120 ;
        RECT 148.740 78.105 149.060 78.120 ;
        RECT 78.640 66.055 146.325 66.290 ;
        RECT 146.560 76.740 149.050 76.995 ;
        RECT 78.640 65.970 143.460 66.055 ;
        RECT 74.485 63.280 74.930 64.605 ;
        RECT 78.640 64.115 79.020 65.970 ;
        RECT 74.460 63.200 143.485 63.280 ;
        RECT 146.560 63.200 146.815 76.740 ;
        RECT 148.730 76.735 149.050 76.740 ;
        RECT 148.645 74.710 149.195 74.765 ;
        RECT 148.625 74.210 149.215 74.710 ;
        RECT 151.675 74.690 152.225 74.745 ;
        RECT 154.685 74.720 155.235 74.775 ;
        RECT 148.645 74.155 149.195 74.210 ;
        RECT 151.655 74.190 152.245 74.690 ;
        RECT 154.665 74.220 155.255 74.720 ;
        RECT 157.715 74.700 158.265 74.755 ;
        RECT 160.685 74.720 161.235 74.775 ;
        RECT 163.725 74.725 164.275 74.780 ;
        RECT 166.725 74.730 167.275 74.785 ;
        RECT 151.675 74.135 152.225 74.190 ;
        RECT 154.685 74.165 155.235 74.220 ;
        RECT 157.695 74.200 158.285 74.700 ;
        RECT 160.665 74.220 161.255 74.720 ;
        RECT 163.705 74.225 164.295 74.725 ;
        RECT 166.705 74.230 167.295 74.730 ;
        RECT 169.755 74.710 170.305 74.765 ;
        RECT 157.715 74.145 158.265 74.200 ;
        RECT 160.685 74.165 161.235 74.220 ;
        RECT 163.725 74.170 164.275 74.225 ;
        RECT 166.725 74.175 167.275 74.230 ;
        RECT 169.735 74.210 170.325 74.710 ;
        RECT 169.755 74.155 170.305 74.210 ;
        RECT 148.660 70.795 149.195 70.850 ;
        RECT 148.640 70.310 149.215 70.795 ;
        RECT 151.690 70.775 152.225 70.830 ;
        RECT 154.700 70.805 155.235 70.860 ;
        RECT 148.660 70.255 149.195 70.310 ;
        RECT 151.670 70.290 152.245 70.775 ;
        RECT 154.680 70.320 155.255 70.805 ;
        RECT 157.730 70.785 158.265 70.840 ;
        RECT 160.700 70.805 161.235 70.860 ;
        RECT 163.740 70.810 164.275 70.865 ;
        RECT 166.740 70.815 167.275 70.870 ;
        RECT 151.690 70.235 152.225 70.290 ;
        RECT 154.700 70.265 155.235 70.320 ;
        RECT 157.710 70.300 158.285 70.785 ;
        RECT 160.680 70.320 161.255 70.805 ;
        RECT 163.720 70.325 164.295 70.810 ;
        RECT 166.720 70.330 167.295 70.815 ;
        RECT 169.770 70.795 170.305 70.850 ;
        RECT 157.730 70.245 158.265 70.300 ;
        RECT 160.700 70.265 161.235 70.320 ;
        RECT 163.740 70.270 164.275 70.325 ;
        RECT 166.740 70.275 167.275 70.330 ;
        RECT 169.750 70.310 170.325 70.795 ;
        RECT 169.770 70.255 170.305 70.310 ;
        RECT 170.065 67.590 170.385 67.640 ;
        RECT 162.285 67.430 170.385 67.590 ;
        RECT 148.695 67.015 149.230 67.070 ;
        RECT 151.725 67.035 152.260 67.090 ;
        RECT 148.675 66.530 149.250 67.015 ;
        RECT 151.705 66.550 152.280 67.035 ;
        RECT 154.735 67.005 155.270 67.060 ;
        RECT 157.765 67.025 158.300 67.080 ;
        RECT 148.695 66.475 149.230 66.530 ;
        RECT 151.725 66.495 152.260 66.550 ;
        RECT 154.715 66.520 155.290 67.005 ;
        RECT 157.745 66.540 158.320 67.025 ;
        RECT 160.735 67.005 161.270 67.060 ;
        RECT 154.735 66.465 155.270 66.520 ;
        RECT 157.765 66.485 158.300 66.540 ;
        RECT 160.715 66.520 161.290 67.005 ;
        RECT 160.735 66.465 161.270 66.520 ;
        RECT 74.460 62.945 146.815 63.200 ;
        RECT 148.680 63.115 149.230 63.170 ;
        RECT 151.710 63.135 152.260 63.190 ;
        RECT 74.460 62.835 143.485 62.945 ;
        RECT 74.485 62.830 74.930 62.835 ;
        RECT 148.660 62.615 149.250 63.115 ;
        RECT 151.690 62.635 152.280 63.135 ;
        RECT 154.720 63.105 155.270 63.160 ;
        RECT 157.750 63.125 158.300 63.180 ;
        RECT 148.680 62.560 149.230 62.615 ;
        RECT 151.710 62.580 152.260 62.635 ;
        RECT 154.700 62.605 155.290 63.105 ;
        RECT 157.730 62.625 158.320 63.125 ;
        RECT 160.720 63.105 161.270 63.160 ;
        RECT 154.720 62.550 155.270 62.605 ;
        RECT 157.750 62.570 158.300 62.625 ;
        RECT 160.700 62.605 161.290 63.105 ;
        RECT 160.720 62.550 161.270 62.605 ;
        RECT 162.285 62.460 162.445 67.430 ;
        RECT 170.065 67.380 170.385 67.430 ;
        RECT 163.765 67.025 164.300 67.080 ;
        RECT 163.745 66.540 164.320 67.025 ;
        RECT 166.775 66.995 167.310 67.050 ;
        RECT 169.805 67.015 170.340 67.070 ;
        RECT 163.765 66.485 164.300 66.540 ;
        RECT 166.755 66.510 167.330 66.995 ;
        RECT 169.785 66.530 170.360 67.015 ;
        RECT 166.775 66.455 167.310 66.510 ;
        RECT 169.805 66.475 170.340 66.530 ;
        RECT 173.115 64.810 173.715 64.895 ;
        RECT 176.540 64.810 177.140 64.895 ;
        RECT 173.115 64.580 177.140 64.810 ;
        RECT 173.115 64.495 173.715 64.580 ;
        RECT 174.805 64.180 175.405 64.580 ;
        RECT 176.540 64.495 177.140 64.580 ;
        RECT 163.750 63.125 164.300 63.180 ;
        RECT 163.730 62.625 164.320 63.125 ;
        RECT 166.760 63.095 167.310 63.150 ;
        RECT 169.790 63.115 170.340 63.170 ;
        RECT 163.750 62.570 164.300 62.625 ;
        RECT 166.740 62.595 167.330 63.095 ;
        RECT 169.770 62.615 170.360 63.115 ;
        RECT 166.760 62.540 167.310 62.595 ;
        RECT 169.790 62.560 170.340 62.615 ;
        RECT 152.045 62.160 152.325 62.255 ;
        RECT 162.205 62.200 162.525 62.460 ;
        RECT 152.045 61.985 156.490 62.160 ;
        RECT 152.045 61.885 152.325 61.985 ;
        RECT 156.315 60.595 156.490 61.985 ;
        RECT 159.935 61.335 160.255 61.595 ;
        RECT 156.275 60.275 156.535 60.595 ;
        RECT 159.375 60.325 159.635 60.645 ;
        RECT 156.235 59.680 156.535 60.030 ;
        RECT 156.200 59.400 156.570 59.680 ;
        RECT 156.235 59.390 156.535 59.400 ;
        RECT 159.425 58.965 159.585 60.325 ;
        RECT 160.015 60.015 160.175 61.335 ;
        RECT 173.115 60.070 173.715 60.155 ;
        RECT 174.805 60.070 175.405 60.470 ;
        RECT 176.540 60.070 177.140 60.155 ;
        RECT 159.965 59.695 160.225 60.015 ;
        RECT 173.115 59.840 177.140 60.070 ;
        RECT 173.115 59.755 173.715 59.840 ;
        RECT 176.540 59.755 177.140 59.840 ;
        RECT 159.375 58.645 159.635 58.965 ;
        RECT 162.115 57.560 162.435 57.820 ;
        RECT 148.795 57.365 149.345 57.420 ;
        RECT 74.485 57.015 74.930 57.020 ;
        RECT 74.460 56.905 143.485 57.015 ;
        RECT 74.460 56.650 146.815 56.905 ;
        RECT 148.775 56.865 149.365 57.365 ;
        RECT 151.825 57.345 152.375 57.400 ;
        RECT 154.835 57.375 155.385 57.430 ;
        RECT 148.795 56.810 149.345 56.865 ;
        RECT 151.805 56.845 152.395 57.345 ;
        RECT 154.815 56.875 155.405 57.375 ;
        RECT 157.865 57.355 158.415 57.410 ;
        RECT 160.835 57.375 161.385 57.430 ;
        RECT 151.825 56.790 152.375 56.845 ;
        RECT 154.835 56.820 155.385 56.875 ;
        RECT 157.845 56.855 158.435 57.355 ;
        RECT 160.815 56.875 161.405 57.375 ;
        RECT 157.865 56.800 158.415 56.855 ;
        RECT 160.835 56.820 161.385 56.875 ;
        RECT 74.460 56.570 143.485 56.650 ;
        RECT 74.485 55.245 74.930 56.570 ;
        RECT 78.640 53.880 79.020 55.735 ;
        RECT 78.640 53.795 143.460 53.880 ;
        RECT 78.640 53.560 146.325 53.795 ;
        RECT 78.640 53.500 143.460 53.560 ;
        RECT 122.535 50.895 122.850 50.925 ;
        RECT 120.725 50.580 122.850 50.895 ;
        RECT 143.075 50.840 143.395 50.860 ;
        RECT 143.075 50.620 145.925 50.840 ;
        RECT 143.075 50.600 143.395 50.620 ;
        RECT 122.535 50.550 122.850 50.580 ;
        RECT 22.785 48.005 23.085 48.395 ;
        RECT 22.840 47.595 23.030 48.005 ;
        RECT 128.605 47.995 128.975 48.015 ;
        RECT 19.940 47.405 48.740 47.595 ;
        RECT 128.550 47.575 129.030 47.995 ;
        RECT 136.635 47.890 136.990 47.915 ;
        RECT 128.605 47.555 128.975 47.575 ;
        RECT 136.610 47.485 140.455 47.890 ;
        RECT 143.120 47.875 143.440 47.880 ;
        RECT 143.120 47.620 145.565 47.875 ;
        RECT 136.635 47.450 136.990 47.485 ;
        RECT 12.415 46.475 12.735 46.510 ;
        RECT 11.870 46.280 12.735 46.475 ;
        RECT 11.870 40.265 12.065 46.280 ;
        RECT 12.415 46.250 12.735 46.280 ;
        RECT 17.065 46.230 17.385 46.490 ;
        RECT 12.750 45.080 13.010 45.400 ;
        RECT 13.915 45.380 14.175 45.410 ;
        RECT 13.885 45.120 14.205 45.380 ;
        RECT 13.915 45.090 14.175 45.120 ;
        RECT 15.095 45.090 15.355 45.410 ;
        RECT 16.285 45.090 16.545 45.410 ;
        RECT 17.455 45.090 17.715 45.410 ;
        RECT 12.785 44.385 12.975 45.080 ;
        RECT 13.950 44.385 14.140 45.090 ;
        RECT 12.785 44.375 14.140 44.385 ;
        RECT 15.130 44.375 15.320 45.090 ;
        RECT 16.320 44.385 16.510 45.090 ;
        RECT 17.490 44.395 17.680 45.090 ;
        RECT 19.940 44.395 20.130 47.405 ;
        RECT 22.030 46.475 22.350 46.510 ;
        RECT 17.490 44.385 20.130 44.395 ;
        RECT 16.320 44.375 20.130 44.385 ;
        RECT 12.785 44.205 20.130 44.375 ;
        RECT 21.485 46.280 22.350 46.475 ;
        RECT 12.785 44.195 17.680 44.205 ;
        RECT 12.785 43.380 12.975 44.195 ;
        RECT 13.950 44.185 16.510 44.195 ;
        RECT 12.750 43.060 13.010 43.380 ;
        RECT 13.950 43.300 14.140 44.185 ;
        RECT 13.915 42.980 14.175 43.300 ;
        RECT 15.130 43.280 15.320 44.185 ;
        RECT 15.095 43.250 15.355 43.280 ;
        RECT 15.065 42.990 15.385 43.250 ;
        RECT 16.320 43.220 16.510 44.185 ;
        RECT 17.490 43.240 17.680 44.195 ;
        RECT 15.095 42.960 15.355 42.990 ;
        RECT 16.285 42.900 16.545 43.220 ;
        RECT 17.455 42.920 17.715 43.240 ;
        RECT 18.020 42.370 18.280 42.430 ;
        RECT 18.020 42.175 18.830 42.370 ;
        RECT 18.020 42.110 18.280 42.175 ;
        RECT 17.100 40.265 17.295 40.270 ;
        RECT 11.870 40.070 17.295 40.265 ;
        RECT 16.380 39.780 16.575 40.070 ;
        RECT 16.350 39.460 16.610 39.780 ;
        RECT 17.100 39.405 17.295 40.070 ;
        RECT 18.635 39.425 18.830 42.175 ;
        RECT 21.485 40.265 21.680 46.280 ;
        RECT 22.030 46.250 22.350 46.280 ;
        RECT 26.680 46.230 27.000 46.490 ;
        RECT 22.365 45.080 22.625 45.400 ;
        RECT 23.530 45.380 23.790 45.410 ;
        RECT 23.500 45.120 23.820 45.380 ;
        RECT 23.530 45.090 23.790 45.120 ;
        RECT 24.710 45.090 24.970 45.410 ;
        RECT 25.900 45.090 26.160 45.410 ;
        RECT 27.070 45.090 27.330 45.410 ;
        RECT 22.400 44.385 22.590 45.080 ;
        RECT 23.565 44.385 23.755 45.090 ;
        RECT 22.400 44.375 23.755 44.385 ;
        RECT 24.745 44.375 24.935 45.090 ;
        RECT 25.935 44.385 26.125 45.090 ;
        RECT 27.105 44.395 27.295 45.090 ;
        RECT 27.105 44.385 29.095 44.395 ;
        RECT 29.490 44.385 29.680 47.405 ;
        RECT 31.645 46.475 31.965 46.510 ;
        RECT 25.935 44.375 29.680 44.385 ;
        RECT 22.400 44.205 29.680 44.375 ;
        RECT 22.400 44.195 27.295 44.205 ;
        RECT 28.900 44.195 29.680 44.205 ;
        RECT 31.100 46.280 31.965 46.475 ;
        RECT 22.400 43.380 22.590 44.195 ;
        RECT 23.565 44.185 26.125 44.195 ;
        RECT 22.365 43.060 22.625 43.380 ;
        RECT 23.565 43.300 23.755 44.185 ;
        RECT 23.530 42.980 23.790 43.300 ;
        RECT 24.745 43.280 24.935 44.185 ;
        RECT 24.710 43.250 24.970 43.280 ;
        RECT 24.680 42.990 25.000 43.250 ;
        RECT 25.935 43.220 26.125 44.185 ;
        RECT 27.105 43.240 27.295 44.195 ;
        RECT 24.710 42.960 24.970 42.990 ;
        RECT 25.900 42.900 26.160 43.220 ;
        RECT 27.070 42.920 27.330 43.240 ;
        RECT 27.635 42.370 27.895 42.430 ;
        RECT 27.635 42.175 28.445 42.370 ;
        RECT 27.635 42.110 27.895 42.175 ;
        RECT 26.715 40.265 26.910 40.270 ;
        RECT 21.485 40.070 26.910 40.265 ;
        RECT 25.995 39.780 26.190 40.070 ;
        RECT 25.965 39.460 26.225 39.780 ;
        RECT 17.100 39.175 17.555 39.405 ;
        RECT 17.235 39.145 17.555 39.175 ;
        RECT 18.605 39.105 18.865 39.425 ;
        RECT 26.715 39.405 26.910 40.070 ;
        RECT 28.250 39.425 28.445 42.175 ;
        RECT 31.100 40.265 31.295 46.280 ;
        RECT 31.645 46.250 31.965 46.280 ;
        RECT 36.295 46.230 36.615 46.490 ;
        RECT 31.980 45.080 32.240 45.400 ;
        RECT 33.145 45.380 33.405 45.410 ;
        RECT 33.115 45.120 33.435 45.380 ;
        RECT 33.145 45.090 33.405 45.120 ;
        RECT 34.325 45.090 34.585 45.410 ;
        RECT 35.515 45.090 35.775 45.410 ;
        RECT 36.685 45.090 36.945 45.410 ;
        RECT 32.015 44.385 32.205 45.080 ;
        RECT 33.180 44.385 33.370 45.090 ;
        RECT 32.015 44.375 33.370 44.385 ;
        RECT 34.360 44.375 34.550 45.090 ;
        RECT 35.550 44.385 35.740 45.090 ;
        RECT 36.720 44.395 36.910 45.090 ;
        RECT 38.910 44.395 39.100 47.405 ;
        RECT 41.260 46.475 41.580 46.510 ;
        RECT 36.720 44.385 39.100 44.395 ;
        RECT 35.550 44.375 39.100 44.385 ;
        RECT 32.015 44.205 39.100 44.375 ;
        RECT 40.715 46.280 41.580 46.475 ;
        RECT 32.015 44.195 36.910 44.205 ;
        RECT 32.015 43.380 32.205 44.195 ;
        RECT 33.180 44.185 35.740 44.195 ;
        RECT 31.980 43.060 32.240 43.380 ;
        RECT 33.180 43.300 33.370 44.185 ;
        RECT 33.145 42.980 33.405 43.300 ;
        RECT 34.360 43.280 34.550 44.185 ;
        RECT 34.325 43.250 34.585 43.280 ;
        RECT 34.295 42.990 34.615 43.250 ;
        RECT 35.550 43.220 35.740 44.185 ;
        RECT 36.720 43.240 36.910 44.195 ;
        RECT 34.325 42.960 34.585 42.990 ;
        RECT 35.515 42.900 35.775 43.220 ;
        RECT 36.685 42.920 36.945 43.240 ;
        RECT 37.250 42.370 37.510 42.430 ;
        RECT 37.250 42.175 38.060 42.370 ;
        RECT 37.250 42.110 37.510 42.175 ;
        RECT 36.330 40.265 36.525 40.270 ;
        RECT 31.100 40.070 36.525 40.265 ;
        RECT 35.610 39.780 35.805 40.070 ;
        RECT 35.580 39.460 35.840 39.780 ;
        RECT 26.715 39.175 27.170 39.405 ;
        RECT 26.850 39.145 27.170 39.175 ;
        RECT 28.220 39.105 28.480 39.425 ;
        RECT 36.330 39.405 36.525 40.070 ;
        RECT 37.865 39.425 38.060 42.175 ;
        RECT 40.715 40.265 40.910 46.280 ;
        RECT 41.260 46.250 41.580 46.280 ;
        RECT 45.910 46.230 46.230 46.490 ;
        RECT 41.595 45.080 41.855 45.400 ;
        RECT 42.760 45.380 43.020 45.410 ;
        RECT 42.730 45.120 43.050 45.380 ;
        RECT 42.760 45.090 43.020 45.120 ;
        RECT 43.940 45.090 44.200 45.410 ;
        RECT 45.130 45.090 45.390 45.410 ;
        RECT 46.300 45.090 46.560 45.410 ;
        RECT 41.630 44.385 41.820 45.080 ;
        RECT 42.795 44.385 42.985 45.090 ;
        RECT 41.630 44.375 42.985 44.385 ;
        RECT 43.975 44.375 44.165 45.090 ;
        RECT 45.165 44.385 45.355 45.090 ;
        RECT 46.335 44.395 46.525 45.090 ;
        RECT 46.335 44.385 48.325 44.395 ;
        RECT 48.550 44.385 48.740 47.405 ;
        RECT 132.700 44.900 133.070 44.920 ;
        RECT 132.645 44.480 133.125 44.900 ;
        RECT 132.700 44.460 133.070 44.480 ;
        RECT 45.165 44.375 48.740 44.385 ;
        RECT 41.630 44.205 48.740 44.375 ;
        RECT 41.630 44.195 46.525 44.205 ;
        RECT 48.160 44.195 48.740 44.205 ;
        RECT 41.630 43.380 41.820 44.195 ;
        RECT 42.795 44.185 45.355 44.195 ;
        RECT 41.595 43.060 41.855 43.380 ;
        RECT 42.795 43.300 42.985 44.185 ;
        RECT 42.760 42.980 43.020 43.300 ;
        RECT 43.975 43.280 44.165 44.185 ;
        RECT 43.940 43.250 44.200 43.280 ;
        RECT 43.910 42.990 44.230 43.250 ;
        RECT 45.165 43.220 45.355 44.185 ;
        RECT 46.335 43.240 46.525 44.195 ;
        RECT 43.940 42.960 44.200 42.990 ;
        RECT 45.130 42.900 45.390 43.220 ;
        RECT 46.300 42.920 46.560 43.240 ;
        RECT 46.865 42.370 47.125 42.430 ;
        RECT 46.865 42.175 47.675 42.370 ;
        RECT 46.865 42.110 47.125 42.175 ;
        RECT 45.945 40.265 46.140 40.270 ;
        RECT 40.715 40.070 46.140 40.265 ;
        RECT 45.225 39.780 45.420 40.070 ;
        RECT 45.195 39.460 45.455 39.780 ;
        RECT 36.330 39.175 36.785 39.405 ;
        RECT 36.465 39.145 36.785 39.175 ;
        RECT 37.835 39.105 38.095 39.425 ;
        RECT 45.945 39.405 46.140 40.070 ;
        RECT 47.480 39.425 47.675 42.175 ;
        RECT 140.050 42.025 140.455 47.485 ;
        RECT 143.035 44.800 143.355 44.810 ;
        RECT 143.035 44.560 145.145 44.800 ;
        RECT 143.035 44.550 143.355 44.560 ;
        RECT 140.020 41.995 140.490 42.025 ;
        RECT 136.610 41.845 139.120 41.875 ;
        RECT 136.590 41.490 139.120 41.845 ;
        RECT 140.020 41.870 143.560 41.995 ;
        RECT 140.020 41.630 144.665 41.870 ;
        RECT 140.020 41.585 143.560 41.630 ;
        RECT 140.020 41.555 140.490 41.585 ;
        RECT 136.610 41.470 139.120 41.490 ;
        RECT 45.945 39.175 46.400 39.405 ;
        RECT 46.080 39.145 46.400 39.175 ;
        RECT 47.450 39.105 47.710 39.425 ;
        RECT 138.715 39.025 139.120 41.470 ;
        RECT 138.715 38.930 143.565 39.025 ;
        RECT 138.715 38.690 144.125 38.930 ;
        RECT 138.715 38.620 143.565 38.690 ;
        RECT 138.710 37.910 139.080 37.930 ;
        RECT 138.655 37.490 139.135 37.910 ;
        RECT 138.680 37.470 139.080 37.490 ;
        RECT 138.680 35.855 139.045 37.470 ;
        RECT 138.680 35.490 143.520 35.855 ;
        RECT 138.725 34.460 139.145 34.940 ;
        RECT 138.775 32.960 139.090 34.460 ;
        RECT 143.150 33.470 143.365 35.490 ;
        RECT 143.885 34.835 144.125 38.690 ;
        RECT 144.425 36.225 144.665 41.630 ;
        RECT 144.905 37.595 145.145 44.560 ;
        RECT 145.310 38.990 145.565 47.620 ;
        RECT 145.705 40.330 145.925 50.620 ;
        RECT 146.090 41.730 146.325 53.560 ;
        RECT 146.560 43.110 146.815 56.650 ;
        RECT 162.195 54.570 162.355 57.560 ;
        RECT 163.865 57.355 164.415 57.410 ;
        RECT 166.875 57.385 167.425 57.440 ;
        RECT 163.845 56.855 164.435 57.355 ;
        RECT 166.855 56.885 167.445 57.385 ;
        RECT 169.905 57.365 170.455 57.420 ;
        RECT 163.865 56.800 164.415 56.855 ;
        RECT 166.875 56.830 167.425 56.885 ;
        RECT 169.885 56.865 170.475 57.365 ;
        RECT 173.115 56.930 173.715 57.015 ;
        RECT 174.805 56.930 175.405 57.330 ;
        RECT 176.540 56.930 177.140 57.015 ;
        RECT 169.905 56.810 170.455 56.865 ;
        RECT 173.115 56.700 177.140 56.930 ;
        RECT 173.115 56.615 173.715 56.700 ;
        RECT 176.540 56.615 177.140 56.700 ;
        RECT 174.975 55.200 175.235 55.520 ;
        RECT 175.025 54.570 175.185 55.200 ;
        RECT 162.195 54.410 175.185 54.570 ;
        RECT 148.810 53.450 149.345 53.505 ;
        RECT 148.790 52.965 149.365 53.450 ;
        RECT 151.840 53.430 152.375 53.485 ;
        RECT 154.850 53.460 155.385 53.515 ;
        RECT 148.810 52.910 149.345 52.965 ;
        RECT 151.820 52.945 152.395 53.430 ;
        RECT 154.830 52.975 155.405 53.460 ;
        RECT 157.880 53.440 158.415 53.495 ;
        RECT 160.850 53.460 161.385 53.515 ;
        RECT 151.840 52.890 152.375 52.945 ;
        RECT 154.850 52.920 155.385 52.975 ;
        RECT 157.860 52.955 158.435 53.440 ;
        RECT 160.830 52.975 161.405 53.460 ;
        RECT 163.880 53.440 164.415 53.495 ;
        RECT 166.890 53.470 167.425 53.525 ;
        RECT 157.880 52.900 158.415 52.955 ;
        RECT 160.850 52.920 161.385 52.975 ;
        RECT 163.860 52.955 164.435 53.440 ;
        RECT 166.870 52.985 167.445 53.470 ;
        RECT 169.920 53.450 170.455 53.505 ;
        RECT 163.880 52.900 164.415 52.955 ;
        RECT 166.890 52.930 167.425 52.985 ;
        RECT 169.900 52.965 170.475 53.450 ;
        RECT 169.920 52.910 170.455 52.965 ;
        RECT 148.775 49.670 149.310 49.725 ;
        RECT 151.805 49.690 152.340 49.745 ;
        RECT 148.755 49.185 149.330 49.670 ;
        RECT 151.785 49.205 152.360 49.690 ;
        RECT 154.815 49.660 155.350 49.715 ;
        RECT 157.845 49.680 158.380 49.735 ;
        RECT 148.775 49.130 149.310 49.185 ;
        RECT 151.805 49.150 152.340 49.205 ;
        RECT 154.795 49.175 155.370 49.660 ;
        RECT 157.825 49.195 158.400 49.680 ;
        RECT 160.815 49.660 161.350 49.715 ;
        RECT 154.815 49.120 155.350 49.175 ;
        RECT 157.845 49.140 158.380 49.195 ;
        RECT 160.795 49.175 161.370 49.660 ;
        RECT 163.855 49.655 164.390 49.710 ;
        RECT 160.815 49.120 161.350 49.175 ;
        RECT 163.835 49.170 164.410 49.655 ;
        RECT 166.855 49.650 167.390 49.705 ;
        RECT 169.885 49.670 170.420 49.725 ;
        RECT 163.855 49.115 164.390 49.170 ;
        RECT 166.835 49.165 167.410 49.650 ;
        RECT 169.865 49.185 170.440 49.670 ;
        RECT 166.855 49.110 167.390 49.165 ;
        RECT 169.885 49.130 170.420 49.185 ;
        RECT 148.760 45.770 149.310 45.825 ;
        RECT 151.790 45.790 152.340 45.845 ;
        RECT 148.740 45.270 149.330 45.770 ;
        RECT 151.770 45.290 152.360 45.790 ;
        RECT 154.800 45.760 155.350 45.815 ;
        RECT 157.830 45.780 158.380 45.835 ;
        RECT 148.760 45.215 149.310 45.270 ;
        RECT 151.790 45.235 152.340 45.290 ;
        RECT 154.780 45.260 155.370 45.760 ;
        RECT 157.810 45.280 158.400 45.780 ;
        RECT 160.800 45.760 161.350 45.815 ;
        RECT 154.800 45.205 155.350 45.260 ;
        RECT 157.830 45.225 158.380 45.280 ;
        RECT 160.780 45.260 161.370 45.760 ;
        RECT 163.840 45.755 164.390 45.810 ;
        RECT 160.800 45.205 161.350 45.260 ;
        RECT 163.820 45.255 164.410 45.755 ;
        RECT 166.840 45.750 167.390 45.805 ;
        RECT 169.870 45.770 170.420 45.825 ;
        RECT 163.840 45.200 164.390 45.255 ;
        RECT 166.820 45.250 167.410 45.750 ;
        RECT 169.850 45.270 170.440 45.770 ;
        RECT 166.840 45.195 167.390 45.250 ;
        RECT 169.870 45.215 170.420 45.270 ;
        RECT 148.730 43.110 149.050 43.115 ;
        RECT 146.560 42.855 149.050 43.110 ;
        RECT 148.740 41.730 149.060 41.745 ;
        RECT 146.090 41.495 149.060 41.730 ;
        RECT 148.740 41.485 149.060 41.495 ;
        RECT 148.760 40.330 149.080 40.350 ;
        RECT 145.705 40.110 149.080 40.330 ;
        RECT 148.760 40.090 149.080 40.110 ;
        RECT 148.760 38.990 149.080 38.995 ;
        RECT 145.310 38.735 149.080 38.990 ;
        RECT 148.735 37.595 149.055 37.605 ;
        RECT 144.905 37.355 149.055 37.595 ;
        RECT 148.735 37.345 149.055 37.355 ;
        RECT 148.730 36.225 149.050 36.235 ;
        RECT 144.425 35.985 149.050 36.225 ;
        RECT 148.730 35.975 149.050 35.985 ;
        RECT 148.765 34.835 149.085 34.845 ;
        RECT 143.885 34.595 149.085 34.835 ;
        RECT 148.765 34.585 149.085 34.595 ;
        RECT 148.750 33.470 149.070 33.495 ;
        RECT 143.150 33.255 149.070 33.470 ;
        RECT 148.750 33.235 149.070 33.255 ;
        RECT 138.775 32.645 143.435 32.960 ;
        RECT 143.170 32.085 143.380 32.645 ;
        RECT 148.760 32.085 149.080 32.110 ;
        RECT 143.170 31.875 149.080 32.085 ;
        RECT 148.760 31.850 149.080 31.875 ;
      LAYER via2 ;
        RECT 138.750 84.965 139.120 85.335 ;
        RECT 138.710 81.965 139.080 82.335 ;
        RECT 136.635 78.005 136.990 78.360 ;
        RECT 132.700 74.975 133.070 75.345 ;
        RECT 128.605 71.880 128.975 72.250 ;
        RECT 136.635 71.980 136.990 72.355 ;
        RECT 22.785 71.500 23.085 71.800 ;
        RECT 120.770 68.955 121.085 69.270 ;
        RECT 74.510 64.155 74.905 64.550 ;
        RECT 78.665 64.170 78.995 64.500 ;
        RECT 148.670 74.210 149.170 74.710 ;
        RECT 151.700 74.190 152.200 74.690 ;
        RECT 154.710 74.220 155.210 74.720 ;
        RECT 157.740 74.200 158.240 74.700 ;
        RECT 160.710 74.220 161.210 74.720 ;
        RECT 163.750 74.225 164.250 74.725 ;
        RECT 166.750 74.230 167.250 74.730 ;
        RECT 169.780 74.210 170.280 74.710 ;
        RECT 148.685 70.310 149.170 70.795 ;
        RECT 151.715 70.290 152.200 70.775 ;
        RECT 154.725 70.320 155.210 70.805 ;
        RECT 157.755 70.300 158.240 70.785 ;
        RECT 160.725 70.320 161.210 70.805 ;
        RECT 163.765 70.325 164.250 70.810 ;
        RECT 166.765 70.330 167.250 70.815 ;
        RECT 169.795 70.310 170.280 70.795 ;
        RECT 148.720 66.530 149.205 67.015 ;
        RECT 151.750 66.550 152.235 67.035 ;
        RECT 154.760 66.520 155.245 67.005 ;
        RECT 157.790 66.540 158.275 67.025 ;
        RECT 160.760 66.520 161.245 67.005 ;
        RECT 148.705 62.615 149.205 63.115 ;
        RECT 151.735 62.635 152.235 63.135 ;
        RECT 154.745 62.605 155.245 63.105 ;
        RECT 157.775 62.625 158.275 63.125 ;
        RECT 160.745 62.605 161.245 63.105 ;
        RECT 163.790 66.540 164.275 67.025 ;
        RECT 166.800 66.510 167.285 66.995 ;
        RECT 169.830 66.530 170.315 67.015 ;
        RECT 163.775 62.625 164.275 63.125 ;
        RECT 166.785 62.595 167.285 63.095 ;
        RECT 169.815 62.615 170.315 63.115 ;
        RECT 152.045 61.930 152.325 62.210 ;
        RECT 156.245 59.400 156.525 59.680 ;
        RECT 148.820 56.865 149.320 57.365 ;
        RECT 151.850 56.845 152.350 57.345 ;
        RECT 154.860 56.875 155.360 57.375 ;
        RECT 157.890 56.855 158.390 57.355 ;
        RECT 160.860 56.875 161.360 57.375 ;
        RECT 74.510 55.300 74.905 55.695 ;
        RECT 78.665 55.350 78.995 55.680 ;
        RECT 120.770 50.580 121.085 50.895 ;
        RECT 22.785 48.050 23.085 48.350 ;
        RECT 128.605 47.600 128.975 47.970 ;
        RECT 136.635 47.495 136.990 47.870 ;
        RECT 132.700 44.505 133.070 44.875 ;
        RECT 136.635 41.490 136.990 41.845 ;
        RECT 138.710 37.515 139.080 37.885 ;
        RECT 138.750 34.515 139.120 34.885 ;
        RECT 163.890 56.855 164.390 57.355 ;
        RECT 166.900 56.885 167.400 57.385 ;
        RECT 169.930 56.865 170.430 57.365 ;
        RECT 148.835 52.965 149.320 53.450 ;
        RECT 151.865 52.945 152.350 53.430 ;
        RECT 154.875 52.975 155.360 53.460 ;
        RECT 157.905 52.955 158.390 53.440 ;
        RECT 160.875 52.975 161.360 53.460 ;
        RECT 163.905 52.955 164.390 53.440 ;
        RECT 166.915 52.985 167.400 53.470 ;
        RECT 169.945 52.965 170.430 53.450 ;
        RECT 148.800 49.185 149.285 49.670 ;
        RECT 151.830 49.205 152.315 49.690 ;
        RECT 154.840 49.175 155.325 49.660 ;
        RECT 157.870 49.195 158.355 49.680 ;
        RECT 160.840 49.175 161.325 49.660 ;
        RECT 163.880 49.170 164.365 49.655 ;
        RECT 166.880 49.165 167.365 49.650 ;
        RECT 169.910 49.185 170.395 49.670 ;
        RECT 148.785 45.270 149.285 45.770 ;
        RECT 151.815 45.290 152.315 45.790 ;
        RECT 154.825 45.260 155.325 45.760 ;
        RECT 157.855 45.280 158.355 45.780 ;
        RECT 160.825 45.260 161.325 45.760 ;
        RECT 163.865 45.255 164.365 45.755 ;
        RECT 166.865 45.250 167.365 45.750 ;
        RECT 169.895 45.270 170.395 45.770 ;
      LAYER met3 ;
        RECT 7.685 87.430 10.115 89.830 ;
        RECT 11.685 87.430 14.115 89.830 ;
        RECT 15.685 87.430 18.115 89.830 ;
        RECT 19.685 87.430 22.115 89.830 ;
        RECT 23.685 87.430 26.115 89.830 ;
        RECT 27.685 87.430 30.115 89.830 ;
        RECT 31.685 87.430 34.115 89.830 ;
        RECT 35.685 87.430 38.115 89.830 ;
        RECT 39.685 87.430 42.115 89.830 ;
        RECT 43.685 87.430 46.115 89.830 ;
        RECT 47.685 87.430 50.115 89.830 ;
        RECT 51.685 87.430 54.115 89.830 ;
        RECT 55.685 87.430 58.115 89.830 ;
        RECT 59.685 87.430 62.115 89.830 ;
        RECT 63.685 87.430 66.115 89.830 ;
        RECT 67.685 87.430 70.115 89.830 ;
        RECT 71.685 87.430 74.115 89.830 ;
        RECT 75.685 87.430 78.115 89.830 ;
        RECT 79.685 87.430 82.115 89.830 ;
        RECT 83.685 87.430 86.115 89.830 ;
        RECT 87.685 87.430 90.115 89.830 ;
        RECT 91.685 87.430 94.115 89.830 ;
        RECT 95.685 87.430 98.115 89.830 ;
        RECT 99.685 87.430 102.115 89.830 ;
        RECT 103.685 87.430 106.115 89.830 ;
        RECT 107.685 87.430 110.115 89.830 ;
        RECT 111.685 87.430 114.115 89.830 ;
        RECT 115.685 87.430 118.115 89.830 ;
        RECT 119.685 87.430 122.115 89.830 ;
        RECT 123.685 87.430 126.115 89.830 ;
        RECT 127.685 87.430 130.115 89.830 ;
        RECT 131.685 87.430 134.115 89.830 ;
        RECT 135.685 87.430 138.115 89.830 ;
        RECT 139.685 87.430 142.115 89.830 ;
        RECT 7.685 84.430 10.115 86.830 ;
        RECT 11.685 85.645 14.115 86.830 ;
        RECT 15.685 85.645 18.115 86.830 ;
        RECT 19.685 85.645 22.115 86.830 ;
        RECT 23.685 85.645 26.115 86.830 ;
        RECT 27.685 85.645 30.115 86.830 ;
        RECT 31.685 85.645 34.115 86.830 ;
        RECT 35.685 85.645 38.115 86.830 ;
        RECT 39.685 85.645 42.115 86.830 ;
        RECT 43.685 85.645 46.115 86.830 ;
        RECT 47.685 85.645 50.115 86.830 ;
        RECT 51.685 85.645 54.115 86.830 ;
        RECT 55.685 85.645 58.115 86.830 ;
        RECT 59.685 85.645 62.115 86.830 ;
        RECT 63.685 85.645 66.115 86.830 ;
        RECT 67.685 85.645 70.115 86.830 ;
        RECT 71.685 85.645 74.115 86.830 ;
        RECT 11.685 85.200 74.115 85.645 ;
        RECT 11.685 84.430 14.115 85.200 ;
        RECT 15.685 84.430 18.115 85.200 ;
        RECT 19.685 84.430 22.115 85.200 ;
        RECT 23.685 84.430 26.115 85.200 ;
        RECT 27.685 84.430 30.115 85.200 ;
        RECT 31.685 84.430 34.115 85.200 ;
        RECT 35.685 84.430 38.115 85.200 ;
        RECT 39.685 84.430 42.115 85.200 ;
        RECT 43.685 84.430 46.115 85.200 ;
        RECT 47.685 84.430 50.115 85.200 ;
        RECT 51.685 84.430 54.115 85.200 ;
        RECT 55.685 84.430 58.115 85.200 ;
        RECT 59.685 84.430 62.115 85.200 ;
        RECT 63.685 84.430 66.115 85.200 ;
        RECT 67.685 84.430 70.115 85.200 ;
        RECT 71.685 84.430 74.115 85.200 ;
        RECT 75.685 85.645 78.115 86.830 ;
        RECT 79.685 85.645 82.115 86.830 ;
        RECT 75.685 85.265 82.115 85.645 ;
        RECT 75.685 84.430 78.115 85.265 ;
        RECT 79.685 84.430 82.115 85.265 ;
        RECT 83.685 85.565 86.115 86.830 ;
        RECT 87.685 85.565 90.115 86.830 ;
        RECT 83.685 85.185 90.115 85.565 ;
        RECT 83.685 84.430 86.115 85.185 ;
        RECT 87.685 84.430 90.115 85.185 ;
        RECT 91.685 85.480 94.115 86.830 ;
        RECT 95.685 85.480 98.115 86.830 ;
        RECT 91.685 85.100 98.115 85.480 ;
        RECT 91.685 84.430 94.115 85.100 ;
        RECT 95.685 84.430 98.115 85.100 ;
        RECT 99.685 85.645 102.115 86.830 ;
        RECT 103.685 85.645 106.115 86.830 ;
        RECT 99.685 85.265 106.115 85.645 ;
        RECT 99.685 84.430 102.115 85.265 ;
        RECT 103.685 84.430 106.115 85.265 ;
        RECT 107.685 85.775 110.115 86.830 ;
        RECT 111.685 85.775 114.115 86.830 ;
        RECT 107.685 85.460 114.115 85.775 ;
        RECT 107.685 84.430 110.115 85.460 ;
        RECT 111.685 84.430 114.115 85.460 ;
        RECT 115.685 85.775 118.115 86.830 ;
        RECT 119.685 85.775 122.115 86.830 ;
        RECT 115.685 85.460 122.115 85.775 ;
        RECT 115.685 84.430 118.115 85.460 ;
        RECT 119.685 84.430 122.115 85.460 ;
        RECT 123.685 85.625 126.115 86.830 ;
        RECT 127.685 85.625 130.115 86.830 ;
        RECT 123.685 85.205 130.115 85.625 ;
        RECT 123.685 84.430 126.115 85.205 ;
        RECT 127.685 84.430 130.115 85.205 ;
        RECT 131.685 84.430 134.115 86.830 ;
        RECT 135.685 85.360 138.115 86.830 ;
        RECT 135.685 84.940 139.145 85.360 ;
        RECT 135.685 84.430 138.115 84.940 ;
        RECT 139.685 84.430 142.115 86.830 ;
        RECT 12.330 83.830 12.775 84.430 ;
        RECT 76.540 83.830 76.920 84.430 ;
        RECT 80.490 83.830 80.870 84.430 ;
        RECT 84.605 83.830 84.985 84.430 ;
        RECT 88.555 83.830 88.935 84.430 ;
        RECT 92.505 83.830 92.885 84.430 ;
        RECT 96.695 83.830 97.075 84.430 ;
        RECT 100.565 83.830 100.945 84.430 ;
        RECT 104.555 83.830 104.935 84.430 ;
        RECT 108.560 83.830 108.875 84.430 ;
        RECT 112.720 83.830 113.035 84.430 ;
        RECT 116.565 83.830 116.880 84.430 ;
        RECT 120.770 83.830 121.085 84.430 ;
        RECT 124.685 83.830 125.105 84.430 ;
        RECT 128.580 83.830 129.000 84.430 ;
        RECT 132.675 83.830 133.095 84.430 ;
        RECT 7.685 81.430 10.115 83.830 ;
        RECT 11.685 82.520 14.115 83.830 ;
        RECT 15.685 82.520 18.115 83.830 ;
        RECT 19.685 82.520 22.115 83.830 ;
        RECT 23.685 82.520 26.115 83.830 ;
        RECT 27.685 82.520 30.115 83.830 ;
        RECT 31.685 82.520 34.115 83.830 ;
        RECT 35.685 82.520 38.115 83.830 ;
        RECT 39.685 82.520 42.115 83.830 ;
        RECT 43.685 82.520 46.115 83.830 ;
        RECT 47.685 82.520 50.115 83.830 ;
        RECT 51.685 82.520 54.115 83.830 ;
        RECT 55.685 82.520 58.115 83.830 ;
        RECT 59.685 82.520 62.115 83.830 ;
        RECT 63.685 82.520 66.115 83.830 ;
        RECT 67.685 82.520 70.115 83.830 ;
        RECT 71.685 82.520 74.115 83.830 ;
        RECT 11.685 82.075 74.115 82.520 ;
        RECT 11.685 81.430 14.115 82.075 ;
        RECT 15.685 81.430 18.115 82.075 ;
        RECT 19.685 81.430 22.115 82.075 ;
        RECT 23.685 81.430 26.115 82.075 ;
        RECT 27.685 81.430 30.115 82.075 ;
        RECT 31.685 81.430 34.115 82.075 ;
        RECT 35.685 81.430 38.115 82.075 ;
        RECT 39.685 81.430 42.115 82.075 ;
        RECT 43.685 81.430 46.115 82.075 ;
        RECT 47.685 81.430 50.115 82.075 ;
        RECT 51.685 81.430 54.115 82.075 ;
        RECT 55.685 81.430 58.115 82.075 ;
        RECT 59.685 81.430 62.115 82.075 ;
        RECT 63.685 81.430 66.115 82.075 ;
        RECT 67.685 81.430 70.115 82.075 ;
        RECT 71.685 81.430 74.115 82.075 ;
        RECT 75.685 81.430 78.115 83.830 ;
        RECT 79.685 81.430 82.115 83.830 ;
        RECT 83.685 81.430 86.115 83.830 ;
        RECT 87.685 81.430 90.115 83.830 ;
        RECT 91.685 81.430 94.115 83.830 ;
        RECT 95.685 81.430 98.115 83.830 ;
        RECT 99.685 81.430 102.115 83.830 ;
        RECT 103.685 81.430 106.115 83.830 ;
        RECT 107.685 81.430 110.115 83.830 ;
        RECT 111.685 81.430 114.115 83.830 ;
        RECT 115.685 81.430 118.115 83.830 ;
        RECT 119.685 81.430 122.115 83.830 ;
        RECT 123.685 81.430 126.115 83.830 ;
        RECT 127.685 81.430 130.115 83.830 ;
        RECT 131.685 81.430 134.115 83.830 ;
        RECT 135.685 82.360 138.115 83.830 ;
        RECT 135.685 81.940 139.105 82.360 ;
        RECT 135.685 81.430 138.115 81.940 ;
        RECT 139.685 81.430 142.115 83.830 ;
        RECT 72.485 80.830 72.930 81.430 ;
        RECT 76.540 80.830 76.920 81.430 ;
        RECT 80.490 80.830 80.870 81.430 ;
        RECT 84.605 80.830 84.985 81.430 ;
        RECT 88.555 80.830 88.935 81.430 ;
        RECT 92.505 80.830 92.885 81.430 ;
        RECT 96.695 80.830 97.075 81.430 ;
        RECT 100.565 80.830 100.945 81.430 ;
        RECT 104.555 80.830 104.935 81.430 ;
        RECT 108.560 80.830 108.875 81.430 ;
        RECT 112.720 80.830 113.035 81.430 ;
        RECT 116.565 80.830 116.880 81.430 ;
        RECT 120.770 80.830 121.085 81.430 ;
        RECT 124.685 80.830 125.105 81.430 ;
        RECT 128.580 80.830 129.000 81.430 ;
        RECT 132.675 80.830 133.095 81.430 ;
        RECT 7.685 78.430 10.115 80.830 ;
        RECT 11.685 79.890 14.115 80.830 ;
        RECT 15.685 79.890 18.115 80.830 ;
        RECT 19.685 79.890 22.115 80.830 ;
        RECT 23.685 79.890 26.115 80.830 ;
        RECT 27.685 79.890 30.115 80.830 ;
        RECT 31.685 79.890 34.115 80.830 ;
        RECT 35.685 79.890 38.115 80.830 ;
        RECT 39.685 79.890 42.115 80.830 ;
        RECT 43.685 79.890 46.115 80.830 ;
        RECT 47.685 79.890 50.115 80.830 ;
        RECT 51.685 79.890 54.115 80.830 ;
        RECT 55.685 79.890 58.115 80.830 ;
        RECT 59.685 79.890 62.115 80.830 ;
        RECT 63.685 79.890 66.115 80.830 ;
        RECT 67.685 79.890 70.115 80.830 ;
        RECT 71.685 79.890 74.115 80.830 ;
        RECT 11.685 79.445 74.115 79.890 ;
        RECT 11.685 78.430 14.115 79.445 ;
        RECT 15.685 78.430 18.115 79.445 ;
        RECT 19.685 78.430 22.115 79.445 ;
        RECT 23.685 78.430 26.115 79.445 ;
        RECT 27.685 78.430 30.115 79.445 ;
        RECT 31.685 78.430 34.115 79.445 ;
        RECT 35.685 78.430 38.115 79.445 ;
        RECT 39.685 78.430 42.115 79.445 ;
        RECT 43.685 78.430 46.115 79.445 ;
        RECT 47.685 78.430 50.115 79.445 ;
        RECT 51.685 78.430 54.115 79.445 ;
        RECT 55.685 78.430 58.115 79.445 ;
        RECT 59.685 78.430 62.115 79.445 ;
        RECT 63.685 78.430 66.115 79.445 ;
        RECT 67.685 78.430 70.115 79.445 ;
        RECT 71.685 78.430 74.115 79.445 ;
        RECT 75.685 78.430 78.115 80.830 ;
        RECT 79.685 78.430 82.115 80.830 ;
        RECT 83.685 78.430 86.115 80.830 ;
        RECT 87.685 78.430 90.115 80.830 ;
        RECT 91.685 78.430 94.115 80.830 ;
        RECT 95.685 78.430 98.115 80.830 ;
        RECT 99.685 78.430 102.115 80.830 ;
        RECT 103.685 78.430 106.115 80.830 ;
        RECT 107.685 78.430 110.115 80.830 ;
        RECT 111.685 78.430 114.115 80.830 ;
        RECT 115.685 78.430 118.115 80.830 ;
        RECT 119.685 78.430 122.115 80.830 ;
        RECT 123.685 78.430 126.115 80.830 ;
        RECT 127.685 78.430 130.115 80.830 ;
        RECT 131.685 78.430 134.115 80.830 ;
        RECT 135.685 78.430 138.115 80.830 ;
        RECT 139.685 78.430 142.115 80.830 ;
        RECT 12.495 77.830 12.940 78.430 ;
        RECT 76.540 77.830 76.920 78.430 ;
        RECT 80.490 77.830 80.870 78.430 ;
        RECT 84.605 77.830 84.985 78.430 ;
        RECT 88.555 77.830 88.935 78.430 ;
        RECT 92.505 77.830 92.885 78.430 ;
        RECT 96.695 77.830 97.075 78.430 ;
        RECT 100.565 77.830 100.945 78.430 ;
        RECT 104.555 77.830 104.935 78.430 ;
        RECT 108.560 77.830 108.875 78.430 ;
        RECT 112.720 77.830 113.035 78.430 ;
        RECT 116.565 77.830 116.880 78.430 ;
        RECT 120.770 77.830 121.085 78.430 ;
        RECT 124.685 77.830 125.105 78.430 ;
        RECT 128.580 77.830 129.000 78.430 ;
        RECT 132.675 77.830 133.095 78.430 ;
        RECT 136.610 77.830 137.015 78.430 ;
        RECT 7.685 75.430 10.115 77.830 ;
        RECT 11.685 76.935 14.115 77.830 ;
        RECT 15.685 76.935 18.115 77.830 ;
        RECT 19.685 76.935 22.115 77.830 ;
        RECT 23.685 76.935 26.115 77.830 ;
        RECT 27.685 76.935 30.115 77.830 ;
        RECT 31.685 76.935 34.115 77.830 ;
        RECT 35.685 76.935 38.115 77.830 ;
        RECT 39.685 76.935 42.115 77.830 ;
        RECT 43.685 76.935 46.115 77.830 ;
        RECT 47.685 76.935 50.115 77.830 ;
        RECT 51.685 76.935 54.115 77.830 ;
        RECT 55.685 76.935 58.115 77.830 ;
        RECT 59.685 76.935 62.115 77.830 ;
        RECT 63.685 76.935 66.115 77.830 ;
        RECT 67.685 76.935 70.115 77.830 ;
        RECT 71.685 76.935 74.115 77.830 ;
        RECT 11.685 76.490 74.115 76.935 ;
        RECT 11.685 75.430 14.115 76.490 ;
        RECT 15.685 75.430 18.115 76.490 ;
        RECT 19.685 75.430 22.115 76.490 ;
        RECT 23.685 75.430 26.115 76.490 ;
        RECT 27.685 75.430 30.115 76.490 ;
        RECT 31.685 75.430 34.115 76.490 ;
        RECT 35.685 75.430 38.115 76.490 ;
        RECT 39.685 75.430 42.115 76.490 ;
        RECT 43.685 75.430 46.115 76.490 ;
        RECT 47.685 75.430 50.115 76.490 ;
        RECT 51.685 75.430 54.115 76.490 ;
        RECT 55.685 75.430 58.115 76.490 ;
        RECT 59.685 75.430 62.115 76.490 ;
        RECT 63.685 75.430 66.115 76.490 ;
        RECT 67.685 75.430 70.115 76.490 ;
        RECT 71.685 75.430 74.115 76.490 ;
        RECT 75.685 75.430 78.115 77.830 ;
        RECT 79.685 75.430 82.115 77.830 ;
        RECT 83.685 75.430 86.115 77.830 ;
        RECT 87.685 75.430 90.115 77.830 ;
        RECT 91.685 75.430 94.115 77.830 ;
        RECT 95.685 75.430 98.115 77.830 ;
        RECT 99.685 75.430 102.115 77.830 ;
        RECT 103.685 75.430 106.115 77.830 ;
        RECT 107.685 75.430 110.115 77.830 ;
        RECT 111.685 75.430 114.115 77.830 ;
        RECT 115.685 75.430 118.115 77.830 ;
        RECT 119.685 75.430 122.115 77.830 ;
        RECT 123.685 75.430 126.115 77.830 ;
        RECT 127.685 75.430 130.115 77.830 ;
        RECT 131.685 75.430 134.115 77.830 ;
        RECT 135.685 75.430 138.115 77.830 ;
        RECT 139.685 75.430 142.115 77.830 ;
        RECT 72.565 74.830 73.010 75.430 ;
        RECT 76.540 74.830 76.920 75.430 ;
        RECT 80.490 74.830 80.870 75.430 ;
        RECT 84.605 74.830 84.985 75.430 ;
        RECT 88.555 74.830 88.935 75.430 ;
        RECT 92.505 74.830 92.885 75.430 ;
        RECT 96.695 74.830 97.075 75.430 ;
        RECT 100.565 74.830 100.945 75.430 ;
        RECT 104.555 74.830 104.935 75.430 ;
        RECT 108.560 74.830 108.875 75.430 ;
        RECT 112.720 74.830 113.035 75.430 ;
        RECT 116.565 74.830 116.880 75.430 ;
        RECT 120.770 74.830 121.085 75.430 ;
        RECT 124.685 74.830 125.105 75.430 ;
        RECT 128.580 74.830 129.000 75.430 ;
        RECT 132.675 74.830 133.095 75.430 ;
        RECT 7.685 72.430 10.115 74.830 ;
        RECT 11.685 73.890 14.115 74.830 ;
        RECT 15.685 73.890 18.115 74.830 ;
        RECT 19.685 73.890 22.115 74.830 ;
        RECT 23.685 73.890 26.115 74.830 ;
        RECT 27.685 73.890 30.115 74.830 ;
        RECT 31.685 73.890 34.115 74.830 ;
        RECT 35.685 73.890 38.115 74.830 ;
        RECT 39.685 73.890 42.115 74.830 ;
        RECT 43.685 73.890 46.115 74.830 ;
        RECT 47.685 73.890 50.115 74.830 ;
        RECT 51.685 73.890 54.115 74.830 ;
        RECT 55.685 73.890 58.115 74.830 ;
        RECT 59.685 73.890 62.115 74.830 ;
        RECT 63.685 73.890 66.115 74.830 ;
        RECT 67.685 73.890 70.115 74.830 ;
        RECT 71.685 73.890 74.115 74.830 ;
        RECT 11.685 73.445 74.115 73.890 ;
        RECT 11.685 72.430 14.115 73.445 ;
        RECT 15.685 72.430 18.115 73.445 ;
        RECT 19.685 72.430 22.115 73.445 ;
        RECT 23.685 72.430 26.115 73.445 ;
        RECT 27.685 72.430 30.115 73.445 ;
        RECT 31.685 72.430 34.115 73.445 ;
        RECT 35.685 72.430 38.115 73.445 ;
        RECT 39.685 72.430 42.115 73.445 ;
        RECT 43.685 72.430 46.115 73.445 ;
        RECT 47.685 72.430 50.115 73.445 ;
        RECT 51.685 72.430 54.115 73.445 ;
        RECT 55.685 72.430 58.115 73.445 ;
        RECT 59.685 72.430 62.115 73.445 ;
        RECT 63.685 72.430 66.115 73.445 ;
        RECT 67.685 72.430 70.115 73.445 ;
        RECT 71.685 72.430 74.115 73.445 ;
        RECT 75.685 72.430 78.115 74.830 ;
        RECT 79.685 72.430 82.115 74.830 ;
        RECT 83.685 72.430 86.115 74.830 ;
        RECT 87.685 72.430 90.115 74.830 ;
        RECT 91.685 72.430 94.115 74.830 ;
        RECT 95.685 72.430 98.115 74.830 ;
        RECT 99.685 72.430 102.115 74.830 ;
        RECT 103.685 72.430 106.115 74.830 ;
        RECT 107.685 72.430 110.115 74.830 ;
        RECT 111.685 72.430 114.115 74.830 ;
        RECT 115.685 72.430 118.115 74.830 ;
        RECT 119.685 72.430 122.115 74.830 ;
        RECT 123.685 72.430 126.115 74.830 ;
        RECT 127.685 72.430 130.115 74.830 ;
        RECT 131.685 72.430 134.115 74.830 ;
        RECT 135.685 72.430 138.115 74.830 ;
        RECT 139.685 72.430 142.115 74.830 ;
        RECT 166.725 74.750 167.275 74.755 ;
        RECT 163.725 74.745 164.275 74.750 ;
        RECT 154.685 74.740 155.235 74.745 ;
        RECT 160.685 74.740 161.235 74.745 ;
        RECT 148.645 74.730 149.195 74.735 ;
        RECT 148.620 74.190 149.220 74.730 ;
        RECT 151.675 74.710 152.225 74.715 ;
        RECT 148.645 74.185 149.195 74.190 ;
        RECT 151.650 74.170 152.250 74.710 ;
        RECT 154.660 74.200 155.260 74.740 ;
        RECT 157.715 74.720 158.265 74.725 ;
        RECT 154.685 74.195 155.235 74.200 ;
        RECT 157.690 74.180 158.290 74.720 ;
        RECT 160.660 74.200 161.260 74.740 ;
        RECT 163.700 74.205 164.300 74.745 ;
        RECT 166.700 74.210 167.300 74.750 ;
        RECT 169.755 74.730 170.305 74.735 ;
        RECT 166.725 74.205 167.275 74.210 ;
        RECT 163.725 74.200 164.275 74.205 ;
        RECT 160.685 74.195 161.235 74.200 ;
        RECT 169.730 74.190 170.330 74.730 ;
        RECT 169.755 74.185 170.305 74.190 ;
        RECT 157.715 74.175 158.265 74.180 ;
        RECT 151.675 74.165 152.225 74.170 ;
        RECT 12.410 71.830 12.855 72.430 ;
        RECT 7.685 69.430 10.115 71.830 ;
        RECT 11.685 70.605 14.115 71.830 ;
        RECT 15.685 70.605 18.115 71.830 ;
        RECT 19.685 70.605 22.115 71.830 ;
        RECT 22.675 71.400 23.175 71.920 ;
        RECT 76.540 71.830 76.920 72.430 ;
        RECT 80.490 71.830 80.870 72.430 ;
        RECT 84.605 71.830 84.985 72.430 ;
        RECT 88.555 71.830 88.935 72.430 ;
        RECT 92.505 71.830 92.885 72.430 ;
        RECT 96.695 71.830 97.075 72.430 ;
        RECT 100.565 71.830 100.945 72.430 ;
        RECT 104.555 71.830 104.935 72.430 ;
        RECT 108.560 71.830 108.875 72.430 ;
        RECT 112.720 71.830 113.035 72.430 ;
        RECT 116.565 71.830 116.880 72.430 ;
        RECT 120.770 71.830 121.085 72.430 ;
        RECT 124.685 71.830 125.105 72.430 ;
        RECT 128.580 71.830 129.000 72.430 ;
        RECT 132.675 71.830 133.095 72.430 ;
        RECT 136.610 71.830 137.015 72.430 ;
        RECT 23.685 70.605 26.115 71.830 ;
        RECT 27.685 70.605 30.115 71.830 ;
        RECT 31.685 70.605 34.115 71.830 ;
        RECT 35.685 70.605 38.115 71.830 ;
        RECT 39.685 70.605 42.115 71.830 ;
        RECT 43.685 70.605 46.115 71.830 ;
        RECT 47.685 70.605 50.115 71.830 ;
        RECT 51.685 70.605 54.115 71.830 ;
        RECT 55.685 70.605 58.115 71.830 ;
        RECT 59.685 70.605 62.115 71.830 ;
        RECT 63.685 70.605 66.115 71.830 ;
        RECT 67.685 70.605 70.115 71.830 ;
        RECT 71.685 70.605 74.115 71.830 ;
        RECT 11.685 70.160 74.115 70.605 ;
        RECT 11.685 69.430 14.115 70.160 ;
        RECT 15.685 69.430 18.115 70.160 ;
        RECT 19.685 69.430 22.115 70.160 ;
        RECT 23.685 69.430 26.115 70.160 ;
        RECT 27.685 69.430 30.115 70.160 ;
        RECT 31.685 69.430 34.115 70.160 ;
        RECT 35.685 69.430 38.115 70.160 ;
        RECT 39.685 69.430 42.115 70.160 ;
        RECT 43.685 69.430 46.115 70.160 ;
        RECT 47.685 69.430 50.115 70.160 ;
        RECT 51.685 69.430 54.115 70.160 ;
        RECT 55.685 69.430 58.115 70.160 ;
        RECT 59.685 69.430 62.115 70.160 ;
        RECT 63.685 69.430 66.115 70.160 ;
        RECT 67.685 69.430 70.115 70.160 ;
        RECT 71.685 69.430 74.115 70.160 ;
        RECT 75.685 69.430 78.115 71.830 ;
        RECT 79.685 69.430 82.115 71.830 ;
        RECT 83.685 69.430 86.115 71.830 ;
        RECT 87.685 69.430 90.115 71.830 ;
        RECT 91.685 69.430 94.115 71.830 ;
        RECT 95.685 69.430 98.115 71.830 ;
        RECT 99.685 69.430 102.115 71.830 ;
        RECT 103.685 69.430 106.115 71.830 ;
        RECT 107.685 69.430 110.115 71.830 ;
        RECT 111.685 69.430 114.115 71.830 ;
        RECT 115.685 69.430 118.115 71.830 ;
        RECT 119.685 69.430 122.115 71.830 ;
        RECT 123.685 69.430 126.115 71.830 ;
        RECT 127.685 69.430 130.115 71.830 ;
        RECT 131.685 69.430 134.115 71.830 ;
        RECT 135.685 69.430 138.115 71.830 ;
        RECT 139.685 69.430 142.115 71.830 ;
        RECT 147.735 71.260 150.135 73.660 ;
        RECT 148.660 70.285 149.195 71.260 ;
        RECT 150.765 71.240 153.165 73.640 ;
        RECT 153.775 71.270 156.175 73.670 ;
        RECT 151.690 70.265 152.225 71.240 ;
        RECT 154.700 70.295 155.235 71.270 ;
        RECT 156.805 71.250 159.205 73.650 ;
        RECT 159.775 71.270 162.175 73.670 ;
        RECT 162.815 71.275 165.215 73.675 ;
        RECT 165.815 71.280 168.215 73.680 ;
        RECT 157.730 70.275 158.265 71.250 ;
        RECT 160.700 70.295 161.235 71.270 ;
        RECT 163.740 70.300 164.275 71.275 ;
        RECT 166.740 70.305 167.275 71.280 ;
        RECT 168.845 71.260 171.245 73.660 ;
        RECT 169.770 70.285 170.305 71.260 ;
        RECT 72.730 68.830 73.175 69.430 ;
        RECT 76.540 68.830 76.920 69.430 ;
        RECT 80.490 68.830 80.870 69.430 ;
        RECT 84.605 68.830 84.985 69.430 ;
        RECT 88.555 68.830 88.935 69.430 ;
        RECT 92.505 68.830 92.885 69.430 ;
        RECT 96.695 68.830 97.075 69.430 ;
        RECT 100.565 68.830 100.945 69.430 ;
        RECT 104.555 68.830 104.935 69.430 ;
        RECT 108.560 68.830 108.875 69.430 ;
        RECT 112.720 68.830 113.035 69.430 ;
        RECT 116.565 68.830 116.880 69.430 ;
        RECT 120.445 68.830 121.420 69.430 ;
        RECT 124.685 68.830 125.105 69.430 ;
        RECT 128.580 68.830 129.000 69.430 ;
        RECT 132.675 68.830 133.095 69.430 ;
        RECT 136.610 68.830 137.015 69.430 ;
        RECT 7.685 66.430 10.115 68.830 ;
        RECT 11.685 67.645 14.115 68.830 ;
        RECT 15.685 67.645 18.115 68.830 ;
        RECT 19.685 67.645 22.115 68.830 ;
        RECT 23.685 67.645 26.115 68.830 ;
        RECT 27.685 67.645 30.115 68.830 ;
        RECT 31.685 67.645 34.115 68.830 ;
        RECT 35.685 67.645 38.115 68.830 ;
        RECT 39.685 67.645 42.115 68.830 ;
        RECT 43.685 67.645 46.115 68.830 ;
        RECT 47.685 67.645 50.115 68.830 ;
        RECT 51.685 67.645 54.115 68.830 ;
        RECT 55.685 67.645 58.115 68.830 ;
        RECT 59.685 67.645 62.115 68.830 ;
        RECT 63.685 67.645 66.115 68.830 ;
        RECT 67.685 67.645 70.115 68.830 ;
        RECT 71.685 67.645 74.115 68.830 ;
        RECT 11.685 67.200 74.115 67.645 ;
        RECT 11.685 66.430 14.115 67.200 ;
        RECT 15.685 66.430 18.115 67.200 ;
        RECT 19.685 66.430 22.115 67.200 ;
        RECT 23.685 66.430 26.115 67.200 ;
        RECT 27.685 66.430 30.115 67.200 ;
        RECT 31.685 66.430 34.115 67.200 ;
        RECT 35.685 66.430 38.115 67.200 ;
        RECT 39.685 66.430 42.115 67.200 ;
        RECT 43.685 66.430 46.115 67.200 ;
        RECT 47.685 66.430 50.115 67.200 ;
        RECT 51.685 66.430 54.115 67.200 ;
        RECT 55.685 66.430 58.115 67.200 ;
        RECT 59.685 66.430 62.115 67.200 ;
        RECT 63.685 66.430 66.115 67.200 ;
        RECT 67.685 66.430 70.115 67.200 ;
        RECT 71.685 66.430 74.115 67.200 ;
        RECT 75.685 66.430 78.115 68.830 ;
        RECT 79.685 66.430 82.115 68.830 ;
        RECT 83.685 66.430 86.115 68.830 ;
        RECT 87.685 66.430 90.115 68.830 ;
        RECT 91.685 66.430 94.115 68.830 ;
        RECT 95.685 66.430 98.115 68.830 ;
        RECT 99.685 66.430 102.115 68.830 ;
        RECT 103.685 66.430 106.115 68.830 ;
        RECT 107.685 66.430 110.115 68.830 ;
        RECT 111.685 66.430 114.115 68.830 ;
        RECT 115.685 66.430 118.115 68.830 ;
        RECT 119.685 66.430 122.115 68.830 ;
        RECT 123.685 66.430 126.115 68.830 ;
        RECT 127.685 66.430 130.115 68.830 ;
        RECT 131.685 66.430 134.115 68.830 ;
        RECT 135.685 66.430 138.115 68.830 ;
        RECT 139.685 66.430 142.115 68.830 ;
        RECT 12.655 65.830 13.100 66.430 ;
        RECT 76.540 65.830 76.920 66.430 ;
        RECT 80.490 65.830 80.870 66.430 ;
        RECT 84.605 65.830 84.985 66.430 ;
        RECT 88.555 65.830 88.935 66.430 ;
        RECT 92.505 65.830 92.885 66.430 ;
        RECT 96.695 65.830 97.075 66.430 ;
        RECT 100.565 65.830 100.945 66.430 ;
        RECT 104.555 65.830 104.935 66.430 ;
        RECT 108.560 65.830 108.875 66.430 ;
        RECT 112.720 65.830 113.035 66.430 ;
        RECT 116.565 65.830 116.880 66.430 ;
        RECT 120.770 65.830 121.085 66.430 ;
        RECT 124.685 65.830 125.105 66.430 ;
        RECT 128.580 65.830 129.000 66.430 ;
        RECT 132.675 65.830 133.095 66.430 ;
        RECT 136.610 65.830 137.015 66.430 ;
        RECT 148.695 66.065 149.230 67.040 ;
        RECT 151.725 66.085 152.260 67.060 ;
        RECT 7.685 63.430 10.115 65.830 ;
        RECT 11.685 64.575 14.115 65.830 ;
        RECT 15.685 64.575 18.115 65.830 ;
        RECT 19.685 64.575 22.115 65.830 ;
        RECT 23.685 64.575 26.115 65.830 ;
        RECT 27.685 64.575 30.115 65.830 ;
        RECT 31.685 64.575 34.115 65.830 ;
        RECT 35.685 64.575 38.115 65.830 ;
        RECT 39.685 64.575 42.115 65.830 ;
        RECT 43.685 64.575 46.115 65.830 ;
        RECT 47.685 64.575 50.115 65.830 ;
        RECT 51.685 64.575 54.115 65.830 ;
        RECT 55.685 64.575 58.115 65.830 ;
        RECT 59.685 64.575 62.115 65.830 ;
        RECT 63.685 64.575 66.115 65.830 ;
        RECT 67.685 64.575 70.115 65.830 ;
        RECT 71.685 64.575 74.115 65.830 ;
        RECT 11.685 64.130 74.930 64.575 ;
        RECT 75.685 64.525 78.115 65.830 ;
        RECT 75.685 64.145 79.020 64.525 ;
        RECT 79.685 64.280 82.115 65.830 ;
        RECT 83.685 64.280 86.115 65.830 ;
        RECT 11.685 63.430 14.115 64.130 ;
        RECT 15.685 63.430 18.115 64.130 ;
        RECT 19.685 63.430 22.115 64.130 ;
        RECT 23.685 63.430 26.115 64.130 ;
        RECT 27.685 63.430 30.115 64.130 ;
        RECT 31.685 63.430 34.115 64.130 ;
        RECT 35.685 63.430 38.115 64.130 ;
        RECT 39.685 63.430 42.115 64.130 ;
        RECT 43.685 63.430 46.115 64.130 ;
        RECT 47.685 63.430 50.115 64.130 ;
        RECT 51.685 63.430 54.115 64.130 ;
        RECT 55.685 63.430 58.115 64.130 ;
        RECT 59.685 63.430 62.115 64.130 ;
        RECT 63.685 63.430 66.115 64.130 ;
        RECT 67.685 63.430 70.115 64.130 ;
        RECT 71.685 63.430 74.115 64.130 ;
        RECT 75.685 63.430 78.115 64.145 ;
        RECT 79.685 63.900 86.115 64.280 ;
        RECT 79.685 63.430 82.115 63.900 ;
        RECT 83.685 63.430 86.115 63.900 ;
        RECT 87.685 64.360 90.115 65.830 ;
        RECT 91.685 64.360 94.115 65.830 ;
        RECT 87.685 63.980 94.115 64.360 ;
        RECT 87.685 63.430 90.115 63.980 ;
        RECT 91.685 63.430 94.115 63.980 ;
        RECT 95.685 64.445 98.115 65.830 ;
        RECT 99.685 64.445 102.115 65.830 ;
        RECT 95.685 64.065 102.115 64.445 ;
        RECT 95.685 63.430 98.115 64.065 ;
        RECT 99.685 63.430 102.115 64.065 ;
        RECT 103.685 63.430 106.115 65.830 ;
        RECT 107.685 63.430 110.115 65.830 ;
        RECT 111.685 64.670 114.115 65.830 ;
        RECT 115.685 64.670 118.115 65.830 ;
        RECT 111.685 64.355 118.115 64.670 ;
        RECT 111.685 63.430 114.115 64.355 ;
        RECT 115.685 63.430 118.115 64.355 ;
        RECT 119.685 63.430 122.115 65.830 ;
        RECT 123.685 64.485 126.115 65.830 ;
        RECT 127.685 64.485 130.115 65.830 ;
        RECT 123.685 64.065 130.115 64.485 ;
        RECT 123.685 63.430 126.115 64.065 ;
        RECT 127.685 63.430 130.115 64.065 ;
        RECT 131.685 63.430 134.115 65.830 ;
        RECT 135.685 63.430 138.115 65.830 ;
        RECT 139.685 63.430 142.115 65.830 ;
        RECT 147.770 63.665 150.170 66.065 ;
        RECT 150.800 63.685 153.200 66.085 ;
        RECT 154.735 66.055 155.270 67.030 ;
        RECT 157.765 66.075 158.300 67.050 ;
        RECT 153.810 63.655 156.210 66.055 ;
        RECT 156.840 63.675 159.240 66.075 ;
        RECT 160.735 66.055 161.270 67.030 ;
        RECT 163.765 66.075 164.300 67.050 ;
        RECT 159.810 63.655 162.210 66.055 ;
        RECT 162.840 63.675 165.240 66.075 ;
        RECT 166.775 66.045 167.310 67.020 ;
        RECT 169.805 66.065 170.340 67.040 ;
        RECT 165.850 63.645 168.250 66.045 ;
        RECT 168.880 63.665 171.280 66.065 ;
        RECT 151.710 63.155 152.260 63.160 ;
        RECT 148.680 63.135 149.230 63.140 ;
        RECT 7.685 60.430 10.115 62.830 ;
        RECT 11.685 60.430 14.115 62.830 ;
        RECT 15.685 60.430 18.115 62.830 ;
        RECT 19.685 60.430 22.115 62.830 ;
        RECT 23.685 60.430 26.115 62.830 ;
        RECT 27.685 60.430 30.115 62.830 ;
        RECT 31.685 60.430 34.115 62.830 ;
        RECT 35.685 60.430 38.115 62.830 ;
        RECT 39.685 60.430 42.115 62.830 ;
        RECT 43.685 60.430 46.115 62.830 ;
        RECT 47.685 60.430 50.115 62.830 ;
        RECT 51.685 60.430 54.115 62.830 ;
        RECT 55.685 60.430 58.115 62.830 ;
        RECT 59.685 60.430 62.115 62.830 ;
        RECT 63.685 60.430 66.115 62.830 ;
        RECT 67.685 60.430 70.115 62.830 ;
        RECT 71.685 60.430 74.115 62.830 ;
        RECT 75.685 60.430 78.115 62.830 ;
        RECT 79.685 60.430 82.115 62.830 ;
        RECT 83.685 60.430 86.115 62.830 ;
        RECT 87.685 60.430 90.115 62.830 ;
        RECT 91.685 60.430 94.115 62.830 ;
        RECT 95.685 60.430 98.115 62.830 ;
        RECT 99.685 60.430 102.115 62.830 ;
        RECT 103.685 60.430 106.115 62.830 ;
        RECT 107.685 60.430 110.115 62.830 ;
        RECT 111.685 60.430 114.115 62.830 ;
        RECT 115.685 60.430 118.115 62.830 ;
        RECT 119.685 60.430 122.115 62.830 ;
        RECT 123.685 60.430 126.115 62.830 ;
        RECT 127.685 60.430 130.115 62.830 ;
        RECT 131.685 60.430 134.115 62.830 ;
        RECT 135.685 60.430 138.115 62.830 ;
        RECT 139.685 60.430 142.115 62.830 ;
        RECT 148.655 62.595 149.255 63.135 ;
        RECT 151.685 62.615 152.285 63.155 ;
        RECT 157.750 63.145 158.300 63.150 ;
        RECT 163.750 63.145 164.300 63.150 ;
        RECT 154.720 63.125 155.270 63.130 ;
        RECT 151.710 62.610 152.260 62.615 ;
        RECT 148.680 62.590 149.230 62.595 ;
        RECT 154.695 62.585 155.295 63.125 ;
        RECT 157.725 62.605 158.325 63.145 ;
        RECT 160.720 63.125 161.270 63.130 ;
        RECT 157.750 62.600 158.300 62.605 ;
        RECT 160.695 62.585 161.295 63.125 ;
        RECT 163.725 62.605 164.325 63.145 ;
        RECT 169.790 63.135 170.340 63.140 ;
        RECT 166.760 63.115 167.310 63.120 ;
        RECT 163.750 62.600 164.300 62.605 ;
        RECT 154.720 62.580 155.270 62.585 ;
        RECT 160.720 62.580 161.270 62.585 ;
        RECT 166.735 62.575 167.335 63.115 ;
        RECT 169.765 62.595 170.365 63.135 ;
        RECT 169.790 62.590 170.340 62.595 ;
        RECT 166.760 62.570 167.310 62.575 ;
        RECT 151.915 61.810 152.405 62.300 ;
        RECT 7.685 57.020 10.115 59.420 ;
        RECT 11.685 57.020 14.115 59.420 ;
        RECT 15.685 57.020 18.115 59.420 ;
        RECT 19.685 57.020 22.115 59.420 ;
        RECT 23.685 57.020 26.115 59.420 ;
        RECT 27.685 57.020 30.115 59.420 ;
        RECT 31.685 57.020 34.115 59.420 ;
        RECT 35.685 57.020 38.115 59.420 ;
        RECT 39.685 57.020 42.115 59.420 ;
        RECT 43.685 57.020 46.115 59.420 ;
        RECT 47.685 57.020 50.115 59.420 ;
        RECT 51.685 57.020 54.115 59.420 ;
        RECT 55.685 57.020 58.115 59.420 ;
        RECT 59.685 57.020 62.115 59.420 ;
        RECT 63.685 57.020 66.115 59.420 ;
        RECT 67.685 57.020 70.115 59.420 ;
        RECT 71.685 57.020 74.115 59.420 ;
        RECT 75.685 57.020 78.115 59.420 ;
        RECT 79.685 57.020 82.115 59.420 ;
        RECT 83.685 57.020 86.115 59.420 ;
        RECT 87.685 57.020 90.115 59.420 ;
        RECT 91.685 57.020 94.115 59.420 ;
        RECT 95.685 57.020 98.115 59.420 ;
        RECT 99.685 57.020 102.115 59.420 ;
        RECT 103.685 57.020 106.115 59.420 ;
        RECT 107.685 57.020 110.115 59.420 ;
        RECT 111.685 57.020 114.115 59.420 ;
        RECT 115.685 57.020 118.115 59.420 ;
        RECT 119.685 57.020 122.115 59.420 ;
        RECT 123.685 57.020 126.115 59.420 ;
        RECT 127.685 57.020 130.115 59.420 ;
        RECT 131.685 57.020 134.115 59.420 ;
        RECT 135.685 57.020 138.115 59.420 ;
        RECT 139.685 57.020 142.115 59.420 ;
        RECT 156.185 59.350 156.565 60.000 ;
        RECT 166.875 57.405 167.425 57.410 ;
        RECT 154.835 57.395 155.385 57.400 ;
        RECT 160.835 57.395 161.385 57.400 ;
        RECT 148.795 57.385 149.345 57.390 ;
        RECT 148.770 56.845 149.370 57.385 ;
        RECT 151.825 57.365 152.375 57.370 ;
        RECT 148.795 56.840 149.345 56.845 ;
        RECT 151.800 56.825 152.400 57.365 ;
        RECT 154.810 56.855 155.410 57.395 ;
        RECT 157.865 57.375 158.415 57.380 ;
        RECT 154.835 56.850 155.385 56.855 ;
        RECT 157.840 56.835 158.440 57.375 ;
        RECT 160.810 56.855 161.410 57.395 ;
        RECT 163.865 57.375 164.415 57.380 ;
        RECT 160.835 56.850 161.385 56.855 ;
        RECT 163.840 56.835 164.440 57.375 ;
        RECT 166.850 56.865 167.450 57.405 ;
        RECT 169.905 57.385 170.455 57.390 ;
        RECT 166.875 56.860 167.425 56.865 ;
        RECT 169.880 56.845 170.480 57.385 ;
        RECT 169.905 56.840 170.455 56.845 ;
        RECT 157.865 56.830 158.415 56.835 ;
        RECT 163.865 56.830 164.415 56.835 ;
        RECT 151.825 56.820 152.375 56.825 ;
        RECT 7.685 54.020 10.115 56.420 ;
        RECT 11.685 55.720 14.115 56.420 ;
        RECT 15.685 55.720 18.115 56.420 ;
        RECT 19.685 55.720 22.115 56.420 ;
        RECT 23.685 55.720 26.115 56.420 ;
        RECT 27.685 55.720 30.115 56.420 ;
        RECT 31.685 55.720 34.115 56.420 ;
        RECT 35.685 55.720 38.115 56.420 ;
        RECT 39.685 55.720 42.115 56.420 ;
        RECT 43.685 55.720 46.115 56.420 ;
        RECT 47.685 55.720 50.115 56.420 ;
        RECT 51.685 55.720 54.115 56.420 ;
        RECT 55.685 55.720 58.115 56.420 ;
        RECT 59.685 55.720 62.115 56.420 ;
        RECT 63.685 55.720 66.115 56.420 ;
        RECT 67.685 55.720 70.115 56.420 ;
        RECT 71.685 55.720 74.115 56.420 ;
        RECT 11.685 55.275 74.930 55.720 ;
        RECT 75.685 55.705 78.115 56.420 ;
        RECT 79.685 55.950 82.115 56.420 ;
        RECT 83.685 55.950 86.115 56.420 ;
        RECT 75.685 55.325 79.020 55.705 ;
        RECT 79.685 55.570 86.115 55.950 ;
        RECT 11.685 54.020 14.115 55.275 ;
        RECT 15.685 54.020 18.115 55.275 ;
        RECT 19.685 54.020 22.115 55.275 ;
        RECT 23.685 54.020 26.115 55.275 ;
        RECT 27.685 54.020 30.115 55.275 ;
        RECT 31.685 54.020 34.115 55.275 ;
        RECT 35.685 54.020 38.115 55.275 ;
        RECT 39.685 54.020 42.115 55.275 ;
        RECT 43.685 54.020 46.115 55.275 ;
        RECT 47.685 54.020 50.115 55.275 ;
        RECT 51.685 54.020 54.115 55.275 ;
        RECT 55.685 54.020 58.115 55.275 ;
        RECT 59.685 54.020 62.115 55.275 ;
        RECT 63.685 54.020 66.115 55.275 ;
        RECT 67.685 54.020 70.115 55.275 ;
        RECT 71.685 54.020 74.115 55.275 ;
        RECT 75.685 54.020 78.115 55.325 ;
        RECT 79.685 54.020 82.115 55.570 ;
        RECT 83.685 54.020 86.115 55.570 ;
        RECT 87.685 55.870 90.115 56.420 ;
        RECT 91.685 55.870 94.115 56.420 ;
        RECT 87.685 55.490 94.115 55.870 ;
        RECT 87.685 54.020 90.115 55.490 ;
        RECT 91.685 54.020 94.115 55.490 ;
        RECT 95.685 55.785 98.115 56.420 ;
        RECT 99.685 55.785 102.115 56.420 ;
        RECT 95.685 55.405 102.115 55.785 ;
        RECT 95.685 54.020 98.115 55.405 ;
        RECT 99.685 54.020 102.115 55.405 ;
        RECT 103.685 54.020 106.115 56.420 ;
        RECT 107.685 54.020 110.115 56.420 ;
        RECT 111.685 55.495 114.115 56.420 ;
        RECT 115.685 55.495 118.115 56.420 ;
        RECT 111.685 55.180 118.115 55.495 ;
        RECT 111.685 54.020 114.115 55.180 ;
        RECT 115.685 54.020 118.115 55.180 ;
        RECT 119.685 54.020 122.115 56.420 ;
        RECT 123.685 55.785 126.115 56.420 ;
        RECT 127.685 55.785 130.115 56.420 ;
        RECT 123.685 55.365 130.115 55.785 ;
        RECT 123.685 54.020 126.115 55.365 ;
        RECT 127.685 54.020 130.115 55.365 ;
        RECT 131.685 54.020 134.115 56.420 ;
        RECT 135.685 54.020 138.115 56.420 ;
        RECT 139.685 54.020 142.115 56.420 ;
        RECT 12.655 53.420 13.100 54.020 ;
        RECT 76.540 53.420 76.920 54.020 ;
        RECT 80.490 53.420 80.870 54.020 ;
        RECT 84.605 53.420 84.985 54.020 ;
        RECT 88.555 53.420 88.935 54.020 ;
        RECT 92.505 53.420 92.885 54.020 ;
        RECT 96.695 53.420 97.075 54.020 ;
        RECT 100.565 53.420 100.945 54.020 ;
        RECT 104.555 53.420 104.935 54.020 ;
        RECT 108.560 53.420 108.875 54.020 ;
        RECT 112.720 53.420 113.035 54.020 ;
        RECT 116.565 53.420 116.880 54.020 ;
        RECT 120.770 53.420 121.085 54.020 ;
        RECT 124.685 53.420 125.105 54.020 ;
        RECT 128.580 53.420 129.000 54.020 ;
        RECT 132.675 53.420 133.095 54.020 ;
        RECT 136.610 53.420 137.015 54.020 ;
        RECT 147.885 53.915 150.285 56.315 ;
        RECT 7.685 51.020 10.115 53.420 ;
        RECT 11.685 52.650 14.115 53.420 ;
        RECT 15.685 52.650 18.115 53.420 ;
        RECT 19.685 52.650 22.115 53.420 ;
        RECT 23.685 52.650 26.115 53.420 ;
        RECT 27.685 52.650 30.115 53.420 ;
        RECT 31.685 52.650 34.115 53.420 ;
        RECT 35.685 52.650 38.115 53.420 ;
        RECT 39.685 52.650 42.115 53.420 ;
        RECT 43.685 52.650 46.115 53.420 ;
        RECT 47.685 52.650 50.115 53.420 ;
        RECT 51.685 52.650 54.115 53.420 ;
        RECT 55.685 52.650 58.115 53.420 ;
        RECT 59.685 52.650 62.115 53.420 ;
        RECT 63.685 52.650 66.115 53.420 ;
        RECT 67.685 52.650 70.115 53.420 ;
        RECT 71.685 52.650 74.115 53.420 ;
        RECT 11.685 52.205 74.115 52.650 ;
        RECT 11.685 51.020 14.115 52.205 ;
        RECT 15.685 51.020 18.115 52.205 ;
        RECT 19.685 51.020 22.115 52.205 ;
        RECT 23.685 51.020 26.115 52.205 ;
        RECT 27.685 51.020 30.115 52.205 ;
        RECT 31.685 51.020 34.115 52.205 ;
        RECT 35.685 51.020 38.115 52.205 ;
        RECT 39.685 51.020 42.115 52.205 ;
        RECT 43.685 51.020 46.115 52.205 ;
        RECT 47.685 51.020 50.115 52.205 ;
        RECT 51.685 51.020 54.115 52.205 ;
        RECT 55.685 51.020 58.115 52.205 ;
        RECT 59.685 51.020 62.115 52.205 ;
        RECT 63.685 51.020 66.115 52.205 ;
        RECT 67.685 51.020 70.115 52.205 ;
        RECT 71.685 51.020 74.115 52.205 ;
        RECT 75.685 51.020 78.115 53.420 ;
        RECT 79.685 51.020 82.115 53.420 ;
        RECT 83.685 51.020 86.115 53.420 ;
        RECT 87.685 51.020 90.115 53.420 ;
        RECT 91.685 51.020 94.115 53.420 ;
        RECT 95.685 51.020 98.115 53.420 ;
        RECT 99.685 51.020 102.115 53.420 ;
        RECT 103.685 51.020 106.115 53.420 ;
        RECT 107.685 51.020 110.115 53.420 ;
        RECT 111.685 51.020 114.115 53.420 ;
        RECT 115.685 51.020 118.115 53.420 ;
        RECT 119.685 51.020 122.115 53.420 ;
        RECT 123.685 51.020 126.115 53.420 ;
        RECT 127.685 51.020 130.115 53.420 ;
        RECT 131.685 51.020 134.115 53.420 ;
        RECT 135.685 51.020 138.115 53.420 ;
        RECT 139.685 51.020 142.115 53.420 ;
        RECT 148.810 52.940 149.345 53.915 ;
        RECT 150.915 53.895 153.315 56.295 ;
        RECT 153.925 53.925 156.325 56.325 ;
        RECT 151.840 52.920 152.375 53.895 ;
        RECT 154.850 52.950 155.385 53.925 ;
        RECT 156.955 53.905 159.355 56.305 ;
        RECT 159.925 53.925 162.325 56.325 ;
        RECT 157.880 52.930 158.415 53.905 ;
        RECT 160.850 52.950 161.385 53.925 ;
        RECT 162.955 53.905 165.355 56.305 ;
        RECT 165.965 53.935 168.365 56.335 ;
        RECT 163.880 52.930 164.415 53.905 ;
        RECT 166.890 52.960 167.425 53.935 ;
        RECT 168.995 53.915 171.395 56.315 ;
        RECT 169.920 52.940 170.455 53.915 ;
        RECT 72.730 50.420 73.175 51.020 ;
        RECT 76.540 50.420 76.920 51.020 ;
        RECT 80.490 50.420 80.870 51.020 ;
        RECT 84.605 50.420 84.985 51.020 ;
        RECT 88.555 50.420 88.935 51.020 ;
        RECT 92.505 50.420 92.885 51.020 ;
        RECT 96.695 50.420 97.075 51.020 ;
        RECT 100.565 50.420 100.945 51.020 ;
        RECT 104.555 50.420 104.935 51.020 ;
        RECT 108.560 50.420 108.875 51.020 ;
        RECT 112.720 50.420 113.035 51.020 ;
        RECT 116.565 50.420 116.880 51.020 ;
        RECT 120.445 50.420 121.420 51.020 ;
        RECT 124.685 50.420 125.105 51.020 ;
        RECT 128.580 50.420 129.000 51.020 ;
        RECT 132.675 50.420 133.095 51.020 ;
        RECT 136.610 50.420 137.015 51.020 ;
        RECT 7.685 48.020 10.115 50.420 ;
        RECT 11.685 49.690 14.115 50.420 ;
        RECT 15.685 49.690 18.115 50.420 ;
        RECT 19.685 49.690 22.115 50.420 ;
        RECT 23.685 49.690 26.115 50.420 ;
        RECT 27.685 49.690 30.115 50.420 ;
        RECT 31.685 49.690 34.115 50.420 ;
        RECT 35.685 49.690 38.115 50.420 ;
        RECT 39.685 49.690 42.115 50.420 ;
        RECT 43.685 49.690 46.115 50.420 ;
        RECT 47.685 49.690 50.115 50.420 ;
        RECT 51.685 49.690 54.115 50.420 ;
        RECT 55.685 49.690 58.115 50.420 ;
        RECT 59.685 49.690 62.115 50.420 ;
        RECT 63.685 49.690 66.115 50.420 ;
        RECT 67.685 49.690 70.115 50.420 ;
        RECT 71.685 49.690 74.115 50.420 ;
        RECT 11.685 49.245 74.115 49.690 ;
        RECT 11.685 48.020 14.115 49.245 ;
        RECT 15.685 48.020 18.115 49.245 ;
        RECT 19.685 48.020 22.115 49.245 ;
        RECT 12.410 47.420 12.855 48.020 ;
        RECT 22.675 47.930 23.175 48.450 ;
        RECT 23.685 48.020 26.115 49.245 ;
        RECT 27.685 48.020 30.115 49.245 ;
        RECT 31.685 48.020 34.115 49.245 ;
        RECT 35.685 48.020 38.115 49.245 ;
        RECT 39.685 48.020 42.115 49.245 ;
        RECT 43.685 48.020 46.115 49.245 ;
        RECT 47.685 48.020 50.115 49.245 ;
        RECT 51.685 48.020 54.115 49.245 ;
        RECT 55.685 48.020 58.115 49.245 ;
        RECT 59.685 48.020 62.115 49.245 ;
        RECT 63.685 48.020 66.115 49.245 ;
        RECT 67.685 48.020 70.115 49.245 ;
        RECT 71.685 48.020 74.115 49.245 ;
        RECT 75.685 48.020 78.115 50.420 ;
        RECT 79.685 48.020 82.115 50.420 ;
        RECT 83.685 48.020 86.115 50.420 ;
        RECT 87.685 48.020 90.115 50.420 ;
        RECT 91.685 48.020 94.115 50.420 ;
        RECT 95.685 48.020 98.115 50.420 ;
        RECT 99.685 48.020 102.115 50.420 ;
        RECT 103.685 48.020 106.115 50.420 ;
        RECT 107.685 48.020 110.115 50.420 ;
        RECT 111.685 48.020 114.115 50.420 ;
        RECT 115.685 48.020 118.115 50.420 ;
        RECT 119.685 48.020 122.115 50.420 ;
        RECT 123.685 48.020 126.115 50.420 ;
        RECT 127.685 48.020 130.115 50.420 ;
        RECT 131.685 48.020 134.115 50.420 ;
        RECT 135.685 48.020 138.115 50.420 ;
        RECT 139.685 48.020 142.115 50.420 ;
        RECT 148.775 48.720 149.310 49.695 ;
        RECT 151.805 48.740 152.340 49.715 ;
        RECT 76.540 47.420 76.920 48.020 ;
        RECT 80.490 47.420 80.870 48.020 ;
        RECT 84.605 47.420 84.985 48.020 ;
        RECT 88.555 47.420 88.935 48.020 ;
        RECT 92.505 47.420 92.885 48.020 ;
        RECT 96.695 47.420 97.075 48.020 ;
        RECT 100.565 47.420 100.945 48.020 ;
        RECT 104.555 47.420 104.935 48.020 ;
        RECT 108.560 47.420 108.875 48.020 ;
        RECT 112.720 47.420 113.035 48.020 ;
        RECT 116.565 47.420 116.880 48.020 ;
        RECT 120.770 47.420 121.085 48.020 ;
        RECT 124.685 47.420 125.105 48.020 ;
        RECT 128.580 47.420 129.000 48.020 ;
        RECT 132.675 47.420 133.095 48.020 ;
        RECT 136.610 47.420 137.015 48.020 ;
        RECT 7.685 45.020 10.115 47.420 ;
        RECT 11.685 46.405 14.115 47.420 ;
        RECT 15.685 46.405 18.115 47.420 ;
        RECT 19.685 46.405 22.115 47.420 ;
        RECT 23.685 46.405 26.115 47.420 ;
        RECT 27.685 46.405 30.115 47.420 ;
        RECT 31.685 46.405 34.115 47.420 ;
        RECT 35.685 46.405 38.115 47.420 ;
        RECT 39.685 46.405 42.115 47.420 ;
        RECT 43.685 46.405 46.115 47.420 ;
        RECT 47.685 46.405 50.115 47.420 ;
        RECT 51.685 46.405 54.115 47.420 ;
        RECT 55.685 46.405 58.115 47.420 ;
        RECT 59.685 46.405 62.115 47.420 ;
        RECT 63.685 46.405 66.115 47.420 ;
        RECT 67.685 46.405 70.115 47.420 ;
        RECT 71.685 46.405 74.115 47.420 ;
        RECT 11.685 45.960 74.115 46.405 ;
        RECT 11.685 45.020 14.115 45.960 ;
        RECT 15.685 45.020 18.115 45.960 ;
        RECT 19.685 45.020 22.115 45.960 ;
        RECT 23.685 45.020 26.115 45.960 ;
        RECT 27.685 45.020 30.115 45.960 ;
        RECT 31.685 45.020 34.115 45.960 ;
        RECT 35.685 45.020 38.115 45.960 ;
        RECT 39.685 45.020 42.115 45.960 ;
        RECT 43.685 45.020 46.115 45.960 ;
        RECT 47.685 45.020 50.115 45.960 ;
        RECT 51.685 45.020 54.115 45.960 ;
        RECT 55.685 45.020 58.115 45.960 ;
        RECT 59.685 45.020 62.115 45.960 ;
        RECT 63.685 45.020 66.115 45.960 ;
        RECT 67.685 45.020 70.115 45.960 ;
        RECT 71.685 45.020 74.115 45.960 ;
        RECT 75.685 45.020 78.115 47.420 ;
        RECT 79.685 45.020 82.115 47.420 ;
        RECT 83.685 45.020 86.115 47.420 ;
        RECT 87.685 45.020 90.115 47.420 ;
        RECT 91.685 45.020 94.115 47.420 ;
        RECT 95.685 45.020 98.115 47.420 ;
        RECT 99.685 45.020 102.115 47.420 ;
        RECT 103.685 45.020 106.115 47.420 ;
        RECT 107.685 45.020 110.115 47.420 ;
        RECT 111.685 45.020 114.115 47.420 ;
        RECT 115.685 45.020 118.115 47.420 ;
        RECT 119.685 45.020 122.115 47.420 ;
        RECT 123.685 45.020 126.115 47.420 ;
        RECT 127.685 45.020 130.115 47.420 ;
        RECT 131.685 45.020 134.115 47.420 ;
        RECT 135.685 45.020 138.115 47.420 ;
        RECT 139.685 45.020 142.115 47.420 ;
        RECT 147.850 46.320 150.250 48.720 ;
        RECT 150.880 46.340 153.280 48.740 ;
        RECT 154.815 48.710 155.350 49.685 ;
        RECT 157.845 48.730 158.380 49.705 ;
        RECT 153.890 46.310 156.290 48.710 ;
        RECT 156.920 46.330 159.320 48.730 ;
        RECT 160.815 48.710 161.350 49.685 ;
        RECT 159.890 46.310 162.290 48.710 ;
        RECT 163.855 48.705 164.390 49.680 ;
        RECT 162.930 46.305 165.330 48.705 ;
        RECT 166.855 48.700 167.390 49.675 ;
        RECT 169.885 48.720 170.420 49.695 ;
        RECT 165.930 46.300 168.330 48.700 ;
        RECT 168.960 46.320 171.360 48.720 ;
        RECT 151.790 45.810 152.340 45.815 ;
        RECT 148.760 45.790 149.310 45.795 ;
        RECT 148.735 45.250 149.335 45.790 ;
        RECT 151.765 45.270 152.365 45.810 ;
        RECT 157.830 45.800 158.380 45.805 ;
        RECT 154.800 45.780 155.350 45.785 ;
        RECT 151.790 45.265 152.340 45.270 ;
        RECT 148.760 45.245 149.310 45.250 ;
        RECT 154.775 45.240 155.375 45.780 ;
        RECT 157.805 45.260 158.405 45.800 ;
        RECT 169.870 45.790 170.420 45.795 ;
        RECT 160.800 45.780 161.350 45.785 ;
        RECT 157.830 45.255 158.380 45.260 ;
        RECT 160.775 45.240 161.375 45.780 ;
        RECT 163.840 45.775 164.390 45.780 ;
        RECT 154.800 45.235 155.350 45.240 ;
        RECT 160.800 45.235 161.350 45.240 ;
        RECT 163.815 45.235 164.415 45.775 ;
        RECT 166.840 45.770 167.390 45.775 ;
        RECT 163.840 45.230 164.390 45.235 ;
        RECT 166.815 45.230 167.415 45.770 ;
        RECT 169.845 45.250 170.445 45.790 ;
        RECT 169.870 45.245 170.420 45.250 ;
        RECT 166.840 45.225 167.390 45.230 ;
        RECT 72.565 44.420 73.010 45.020 ;
        RECT 76.540 44.420 76.920 45.020 ;
        RECT 80.490 44.420 80.870 45.020 ;
        RECT 84.605 44.420 84.985 45.020 ;
        RECT 88.555 44.420 88.935 45.020 ;
        RECT 92.505 44.420 92.885 45.020 ;
        RECT 96.695 44.420 97.075 45.020 ;
        RECT 100.565 44.420 100.945 45.020 ;
        RECT 104.555 44.420 104.935 45.020 ;
        RECT 108.560 44.420 108.875 45.020 ;
        RECT 112.720 44.420 113.035 45.020 ;
        RECT 116.565 44.420 116.880 45.020 ;
        RECT 120.770 44.420 121.085 45.020 ;
        RECT 124.685 44.420 125.105 45.020 ;
        RECT 128.580 44.420 129.000 45.020 ;
        RECT 132.675 44.420 133.095 45.020 ;
        RECT 7.685 42.020 10.115 44.420 ;
        RECT 11.685 43.360 14.115 44.420 ;
        RECT 15.685 43.360 18.115 44.420 ;
        RECT 19.685 43.360 22.115 44.420 ;
        RECT 23.685 43.360 26.115 44.420 ;
        RECT 27.685 43.360 30.115 44.420 ;
        RECT 31.685 43.360 34.115 44.420 ;
        RECT 35.685 43.360 38.115 44.420 ;
        RECT 39.685 43.360 42.115 44.420 ;
        RECT 43.685 43.360 46.115 44.420 ;
        RECT 47.685 43.360 50.115 44.420 ;
        RECT 51.685 43.360 54.115 44.420 ;
        RECT 55.685 43.360 58.115 44.420 ;
        RECT 59.685 43.360 62.115 44.420 ;
        RECT 63.685 43.360 66.115 44.420 ;
        RECT 67.685 43.360 70.115 44.420 ;
        RECT 71.685 43.360 74.115 44.420 ;
        RECT 11.685 42.915 74.115 43.360 ;
        RECT 11.685 42.020 14.115 42.915 ;
        RECT 15.685 42.020 18.115 42.915 ;
        RECT 19.685 42.020 22.115 42.915 ;
        RECT 23.685 42.020 26.115 42.915 ;
        RECT 27.685 42.020 30.115 42.915 ;
        RECT 31.685 42.020 34.115 42.915 ;
        RECT 35.685 42.020 38.115 42.915 ;
        RECT 39.685 42.020 42.115 42.915 ;
        RECT 43.685 42.020 46.115 42.915 ;
        RECT 47.685 42.020 50.115 42.915 ;
        RECT 51.685 42.020 54.115 42.915 ;
        RECT 55.685 42.020 58.115 42.915 ;
        RECT 59.685 42.020 62.115 42.915 ;
        RECT 63.685 42.020 66.115 42.915 ;
        RECT 67.685 42.020 70.115 42.915 ;
        RECT 71.685 42.020 74.115 42.915 ;
        RECT 75.685 42.020 78.115 44.420 ;
        RECT 79.685 42.020 82.115 44.420 ;
        RECT 83.685 42.020 86.115 44.420 ;
        RECT 87.685 42.020 90.115 44.420 ;
        RECT 91.685 42.020 94.115 44.420 ;
        RECT 95.685 42.020 98.115 44.420 ;
        RECT 99.685 42.020 102.115 44.420 ;
        RECT 103.685 42.020 106.115 44.420 ;
        RECT 107.685 42.020 110.115 44.420 ;
        RECT 111.685 42.020 114.115 44.420 ;
        RECT 115.685 42.020 118.115 44.420 ;
        RECT 119.685 42.020 122.115 44.420 ;
        RECT 123.685 42.020 126.115 44.420 ;
        RECT 127.685 42.020 130.115 44.420 ;
        RECT 131.685 42.020 134.115 44.420 ;
        RECT 135.685 42.020 138.115 44.420 ;
        RECT 139.685 42.020 142.115 44.420 ;
        RECT 12.495 41.420 12.940 42.020 ;
        RECT 76.540 41.420 76.920 42.020 ;
        RECT 80.490 41.420 80.870 42.020 ;
        RECT 84.605 41.420 84.985 42.020 ;
        RECT 88.555 41.420 88.935 42.020 ;
        RECT 92.505 41.420 92.885 42.020 ;
        RECT 96.695 41.420 97.075 42.020 ;
        RECT 100.565 41.420 100.945 42.020 ;
        RECT 104.555 41.420 104.935 42.020 ;
        RECT 108.560 41.420 108.875 42.020 ;
        RECT 112.720 41.420 113.035 42.020 ;
        RECT 116.565 41.420 116.880 42.020 ;
        RECT 120.770 41.420 121.085 42.020 ;
        RECT 124.685 41.420 125.105 42.020 ;
        RECT 128.580 41.420 129.000 42.020 ;
        RECT 132.675 41.420 133.095 42.020 ;
        RECT 136.610 41.420 137.015 42.020 ;
        RECT 7.685 39.020 10.115 41.420 ;
        RECT 11.685 40.405 14.115 41.420 ;
        RECT 15.685 40.405 18.115 41.420 ;
        RECT 19.685 40.405 22.115 41.420 ;
        RECT 23.685 40.405 26.115 41.420 ;
        RECT 27.685 40.405 30.115 41.420 ;
        RECT 31.685 40.405 34.115 41.420 ;
        RECT 35.685 40.405 38.115 41.420 ;
        RECT 39.685 40.405 42.115 41.420 ;
        RECT 43.685 40.405 46.115 41.420 ;
        RECT 47.685 40.405 50.115 41.420 ;
        RECT 51.685 40.405 54.115 41.420 ;
        RECT 55.685 40.405 58.115 41.420 ;
        RECT 59.685 40.405 62.115 41.420 ;
        RECT 63.685 40.405 66.115 41.420 ;
        RECT 67.685 40.405 70.115 41.420 ;
        RECT 71.685 40.405 74.115 41.420 ;
        RECT 11.685 39.960 74.115 40.405 ;
        RECT 11.685 39.020 14.115 39.960 ;
        RECT 15.685 39.020 18.115 39.960 ;
        RECT 19.685 39.020 22.115 39.960 ;
        RECT 23.685 39.020 26.115 39.960 ;
        RECT 27.685 39.020 30.115 39.960 ;
        RECT 31.685 39.020 34.115 39.960 ;
        RECT 35.685 39.020 38.115 39.960 ;
        RECT 39.685 39.020 42.115 39.960 ;
        RECT 43.685 39.020 46.115 39.960 ;
        RECT 47.685 39.020 50.115 39.960 ;
        RECT 51.685 39.020 54.115 39.960 ;
        RECT 55.685 39.020 58.115 39.960 ;
        RECT 59.685 39.020 62.115 39.960 ;
        RECT 63.685 39.020 66.115 39.960 ;
        RECT 67.685 39.020 70.115 39.960 ;
        RECT 71.685 39.020 74.115 39.960 ;
        RECT 75.685 39.020 78.115 41.420 ;
        RECT 79.685 39.020 82.115 41.420 ;
        RECT 83.685 39.020 86.115 41.420 ;
        RECT 87.685 39.020 90.115 41.420 ;
        RECT 91.685 39.020 94.115 41.420 ;
        RECT 95.685 39.020 98.115 41.420 ;
        RECT 99.685 39.020 102.115 41.420 ;
        RECT 103.685 39.020 106.115 41.420 ;
        RECT 107.685 39.020 110.115 41.420 ;
        RECT 111.685 39.020 114.115 41.420 ;
        RECT 115.685 39.020 118.115 41.420 ;
        RECT 119.685 39.020 122.115 41.420 ;
        RECT 123.685 39.020 126.115 41.420 ;
        RECT 127.685 39.020 130.115 41.420 ;
        RECT 131.685 39.020 134.115 41.420 ;
        RECT 135.685 39.020 138.115 41.420 ;
        RECT 139.685 39.020 142.115 41.420 ;
        RECT 72.485 38.420 72.930 39.020 ;
        RECT 76.540 38.420 76.920 39.020 ;
        RECT 80.490 38.420 80.870 39.020 ;
        RECT 84.605 38.420 84.985 39.020 ;
        RECT 88.555 38.420 88.935 39.020 ;
        RECT 92.505 38.420 92.885 39.020 ;
        RECT 96.695 38.420 97.075 39.020 ;
        RECT 100.565 38.420 100.945 39.020 ;
        RECT 104.555 38.420 104.935 39.020 ;
        RECT 108.560 38.420 108.875 39.020 ;
        RECT 112.720 38.420 113.035 39.020 ;
        RECT 116.565 38.420 116.880 39.020 ;
        RECT 120.770 38.420 121.085 39.020 ;
        RECT 124.685 38.420 125.105 39.020 ;
        RECT 128.580 38.420 129.000 39.020 ;
        RECT 132.675 38.420 133.095 39.020 ;
        RECT 7.685 36.020 10.115 38.420 ;
        RECT 11.685 37.775 14.115 38.420 ;
        RECT 15.685 37.775 18.115 38.420 ;
        RECT 19.685 37.775 22.115 38.420 ;
        RECT 23.685 37.775 26.115 38.420 ;
        RECT 27.685 37.775 30.115 38.420 ;
        RECT 31.685 37.775 34.115 38.420 ;
        RECT 35.685 37.775 38.115 38.420 ;
        RECT 39.685 37.775 42.115 38.420 ;
        RECT 43.685 37.775 46.115 38.420 ;
        RECT 47.685 37.775 50.115 38.420 ;
        RECT 51.685 37.775 54.115 38.420 ;
        RECT 55.685 37.775 58.115 38.420 ;
        RECT 59.685 37.775 62.115 38.420 ;
        RECT 63.685 37.775 66.115 38.420 ;
        RECT 67.685 37.775 70.115 38.420 ;
        RECT 71.685 37.775 74.115 38.420 ;
        RECT 11.685 37.330 74.115 37.775 ;
        RECT 11.685 36.020 14.115 37.330 ;
        RECT 15.685 36.020 18.115 37.330 ;
        RECT 19.685 36.020 22.115 37.330 ;
        RECT 23.685 36.020 26.115 37.330 ;
        RECT 27.685 36.020 30.115 37.330 ;
        RECT 31.685 36.020 34.115 37.330 ;
        RECT 35.685 36.020 38.115 37.330 ;
        RECT 39.685 36.020 42.115 37.330 ;
        RECT 43.685 36.020 46.115 37.330 ;
        RECT 47.685 36.020 50.115 37.330 ;
        RECT 51.685 36.020 54.115 37.330 ;
        RECT 55.685 36.020 58.115 37.330 ;
        RECT 59.685 36.020 62.115 37.330 ;
        RECT 63.685 36.020 66.115 37.330 ;
        RECT 67.685 36.020 70.115 37.330 ;
        RECT 71.685 36.020 74.115 37.330 ;
        RECT 75.685 36.020 78.115 38.420 ;
        RECT 79.685 36.020 82.115 38.420 ;
        RECT 83.685 36.020 86.115 38.420 ;
        RECT 87.685 36.020 90.115 38.420 ;
        RECT 91.685 36.020 94.115 38.420 ;
        RECT 95.685 36.020 98.115 38.420 ;
        RECT 99.685 36.020 102.115 38.420 ;
        RECT 103.685 36.020 106.115 38.420 ;
        RECT 107.685 36.020 110.115 38.420 ;
        RECT 111.685 36.020 114.115 38.420 ;
        RECT 115.685 36.020 118.115 38.420 ;
        RECT 119.685 36.020 122.115 38.420 ;
        RECT 123.685 36.020 126.115 38.420 ;
        RECT 127.685 36.020 130.115 38.420 ;
        RECT 131.685 36.020 134.115 38.420 ;
        RECT 135.685 37.910 138.115 38.420 ;
        RECT 135.685 37.490 139.105 37.910 ;
        RECT 135.685 36.020 138.115 37.490 ;
        RECT 139.685 36.020 142.115 38.420 ;
        RECT 12.330 35.420 12.775 36.020 ;
        RECT 76.540 35.420 76.920 36.020 ;
        RECT 80.490 35.420 80.870 36.020 ;
        RECT 84.605 35.420 84.985 36.020 ;
        RECT 88.555 35.420 88.935 36.020 ;
        RECT 92.505 35.420 92.885 36.020 ;
        RECT 96.695 35.420 97.075 36.020 ;
        RECT 100.565 35.420 100.945 36.020 ;
        RECT 104.555 35.420 104.935 36.020 ;
        RECT 108.560 35.420 108.875 36.020 ;
        RECT 112.720 35.420 113.035 36.020 ;
        RECT 116.565 35.420 116.880 36.020 ;
        RECT 120.770 35.420 121.085 36.020 ;
        RECT 124.685 35.420 125.105 36.020 ;
        RECT 128.580 35.420 129.000 36.020 ;
        RECT 132.675 35.420 133.095 36.020 ;
        RECT 7.685 33.020 10.115 35.420 ;
        RECT 11.685 34.650 14.115 35.420 ;
        RECT 15.685 34.650 18.115 35.420 ;
        RECT 19.685 34.650 22.115 35.420 ;
        RECT 23.685 34.650 26.115 35.420 ;
        RECT 27.685 34.650 30.115 35.420 ;
        RECT 31.685 34.650 34.115 35.420 ;
        RECT 35.685 34.650 38.115 35.420 ;
        RECT 39.685 34.650 42.115 35.420 ;
        RECT 43.685 34.650 46.115 35.420 ;
        RECT 47.685 34.650 50.115 35.420 ;
        RECT 51.685 34.650 54.115 35.420 ;
        RECT 55.685 34.650 58.115 35.420 ;
        RECT 59.685 34.650 62.115 35.420 ;
        RECT 63.685 34.650 66.115 35.420 ;
        RECT 67.685 34.650 70.115 35.420 ;
        RECT 71.685 34.650 74.115 35.420 ;
        RECT 11.685 34.205 74.115 34.650 ;
        RECT 11.685 33.020 14.115 34.205 ;
        RECT 15.685 33.020 18.115 34.205 ;
        RECT 19.685 33.020 22.115 34.205 ;
        RECT 23.685 33.020 26.115 34.205 ;
        RECT 27.685 33.020 30.115 34.205 ;
        RECT 31.685 33.020 34.115 34.205 ;
        RECT 35.685 33.020 38.115 34.205 ;
        RECT 39.685 33.020 42.115 34.205 ;
        RECT 43.685 33.020 46.115 34.205 ;
        RECT 47.685 33.020 50.115 34.205 ;
        RECT 51.685 33.020 54.115 34.205 ;
        RECT 55.685 33.020 58.115 34.205 ;
        RECT 59.685 33.020 62.115 34.205 ;
        RECT 63.685 33.020 66.115 34.205 ;
        RECT 67.685 33.020 70.115 34.205 ;
        RECT 71.685 33.020 74.115 34.205 ;
        RECT 75.685 34.585 78.115 35.420 ;
        RECT 79.685 34.585 82.115 35.420 ;
        RECT 75.685 34.205 82.115 34.585 ;
        RECT 75.685 33.020 78.115 34.205 ;
        RECT 79.685 33.020 82.115 34.205 ;
        RECT 83.685 34.665 86.115 35.420 ;
        RECT 87.685 34.665 90.115 35.420 ;
        RECT 83.685 34.285 90.115 34.665 ;
        RECT 83.685 33.020 86.115 34.285 ;
        RECT 87.685 33.020 90.115 34.285 ;
        RECT 91.685 34.750 94.115 35.420 ;
        RECT 95.685 34.750 98.115 35.420 ;
        RECT 91.685 34.370 98.115 34.750 ;
        RECT 91.685 33.020 94.115 34.370 ;
        RECT 95.685 33.020 98.115 34.370 ;
        RECT 99.685 34.585 102.115 35.420 ;
        RECT 103.685 34.585 106.115 35.420 ;
        RECT 99.685 34.205 106.115 34.585 ;
        RECT 99.685 33.020 102.115 34.205 ;
        RECT 103.685 33.020 106.115 34.205 ;
        RECT 107.685 34.390 110.115 35.420 ;
        RECT 111.685 34.390 114.115 35.420 ;
        RECT 107.685 34.075 114.115 34.390 ;
        RECT 107.685 33.020 110.115 34.075 ;
        RECT 111.685 33.020 114.115 34.075 ;
        RECT 115.685 34.390 118.115 35.420 ;
        RECT 119.685 34.390 122.115 35.420 ;
        RECT 115.685 34.075 122.115 34.390 ;
        RECT 115.685 33.020 118.115 34.075 ;
        RECT 119.685 33.020 122.115 34.075 ;
        RECT 123.685 34.645 126.115 35.420 ;
        RECT 127.685 34.645 130.115 35.420 ;
        RECT 123.685 34.225 130.115 34.645 ;
        RECT 123.685 33.020 126.115 34.225 ;
        RECT 127.685 33.020 130.115 34.225 ;
        RECT 131.685 33.020 134.115 35.420 ;
        RECT 135.685 34.910 138.115 35.420 ;
        RECT 135.685 34.490 139.145 34.910 ;
        RECT 135.685 33.020 138.115 34.490 ;
        RECT 139.685 33.020 142.115 35.420 ;
        RECT 7.685 30.020 10.115 32.420 ;
        RECT 11.685 30.020 14.115 32.420 ;
        RECT 15.685 30.020 18.115 32.420 ;
        RECT 19.685 30.020 22.115 32.420 ;
        RECT 23.685 30.020 26.115 32.420 ;
        RECT 27.685 30.020 30.115 32.420 ;
        RECT 31.685 30.020 34.115 32.420 ;
        RECT 35.685 30.020 38.115 32.420 ;
        RECT 39.685 30.020 42.115 32.420 ;
        RECT 43.685 30.020 46.115 32.420 ;
        RECT 47.685 30.020 50.115 32.420 ;
        RECT 51.685 30.020 54.115 32.420 ;
        RECT 55.685 30.020 58.115 32.420 ;
        RECT 59.685 30.020 62.115 32.420 ;
        RECT 63.685 30.020 66.115 32.420 ;
        RECT 67.685 30.020 70.115 32.420 ;
        RECT 71.685 30.020 74.115 32.420 ;
        RECT 75.685 30.020 78.115 32.420 ;
        RECT 79.685 30.020 82.115 32.420 ;
        RECT 83.685 30.020 86.115 32.420 ;
        RECT 87.685 30.020 90.115 32.420 ;
        RECT 91.685 30.020 94.115 32.420 ;
        RECT 95.685 30.020 98.115 32.420 ;
        RECT 99.685 30.020 102.115 32.420 ;
        RECT 103.685 30.020 106.115 32.420 ;
        RECT 107.685 30.020 110.115 32.420 ;
        RECT 111.685 30.020 114.115 32.420 ;
        RECT 115.685 30.020 118.115 32.420 ;
        RECT 119.685 30.020 122.115 32.420 ;
        RECT 123.685 30.020 126.115 32.420 ;
        RECT 127.685 30.020 130.115 32.420 ;
        RECT 131.685 30.020 134.115 32.420 ;
        RECT 135.685 30.020 138.115 32.420 ;
        RECT 139.685 30.020 142.115 32.420 ;
      LAYER via3 ;
        RECT 148.650 74.190 149.190 74.730 ;
        RECT 151.680 74.170 152.220 74.710 ;
        RECT 154.690 74.200 155.230 74.740 ;
        RECT 157.720 74.180 158.260 74.720 ;
        RECT 160.690 74.200 161.230 74.740 ;
        RECT 163.730 74.205 164.270 74.745 ;
        RECT 166.730 74.210 167.270 74.750 ;
        RECT 169.760 74.190 170.300 74.730 ;
        RECT 22.760 71.475 23.110 71.825 ;
        RECT 148.685 62.595 149.225 63.135 ;
        RECT 151.715 62.615 152.255 63.155 ;
        RECT 154.725 62.585 155.265 63.125 ;
        RECT 157.755 62.605 158.295 63.145 ;
        RECT 160.725 62.585 161.265 63.125 ;
        RECT 163.755 62.605 164.295 63.145 ;
        RECT 166.765 62.575 167.305 63.115 ;
        RECT 169.795 62.595 170.335 63.135 ;
        RECT 152.025 61.910 152.345 62.230 ;
        RECT 156.225 59.380 156.545 59.700 ;
        RECT 148.800 56.845 149.340 57.385 ;
        RECT 151.830 56.825 152.370 57.365 ;
        RECT 154.840 56.855 155.380 57.395 ;
        RECT 157.870 56.835 158.410 57.375 ;
        RECT 160.840 56.855 161.380 57.395 ;
        RECT 163.870 56.835 164.410 57.375 ;
        RECT 166.880 56.865 167.420 57.405 ;
        RECT 169.910 56.845 170.450 57.385 ;
        RECT 22.760 48.025 23.110 48.375 ;
        RECT 148.765 45.250 149.305 45.790 ;
        RECT 151.795 45.270 152.335 45.810 ;
        RECT 154.805 45.240 155.345 45.780 ;
        RECT 157.835 45.260 158.375 45.800 ;
        RECT 160.805 45.240 161.345 45.780 ;
        RECT 163.845 45.235 164.385 45.775 ;
        RECT 166.845 45.230 167.385 45.770 ;
        RECT 169.875 45.250 170.415 45.790 ;
      LAYER met4 ;
        RECT 8.080 88.800 9.690 89.435 ;
        RECT 12.080 88.800 13.690 89.435 ;
        RECT 16.080 88.800 17.690 89.435 ;
        RECT 20.080 88.800 21.690 89.435 ;
        RECT 24.080 88.800 25.690 89.435 ;
        RECT 28.080 88.800 29.690 89.435 ;
        RECT 32.080 88.800 33.690 89.435 ;
        RECT 36.080 88.800 37.690 89.435 ;
        RECT 40.080 88.800 41.690 89.435 ;
        RECT 44.080 88.800 45.690 89.435 ;
        RECT 48.080 88.800 49.690 89.435 ;
        RECT 52.080 88.800 53.690 89.435 ;
        RECT 56.080 88.800 57.690 89.435 ;
        RECT 60.080 88.800 61.690 89.435 ;
        RECT 64.080 88.800 65.690 89.435 ;
        RECT 68.080 88.800 69.690 89.435 ;
        RECT 72.080 88.800 73.690 89.435 ;
        RECT 76.080 88.800 77.690 89.435 ;
        RECT 80.080 88.800 81.690 89.435 ;
        RECT 84.080 88.800 85.690 89.435 ;
        RECT 88.080 88.800 89.690 89.435 ;
        RECT 92.080 88.800 93.690 89.435 ;
        RECT 96.080 88.800 97.690 89.435 ;
        RECT 100.080 88.800 101.690 89.435 ;
        RECT 104.080 88.800 105.690 89.435 ;
        RECT 108.080 88.800 109.690 89.435 ;
        RECT 112.080 88.800 113.690 89.435 ;
        RECT 116.080 88.800 117.690 89.435 ;
        RECT 120.080 88.800 121.690 89.435 ;
        RECT 124.080 88.800 125.690 89.435 ;
        RECT 128.080 88.800 129.690 89.435 ;
        RECT 132.080 88.800 133.690 89.435 ;
        RECT 136.080 88.800 137.690 89.435 ;
        RECT 140.080 88.800 141.690 89.435 ;
        RECT 8.080 88.500 141.690 88.800 ;
        RECT 8.080 87.825 9.690 88.500 ;
        RECT 12.080 87.825 13.690 88.500 ;
        RECT 16.080 87.825 17.690 88.500 ;
        RECT 20.080 87.825 21.690 88.500 ;
        RECT 24.080 87.825 25.690 88.500 ;
        RECT 28.080 87.825 29.690 88.500 ;
        RECT 32.080 87.825 33.690 88.500 ;
        RECT 36.080 87.825 37.690 88.500 ;
        RECT 40.080 87.825 41.690 88.500 ;
        RECT 44.080 87.825 45.690 88.500 ;
        RECT 48.080 87.825 49.690 88.500 ;
        RECT 52.080 87.825 53.690 88.500 ;
        RECT 56.080 87.825 57.690 88.500 ;
        RECT 60.080 87.825 61.690 88.500 ;
        RECT 64.080 87.825 65.690 88.500 ;
        RECT 68.080 87.825 69.690 88.500 ;
        RECT 72.080 87.825 73.690 88.500 ;
        RECT 76.080 87.825 77.690 88.500 ;
        RECT 80.080 87.825 81.690 88.500 ;
        RECT 84.080 87.825 85.690 88.500 ;
        RECT 88.080 87.825 89.690 88.500 ;
        RECT 92.080 87.825 93.690 88.500 ;
        RECT 96.080 87.825 97.690 88.500 ;
        RECT 100.080 87.825 101.690 88.500 ;
        RECT 104.080 87.825 105.690 88.500 ;
        RECT 108.080 87.825 109.690 88.500 ;
        RECT 112.080 87.825 113.690 88.500 ;
        RECT 116.080 87.825 117.690 88.500 ;
        RECT 120.080 87.825 121.690 88.500 ;
        RECT 124.080 87.825 125.690 88.500 ;
        RECT 128.080 87.825 129.690 88.500 ;
        RECT 132.080 87.825 133.690 88.500 ;
        RECT 136.080 87.825 137.690 88.500 ;
        RECT 140.080 87.825 141.690 88.500 ;
        RECT 8.660 86.435 8.960 87.825 ;
        RECT 140.790 86.435 141.090 87.825 ;
        RECT 8.080 86.140 9.690 86.435 ;
        RECT 12.080 86.140 13.690 86.435 ;
        RECT 16.080 86.140 17.690 86.435 ;
        RECT 20.080 86.140 21.690 86.435 ;
        RECT 24.080 86.140 25.690 86.435 ;
        RECT 28.080 86.140 29.690 86.435 ;
        RECT 32.080 86.140 33.690 86.435 ;
        RECT 36.080 86.140 37.690 86.435 ;
        RECT 40.080 86.140 41.690 86.435 ;
        RECT 44.080 86.140 45.690 86.435 ;
        RECT 48.080 86.140 49.690 86.435 ;
        RECT 52.080 86.140 53.690 86.435 ;
        RECT 56.080 86.140 57.690 86.435 ;
        RECT 60.080 86.140 61.690 86.435 ;
        RECT 64.080 86.140 65.690 86.435 ;
        RECT 68.080 86.140 69.690 86.435 ;
        RECT 72.080 86.140 73.690 86.435 ;
        RECT 76.080 86.140 77.690 86.435 ;
        RECT 80.080 86.140 81.690 86.435 ;
        RECT 84.080 86.140 85.690 86.435 ;
        RECT 88.080 86.140 89.690 86.435 ;
        RECT 92.080 86.140 93.690 86.435 ;
        RECT 96.080 86.140 97.690 86.435 ;
        RECT 100.080 86.140 101.690 86.435 ;
        RECT 104.080 86.140 105.690 86.435 ;
        RECT 108.080 86.140 109.690 86.435 ;
        RECT 112.080 86.140 113.690 86.435 ;
        RECT 116.080 86.140 117.690 86.435 ;
        RECT 120.080 86.140 121.690 86.435 ;
        RECT 124.080 86.140 125.690 86.435 ;
        RECT 128.080 86.140 129.690 86.435 ;
        RECT 132.080 86.140 133.690 86.435 ;
        RECT 136.080 86.140 137.690 86.435 ;
        RECT 8.080 85.840 137.690 86.140 ;
        RECT 8.080 84.825 9.690 85.840 ;
        RECT 12.080 84.825 13.690 85.840 ;
        RECT 16.080 84.825 17.690 85.840 ;
        RECT 20.080 84.825 21.690 85.840 ;
        RECT 24.080 84.825 25.690 85.840 ;
        RECT 28.080 84.825 29.690 85.840 ;
        RECT 32.080 84.825 33.690 85.840 ;
        RECT 36.080 84.825 37.690 85.840 ;
        RECT 40.080 84.825 41.690 85.840 ;
        RECT 44.080 84.825 45.690 85.840 ;
        RECT 48.080 84.825 49.690 85.840 ;
        RECT 52.080 84.825 53.690 85.840 ;
        RECT 56.080 84.825 57.690 85.840 ;
        RECT 60.080 84.825 61.690 85.840 ;
        RECT 64.080 84.825 65.690 85.840 ;
        RECT 68.080 84.825 69.690 85.840 ;
        RECT 72.080 84.825 73.690 85.840 ;
        RECT 76.080 84.825 77.690 85.840 ;
        RECT 80.080 84.825 81.690 85.840 ;
        RECT 84.080 84.825 85.690 85.840 ;
        RECT 88.080 84.825 89.690 85.840 ;
        RECT 92.080 84.825 93.690 85.840 ;
        RECT 96.080 84.825 97.690 85.840 ;
        RECT 100.080 84.825 101.690 85.840 ;
        RECT 104.080 84.825 105.690 85.840 ;
        RECT 108.080 84.825 109.690 85.840 ;
        RECT 112.080 84.825 113.690 85.840 ;
        RECT 116.080 84.825 117.690 85.840 ;
        RECT 120.080 84.825 121.690 85.840 ;
        RECT 124.080 84.825 125.690 85.840 ;
        RECT 128.080 84.825 129.690 85.840 ;
        RECT 132.080 84.825 133.690 85.840 ;
        RECT 136.080 84.825 137.690 85.840 ;
        RECT 140.080 84.825 141.690 86.435 ;
        RECT 8.660 83.435 8.960 84.825 ;
        RECT 140.790 83.435 141.090 84.825 ;
        RECT 8.080 83.140 9.690 83.435 ;
        RECT 12.080 83.140 13.690 83.435 ;
        RECT 16.080 83.140 17.690 83.435 ;
        RECT 20.080 83.140 21.690 83.435 ;
        RECT 24.080 83.140 25.690 83.435 ;
        RECT 28.080 83.140 29.690 83.435 ;
        RECT 32.080 83.140 33.690 83.435 ;
        RECT 36.080 83.140 37.690 83.435 ;
        RECT 40.080 83.140 41.690 83.435 ;
        RECT 44.080 83.140 45.690 83.435 ;
        RECT 48.080 83.140 49.690 83.435 ;
        RECT 52.080 83.140 53.690 83.435 ;
        RECT 56.080 83.140 57.690 83.435 ;
        RECT 60.080 83.140 61.690 83.435 ;
        RECT 64.080 83.140 65.690 83.435 ;
        RECT 68.080 83.140 69.690 83.435 ;
        RECT 72.080 83.140 73.690 83.435 ;
        RECT 76.080 83.140 77.690 83.435 ;
        RECT 80.080 83.140 81.690 83.435 ;
        RECT 84.080 83.140 85.690 83.435 ;
        RECT 88.080 83.140 89.690 83.435 ;
        RECT 92.080 83.140 93.690 83.435 ;
        RECT 96.080 83.140 97.690 83.435 ;
        RECT 100.080 83.140 101.690 83.435 ;
        RECT 104.080 83.140 105.690 83.435 ;
        RECT 108.080 83.140 109.690 83.435 ;
        RECT 112.080 83.140 113.690 83.435 ;
        RECT 116.080 83.140 117.690 83.435 ;
        RECT 120.080 83.140 121.690 83.435 ;
        RECT 124.080 83.140 125.690 83.435 ;
        RECT 128.080 83.140 129.690 83.435 ;
        RECT 132.080 83.140 133.690 83.435 ;
        RECT 136.080 83.140 137.690 83.435 ;
        RECT 8.080 82.840 137.690 83.140 ;
        RECT 8.080 81.825 9.690 82.840 ;
        RECT 12.080 81.825 13.690 82.840 ;
        RECT 16.080 81.825 17.690 82.840 ;
        RECT 20.080 81.825 21.690 82.840 ;
        RECT 24.080 81.825 25.690 82.840 ;
        RECT 28.080 81.825 29.690 82.840 ;
        RECT 32.080 81.825 33.690 82.840 ;
        RECT 36.080 81.825 37.690 82.840 ;
        RECT 40.080 81.825 41.690 82.840 ;
        RECT 44.080 81.825 45.690 82.840 ;
        RECT 48.080 81.825 49.690 82.840 ;
        RECT 52.080 81.825 53.690 82.840 ;
        RECT 56.080 81.825 57.690 82.840 ;
        RECT 60.080 81.825 61.690 82.840 ;
        RECT 64.080 81.825 65.690 82.840 ;
        RECT 68.080 81.825 69.690 82.840 ;
        RECT 72.080 81.825 73.690 82.840 ;
        RECT 76.080 81.825 77.690 82.840 ;
        RECT 80.080 81.825 81.690 82.840 ;
        RECT 84.080 81.825 85.690 82.840 ;
        RECT 88.080 81.825 89.690 82.840 ;
        RECT 92.080 81.825 93.690 82.840 ;
        RECT 96.080 81.825 97.690 82.840 ;
        RECT 100.080 81.825 101.690 82.840 ;
        RECT 104.080 81.825 105.690 82.840 ;
        RECT 108.080 81.825 109.690 82.840 ;
        RECT 112.080 81.825 113.690 82.840 ;
        RECT 116.080 81.825 117.690 82.840 ;
        RECT 120.080 81.825 121.690 82.840 ;
        RECT 124.080 81.825 125.690 82.840 ;
        RECT 128.080 81.825 129.690 82.840 ;
        RECT 132.080 81.825 133.690 82.840 ;
        RECT 136.080 81.825 137.690 82.840 ;
        RECT 140.080 81.825 141.690 83.435 ;
        RECT 8.660 80.435 8.960 81.825 ;
        RECT 140.790 80.435 141.090 81.825 ;
        RECT 8.080 80.090 9.690 80.435 ;
        RECT 12.080 80.090 13.690 80.435 ;
        RECT 16.080 80.090 17.690 80.435 ;
        RECT 20.080 80.090 21.690 80.435 ;
        RECT 24.080 80.090 25.690 80.435 ;
        RECT 28.080 80.090 29.690 80.435 ;
        RECT 32.080 80.090 33.690 80.435 ;
        RECT 36.080 80.090 37.690 80.435 ;
        RECT 40.080 80.090 41.690 80.435 ;
        RECT 44.080 80.090 45.690 80.435 ;
        RECT 48.080 80.090 49.690 80.435 ;
        RECT 52.080 80.090 53.690 80.435 ;
        RECT 56.080 80.090 57.690 80.435 ;
        RECT 60.080 80.090 61.690 80.435 ;
        RECT 64.080 80.090 65.690 80.435 ;
        RECT 68.080 80.090 69.690 80.435 ;
        RECT 72.080 80.090 73.690 80.435 ;
        RECT 76.080 80.090 77.690 80.435 ;
        RECT 80.080 80.090 81.690 80.435 ;
        RECT 84.080 80.090 85.690 80.435 ;
        RECT 88.080 80.090 89.690 80.435 ;
        RECT 92.080 80.090 93.690 80.435 ;
        RECT 96.080 80.090 97.690 80.435 ;
        RECT 100.080 80.090 101.690 80.435 ;
        RECT 104.080 80.090 105.690 80.435 ;
        RECT 108.080 80.090 109.690 80.435 ;
        RECT 112.080 80.090 113.690 80.435 ;
        RECT 116.080 80.090 117.690 80.435 ;
        RECT 120.080 80.090 121.690 80.435 ;
        RECT 124.080 80.090 125.690 80.435 ;
        RECT 128.080 80.090 129.690 80.435 ;
        RECT 132.080 80.090 133.690 80.435 ;
        RECT 136.080 80.090 137.690 80.435 ;
        RECT 8.080 79.790 137.690 80.090 ;
        RECT 8.080 78.825 9.690 79.790 ;
        RECT 12.080 78.825 13.690 79.790 ;
        RECT 16.080 78.825 17.690 79.790 ;
        RECT 20.080 78.825 21.690 79.790 ;
        RECT 24.080 78.825 25.690 79.790 ;
        RECT 28.080 78.825 29.690 79.790 ;
        RECT 32.080 78.825 33.690 79.790 ;
        RECT 36.080 78.825 37.690 79.790 ;
        RECT 40.080 78.825 41.690 79.790 ;
        RECT 44.080 78.825 45.690 79.790 ;
        RECT 48.080 78.825 49.690 79.790 ;
        RECT 52.080 78.825 53.690 79.790 ;
        RECT 56.080 78.825 57.690 79.790 ;
        RECT 60.080 78.825 61.690 79.790 ;
        RECT 64.080 78.825 65.690 79.790 ;
        RECT 68.080 78.825 69.690 79.790 ;
        RECT 72.080 78.825 73.690 79.790 ;
        RECT 76.080 78.825 77.690 79.790 ;
        RECT 80.080 78.825 81.690 79.790 ;
        RECT 84.080 78.825 85.690 79.790 ;
        RECT 88.080 78.825 89.690 79.790 ;
        RECT 92.080 78.825 93.690 79.790 ;
        RECT 96.080 78.825 97.690 79.790 ;
        RECT 100.080 78.825 101.690 79.790 ;
        RECT 104.080 78.825 105.690 79.790 ;
        RECT 108.080 78.825 109.690 79.790 ;
        RECT 112.080 78.825 113.690 79.790 ;
        RECT 116.080 78.825 117.690 79.790 ;
        RECT 120.080 78.825 121.690 79.790 ;
        RECT 124.080 78.825 125.690 79.790 ;
        RECT 128.080 78.825 129.690 79.790 ;
        RECT 132.080 78.825 133.690 79.790 ;
        RECT 136.080 78.825 137.690 79.790 ;
        RECT 140.080 78.825 141.690 80.435 ;
        RECT 8.660 77.435 8.960 78.825 ;
        RECT 140.790 77.435 141.090 78.825 ;
        RECT 8.080 77.180 9.690 77.435 ;
        RECT 12.080 77.180 13.690 77.435 ;
        RECT 16.080 77.180 17.690 77.435 ;
        RECT 20.080 77.180 21.690 77.435 ;
        RECT 24.080 77.180 25.690 77.435 ;
        RECT 28.080 77.180 29.690 77.435 ;
        RECT 32.080 77.180 33.690 77.435 ;
        RECT 36.080 77.180 37.690 77.435 ;
        RECT 40.080 77.180 41.690 77.435 ;
        RECT 44.080 77.180 45.690 77.435 ;
        RECT 48.080 77.180 49.690 77.435 ;
        RECT 52.080 77.180 53.690 77.435 ;
        RECT 56.080 77.180 57.690 77.435 ;
        RECT 60.080 77.180 61.690 77.435 ;
        RECT 64.080 77.180 65.690 77.435 ;
        RECT 68.080 77.180 69.690 77.435 ;
        RECT 72.080 77.180 73.690 77.435 ;
        RECT 76.080 77.180 77.690 77.435 ;
        RECT 80.080 77.180 81.690 77.435 ;
        RECT 84.080 77.180 85.690 77.435 ;
        RECT 88.080 77.180 89.690 77.435 ;
        RECT 92.080 77.180 93.690 77.435 ;
        RECT 96.080 77.180 97.690 77.435 ;
        RECT 100.080 77.180 101.690 77.435 ;
        RECT 104.080 77.180 105.690 77.435 ;
        RECT 108.080 77.180 109.690 77.435 ;
        RECT 112.080 77.180 113.690 77.435 ;
        RECT 116.080 77.180 117.690 77.435 ;
        RECT 120.080 77.180 121.690 77.435 ;
        RECT 124.080 77.180 125.690 77.435 ;
        RECT 128.080 77.180 129.690 77.435 ;
        RECT 132.080 77.180 133.690 77.435 ;
        RECT 136.080 77.180 137.690 77.435 ;
        RECT 8.080 76.880 137.690 77.180 ;
        RECT 8.080 75.825 9.690 76.880 ;
        RECT 12.080 75.825 13.690 76.880 ;
        RECT 16.080 75.825 17.690 76.880 ;
        RECT 20.080 75.825 21.690 76.880 ;
        RECT 24.080 75.825 25.690 76.880 ;
        RECT 28.080 75.825 29.690 76.880 ;
        RECT 32.080 75.825 33.690 76.880 ;
        RECT 36.080 75.825 37.690 76.880 ;
        RECT 40.080 75.825 41.690 76.880 ;
        RECT 44.080 75.825 45.690 76.880 ;
        RECT 48.080 75.825 49.690 76.880 ;
        RECT 52.080 75.825 53.690 76.880 ;
        RECT 56.080 75.825 57.690 76.880 ;
        RECT 60.080 75.825 61.690 76.880 ;
        RECT 64.080 75.825 65.690 76.880 ;
        RECT 68.080 75.825 69.690 76.880 ;
        RECT 72.080 75.825 73.690 76.880 ;
        RECT 76.080 75.825 77.690 76.880 ;
        RECT 80.080 75.825 81.690 76.880 ;
        RECT 84.080 75.825 85.690 76.880 ;
        RECT 88.080 75.825 89.690 76.880 ;
        RECT 92.080 75.825 93.690 76.880 ;
        RECT 96.080 75.825 97.690 76.880 ;
        RECT 100.080 75.825 101.690 76.880 ;
        RECT 104.080 75.825 105.690 76.880 ;
        RECT 108.080 75.825 109.690 76.880 ;
        RECT 112.080 75.825 113.690 76.880 ;
        RECT 116.080 75.825 117.690 76.880 ;
        RECT 120.080 75.825 121.690 76.880 ;
        RECT 124.080 75.825 125.690 76.880 ;
        RECT 128.080 75.825 129.690 76.880 ;
        RECT 132.080 75.825 133.690 76.880 ;
        RECT 136.080 75.825 137.690 76.880 ;
        RECT 140.080 75.825 141.690 77.435 ;
        RECT 8.660 74.435 8.960 75.825 ;
        RECT 140.790 74.435 141.090 75.825 ;
        RECT 8.080 74.180 9.690 74.435 ;
        RECT 12.080 74.180 13.690 74.435 ;
        RECT 16.080 74.180 17.690 74.435 ;
        RECT 20.080 74.180 21.690 74.435 ;
        RECT 24.080 74.180 25.690 74.435 ;
        RECT 28.080 74.180 29.690 74.435 ;
        RECT 32.080 74.180 33.690 74.435 ;
        RECT 36.080 74.180 37.690 74.435 ;
        RECT 40.080 74.180 41.690 74.435 ;
        RECT 44.080 74.180 45.690 74.435 ;
        RECT 48.080 74.180 49.690 74.435 ;
        RECT 52.080 74.180 53.690 74.435 ;
        RECT 56.080 74.180 57.690 74.435 ;
        RECT 60.080 74.180 61.690 74.435 ;
        RECT 64.080 74.180 65.690 74.435 ;
        RECT 68.080 74.180 69.690 74.435 ;
        RECT 72.080 74.180 73.690 74.435 ;
        RECT 76.080 74.180 77.690 74.435 ;
        RECT 80.080 74.180 81.690 74.435 ;
        RECT 84.080 74.180 85.690 74.435 ;
        RECT 88.080 74.180 89.690 74.435 ;
        RECT 92.080 74.180 93.690 74.435 ;
        RECT 96.080 74.180 97.690 74.435 ;
        RECT 100.080 74.180 101.690 74.435 ;
        RECT 104.080 74.180 105.690 74.435 ;
        RECT 108.080 74.180 109.690 74.435 ;
        RECT 112.080 74.180 113.690 74.435 ;
        RECT 116.080 74.180 117.690 74.435 ;
        RECT 120.080 74.180 121.690 74.435 ;
        RECT 124.080 74.180 125.690 74.435 ;
        RECT 128.080 74.180 129.690 74.435 ;
        RECT 132.080 74.180 133.690 74.435 ;
        RECT 136.080 74.180 137.690 74.435 ;
        RECT 8.080 73.880 137.690 74.180 ;
        RECT 8.080 72.825 9.690 73.880 ;
        RECT 12.080 72.825 13.690 73.880 ;
        RECT 16.080 72.825 17.690 73.880 ;
        RECT 20.080 72.825 21.690 73.880 ;
        RECT 24.080 72.825 25.690 73.880 ;
        RECT 28.080 72.825 29.690 73.880 ;
        RECT 32.080 72.825 33.690 73.880 ;
        RECT 36.080 72.825 37.690 73.880 ;
        RECT 40.080 72.825 41.690 73.880 ;
        RECT 44.080 72.825 45.690 73.880 ;
        RECT 48.080 72.825 49.690 73.880 ;
        RECT 52.080 72.825 53.690 73.880 ;
        RECT 56.080 72.825 57.690 73.880 ;
        RECT 60.080 72.825 61.690 73.880 ;
        RECT 64.080 72.825 65.690 73.880 ;
        RECT 68.080 72.825 69.690 73.880 ;
        RECT 72.080 72.825 73.690 73.880 ;
        RECT 76.080 72.825 77.690 73.880 ;
        RECT 80.080 72.825 81.690 73.880 ;
        RECT 84.080 72.825 85.690 73.880 ;
        RECT 88.080 72.825 89.690 73.880 ;
        RECT 92.080 72.825 93.690 73.880 ;
        RECT 96.080 72.825 97.690 73.880 ;
        RECT 100.080 72.825 101.690 73.880 ;
        RECT 104.080 72.825 105.690 73.880 ;
        RECT 108.080 72.825 109.690 73.880 ;
        RECT 112.080 72.825 113.690 73.880 ;
        RECT 116.080 72.825 117.690 73.880 ;
        RECT 120.080 72.825 121.690 73.880 ;
        RECT 124.080 72.825 125.690 73.880 ;
        RECT 128.080 72.825 129.690 73.880 ;
        RECT 132.080 72.825 133.690 73.880 ;
        RECT 136.080 72.825 137.690 73.880 ;
        RECT 140.080 72.825 141.690 74.435 ;
        RECT 148.645 73.265 149.195 74.735 ;
        RECT 8.660 71.435 8.960 72.825 ;
        RECT 22.755 71.470 23.115 71.830 ;
        RECT 8.080 71.080 9.690 71.435 ;
        RECT 12.080 71.080 13.690 71.435 ;
        RECT 16.080 71.080 17.690 71.435 ;
        RECT 20.080 71.080 21.690 71.435 ;
        RECT 22.785 71.080 23.085 71.470 ;
        RECT 140.790 71.435 141.090 72.825 ;
        RECT 148.130 71.655 149.740 73.265 ;
        RECT 151.675 73.245 152.225 74.715 ;
        RECT 154.685 73.275 155.235 74.745 ;
        RECT 151.160 71.635 152.770 73.245 ;
        RECT 154.170 71.665 155.780 73.275 ;
        RECT 157.715 73.255 158.265 74.725 ;
        RECT 160.685 73.275 161.235 74.745 ;
        RECT 163.725 73.280 164.275 74.750 ;
        RECT 166.725 73.285 167.275 74.755 ;
        RECT 157.200 71.645 158.810 73.255 ;
        RECT 160.170 71.665 161.780 73.275 ;
        RECT 163.210 71.670 164.820 73.280 ;
        RECT 166.210 71.675 167.820 73.285 ;
        RECT 169.755 73.265 170.305 74.735 ;
        RECT 169.240 71.655 170.850 73.265 ;
        RECT 24.080 71.080 25.690 71.435 ;
        RECT 28.080 71.080 29.690 71.435 ;
        RECT 32.080 71.080 33.690 71.435 ;
        RECT 36.080 71.080 37.690 71.435 ;
        RECT 40.080 71.080 41.690 71.435 ;
        RECT 44.080 71.080 45.690 71.435 ;
        RECT 48.080 71.080 49.690 71.435 ;
        RECT 52.080 71.080 53.690 71.435 ;
        RECT 56.080 71.080 57.690 71.435 ;
        RECT 60.080 71.080 61.690 71.435 ;
        RECT 64.080 71.080 65.690 71.435 ;
        RECT 68.080 71.080 69.690 71.435 ;
        RECT 72.080 71.080 73.690 71.435 ;
        RECT 76.080 71.080 77.690 71.435 ;
        RECT 80.080 71.080 81.690 71.435 ;
        RECT 84.080 71.080 85.690 71.435 ;
        RECT 88.080 71.080 89.690 71.435 ;
        RECT 92.080 71.080 93.690 71.435 ;
        RECT 96.080 71.080 97.690 71.435 ;
        RECT 100.080 71.080 101.690 71.435 ;
        RECT 104.080 71.080 105.690 71.435 ;
        RECT 108.080 71.080 109.690 71.435 ;
        RECT 112.080 71.080 113.690 71.435 ;
        RECT 116.080 71.080 117.690 71.435 ;
        RECT 120.080 71.080 121.690 71.435 ;
        RECT 124.080 71.080 125.690 71.435 ;
        RECT 128.080 71.080 129.690 71.435 ;
        RECT 132.080 71.080 133.690 71.435 ;
        RECT 136.080 71.080 137.690 71.435 ;
        RECT 8.080 70.780 137.690 71.080 ;
        RECT 8.080 69.825 9.690 70.780 ;
        RECT 12.080 69.825 13.690 70.780 ;
        RECT 16.080 69.825 17.690 70.780 ;
        RECT 20.080 69.825 21.690 70.780 ;
        RECT 24.080 69.825 25.690 70.780 ;
        RECT 28.080 69.825 29.690 70.780 ;
        RECT 32.080 69.825 33.690 70.780 ;
        RECT 36.080 69.825 37.690 70.780 ;
        RECT 40.080 69.825 41.690 70.780 ;
        RECT 44.080 69.825 45.690 70.780 ;
        RECT 48.080 69.825 49.690 70.780 ;
        RECT 52.080 69.825 53.690 70.780 ;
        RECT 56.080 69.825 57.690 70.780 ;
        RECT 60.080 69.825 61.690 70.780 ;
        RECT 64.080 69.825 65.690 70.780 ;
        RECT 68.080 69.825 69.690 70.780 ;
        RECT 72.080 69.825 73.690 70.780 ;
        RECT 76.080 69.825 77.690 70.780 ;
        RECT 80.080 69.825 81.690 70.780 ;
        RECT 84.080 69.825 85.690 70.780 ;
        RECT 88.080 69.825 89.690 70.780 ;
        RECT 92.080 69.825 93.690 70.780 ;
        RECT 96.080 69.825 97.690 70.780 ;
        RECT 100.080 69.825 101.690 70.780 ;
        RECT 104.080 69.825 105.690 70.780 ;
        RECT 108.080 69.825 109.690 70.780 ;
        RECT 112.080 69.825 113.690 70.780 ;
        RECT 116.080 69.825 117.690 70.780 ;
        RECT 120.080 69.825 121.690 70.780 ;
        RECT 124.080 69.825 125.690 70.780 ;
        RECT 128.080 69.825 129.690 70.780 ;
        RECT 132.080 69.825 133.690 70.780 ;
        RECT 136.080 69.825 137.690 70.780 ;
        RECT 140.080 69.825 141.690 71.435 ;
        RECT 8.660 68.435 8.960 69.825 ;
        RECT 140.790 68.435 141.090 69.825 ;
        RECT 8.080 68.240 9.690 68.435 ;
        RECT 12.080 68.240 13.690 68.435 ;
        RECT 16.080 68.240 17.690 68.435 ;
        RECT 20.080 68.240 21.690 68.435 ;
        RECT 24.080 68.240 25.690 68.435 ;
        RECT 28.080 68.240 29.690 68.435 ;
        RECT 32.080 68.240 33.690 68.435 ;
        RECT 36.080 68.240 37.690 68.435 ;
        RECT 40.080 68.240 41.690 68.435 ;
        RECT 44.080 68.240 45.690 68.435 ;
        RECT 48.080 68.240 49.690 68.435 ;
        RECT 52.080 68.240 53.690 68.435 ;
        RECT 56.080 68.240 57.690 68.435 ;
        RECT 60.080 68.240 61.690 68.435 ;
        RECT 64.080 68.240 65.690 68.435 ;
        RECT 68.080 68.240 69.690 68.435 ;
        RECT 72.080 68.240 73.690 68.435 ;
        RECT 76.080 68.240 77.690 68.435 ;
        RECT 80.080 68.240 81.690 68.435 ;
        RECT 84.080 68.240 85.690 68.435 ;
        RECT 88.080 68.240 89.690 68.435 ;
        RECT 92.080 68.240 93.690 68.435 ;
        RECT 96.080 68.240 97.690 68.435 ;
        RECT 100.080 68.240 101.690 68.435 ;
        RECT 104.080 68.240 105.690 68.435 ;
        RECT 108.080 68.240 109.690 68.435 ;
        RECT 112.080 68.240 113.690 68.435 ;
        RECT 116.080 68.240 117.690 68.435 ;
        RECT 120.080 68.240 121.690 68.435 ;
        RECT 124.080 68.240 125.690 68.435 ;
        RECT 128.080 68.240 129.690 68.435 ;
        RECT 132.080 68.240 133.690 68.435 ;
        RECT 136.080 68.240 137.690 68.435 ;
        RECT 8.080 67.940 137.690 68.240 ;
        RECT 8.080 66.825 9.690 67.940 ;
        RECT 12.080 66.825 13.690 67.940 ;
        RECT 16.080 66.825 17.690 67.940 ;
        RECT 20.080 66.825 21.690 67.940 ;
        RECT 24.080 66.825 25.690 67.940 ;
        RECT 28.080 66.825 29.690 67.940 ;
        RECT 32.080 66.825 33.690 67.940 ;
        RECT 36.080 66.825 37.690 67.940 ;
        RECT 40.080 66.825 41.690 67.940 ;
        RECT 44.080 66.825 45.690 67.940 ;
        RECT 48.080 66.825 49.690 67.940 ;
        RECT 52.080 66.825 53.690 67.940 ;
        RECT 56.080 66.825 57.690 67.940 ;
        RECT 60.080 66.825 61.690 67.940 ;
        RECT 64.080 66.825 65.690 67.940 ;
        RECT 68.080 66.825 69.690 67.940 ;
        RECT 72.080 66.825 73.690 67.940 ;
        RECT 76.080 66.825 77.690 67.940 ;
        RECT 80.080 66.825 81.690 67.940 ;
        RECT 84.080 66.825 85.690 67.940 ;
        RECT 88.080 66.825 89.690 67.940 ;
        RECT 92.080 66.825 93.690 67.940 ;
        RECT 96.080 66.825 97.690 67.940 ;
        RECT 100.080 66.825 101.690 67.940 ;
        RECT 104.080 66.825 105.690 67.940 ;
        RECT 108.080 66.825 109.690 67.940 ;
        RECT 112.080 66.825 113.690 67.940 ;
        RECT 116.080 66.825 117.690 67.940 ;
        RECT 120.080 66.825 121.690 67.940 ;
        RECT 124.080 66.825 125.690 67.940 ;
        RECT 128.080 66.825 129.690 67.940 ;
        RECT 132.080 66.825 133.690 67.940 ;
        RECT 136.080 66.825 137.690 67.940 ;
        RECT 140.080 66.825 141.690 68.435 ;
        RECT 8.660 65.435 8.960 66.825 ;
        RECT 140.790 65.435 141.090 66.825 ;
        RECT 8.080 65.170 9.690 65.435 ;
        RECT 12.080 65.170 13.690 65.435 ;
        RECT 16.080 65.170 17.690 65.435 ;
        RECT 20.080 65.170 21.690 65.435 ;
        RECT 24.080 65.170 25.690 65.435 ;
        RECT 28.080 65.170 29.690 65.435 ;
        RECT 32.080 65.170 33.690 65.435 ;
        RECT 36.080 65.170 37.690 65.435 ;
        RECT 40.080 65.170 41.690 65.435 ;
        RECT 44.080 65.170 45.690 65.435 ;
        RECT 48.080 65.170 49.690 65.435 ;
        RECT 52.080 65.170 53.690 65.435 ;
        RECT 56.080 65.170 57.690 65.435 ;
        RECT 60.080 65.170 61.690 65.435 ;
        RECT 64.080 65.170 65.690 65.435 ;
        RECT 68.080 65.170 69.690 65.435 ;
        RECT 72.080 65.170 73.690 65.435 ;
        RECT 76.080 65.170 77.690 65.435 ;
        RECT 80.080 65.170 81.690 65.435 ;
        RECT 84.080 65.170 85.690 65.435 ;
        RECT 88.080 65.170 89.690 65.435 ;
        RECT 92.080 65.170 93.690 65.435 ;
        RECT 96.080 65.170 97.690 65.435 ;
        RECT 100.080 65.170 101.690 65.435 ;
        RECT 104.080 65.170 105.690 65.435 ;
        RECT 108.080 65.170 109.690 65.435 ;
        RECT 112.080 65.170 113.690 65.435 ;
        RECT 116.080 65.170 117.690 65.435 ;
        RECT 120.080 65.170 121.690 65.435 ;
        RECT 124.080 65.170 125.690 65.435 ;
        RECT 128.080 65.170 129.690 65.435 ;
        RECT 132.080 65.170 133.690 65.435 ;
        RECT 136.080 65.170 137.690 65.435 ;
        RECT 8.080 64.870 137.690 65.170 ;
        RECT 8.080 63.825 9.690 64.870 ;
        RECT 12.080 63.825 13.690 64.870 ;
        RECT 16.080 63.825 17.690 64.870 ;
        RECT 20.080 63.825 21.690 64.870 ;
        RECT 24.080 63.825 25.690 64.870 ;
        RECT 28.080 63.825 29.690 64.870 ;
        RECT 32.080 63.825 33.690 64.870 ;
        RECT 36.080 63.825 37.690 64.870 ;
        RECT 40.080 63.825 41.690 64.870 ;
        RECT 44.080 63.825 45.690 64.870 ;
        RECT 48.080 63.825 49.690 64.870 ;
        RECT 52.080 63.825 53.690 64.870 ;
        RECT 56.080 63.825 57.690 64.870 ;
        RECT 60.080 63.825 61.690 64.870 ;
        RECT 64.080 63.825 65.690 64.870 ;
        RECT 68.080 63.825 69.690 64.870 ;
        RECT 72.080 63.825 73.690 64.870 ;
        RECT 76.080 63.825 77.690 64.870 ;
        RECT 80.080 63.825 81.690 64.870 ;
        RECT 84.080 63.825 85.690 64.870 ;
        RECT 88.080 63.825 89.690 64.870 ;
        RECT 92.080 63.825 93.690 64.870 ;
        RECT 96.080 63.825 97.690 64.870 ;
        RECT 100.080 63.825 101.690 64.870 ;
        RECT 104.080 63.825 105.690 64.870 ;
        RECT 108.080 63.825 109.690 64.870 ;
        RECT 112.080 63.825 113.690 64.870 ;
        RECT 116.080 63.825 117.690 64.870 ;
        RECT 120.080 63.825 121.690 64.870 ;
        RECT 124.080 63.825 125.690 64.870 ;
        RECT 128.080 63.825 129.690 64.870 ;
        RECT 132.080 63.825 133.690 64.870 ;
        RECT 136.080 63.825 137.690 64.870 ;
        RECT 140.080 63.825 141.690 65.435 ;
        RECT 148.165 64.060 149.775 65.670 ;
        RECT 151.195 64.080 152.805 65.690 ;
        RECT 8.660 62.435 8.960 63.825 ;
        RECT 140.790 62.435 141.090 63.825 ;
        RECT 148.680 62.590 149.230 64.060 ;
        RECT 151.710 62.610 152.260 64.080 ;
        RECT 154.205 64.050 155.815 65.660 ;
        RECT 157.235 64.070 158.845 65.680 ;
        RECT 154.720 62.580 155.270 64.050 ;
        RECT 157.750 62.600 158.300 64.070 ;
        RECT 160.205 64.050 161.815 65.660 ;
        RECT 163.235 64.070 164.845 65.680 ;
        RECT 160.720 62.580 161.270 64.050 ;
        RECT 163.750 62.600 164.300 64.070 ;
        RECT 166.245 64.040 167.855 65.650 ;
        RECT 169.275 64.060 170.885 65.670 ;
        RECT 166.760 62.570 167.310 64.040 ;
        RECT 169.790 62.590 170.340 64.060 ;
        RECT 8.080 61.840 9.690 62.435 ;
        RECT 12.080 61.840 13.690 62.435 ;
        RECT 16.080 61.840 17.690 62.435 ;
        RECT 20.080 61.840 21.690 62.435 ;
        RECT 24.080 61.840 25.690 62.435 ;
        RECT 28.080 61.840 29.690 62.435 ;
        RECT 32.080 61.840 33.690 62.435 ;
        RECT 36.080 61.840 37.690 62.435 ;
        RECT 40.080 61.840 41.690 62.435 ;
        RECT 44.080 61.840 45.690 62.435 ;
        RECT 48.080 61.840 49.690 62.435 ;
        RECT 52.080 61.840 53.690 62.435 ;
        RECT 56.080 61.840 57.690 62.435 ;
        RECT 60.080 61.840 61.690 62.435 ;
        RECT 64.080 61.840 65.690 62.435 ;
        RECT 68.080 61.840 69.690 62.435 ;
        RECT 72.080 61.840 73.690 62.435 ;
        RECT 76.080 61.840 77.690 62.435 ;
        RECT 80.080 61.840 81.690 62.435 ;
        RECT 84.080 61.840 85.690 62.435 ;
        RECT 88.080 61.840 89.690 62.435 ;
        RECT 92.080 61.840 93.690 62.435 ;
        RECT 96.080 61.840 97.690 62.435 ;
        RECT 100.080 61.840 101.690 62.435 ;
        RECT 104.080 61.840 105.690 62.435 ;
        RECT 108.080 61.840 109.690 62.435 ;
        RECT 112.080 61.840 113.690 62.435 ;
        RECT 116.080 61.840 117.690 62.435 ;
        RECT 120.080 61.840 121.690 62.435 ;
        RECT 124.080 61.840 125.690 62.435 ;
        RECT 128.080 61.840 129.690 62.435 ;
        RECT 132.080 61.840 133.690 62.435 ;
        RECT 136.080 61.840 137.690 62.435 ;
        RECT 140.080 61.840 141.690 62.435 ;
        RECT 152.020 61.905 152.350 62.235 ;
        RECT 8.080 61.540 141.690 61.840 ;
        RECT 8.080 60.825 9.690 61.540 ;
        RECT 12.080 60.825 13.690 61.540 ;
        RECT 16.080 60.825 17.690 61.540 ;
        RECT 20.080 60.825 21.690 61.540 ;
        RECT 24.080 60.825 25.690 61.540 ;
        RECT 28.080 60.825 29.690 61.540 ;
        RECT 32.080 60.825 33.690 61.540 ;
        RECT 36.080 60.825 37.690 61.540 ;
        RECT 40.080 60.825 41.690 61.540 ;
        RECT 44.080 60.825 45.690 61.540 ;
        RECT 48.080 60.825 49.690 61.540 ;
        RECT 52.080 60.825 53.690 61.540 ;
        RECT 56.080 60.825 57.690 61.540 ;
        RECT 60.080 60.825 61.690 61.540 ;
        RECT 64.080 60.825 65.690 61.540 ;
        RECT 68.080 60.825 69.690 61.540 ;
        RECT 72.080 60.825 73.690 61.540 ;
        RECT 76.080 60.825 77.690 61.540 ;
        RECT 80.080 60.825 81.690 61.540 ;
        RECT 84.080 60.825 85.690 61.540 ;
        RECT 88.080 60.825 89.690 61.540 ;
        RECT 92.080 60.825 93.690 61.540 ;
        RECT 96.080 60.825 97.690 61.540 ;
        RECT 100.080 60.825 101.690 61.540 ;
        RECT 104.080 60.825 105.690 61.540 ;
        RECT 108.080 60.825 109.690 61.540 ;
        RECT 112.080 60.825 113.690 61.540 ;
        RECT 116.080 60.825 117.690 61.540 ;
        RECT 120.080 60.825 121.690 61.540 ;
        RECT 124.080 60.825 125.690 61.540 ;
        RECT 128.080 60.825 129.690 61.540 ;
        RECT 132.080 60.825 133.690 61.540 ;
        RECT 136.080 60.825 137.690 61.540 ;
        RECT 138.965 60.400 139.265 61.540 ;
        RECT 140.080 60.825 141.690 61.540 ;
        RECT 152.035 60.400 152.335 61.905 ;
        RECT 138.965 60.100 152.345 60.400 ;
        RECT 156.220 59.690 156.550 59.705 ;
        RECT 138.965 59.390 156.550 59.690 ;
        RECT 8.080 58.310 9.690 59.025 ;
        RECT 12.080 58.310 13.690 59.025 ;
        RECT 16.080 58.310 17.690 59.025 ;
        RECT 20.080 58.310 21.690 59.025 ;
        RECT 24.080 58.310 25.690 59.025 ;
        RECT 28.080 58.310 29.690 59.025 ;
        RECT 32.080 58.310 33.690 59.025 ;
        RECT 36.080 58.310 37.690 59.025 ;
        RECT 40.080 58.310 41.690 59.025 ;
        RECT 44.080 58.310 45.690 59.025 ;
        RECT 48.080 58.310 49.690 59.025 ;
        RECT 52.080 58.310 53.690 59.025 ;
        RECT 56.080 58.310 57.690 59.025 ;
        RECT 60.080 58.310 61.690 59.025 ;
        RECT 64.080 58.310 65.690 59.025 ;
        RECT 68.080 58.310 69.690 59.025 ;
        RECT 72.080 58.310 73.690 59.025 ;
        RECT 76.080 58.310 77.690 59.025 ;
        RECT 80.080 58.310 81.690 59.025 ;
        RECT 84.080 58.310 85.690 59.025 ;
        RECT 88.080 58.310 89.690 59.025 ;
        RECT 92.080 58.310 93.690 59.025 ;
        RECT 96.080 58.310 97.690 59.025 ;
        RECT 100.080 58.310 101.690 59.025 ;
        RECT 104.080 58.310 105.690 59.025 ;
        RECT 108.080 58.310 109.690 59.025 ;
        RECT 112.080 58.310 113.690 59.025 ;
        RECT 116.080 58.310 117.690 59.025 ;
        RECT 120.080 58.310 121.690 59.025 ;
        RECT 124.080 58.310 125.690 59.025 ;
        RECT 128.080 58.310 129.690 59.025 ;
        RECT 132.080 58.310 133.690 59.025 ;
        RECT 136.080 58.310 137.690 59.025 ;
        RECT 138.965 58.310 139.265 59.390 ;
        RECT 156.220 59.375 156.550 59.390 ;
        RECT 140.080 58.310 141.690 59.025 ;
        RECT 8.080 58.010 141.690 58.310 ;
        RECT 8.080 57.415 9.690 58.010 ;
        RECT 12.080 57.415 13.690 58.010 ;
        RECT 16.080 57.415 17.690 58.010 ;
        RECT 20.080 57.415 21.690 58.010 ;
        RECT 24.080 57.415 25.690 58.010 ;
        RECT 28.080 57.415 29.690 58.010 ;
        RECT 32.080 57.415 33.690 58.010 ;
        RECT 36.080 57.415 37.690 58.010 ;
        RECT 40.080 57.415 41.690 58.010 ;
        RECT 44.080 57.415 45.690 58.010 ;
        RECT 48.080 57.415 49.690 58.010 ;
        RECT 52.080 57.415 53.690 58.010 ;
        RECT 56.080 57.415 57.690 58.010 ;
        RECT 60.080 57.415 61.690 58.010 ;
        RECT 64.080 57.415 65.690 58.010 ;
        RECT 68.080 57.415 69.690 58.010 ;
        RECT 72.080 57.415 73.690 58.010 ;
        RECT 76.080 57.415 77.690 58.010 ;
        RECT 80.080 57.415 81.690 58.010 ;
        RECT 84.080 57.415 85.690 58.010 ;
        RECT 88.080 57.415 89.690 58.010 ;
        RECT 92.080 57.415 93.690 58.010 ;
        RECT 96.080 57.415 97.690 58.010 ;
        RECT 100.080 57.415 101.690 58.010 ;
        RECT 104.080 57.415 105.690 58.010 ;
        RECT 108.080 57.415 109.690 58.010 ;
        RECT 112.080 57.415 113.690 58.010 ;
        RECT 116.080 57.415 117.690 58.010 ;
        RECT 120.080 57.415 121.690 58.010 ;
        RECT 124.080 57.415 125.690 58.010 ;
        RECT 128.080 57.415 129.690 58.010 ;
        RECT 132.080 57.415 133.690 58.010 ;
        RECT 136.080 57.415 137.690 58.010 ;
        RECT 140.080 57.415 141.690 58.010 ;
        RECT 8.660 56.025 8.960 57.415 ;
        RECT 140.790 56.025 141.090 57.415 ;
        RECT 8.080 54.980 9.690 56.025 ;
        RECT 12.080 54.980 13.690 56.025 ;
        RECT 16.080 54.980 17.690 56.025 ;
        RECT 20.080 54.980 21.690 56.025 ;
        RECT 24.080 54.980 25.690 56.025 ;
        RECT 28.080 54.980 29.690 56.025 ;
        RECT 32.080 54.980 33.690 56.025 ;
        RECT 36.080 54.980 37.690 56.025 ;
        RECT 40.080 54.980 41.690 56.025 ;
        RECT 44.080 54.980 45.690 56.025 ;
        RECT 48.080 54.980 49.690 56.025 ;
        RECT 52.080 54.980 53.690 56.025 ;
        RECT 56.080 54.980 57.690 56.025 ;
        RECT 60.080 54.980 61.690 56.025 ;
        RECT 64.080 54.980 65.690 56.025 ;
        RECT 68.080 54.980 69.690 56.025 ;
        RECT 72.080 54.980 73.690 56.025 ;
        RECT 76.080 54.980 77.690 56.025 ;
        RECT 80.080 54.980 81.690 56.025 ;
        RECT 84.080 54.980 85.690 56.025 ;
        RECT 88.080 54.980 89.690 56.025 ;
        RECT 92.080 54.980 93.690 56.025 ;
        RECT 96.080 54.980 97.690 56.025 ;
        RECT 100.080 54.980 101.690 56.025 ;
        RECT 104.080 54.980 105.690 56.025 ;
        RECT 108.080 54.980 109.690 56.025 ;
        RECT 112.080 54.980 113.690 56.025 ;
        RECT 116.080 54.980 117.690 56.025 ;
        RECT 120.080 54.980 121.690 56.025 ;
        RECT 124.080 54.980 125.690 56.025 ;
        RECT 128.080 54.980 129.690 56.025 ;
        RECT 132.080 54.980 133.690 56.025 ;
        RECT 136.080 54.980 137.690 56.025 ;
        RECT 8.080 54.680 137.690 54.980 ;
        RECT 8.080 54.415 9.690 54.680 ;
        RECT 12.080 54.415 13.690 54.680 ;
        RECT 16.080 54.415 17.690 54.680 ;
        RECT 20.080 54.415 21.690 54.680 ;
        RECT 24.080 54.415 25.690 54.680 ;
        RECT 28.080 54.415 29.690 54.680 ;
        RECT 32.080 54.415 33.690 54.680 ;
        RECT 36.080 54.415 37.690 54.680 ;
        RECT 40.080 54.415 41.690 54.680 ;
        RECT 44.080 54.415 45.690 54.680 ;
        RECT 48.080 54.415 49.690 54.680 ;
        RECT 52.080 54.415 53.690 54.680 ;
        RECT 56.080 54.415 57.690 54.680 ;
        RECT 60.080 54.415 61.690 54.680 ;
        RECT 64.080 54.415 65.690 54.680 ;
        RECT 68.080 54.415 69.690 54.680 ;
        RECT 72.080 54.415 73.690 54.680 ;
        RECT 76.080 54.415 77.690 54.680 ;
        RECT 80.080 54.415 81.690 54.680 ;
        RECT 84.080 54.415 85.690 54.680 ;
        RECT 88.080 54.415 89.690 54.680 ;
        RECT 92.080 54.415 93.690 54.680 ;
        RECT 96.080 54.415 97.690 54.680 ;
        RECT 100.080 54.415 101.690 54.680 ;
        RECT 104.080 54.415 105.690 54.680 ;
        RECT 108.080 54.415 109.690 54.680 ;
        RECT 112.080 54.415 113.690 54.680 ;
        RECT 116.080 54.415 117.690 54.680 ;
        RECT 120.080 54.415 121.690 54.680 ;
        RECT 124.080 54.415 125.690 54.680 ;
        RECT 128.080 54.415 129.690 54.680 ;
        RECT 132.080 54.415 133.690 54.680 ;
        RECT 136.080 54.415 137.690 54.680 ;
        RECT 140.080 54.415 141.690 56.025 ;
        RECT 148.795 55.920 149.345 57.390 ;
        RECT 8.660 53.025 8.960 54.415 ;
        RECT 140.790 53.025 141.090 54.415 ;
        RECT 148.280 54.310 149.890 55.920 ;
        RECT 151.825 55.900 152.375 57.370 ;
        RECT 154.835 55.930 155.385 57.400 ;
        RECT 151.310 54.290 152.920 55.900 ;
        RECT 154.320 54.320 155.930 55.930 ;
        RECT 157.865 55.910 158.415 57.380 ;
        RECT 160.835 55.930 161.385 57.400 ;
        RECT 157.350 54.300 158.960 55.910 ;
        RECT 160.320 54.320 161.930 55.930 ;
        RECT 163.865 55.910 164.415 57.380 ;
        RECT 166.875 55.940 167.425 57.410 ;
        RECT 163.350 54.300 164.960 55.910 ;
        RECT 166.360 54.330 167.970 55.940 ;
        RECT 169.905 55.920 170.455 57.390 ;
        RECT 169.390 54.310 171.000 55.920 ;
        RECT 8.080 51.910 9.690 53.025 ;
        RECT 12.080 51.910 13.690 53.025 ;
        RECT 16.080 51.910 17.690 53.025 ;
        RECT 20.080 51.910 21.690 53.025 ;
        RECT 24.080 51.910 25.690 53.025 ;
        RECT 28.080 51.910 29.690 53.025 ;
        RECT 32.080 51.910 33.690 53.025 ;
        RECT 36.080 51.910 37.690 53.025 ;
        RECT 40.080 51.910 41.690 53.025 ;
        RECT 44.080 51.910 45.690 53.025 ;
        RECT 48.080 51.910 49.690 53.025 ;
        RECT 52.080 51.910 53.690 53.025 ;
        RECT 56.080 51.910 57.690 53.025 ;
        RECT 60.080 51.910 61.690 53.025 ;
        RECT 64.080 51.910 65.690 53.025 ;
        RECT 68.080 51.910 69.690 53.025 ;
        RECT 72.080 51.910 73.690 53.025 ;
        RECT 76.080 51.910 77.690 53.025 ;
        RECT 80.080 51.910 81.690 53.025 ;
        RECT 84.080 51.910 85.690 53.025 ;
        RECT 88.080 51.910 89.690 53.025 ;
        RECT 92.080 51.910 93.690 53.025 ;
        RECT 96.080 51.910 97.690 53.025 ;
        RECT 100.080 51.910 101.690 53.025 ;
        RECT 104.080 51.910 105.690 53.025 ;
        RECT 108.080 51.910 109.690 53.025 ;
        RECT 112.080 51.910 113.690 53.025 ;
        RECT 116.080 51.910 117.690 53.025 ;
        RECT 120.080 51.910 121.690 53.025 ;
        RECT 124.080 51.910 125.690 53.025 ;
        RECT 128.080 51.910 129.690 53.025 ;
        RECT 132.080 51.910 133.690 53.025 ;
        RECT 136.080 51.910 137.690 53.025 ;
        RECT 8.080 51.610 137.690 51.910 ;
        RECT 8.080 51.415 9.690 51.610 ;
        RECT 12.080 51.415 13.690 51.610 ;
        RECT 16.080 51.415 17.690 51.610 ;
        RECT 20.080 51.415 21.690 51.610 ;
        RECT 24.080 51.415 25.690 51.610 ;
        RECT 28.080 51.415 29.690 51.610 ;
        RECT 32.080 51.415 33.690 51.610 ;
        RECT 36.080 51.415 37.690 51.610 ;
        RECT 40.080 51.415 41.690 51.610 ;
        RECT 44.080 51.415 45.690 51.610 ;
        RECT 48.080 51.415 49.690 51.610 ;
        RECT 52.080 51.415 53.690 51.610 ;
        RECT 56.080 51.415 57.690 51.610 ;
        RECT 60.080 51.415 61.690 51.610 ;
        RECT 64.080 51.415 65.690 51.610 ;
        RECT 68.080 51.415 69.690 51.610 ;
        RECT 72.080 51.415 73.690 51.610 ;
        RECT 76.080 51.415 77.690 51.610 ;
        RECT 80.080 51.415 81.690 51.610 ;
        RECT 84.080 51.415 85.690 51.610 ;
        RECT 88.080 51.415 89.690 51.610 ;
        RECT 92.080 51.415 93.690 51.610 ;
        RECT 96.080 51.415 97.690 51.610 ;
        RECT 100.080 51.415 101.690 51.610 ;
        RECT 104.080 51.415 105.690 51.610 ;
        RECT 108.080 51.415 109.690 51.610 ;
        RECT 112.080 51.415 113.690 51.610 ;
        RECT 116.080 51.415 117.690 51.610 ;
        RECT 120.080 51.415 121.690 51.610 ;
        RECT 124.080 51.415 125.690 51.610 ;
        RECT 128.080 51.415 129.690 51.610 ;
        RECT 132.080 51.415 133.690 51.610 ;
        RECT 136.080 51.415 137.690 51.610 ;
        RECT 140.080 51.415 141.690 53.025 ;
        RECT 8.660 50.025 8.960 51.415 ;
        RECT 140.790 50.025 141.090 51.415 ;
        RECT 8.080 49.070 9.690 50.025 ;
        RECT 12.080 49.070 13.690 50.025 ;
        RECT 16.080 49.070 17.690 50.025 ;
        RECT 20.080 49.070 21.690 50.025 ;
        RECT 24.080 49.070 25.690 50.025 ;
        RECT 28.080 49.070 29.690 50.025 ;
        RECT 32.080 49.070 33.690 50.025 ;
        RECT 36.080 49.070 37.690 50.025 ;
        RECT 40.080 49.070 41.690 50.025 ;
        RECT 44.080 49.070 45.690 50.025 ;
        RECT 48.080 49.070 49.690 50.025 ;
        RECT 52.080 49.070 53.690 50.025 ;
        RECT 56.080 49.070 57.690 50.025 ;
        RECT 60.080 49.070 61.690 50.025 ;
        RECT 64.080 49.070 65.690 50.025 ;
        RECT 68.080 49.070 69.690 50.025 ;
        RECT 72.080 49.070 73.690 50.025 ;
        RECT 76.080 49.070 77.690 50.025 ;
        RECT 80.080 49.070 81.690 50.025 ;
        RECT 84.080 49.070 85.690 50.025 ;
        RECT 88.080 49.070 89.690 50.025 ;
        RECT 92.080 49.070 93.690 50.025 ;
        RECT 96.080 49.070 97.690 50.025 ;
        RECT 100.080 49.070 101.690 50.025 ;
        RECT 104.080 49.070 105.690 50.025 ;
        RECT 108.080 49.070 109.690 50.025 ;
        RECT 112.080 49.070 113.690 50.025 ;
        RECT 116.080 49.070 117.690 50.025 ;
        RECT 120.080 49.070 121.690 50.025 ;
        RECT 124.080 49.070 125.690 50.025 ;
        RECT 128.080 49.070 129.690 50.025 ;
        RECT 132.080 49.070 133.690 50.025 ;
        RECT 136.080 49.070 137.690 50.025 ;
        RECT 8.080 48.770 137.690 49.070 ;
        RECT 8.080 48.415 9.690 48.770 ;
        RECT 12.080 48.415 13.690 48.770 ;
        RECT 16.080 48.415 17.690 48.770 ;
        RECT 20.080 48.415 21.690 48.770 ;
        RECT 8.660 47.025 8.960 48.415 ;
        RECT 22.785 48.380 23.085 48.770 ;
        RECT 24.080 48.415 25.690 48.770 ;
        RECT 28.080 48.415 29.690 48.770 ;
        RECT 32.080 48.415 33.690 48.770 ;
        RECT 36.080 48.415 37.690 48.770 ;
        RECT 40.080 48.415 41.690 48.770 ;
        RECT 44.080 48.415 45.690 48.770 ;
        RECT 48.080 48.415 49.690 48.770 ;
        RECT 52.080 48.415 53.690 48.770 ;
        RECT 56.080 48.415 57.690 48.770 ;
        RECT 60.080 48.415 61.690 48.770 ;
        RECT 64.080 48.415 65.690 48.770 ;
        RECT 68.080 48.415 69.690 48.770 ;
        RECT 72.080 48.415 73.690 48.770 ;
        RECT 76.080 48.415 77.690 48.770 ;
        RECT 80.080 48.415 81.690 48.770 ;
        RECT 84.080 48.415 85.690 48.770 ;
        RECT 88.080 48.415 89.690 48.770 ;
        RECT 92.080 48.415 93.690 48.770 ;
        RECT 96.080 48.415 97.690 48.770 ;
        RECT 100.080 48.415 101.690 48.770 ;
        RECT 104.080 48.415 105.690 48.770 ;
        RECT 108.080 48.415 109.690 48.770 ;
        RECT 112.080 48.415 113.690 48.770 ;
        RECT 116.080 48.415 117.690 48.770 ;
        RECT 120.080 48.415 121.690 48.770 ;
        RECT 124.080 48.415 125.690 48.770 ;
        RECT 128.080 48.415 129.690 48.770 ;
        RECT 132.080 48.415 133.690 48.770 ;
        RECT 136.080 48.415 137.690 48.770 ;
        RECT 140.080 48.415 141.690 50.025 ;
        RECT 22.755 48.020 23.115 48.380 ;
        RECT 140.790 47.025 141.090 48.415 ;
        RECT 8.080 45.970 9.690 47.025 ;
        RECT 12.080 45.970 13.690 47.025 ;
        RECT 16.080 45.970 17.690 47.025 ;
        RECT 20.080 45.970 21.690 47.025 ;
        RECT 24.080 45.970 25.690 47.025 ;
        RECT 28.080 45.970 29.690 47.025 ;
        RECT 32.080 45.970 33.690 47.025 ;
        RECT 36.080 45.970 37.690 47.025 ;
        RECT 40.080 45.970 41.690 47.025 ;
        RECT 44.080 45.970 45.690 47.025 ;
        RECT 48.080 45.970 49.690 47.025 ;
        RECT 52.080 45.970 53.690 47.025 ;
        RECT 56.080 45.970 57.690 47.025 ;
        RECT 60.080 45.970 61.690 47.025 ;
        RECT 64.080 45.970 65.690 47.025 ;
        RECT 68.080 45.970 69.690 47.025 ;
        RECT 72.080 45.970 73.690 47.025 ;
        RECT 76.080 45.970 77.690 47.025 ;
        RECT 80.080 45.970 81.690 47.025 ;
        RECT 84.080 45.970 85.690 47.025 ;
        RECT 88.080 45.970 89.690 47.025 ;
        RECT 92.080 45.970 93.690 47.025 ;
        RECT 96.080 45.970 97.690 47.025 ;
        RECT 100.080 45.970 101.690 47.025 ;
        RECT 104.080 45.970 105.690 47.025 ;
        RECT 108.080 45.970 109.690 47.025 ;
        RECT 112.080 45.970 113.690 47.025 ;
        RECT 116.080 45.970 117.690 47.025 ;
        RECT 120.080 45.970 121.690 47.025 ;
        RECT 124.080 45.970 125.690 47.025 ;
        RECT 128.080 45.970 129.690 47.025 ;
        RECT 132.080 45.970 133.690 47.025 ;
        RECT 136.080 45.970 137.690 47.025 ;
        RECT 8.080 45.670 137.690 45.970 ;
        RECT 8.080 45.415 9.690 45.670 ;
        RECT 12.080 45.415 13.690 45.670 ;
        RECT 16.080 45.415 17.690 45.670 ;
        RECT 20.080 45.415 21.690 45.670 ;
        RECT 24.080 45.415 25.690 45.670 ;
        RECT 28.080 45.415 29.690 45.670 ;
        RECT 32.080 45.415 33.690 45.670 ;
        RECT 36.080 45.415 37.690 45.670 ;
        RECT 40.080 45.415 41.690 45.670 ;
        RECT 44.080 45.415 45.690 45.670 ;
        RECT 48.080 45.415 49.690 45.670 ;
        RECT 52.080 45.415 53.690 45.670 ;
        RECT 56.080 45.415 57.690 45.670 ;
        RECT 60.080 45.415 61.690 45.670 ;
        RECT 64.080 45.415 65.690 45.670 ;
        RECT 68.080 45.415 69.690 45.670 ;
        RECT 72.080 45.415 73.690 45.670 ;
        RECT 76.080 45.415 77.690 45.670 ;
        RECT 80.080 45.415 81.690 45.670 ;
        RECT 84.080 45.415 85.690 45.670 ;
        RECT 88.080 45.415 89.690 45.670 ;
        RECT 92.080 45.415 93.690 45.670 ;
        RECT 96.080 45.415 97.690 45.670 ;
        RECT 100.080 45.415 101.690 45.670 ;
        RECT 104.080 45.415 105.690 45.670 ;
        RECT 108.080 45.415 109.690 45.670 ;
        RECT 112.080 45.415 113.690 45.670 ;
        RECT 116.080 45.415 117.690 45.670 ;
        RECT 120.080 45.415 121.690 45.670 ;
        RECT 124.080 45.415 125.690 45.670 ;
        RECT 128.080 45.415 129.690 45.670 ;
        RECT 132.080 45.415 133.690 45.670 ;
        RECT 136.080 45.415 137.690 45.670 ;
        RECT 140.080 45.415 141.690 47.025 ;
        RECT 148.245 46.715 149.855 48.325 ;
        RECT 151.275 46.735 152.885 48.345 ;
        RECT 8.660 44.025 8.960 45.415 ;
        RECT 140.790 44.025 141.090 45.415 ;
        RECT 148.760 45.245 149.310 46.715 ;
        RECT 151.790 45.265 152.340 46.735 ;
        RECT 154.285 46.705 155.895 48.315 ;
        RECT 157.315 46.725 158.925 48.335 ;
        RECT 154.800 45.235 155.350 46.705 ;
        RECT 157.830 45.255 158.380 46.725 ;
        RECT 160.285 46.705 161.895 48.315 ;
        RECT 160.800 45.235 161.350 46.705 ;
        RECT 163.325 46.700 164.935 48.310 ;
        RECT 163.840 45.230 164.390 46.700 ;
        RECT 166.325 46.695 167.935 48.305 ;
        RECT 169.355 46.715 170.965 48.325 ;
        RECT 166.840 45.225 167.390 46.695 ;
        RECT 169.870 45.245 170.420 46.715 ;
        RECT 8.080 42.970 9.690 44.025 ;
        RECT 12.080 42.970 13.690 44.025 ;
        RECT 16.080 42.970 17.690 44.025 ;
        RECT 20.080 42.970 21.690 44.025 ;
        RECT 24.080 42.970 25.690 44.025 ;
        RECT 28.080 42.970 29.690 44.025 ;
        RECT 32.080 42.970 33.690 44.025 ;
        RECT 36.080 42.970 37.690 44.025 ;
        RECT 40.080 42.970 41.690 44.025 ;
        RECT 44.080 42.970 45.690 44.025 ;
        RECT 48.080 42.970 49.690 44.025 ;
        RECT 52.080 42.970 53.690 44.025 ;
        RECT 56.080 42.970 57.690 44.025 ;
        RECT 60.080 42.970 61.690 44.025 ;
        RECT 64.080 42.970 65.690 44.025 ;
        RECT 68.080 42.970 69.690 44.025 ;
        RECT 72.080 42.970 73.690 44.025 ;
        RECT 76.080 42.970 77.690 44.025 ;
        RECT 80.080 42.970 81.690 44.025 ;
        RECT 84.080 42.970 85.690 44.025 ;
        RECT 88.080 42.970 89.690 44.025 ;
        RECT 92.080 42.970 93.690 44.025 ;
        RECT 96.080 42.970 97.690 44.025 ;
        RECT 100.080 42.970 101.690 44.025 ;
        RECT 104.080 42.970 105.690 44.025 ;
        RECT 108.080 42.970 109.690 44.025 ;
        RECT 112.080 42.970 113.690 44.025 ;
        RECT 116.080 42.970 117.690 44.025 ;
        RECT 120.080 42.970 121.690 44.025 ;
        RECT 124.080 42.970 125.690 44.025 ;
        RECT 128.080 42.970 129.690 44.025 ;
        RECT 132.080 42.970 133.690 44.025 ;
        RECT 136.080 42.970 137.690 44.025 ;
        RECT 8.080 42.670 137.690 42.970 ;
        RECT 8.080 42.415 9.690 42.670 ;
        RECT 12.080 42.415 13.690 42.670 ;
        RECT 16.080 42.415 17.690 42.670 ;
        RECT 20.080 42.415 21.690 42.670 ;
        RECT 24.080 42.415 25.690 42.670 ;
        RECT 28.080 42.415 29.690 42.670 ;
        RECT 32.080 42.415 33.690 42.670 ;
        RECT 36.080 42.415 37.690 42.670 ;
        RECT 40.080 42.415 41.690 42.670 ;
        RECT 44.080 42.415 45.690 42.670 ;
        RECT 48.080 42.415 49.690 42.670 ;
        RECT 52.080 42.415 53.690 42.670 ;
        RECT 56.080 42.415 57.690 42.670 ;
        RECT 60.080 42.415 61.690 42.670 ;
        RECT 64.080 42.415 65.690 42.670 ;
        RECT 68.080 42.415 69.690 42.670 ;
        RECT 72.080 42.415 73.690 42.670 ;
        RECT 76.080 42.415 77.690 42.670 ;
        RECT 80.080 42.415 81.690 42.670 ;
        RECT 84.080 42.415 85.690 42.670 ;
        RECT 88.080 42.415 89.690 42.670 ;
        RECT 92.080 42.415 93.690 42.670 ;
        RECT 96.080 42.415 97.690 42.670 ;
        RECT 100.080 42.415 101.690 42.670 ;
        RECT 104.080 42.415 105.690 42.670 ;
        RECT 108.080 42.415 109.690 42.670 ;
        RECT 112.080 42.415 113.690 42.670 ;
        RECT 116.080 42.415 117.690 42.670 ;
        RECT 120.080 42.415 121.690 42.670 ;
        RECT 124.080 42.415 125.690 42.670 ;
        RECT 128.080 42.415 129.690 42.670 ;
        RECT 132.080 42.415 133.690 42.670 ;
        RECT 136.080 42.415 137.690 42.670 ;
        RECT 140.080 42.415 141.690 44.025 ;
        RECT 8.660 41.025 8.960 42.415 ;
        RECT 140.790 41.025 141.090 42.415 ;
        RECT 8.080 40.060 9.690 41.025 ;
        RECT 12.080 40.060 13.690 41.025 ;
        RECT 16.080 40.060 17.690 41.025 ;
        RECT 20.080 40.060 21.690 41.025 ;
        RECT 24.080 40.060 25.690 41.025 ;
        RECT 28.080 40.060 29.690 41.025 ;
        RECT 32.080 40.060 33.690 41.025 ;
        RECT 36.080 40.060 37.690 41.025 ;
        RECT 40.080 40.060 41.690 41.025 ;
        RECT 44.080 40.060 45.690 41.025 ;
        RECT 48.080 40.060 49.690 41.025 ;
        RECT 52.080 40.060 53.690 41.025 ;
        RECT 56.080 40.060 57.690 41.025 ;
        RECT 60.080 40.060 61.690 41.025 ;
        RECT 64.080 40.060 65.690 41.025 ;
        RECT 68.080 40.060 69.690 41.025 ;
        RECT 72.080 40.060 73.690 41.025 ;
        RECT 76.080 40.060 77.690 41.025 ;
        RECT 80.080 40.060 81.690 41.025 ;
        RECT 84.080 40.060 85.690 41.025 ;
        RECT 88.080 40.060 89.690 41.025 ;
        RECT 92.080 40.060 93.690 41.025 ;
        RECT 96.080 40.060 97.690 41.025 ;
        RECT 100.080 40.060 101.690 41.025 ;
        RECT 104.080 40.060 105.690 41.025 ;
        RECT 108.080 40.060 109.690 41.025 ;
        RECT 112.080 40.060 113.690 41.025 ;
        RECT 116.080 40.060 117.690 41.025 ;
        RECT 120.080 40.060 121.690 41.025 ;
        RECT 124.080 40.060 125.690 41.025 ;
        RECT 128.080 40.060 129.690 41.025 ;
        RECT 132.080 40.060 133.690 41.025 ;
        RECT 136.080 40.060 137.690 41.025 ;
        RECT 8.080 39.760 137.690 40.060 ;
        RECT 8.080 39.415 9.690 39.760 ;
        RECT 12.080 39.415 13.690 39.760 ;
        RECT 16.080 39.415 17.690 39.760 ;
        RECT 20.080 39.415 21.690 39.760 ;
        RECT 24.080 39.415 25.690 39.760 ;
        RECT 28.080 39.415 29.690 39.760 ;
        RECT 32.080 39.415 33.690 39.760 ;
        RECT 36.080 39.415 37.690 39.760 ;
        RECT 40.080 39.415 41.690 39.760 ;
        RECT 44.080 39.415 45.690 39.760 ;
        RECT 48.080 39.415 49.690 39.760 ;
        RECT 52.080 39.415 53.690 39.760 ;
        RECT 56.080 39.415 57.690 39.760 ;
        RECT 60.080 39.415 61.690 39.760 ;
        RECT 64.080 39.415 65.690 39.760 ;
        RECT 68.080 39.415 69.690 39.760 ;
        RECT 72.080 39.415 73.690 39.760 ;
        RECT 76.080 39.415 77.690 39.760 ;
        RECT 80.080 39.415 81.690 39.760 ;
        RECT 84.080 39.415 85.690 39.760 ;
        RECT 88.080 39.415 89.690 39.760 ;
        RECT 92.080 39.415 93.690 39.760 ;
        RECT 96.080 39.415 97.690 39.760 ;
        RECT 100.080 39.415 101.690 39.760 ;
        RECT 104.080 39.415 105.690 39.760 ;
        RECT 108.080 39.415 109.690 39.760 ;
        RECT 112.080 39.415 113.690 39.760 ;
        RECT 116.080 39.415 117.690 39.760 ;
        RECT 120.080 39.415 121.690 39.760 ;
        RECT 124.080 39.415 125.690 39.760 ;
        RECT 128.080 39.415 129.690 39.760 ;
        RECT 132.080 39.415 133.690 39.760 ;
        RECT 136.080 39.415 137.690 39.760 ;
        RECT 140.080 39.415 141.690 41.025 ;
        RECT 8.660 38.025 8.960 39.415 ;
        RECT 140.790 38.025 141.090 39.415 ;
        RECT 8.080 37.010 9.690 38.025 ;
        RECT 12.080 37.010 13.690 38.025 ;
        RECT 16.080 37.010 17.690 38.025 ;
        RECT 20.080 37.010 21.690 38.025 ;
        RECT 24.080 37.010 25.690 38.025 ;
        RECT 28.080 37.010 29.690 38.025 ;
        RECT 32.080 37.010 33.690 38.025 ;
        RECT 36.080 37.010 37.690 38.025 ;
        RECT 40.080 37.010 41.690 38.025 ;
        RECT 44.080 37.010 45.690 38.025 ;
        RECT 48.080 37.010 49.690 38.025 ;
        RECT 52.080 37.010 53.690 38.025 ;
        RECT 56.080 37.010 57.690 38.025 ;
        RECT 60.080 37.010 61.690 38.025 ;
        RECT 64.080 37.010 65.690 38.025 ;
        RECT 68.080 37.010 69.690 38.025 ;
        RECT 72.080 37.010 73.690 38.025 ;
        RECT 76.080 37.010 77.690 38.025 ;
        RECT 80.080 37.010 81.690 38.025 ;
        RECT 84.080 37.010 85.690 38.025 ;
        RECT 88.080 37.010 89.690 38.025 ;
        RECT 92.080 37.010 93.690 38.025 ;
        RECT 96.080 37.010 97.690 38.025 ;
        RECT 100.080 37.010 101.690 38.025 ;
        RECT 104.080 37.010 105.690 38.025 ;
        RECT 108.080 37.010 109.690 38.025 ;
        RECT 112.080 37.010 113.690 38.025 ;
        RECT 116.080 37.010 117.690 38.025 ;
        RECT 120.080 37.010 121.690 38.025 ;
        RECT 124.080 37.010 125.690 38.025 ;
        RECT 128.080 37.010 129.690 38.025 ;
        RECT 132.080 37.010 133.690 38.025 ;
        RECT 136.080 37.010 137.690 38.025 ;
        RECT 8.080 36.710 137.690 37.010 ;
        RECT 8.080 36.415 9.690 36.710 ;
        RECT 12.080 36.415 13.690 36.710 ;
        RECT 16.080 36.415 17.690 36.710 ;
        RECT 20.080 36.415 21.690 36.710 ;
        RECT 24.080 36.415 25.690 36.710 ;
        RECT 28.080 36.415 29.690 36.710 ;
        RECT 32.080 36.415 33.690 36.710 ;
        RECT 36.080 36.415 37.690 36.710 ;
        RECT 40.080 36.415 41.690 36.710 ;
        RECT 44.080 36.415 45.690 36.710 ;
        RECT 48.080 36.415 49.690 36.710 ;
        RECT 52.080 36.415 53.690 36.710 ;
        RECT 56.080 36.415 57.690 36.710 ;
        RECT 60.080 36.415 61.690 36.710 ;
        RECT 64.080 36.415 65.690 36.710 ;
        RECT 68.080 36.415 69.690 36.710 ;
        RECT 72.080 36.415 73.690 36.710 ;
        RECT 76.080 36.415 77.690 36.710 ;
        RECT 80.080 36.415 81.690 36.710 ;
        RECT 84.080 36.415 85.690 36.710 ;
        RECT 88.080 36.415 89.690 36.710 ;
        RECT 92.080 36.415 93.690 36.710 ;
        RECT 96.080 36.415 97.690 36.710 ;
        RECT 100.080 36.415 101.690 36.710 ;
        RECT 104.080 36.415 105.690 36.710 ;
        RECT 108.080 36.415 109.690 36.710 ;
        RECT 112.080 36.415 113.690 36.710 ;
        RECT 116.080 36.415 117.690 36.710 ;
        RECT 120.080 36.415 121.690 36.710 ;
        RECT 124.080 36.415 125.690 36.710 ;
        RECT 128.080 36.415 129.690 36.710 ;
        RECT 132.080 36.415 133.690 36.710 ;
        RECT 136.080 36.415 137.690 36.710 ;
        RECT 140.080 36.415 141.690 38.025 ;
        RECT 8.660 35.025 8.960 36.415 ;
        RECT 140.790 35.025 141.090 36.415 ;
        RECT 8.080 34.010 9.690 35.025 ;
        RECT 12.080 34.010 13.690 35.025 ;
        RECT 16.080 34.010 17.690 35.025 ;
        RECT 20.080 34.010 21.690 35.025 ;
        RECT 24.080 34.010 25.690 35.025 ;
        RECT 28.080 34.010 29.690 35.025 ;
        RECT 32.080 34.010 33.690 35.025 ;
        RECT 36.080 34.010 37.690 35.025 ;
        RECT 40.080 34.010 41.690 35.025 ;
        RECT 44.080 34.010 45.690 35.025 ;
        RECT 48.080 34.010 49.690 35.025 ;
        RECT 52.080 34.010 53.690 35.025 ;
        RECT 56.080 34.010 57.690 35.025 ;
        RECT 60.080 34.010 61.690 35.025 ;
        RECT 64.080 34.010 65.690 35.025 ;
        RECT 68.080 34.010 69.690 35.025 ;
        RECT 72.080 34.010 73.690 35.025 ;
        RECT 76.080 34.010 77.690 35.025 ;
        RECT 80.080 34.010 81.690 35.025 ;
        RECT 84.080 34.010 85.690 35.025 ;
        RECT 88.080 34.010 89.690 35.025 ;
        RECT 92.080 34.010 93.690 35.025 ;
        RECT 96.080 34.010 97.690 35.025 ;
        RECT 100.080 34.010 101.690 35.025 ;
        RECT 104.080 34.010 105.690 35.025 ;
        RECT 108.080 34.010 109.690 35.025 ;
        RECT 112.080 34.010 113.690 35.025 ;
        RECT 116.080 34.010 117.690 35.025 ;
        RECT 120.080 34.010 121.690 35.025 ;
        RECT 124.080 34.010 125.690 35.025 ;
        RECT 128.080 34.010 129.690 35.025 ;
        RECT 132.080 34.010 133.690 35.025 ;
        RECT 136.080 34.010 137.690 35.025 ;
        RECT 8.080 33.710 137.690 34.010 ;
        RECT 8.080 33.415 9.690 33.710 ;
        RECT 12.080 33.415 13.690 33.710 ;
        RECT 16.080 33.415 17.690 33.710 ;
        RECT 20.080 33.415 21.690 33.710 ;
        RECT 24.080 33.415 25.690 33.710 ;
        RECT 28.080 33.415 29.690 33.710 ;
        RECT 32.080 33.415 33.690 33.710 ;
        RECT 36.080 33.415 37.690 33.710 ;
        RECT 40.080 33.415 41.690 33.710 ;
        RECT 44.080 33.415 45.690 33.710 ;
        RECT 48.080 33.415 49.690 33.710 ;
        RECT 52.080 33.415 53.690 33.710 ;
        RECT 56.080 33.415 57.690 33.710 ;
        RECT 60.080 33.415 61.690 33.710 ;
        RECT 64.080 33.415 65.690 33.710 ;
        RECT 68.080 33.415 69.690 33.710 ;
        RECT 72.080 33.415 73.690 33.710 ;
        RECT 76.080 33.415 77.690 33.710 ;
        RECT 80.080 33.415 81.690 33.710 ;
        RECT 84.080 33.415 85.690 33.710 ;
        RECT 88.080 33.415 89.690 33.710 ;
        RECT 92.080 33.415 93.690 33.710 ;
        RECT 96.080 33.415 97.690 33.710 ;
        RECT 100.080 33.415 101.690 33.710 ;
        RECT 104.080 33.415 105.690 33.710 ;
        RECT 108.080 33.415 109.690 33.710 ;
        RECT 112.080 33.415 113.690 33.710 ;
        RECT 116.080 33.415 117.690 33.710 ;
        RECT 120.080 33.415 121.690 33.710 ;
        RECT 124.080 33.415 125.690 33.710 ;
        RECT 128.080 33.415 129.690 33.710 ;
        RECT 132.080 33.415 133.690 33.710 ;
        RECT 136.080 33.415 137.690 33.710 ;
        RECT 140.080 33.415 141.690 35.025 ;
        RECT 8.660 32.025 8.960 33.415 ;
        RECT 140.790 32.025 141.090 33.415 ;
        RECT 8.080 31.350 9.690 32.025 ;
        RECT 12.080 31.350 13.690 32.025 ;
        RECT 16.080 31.350 17.690 32.025 ;
        RECT 20.080 31.350 21.690 32.025 ;
        RECT 24.080 31.350 25.690 32.025 ;
        RECT 28.080 31.350 29.690 32.025 ;
        RECT 32.080 31.350 33.690 32.025 ;
        RECT 36.080 31.350 37.690 32.025 ;
        RECT 40.080 31.350 41.690 32.025 ;
        RECT 44.080 31.350 45.690 32.025 ;
        RECT 48.080 31.350 49.690 32.025 ;
        RECT 52.080 31.350 53.690 32.025 ;
        RECT 56.080 31.350 57.690 32.025 ;
        RECT 60.080 31.350 61.690 32.025 ;
        RECT 64.080 31.350 65.690 32.025 ;
        RECT 68.080 31.350 69.690 32.025 ;
        RECT 72.080 31.350 73.690 32.025 ;
        RECT 76.080 31.350 77.690 32.025 ;
        RECT 80.080 31.350 81.690 32.025 ;
        RECT 84.080 31.350 85.690 32.025 ;
        RECT 88.080 31.350 89.690 32.025 ;
        RECT 92.080 31.350 93.690 32.025 ;
        RECT 96.080 31.350 97.690 32.025 ;
        RECT 100.080 31.350 101.690 32.025 ;
        RECT 104.080 31.350 105.690 32.025 ;
        RECT 108.080 31.350 109.690 32.025 ;
        RECT 112.080 31.350 113.690 32.025 ;
        RECT 116.080 31.350 117.690 32.025 ;
        RECT 120.080 31.350 121.690 32.025 ;
        RECT 124.080 31.350 125.690 32.025 ;
        RECT 128.080 31.350 129.690 32.025 ;
        RECT 132.080 31.350 133.690 32.025 ;
        RECT 136.080 31.350 137.690 32.025 ;
        RECT 140.080 31.350 141.690 32.025 ;
        RECT 8.080 31.050 141.690 31.350 ;
        RECT 8.080 30.415 9.690 31.050 ;
        RECT 12.080 30.415 13.690 31.050 ;
        RECT 16.080 30.415 17.690 31.050 ;
        RECT 20.080 30.415 21.690 31.050 ;
        RECT 24.080 30.415 25.690 31.050 ;
        RECT 28.080 30.415 29.690 31.050 ;
        RECT 32.080 30.415 33.690 31.050 ;
        RECT 36.080 30.415 37.690 31.050 ;
        RECT 40.080 30.415 41.690 31.050 ;
        RECT 44.080 30.415 45.690 31.050 ;
        RECT 48.080 30.415 49.690 31.050 ;
        RECT 52.080 30.415 53.690 31.050 ;
        RECT 56.080 30.415 57.690 31.050 ;
        RECT 60.080 30.415 61.690 31.050 ;
        RECT 64.080 30.415 65.690 31.050 ;
        RECT 68.080 30.415 69.690 31.050 ;
        RECT 72.080 30.415 73.690 31.050 ;
        RECT 76.080 30.415 77.690 31.050 ;
        RECT 80.080 30.415 81.690 31.050 ;
        RECT 84.080 30.415 85.690 31.050 ;
        RECT 88.080 30.415 89.690 31.050 ;
        RECT 92.080 30.415 93.690 31.050 ;
        RECT 96.080 30.415 97.690 31.050 ;
        RECT 100.080 30.415 101.690 31.050 ;
        RECT 104.080 30.415 105.690 31.050 ;
        RECT 108.080 30.415 109.690 31.050 ;
        RECT 112.080 30.415 113.690 31.050 ;
        RECT 116.080 30.415 117.690 31.050 ;
        RECT 120.080 30.415 121.690 31.050 ;
        RECT 124.080 30.415 125.690 31.050 ;
        RECT 128.080 30.415 129.690 31.050 ;
        RECT 132.080 30.415 133.690 31.050 ;
        RECT 136.080 30.415 137.690 31.050 ;
        RECT 140.080 30.415 141.690 31.050 ;
  END
END sar_analog
END LIBRARY

