VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC
  CLASS BLOCK ;
  FOREIGN DAC ;
  ORIGIN 14.155 4.275 ;
  SIZE 249.630 BY 20.910 ;
  PIN enb
    ANTENNAGATEAREA 3.990000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 223.185 47.650 223.355 47.980 ;
        RECT 223.185 47.060 223.355 47.390 ;
        RECT 223.185 46.470 223.355 46.800 ;
        RECT 231.450 46.335 231.700 47.965 ;
        RECT 223.185 45.880 223.355 46.210 ;
        RECT 231.090 45.835 232.050 46.100 ;
        RECT 231.090 45.665 231.280 45.835 ;
        RECT 223.185 45.290 223.355 45.620 ;
        RECT 230.310 45.335 231.280 45.665 ;
        RECT 223.185 44.700 223.355 45.030 ;
        RECT 231.110 44.825 231.280 45.335 ;
        RECT 230.310 44.495 231.280 44.825 ;
        RECT 231.870 45.665 232.050 45.835 ;
        RECT 231.870 45.335 232.520 45.665 ;
        RECT 231.870 44.825 232.050 45.335 ;
        RECT 231.870 44.495 232.520 44.825 ;
        RECT 223.185 44.110 223.355 44.440 ;
        RECT 223.185 43.520 223.355 43.850 ;
        RECT 223.185 42.930 223.355 43.260 ;
        RECT 223.185 42.340 223.355 42.670 ;
      LAYER mcon ;
        RECT 223.185 47.730 223.355 47.900 ;
        RECT 223.185 47.140 223.355 47.310 ;
        RECT 223.185 46.550 223.355 46.720 ;
        RECT 231.490 46.500 231.660 46.670 ;
        RECT 223.185 45.960 223.355 46.130 ;
        RECT 231.160 45.915 231.330 46.085 ;
        RECT 223.185 45.370 223.355 45.540 ;
        RECT 223.185 44.780 223.355 44.950 ;
        RECT 223.185 44.190 223.355 44.360 ;
        RECT 223.185 43.600 223.355 43.770 ;
        RECT 223.185 43.010 223.355 43.180 ;
        RECT 223.185 42.420 223.355 42.590 ;
      LAYER met1 ;
        RECT 223.155 49.220 223.855 49.520 ;
        RECT 223.155 42.360 223.385 49.220 ;
        RECT 231.425 46.150 231.725 46.765 ;
        RECT 231.085 45.850 231.725 46.150 ;
      LAYER via ;
        RECT 223.215 49.240 223.475 49.500 ;
        RECT 223.535 49.240 223.795 49.500 ;
        RECT 231.115 45.870 231.375 46.130 ;
      LAYER met2 ;
        RECT 223.205 49.520 223.805 49.570 ;
        RECT 223.205 49.220 229.670 49.520 ;
        RECT 223.205 49.170 223.805 49.220 ;
        RECT 229.370 46.150 229.670 49.220 ;
        RECT 231.115 46.150 231.375 46.160 ;
        RECT 229.370 45.850 231.410 46.150 ;
        RECT 231.115 45.840 231.375 45.850 ;
    END
    PORT
      LAYER li1 ;
        RECT 223.185 26.490 223.355 26.820 ;
        RECT 223.185 25.900 223.355 26.230 ;
        RECT 223.185 25.310 223.355 25.640 ;
        RECT 231.450 25.175 231.700 26.805 ;
        RECT 223.185 24.720 223.355 25.050 ;
        RECT 231.090 24.675 232.050 24.940 ;
        RECT 231.090 24.505 231.280 24.675 ;
        RECT 223.185 24.130 223.355 24.460 ;
        RECT 230.310 24.175 231.280 24.505 ;
        RECT 223.185 23.540 223.355 23.870 ;
        RECT 231.110 23.665 231.280 24.175 ;
        RECT 230.310 23.335 231.280 23.665 ;
        RECT 231.870 24.505 232.050 24.675 ;
        RECT 231.870 24.175 232.520 24.505 ;
        RECT 231.870 23.665 232.050 24.175 ;
        RECT 231.870 23.335 232.520 23.665 ;
        RECT 223.185 22.950 223.355 23.280 ;
        RECT 223.185 22.360 223.355 22.690 ;
        RECT 223.185 21.770 223.355 22.100 ;
        RECT 223.185 21.180 223.355 21.510 ;
      LAYER mcon ;
        RECT 223.185 26.570 223.355 26.740 ;
        RECT 223.185 25.980 223.355 26.150 ;
        RECT 223.185 25.390 223.355 25.560 ;
        RECT 231.490 25.340 231.660 25.510 ;
        RECT 223.185 24.800 223.355 24.970 ;
        RECT 231.160 24.755 231.330 24.925 ;
        RECT 223.185 24.210 223.355 24.380 ;
        RECT 223.185 23.620 223.355 23.790 ;
        RECT 223.185 23.030 223.355 23.200 ;
        RECT 223.185 22.440 223.355 22.610 ;
        RECT 223.185 21.850 223.355 22.020 ;
        RECT 223.185 21.260 223.355 21.430 ;
      LAYER met1 ;
        RECT 223.155 28.060 223.855 28.360 ;
        RECT 223.155 21.200 223.385 28.060 ;
        RECT 231.425 24.990 231.725 25.605 ;
        RECT 231.085 24.690 231.725 24.990 ;
      LAYER via ;
        RECT 223.215 28.080 223.475 28.340 ;
        RECT 223.535 28.080 223.795 28.340 ;
        RECT 231.115 24.710 231.375 24.970 ;
      LAYER met2 ;
        RECT 223.205 28.360 223.805 28.410 ;
        RECT 223.205 28.060 229.670 28.360 ;
        RECT 223.205 28.010 223.805 28.060 ;
        RECT 229.370 24.990 229.670 28.060 ;
        RECT 231.115 24.990 231.375 25.000 ;
        RECT 229.370 24.690 231.410 24.990 ;
        RECT 231.115 24.680 231.375 24.690 ;
    END
  END enb
  PIN en_buf
    ANTENNAGATEAREA 3.000000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 231.090 48.135 232.050 48.400 ;
        RECT 228.640 47.650 228.810 47.980 ;
        RECT 231.090 47.965 231.280 48.135 ;
        RECT 230.310 47.635 231.280 47.965 ;
        RECT 228.640 47.060 228.810 47.390 ;
        RECT 231.110 47.125 231.280 47.635 ;
        RECT 228.640 46.470 228.810 46.800 ;
        RECT 230.310 46.795 231.280 47.125 ;
        RECT 231.870 47.965 232.050 48.135 ;
        RECT 231.870 47.635 232.520 47.965 ;
        RECT 231.870 47.125 232.050 47.635 ;
        RECT 231.870 46.795 232.520 47.125 ;
        RECT 228.640 45.880 228.810 46.210 ;
        RECT 228.640 45.290 228.810 45.620 ;
        RECT 228.640 44.700 228.810 45.030 ;
        RECT 228.640 44.110 228.810 44.440 ;
        RECT 228.640 43.520 228.810 43.850 ;
        RECT 228.640 42.930 228.810 43.260 ;
        RECT 228.640 42.340 228.810 42.670 ;
      LAYER mcon ;
        RECT 231.160 48.215 231.330 48.385 ;
        RECT 228.640 47.730 228.810 47.900 ;
        RECT 228.640 47.140 228.810 47.310 ;
        RECT 228.640 46.550 228.810 46.720 ;
        RECT 228.640 45.960 228.810 46.130 ;
        RECT 228.640 45.370 228.810 45.540 ;
        RECT 228.640 44.780 228.810 44.950 ;
        RECT 228.640 44.190 228.810 44.360 ;
        RECT 228.640 43.600 228.810 43.770 ;
        RECT 228.640 43.010 228.810 43.180 ;
        RECT 228.640 42.420 228.810 42.590 ;
      LAYER met1 ;
        RECT 231.085 48.170 231.405 48.430 ;
        RECT 228.610 45.510 228.840 47.960 ;
        RECT 228.610 44.810 228.910 45.510 ;
        RECT 228.610 42.360 228.840 44.810 ;
      LAYER via ;
        RECT 231.115 48.170 231.375 48.430 ;
        RECT 228.630 45.190 228.890 45.450 ;
        RECT 228.630 44.870 228.890 45.130 ;
      LAYER met2 ;
        RECT 231.115 48.450 231.375 48.460 ;
        RECT 231.115 48.150 232.215 48.450 ;
        RECT 231.115 48.140 231.375 48.150 ;
        RECT 228.560 45.310 228.960 45.460 ;
        RECT 231.915 45.310 232.215 48.150 ;
        RECT 228.560 45.010 232.215 45.310 ;
        RECT 228.560 44.860 228.960 45.010 ;
    END
    PORT
      LAYER li1 ;
        RECT 231.090 26.975 232.050 27.240 ;
        RECT 228.640 26.490 228.810 26.820 ;
        RECT 231.090 26.805 231.280 26.975 ;
        RECT 230.310 26.475 231.280 26.805 ;
        RECT 228.640 25.900 228.810 26.230 ;
        RECT 231.110 25.965 231.280 26.475 ;
        RECT 228.640 25.310 228.810 25.640 ;
        RECT 230.310 25.635 231.280 25.965 ;
        RECT 231.870 26.805 232.050 26.975 ;
        RECT 231.870 26.475 232.520 26.805 ;
        RECT 231.870 25.965 232.050 26.475 ;
        RECT 231.870 25.635 232.520 25.965 ;
        RECT 228.640 24.720 228.810 25.050 ;
        RECT 228.640 24.130 228.810 24.460 ;
        RECT 228.640 23.540 228.810 23.870 ;
        RECT 228.640 22.950 228.810 23.280 ;
        RECT 228.640 22.360 228.810 22.690 ;
        RECT 228.640 21.770 228.810 22.100 ;
        RECT 228.640 21.180 228.810 21.510 ;
      LAYER mcon ;
        RECT 231.160 27.055 231.330 27.225 ;
        RECT 228.640 26.570 228.810 26.740 ;
        RECT 228.640 25.980 228.810 26.150 ;
        RECT 228.640 25.390 228.810 25.560 ;
        RECT 228.640 24.800 228.810 24.970 ;
        RECT 228.640 24.210 228.810 24.380 ;
        RECT 228.640 23.620 228.810 23.790 ;
        RECT 228.640 23.030 228.810 23.200 ;
        RECT 228.640 22.440 228.810 22.610 ;
        RECT 228.640 21.850 228.810 22.020 ;
        RECT 228.640 21.260 228.810 21.430 ;
      LAYER met1 ;
        RECT 231.085 27.010 231.405 27.270 ;
        RECT 228.610 24.350 228.840 26.800 ;
        RECT 228.610 23.650 228.910 24.350 ;
        RECT 228.610 21.200 228.840 23.650 ;
      LAYER via ;
        RECT 231.115 27.010 231.375 27.270 ;
        RECT 228.630 24.030 228.890 24.290 ;
        RECT 228.630 23.710 228.890 23.970 ;
      LAYER met2 ;
        RECT 231.115 27.290 231.375 27.300 ;
        RECT 231.115 26.990 232.215 27.290 ;
        RECT 231.115 26.980 231.375 26.990 ;
        RECT 228.560 24.150 228.960 24.300 ;
        RECT 231.915 24.150 232.215 26.990 ;
        RECT 228.560 23.850 232.215 24.150 ;
        RECT 228.560 23.700 228.960 23.850 ;
    END
  END en_buf
  PIN ctl1
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 5.790 -10.185 6.120 ;
      LAYER mcon ;
        RECT -10.400 5.910 -10.230 6.080 ;
      LAYER met1 ;
        RECT -10.445 5.835 -10.185 6.155 ;
      LAYER via ;
        RECT -10.445 5.865 -10.185 6.125 ;
      LAYER met2 ;
        RECT -14.155 5.795 -10.105 6.195 ;
    END
  END ctl1
  PIN ctl0
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 4.410 -10.185 4.740 ;
      LAYER mcon ;
        RECT -10.400 4.530 -10.230 4.700 ;
      LAYER met1 ;
        RECT -10.445 4.455 -10.185 4.775 ;
      LAYER via ;
        RECT -10.445 4.485 -10.185 4.745 ;
      LAYER met2 ;
        RECT -14.155 4.415 -10.105 4.815 ;
    END
  END ctl0
  PIN dum
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 3.030 -10.185 3.360 ;
      LAYER mcon ;
        RECT -10.400 3.150 -10.230 3.320 ;
      LAYER met1 ;
        RECT -10.445 3.075 -10.185 3.395 ;
      LAYER via ;
        RECT -10.445 3.105 -10.185 3.365 ;
      LAYER met2 ;
        RECT -14.155 3.035 -10.105 3.435 ;
    END
  END dum
  PIN ctl3
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 12.690 -10.185 13.020 ;
      LAYER mcon ;
        RECT -10.400 12.810 -10.230 12.980 ;
      LAYER met1 ;
        RECT -10.445 12.735 -10.185 13.055 ;
      LAYER via ;
        RECT -10.445 12.765 -10.185 13.025 ;
      LAYER met2 ;
        RECT -14.155 12.695 -10.105 13.095 ;
    END
  END ctl3
  PIN ctl4
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 11.310 -10.185 11.640 ;
      LAYER mcon ;
        RECT -10.400 11.430 -10.230 11.600 ;
      LAYER met1 ;
        RECT -10.445 11.355 -10.185 11.675 ;
      LAYER via ;
        RECT -10.445 11.385 -10.185 11.645 ;
      LAYER met2 ;
        RECT -14.155 11.315 -10.105 11.715 ;
    END
  END ctl4
  PIN ctl5
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 9.930 -10.185 10.260 ;
      LAYER mcon ;
        RECT -10.400 10.050 -10.230 10.220 ;
      LAYER met1 ;
        RECT -10.445 9.975 -10.185 10.295 ;
      LAYER via ;
        RECT -10.445 10.005 -10.185 10.265 ;
      LAYER met2 ;
        RECT -14.155 9.935 -10.105 10.335 ;
    END
  END ctl5
  PIN ctl6
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 8.550 -10.185 8.880 ;
      LAYER mcon ;
        RECT -10.400 8.670 -10.230 8.840 ;
      LAYER met1 ;
        RECT -10.445 8.595 -10.185 8.915 ;
      LAYER via ;
        RECT -10.445 8.625 -10.185 8.885 ;
      LAYER met2 ;
        RECT -14.155 8.555 -10.105 8.955 ;
    END
  END ctl6
  PIN ctl7
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 7.170 -10.185 7.500 ;
      LAYER mcon ;
        RECT -10.400 7.290 -10.230 7.460 ;
      LAYER met1 ;
        RECT -10.445 7.215 -10.185 7.535 ;
      LAYER via ;
        RECT -10.445 7.245 -10.185 7.505 ;
      LAYER met2 ;
        RECT -14.155 7.175 -10.105 7.575 ;
    END
  END ctl7
  PIN ctl2
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -10.435 14.070 -10.185 14.400 ;
      LAYER mcon ;
        RECT -10.400 14.190 -10.230 14.360 ;
      LAYER met1 ;
        RECT -10.445 14.115 -10.185 14.435 ;
      LAYER via ;
        RECT -10.445 14.145 -10.185 14.405 ;
      LAYER met2 ;
        RECT -14.155 14.075 -10.105 14.475 ;
    END
  END ctl2
  PIN vdd
    ANTENNAGATEAREA 7.656000 ;
    ANTENNADIFFAREA 24.308949 ;
    PORT
      LAYER nwell ;
        RECT 222.490 41.375 225.330 48.945 ;
        RECT 222.490 30.795 225.330 38.365 ;
        RECT 222.490 20.215 225.330 27.785 ;
        RECT 222.490 9.635 225.330 17.205 ;
        RECT 229.865 8.320 231.470 50.100 ;
      LAYER li1 ;
        RECT 229.970 49.825 230.140 49.910 ;
        RECT 229.970 49.305 231.770 49.825 ;
        RECT 222.670 48.595 225.150 48.765 ;
        RECT 222.670 41.725 222.840 48.595 ;
        RECT 224.980 41.725 225.150 48.595 ;
        RECT 222.670 41.555 225.150 41.725 ;
        RECT 229.970 48.615 231.230 49.305 ;
        RECT 229.970 48.345 230.140 48.615 ;
        RECT 229.970 48.135 230.600 48.345 ;
        RECT 229.970 47.465 230.140 48.135 ;
        RECT 229.970 47.295 230.940 47.465 ;
        RECT 229.970 46.625 230.140 47.295 ;
        RECT 229.970 46.360 231.280 46.625 ;
        RECT 229.970 46.045 230.140 46.360 ;
        RECT 229.970 45.835 230.600 46.045 ;
        RECT 229.970 45.165 230.140 45.835 ;
        RECT 229.970 44.995 230.940 45.165 ;
        RECT 229.970 44.325 230.140 44.995 ;
        RECT 229.970 44.060 231.280 44.325 ;
        RECT 229.970 43.845 230.140 44.060 ;
        RECT 229.970 42.155 231.750 43.845 ;
        RECT 229.970 40.335 231.230 42.155 ;
        RECT 229.970 40.165 230.140 40.335 ;
        RECT 229.970 39.415 231.305 40.165 ;
        RECT 229.970 39.245 230.140 39.415 ;
        RECT 229.970 38.725 231.770 39.245 ;
        RECT 222.670 38.015 225.150 38.185 ;
        RECT 222.670 31.145 222.840 38.015 ;
        RECT 224.980 31.145 225.150 38.015 ;
        RECT 222.670 30.975 225.150 31.145 ;
        RECT 229.970 38.035 231.230 38.725 ;
        RECT 229.970 37.765 230.140 38.035 ;
        RECT 229.970 37.555 230.600 37.765 ;
        RECT 229.970 36.885 230.140 37.555 ;
        RECT 229.970 36.715 230.940 36.885 ;
        RECT 229.970 36.045 230.140 36.715 ;
        RECT 229.970 35.780 231.280 36.045 ;
        RECT 229.970 35.465 230.140 35.780 ;
        RECT 229.970 35.255 230.600 35.465 ;
        RECT 229.970 34.585 230.140 35.255 ;
        RECT 229.970 34.415 230.940 34.585 ;
        RECT 229.970 33.745 230.140 34.415 ;
        RECT 229.970 33.480 231.280 33.745 ;
        RECT 229.970 33.265 230.140 33.480 ;
        RECT 229.970 31.575 231.750 33.265 ;
        RECT 229.970 29.755 231.230 31.575 ;
        RECT 229.970 29.585 230.140 29.755 ;
        RECT 229.970 28.835 231.305 29.585 ;
        RECT 229.970 28.665 230.140 28.835 ;
        RECT 229.970 28.145 231.770 28.665 ;
        RECT 222.670 27.435 225.150 27.605 ;
        RECT 222.670 20.565 222.840 27.435 ;
        RECT 224.980 20.565 225.150 27.435 ;
        RECT 222.670 20.395 225.150 20.565 ;
        RECT 229.970 27.455 231.230 28.145 ;
        RECT 229.970 27.185 230.140 27.455 ;
        RECT 229.970 26.975 230.600 27.185 ;
        RECT 229.970 26.305 230.140 26.975 ;
        RECT 229.970 26.135 230.940 26.305 ;
        RECT 229.970 25.465 230.140 26.135 ;
        RECT 229.970 25.200 231.280 25.465 ;
        RECT 229.970 24.885 230.140 25.200 ;
        RECT 229.970 24.675 230.600 24.885 ;
        RECT 229.970 24.005 230.140 24.675 ;
        RECT 229.970 23.835 230.940 24.005 ;
        RECT 229.970 23.165 230.140 23.835 ;
        RECT 229.970 22.900 231.280 23.165 ;
        RECT 229.970 22.685 230.140 22.900 ;
        RECT 229.970 20.995 231.750 22.685 ;
        RECT 229.970 19.175 231.230 20.995 ;
        RECT 229.970 19.005 230.140 19.175 ;
        RECT 229.970 18.255 231.305 19.005 ;
        RECT 229.970 18.085 230.140 18.255 ;
        RECT 229.970 17.565 231.770 18.085 ;
        RECT 222.670 16.855 225.150 17.025 ;
        RECT 222.670 9.985 222.840 16.855 ;
        RECT 224.980 9.985 225.150 16.855 ;
        RECT 222.670 9.815 225.150 9.985 ;
        RECT 229.970 16.875 231.230 17.565 ;
        RECT 229.970 16.605 230.140 16.875 ;
        RECT 229.970 16.395 230.600 16.605 ;
        RECT 229.970 15.725 230.140 16.395 ;
        RECT 229.970 15.555 230.940 15.725 ;
        RECT 229.970 14.885 230.140 15.555 ;
        RECT 229.970 14.620 231.280 14.885 ;
        RECT 229.970 14.305 230.140 14.620 ;
        RECT 229.970 14.095 230.600 14.305 ;
        RECT 229.970 13.425 230.140 14.095 ;
        RECT 229.970 13.255 230.940 13.425 ;
        RECT 229.970 12.585 230.140 13.255 ;
        RECT 229.970 12.320 231.280 12.585 ;
        RECT 229.970 12.105 230.140 12.320 ;
        RECT 229.970 10.415 231.750 12.105 ;
        RECT 229.970 8.595 231.230 10.415 ;
        RECT 229.970 8.510 230.140 8.595 ;
      LAYER mcon ;
        RECT 229.970 49.595 230.140 49.765 ;
        RECT 229.970 49.135 230.140 49.305 ;
        RECT 223.305 41.555 223.475 41.725 ;
        RECT 223.665 41.555 223.835 41.725 ;
        RECT 224.025 41.555 224.195 41.725 ;
        RECT 224.385 41.555 224.555 41.725 ;
        RECT 229.970 48.675 230.140 48.845 ;
        RECT 229.970 48.215 230.140 48.385 ;
        RECT 229.970 47.755 230.140 47.925 ;
        RECT 229.970 46.835 230.140 47.005 ;
        RECT 229.970 46.375 230.140 46.545 ;
        RECT 229.970 45.915 230.140 46.085 ;
        RECT 229.970 45.455 230.140 45.625 ;
        RECT 229.970 44.535 230.140 44.705 ;
        RECT 229.970 44.075 230.140 44.245 ;
        RECT 229.970 43.615 230.140 43.785 ;
        RECT 229.970 43.155 230.140 43.325 ;
        RECT 229.970 42.695 230.140 42.865 ;
        RECT 229.970 42.235 230.140 42.405 ;
        RECT 229.970 41.775 230.140 41.945 ;
        RECT 229.970 41.315 230.140 41.485 ;
        RECT 229.970 40.855 230.140 41.025 ;
        RECT 229.970 40.395 230.140 40.565 ;
        RECT 229.970 39.935 230.140 40.105 ;
        RECT 229.970 39.475 230.140 39.645 ;
        RECT 229.970 39.015 230.140 39.185 ;
        RECT 229.970 38.555 230.140 38.725 ;
        RECT 223.305 30.975 223.475 31.145 ;
        RECT 223.665 30.975 223.835 31.145 ;
        RECT 224.025 30.975 224.195 31.145 ;
        RECT 224.385 30.975 224.555 31.145 ;
        RECT 229.970 38.095 230.140 38.265 ;
        RECT 229.970 37.635 230.140 37.805 ;
        RECT 229.970 37.175 230.140 37.345 ;
        RECT 229.970 36.255 230.140 36.425 ;
        RECT 229.970 35.795 230.140 35.965 ;
        RECT 229.970 35.335 230.140 35.505 ;
        RECT 229.970 34.875 230.140 35.045 ;
        RECT 229.970 33.955 230.140 34.125 ;
        RECT 229.970 33.495 230.140 33.665 ;
        RECT 229.970 33.035 230.140 33.205 ;
        RECT 229.970 32.575 230.140 32.745 ;
        RECT 229.970 32.115 230.140 32.285 ;
        RECT 229.970 31.655 230.140 31.825 ;
        RECT 229.970 31.195 230.140 31.365 ;
        RECT 229.970 30.735 230.140 30.905 ;
        RECT 229.970 30.275 230.140 30.445 ;
        RECT 229.970 29.815 230.140 29.985 ;
        RECT 229.970 29.355 230.140 29.525 ;
        RECT 229.970 28.895 230.140 29.065 ;
        RECT 229.970 28.435 230.140 28.605 ;
        RECT 229.970 27.975 230.140 28.145 ;
        RECT 223.305 20.395 223.475 20.565 ;
        RECT 223.665 20.395 223.835 20.565 ;
        RECT 224.025 20.395 224.195 20.565 ;
        RECT 224.385 20.395 224.555 20.565 ;
        RECT 229.970 27.515 230.140 27.685 ;
        RECT 229.970 27.055 230.140 27.225 ;
        RECT 229.970 26.595 230.140 26.765 ;
        RECT 229.970 25.675 230.140 25.845 ;
        RECT 229.970 25.215 230.140 25.385 ;
        RECT 229.970 24.755 230.140 24.925 ;
        RECT 229.970 24.295 230.140 24.465 ;
        RECT 229.970 23.375 230.140 23.545 ;
        RECT 229.970 22.915 230.140 23.085 ;
        RECT 229.970 22.455 230.140 22.625 ;
        RECT 229.970 21.995 230.140 22.165 ;
        RECT 229.970 21.535 230.140 21.705 ;
        RECT 229.970 21.075 230.140 21.245 ;
        RECT 229.970 20.615 230.140 20.785 ;
        RECT 229.970 20.155 230.140 20.325 ;
        RECT 229.970 19.695 230.140 19.865 ;
        RECT 229.970 19.235 230.140 19.405 ;
        RECT 229.970 18.775 230.140 18.945 ;
        RECT 229.970 18.315 230.140 18.485 ;
        RECT 229.970 17.855 230.140 18.025 ;
        RECT 229.970 17.395 230.140 17.565 ;
        RECT 223.305 9.815 223.475 9.985 ;
        RECT 223.665 9.815 223.835 9.985 ;
        RECT 224.025 9.815 224.195 9.985 ;
        RECT 224.385 9.815 224.555 9.985 ;
        RECT 229.970 16.935 230.140 17.105 ;
        RECT 229.970 16.475 230.140 16.645 ;
        RECT 229.970 16.015 230.140 16.185 ;
        RECT 229.970 15.095 230.140 15.265 ;
        RECT 229.970 14.635 230.140 14.805 ;
        RECT 229.970 14.175 230.140 14.345 ;
        RECT 229.970 13.715 230.140 13.885 ;
        RECT 229.970 12.795 230.140 12.965 ;
        RECT 229.970 12.335 230.140 12.505 ;
        RECT 229.970 11.875 230.140 12.045 ;
        RECT 229.970 11.415 230.140 11.585 ;
        RECT 229.970 10.955 230.140 11.125 ;
        RECT 229.970 10.495 230.140 10.665 ;
        RECT 229.970 10.035 230.140 10.205 ;
        RECT 229.970 9.575 230.140 9.745 ;
        RECT 229.970 9.115 230.140 9.285 ;
        RECT 229.970 8.655 230.140 8.825 ;
      LAYER met1 ;
        RECT 223.070 41.525 224.745 41.755 ;
        RECT 224.045 41.000 224.745 41.525 ;
        RECT 229.815 41.000 230.295 49.910 ;
        RECT 224.045 40.700 230.295 41.000 ;
        RECT 223.070 30.945 224.745 31.175 ;
        RECT 224.045 30.420 224.745 30.945 ;
        RECT 229.815 30.420 230.295 40.700 ;
        RECT 224.045 30.120 230.295 30.420 ;
        RECT 223.070 20.365 224.745 20.595 ;
        RECT 224.045 19.840 224.745 20.365 ;
        RECT 229.815 19.840 230.295 30.120 ;
        RECT 224.045 19.540 230.295 19.840 ;
        RECT 223.070 9.785 224.745 10.015 ;
        RECT 224.045 9.260 224.745 9.785 ;
        RECT 229.815 9.260 230.295 19.540 ;
        RECT 224.045 8.960 230.295 9.260 ;
        RECT 229.815 -3.375 230.295 8.960 ;
        RECT 229.425 -4.075 230.685 -3.375 ;
      LAYER via ;
        RECT 229.445 -3.695 229.705 -3.435 ;
        RECT 229.765 -3.695 230.025 -3.435 ;
        RECT 230.085 -3.695 230.345 -3.435 ;
        RECT 230.405 -3.695 230.665 -3.435 ;
        RECT 229.445 -4.015 229.705 -3.755 ;
        RECT 229.765 -4.015 230.025 -3.755 ;
        RECT 230.085 -4.015 230.345 -3.755 ;
        RECT 230.405 -4.015 230.665 -3.755 ;
      LAYER met2 ;
        RECT 229.235 -4.225 230.835 -3.225 ;
      LAYER via2 ;
        RECT 229.295 -4.065 230.775 -3.385 ;
      LAYER met3 ;
        RECT 229.260 -4.275 235.475 -3.175 ;
    END
    PORT
      LAYER nwell ;
        RECT -10.205 0.975 -8.600 15.615 ;
      LAYER li1 ;
        RECT -8.875 15.340 -8.705 15.425 ;
        RECT -10.040 14.590 -8.705 15.340 ;
        RECT -8.875 14.380 -8.705 14.590 ;
        RECT -10.015 14.150 -8.705 14.380 ;
        RECT -8.875 13.480 -8.705 14.150 ;
        RECT -10.015 13.270 -8.705 13.480 ;
        RECT -8.875 13.000 -8.705 13.270 ;
        RECT -10.015 12.770 -8.705 13.000 ;
        RECT -8.875 12.100 -8.705 12.770 ;
        RECT -10.015 11.890 -8.705 12.100 ;
        RECT -8.875 11.620 -8.705 11.890 ;
        RECT -10.015 11.390 -8.705 11.620 ;
        RECT -8.875 10.720 -8.705 11.390 ;
        RECT -10.015 10.510 -8.705 10.720 ;
        RECT -8.875 10.240 -8.705 10.510 ;
        RECT -10.015 10.010 -8.705 10.240 ;
        RECT -8.875 9.340 -8.705 10.010 ;
        RECT -10.015 9.130 -8.705 9.340 ;
        RECT -8.875 8.860 -8.705 9.130 ;
        RECT -10.015 8.630 -8.705 8.860 ;
        RECT -8.875 7.960 -8.705 8.630 ;
        RECT -10.015 7.750 -8.705 7.960 ;
        RECT -8.875 7.480 -8.705 7.750 ;
        RECT -10.015 7.250 -8.705 7.480 ;
        RECT -8.875 6.580 -8.705 7.250 ;
        RECT -10.015 6.370 -8.705 6.580 ;
        RECT -8.875 6.100 -8.705 6.370 ;
        RECT -10.015 5.870 -8.705 6.100 ;
        RECT -8.875 5.200 -8.705 5.870 ;
        RECT -10.015 4.990 -8.705 5.200 ;
        RECT -8.875 4.720 -8.705 4.990 ;
        RECT -10.015 4.490 -8.705 4.720 ;
        RECT -8.875 3.820 -8.705 4.490 ;
        RECT -10.015 3.610 -8.705 3.820 ;
        RECT -8.875 3.340 -8.705 3.610 ;
        RECT -10.015 3.110 -8.705 3.340 ;
        RECT -8.875 2.440 -8.705 3.110 ;
        RECT -10.015 2.230 -8.705 2.440 ;
        RECT -8.875 2.000 -8.705 2.230 ;
        RECT -10.040 1.250 -8.705 2.000 ;
        RECT -8.875 1.165 -8.705 1.250 ;
      LAYER mcon ;
        RECT -8.875 15.110 -8.705 15.280 ;
        RECT -8.875 14.650 -8.705 14.820 ;
        RECT -8.875 14.190 -8.705 14.360 ;
        RECT -8.875 13.730 -8.705 13.900 ;
        RECT -8.875 13.270 -8.705 13.440 ;
        RECT -8.875 12.810 -8.705 12.980 ;
        RECT -8.875 12.350 -8.705 12.520 ;
        RECT -8.875 11.890 -8.705 12.060 ;
        RECT -8.875 11.430 -8.705 11.600 ;
        RECT -8.875 10.970 -8.705 11.140 ;
        RECT -8.875 10.510 -8.705 10.680 ;
        RECT -8.875 10.050 -8.705 10.220 ;
        RECT -8.875 9.590 -8.705 9.760 ;
        RECT -8.875 9.130 -8.705 9.300 ;
        RECT -8.875 8.670 -8.705 8.840 ;
        RECT -8.875 8.210 -8.705 8.380 ;
        RECT -8.875 7.750 -8.705 7.920 ;
        RECT -8.875 7.290 -8.705 7.460 ;
        RECT -8.875 6.830 -8.705 7.000 ;
        RECT -8.875 6.370 -8.705 6.540 ;
        RECT -8.875 5.910 -8.705 6.080 ;
        RECT -8.875 5.450 -8.705 5.620 ;
        RECT -8.875 4.990 -8.705 5.160 ;
        RECT -8.875 4.530 -8.705 4.700 ;
        RECT -8.875 4.070 -8.705 4.240 ;
        RECT -8.875 3.610 -8.705 3.780 ;
        RECT -8.875 3.150 -8.705 3.320 ;
        RECT -8.875 2.690 -8.705 2.860 ;
        RECT -8.875 2.230 -8.705 2.400 ;
        RECT -8.875 1.770 -8.705 1.940 ;
        RECT -8.875 1.310 -8.705 1.480 ;
      LAYER met1 ;
        RECT -9.030 -3.375 -8.550 15.425 ;
        RECT -9.420 -4.075 -8.160 -3.375 ;
      LAYER via ;
        RECT -9.400 -3.695 -9.140 -3.435 ;
        RECT -9.080 -3.695 -8.820 -3.435 ;
        RECT -8.760 -3.695 -8.500 -3.435 ;
        RECT -8.440 -3.695 -8.180 -3.435 ;
        RECT -9.400 -4.015 -9.140 -3.755 ;
        RECT -9.080 -4.015 -8.820 -3.755 ;
        RECT -8.760 -4.015 -8.500 -3.755 ;
        RECT -8.440 -4.015 -8.180 -3.755 ;
      LAYER met2 ;
        RECT -9.610 -4.225 -8.010 -3.225 ;
      LAYER via2 ;
        RECT -9.550 -4.065 -8.070 -3.385 ;
      LAYER met3 ;
        RECT -14.160 -4.275 -7.190 -3.175 ;
    END
  END vdd
  PIN vss
    ANTENNAGATEAREA 12.110399 ;
    ANTENNADIFFAREA 20.036249 ;
    PORT
      LAYER pwell ;
        RECT 226.760 41.425 229.450 48.895 ;
        RECT 231.800 39.345 232.585 40.235 ;
        RECT 226.760 30.845 229.450 38.315 ;
        RECT 231.800 28.765 232.585 29.655 ;
        RECT 226.760 20.265 229.450 27.735 ;
        RECT 231.800 18.185 232.585 19.075 ;
        RECT 226.760 9.685 229.450 17.155 ;
      LAYER li1 ;
        RECT 232.690 49.825 232.860 49.910 ;
        RECT 231.940 49.135 232.860 49.825 ;
        RECT 226.890 48.595 229.320 48.765 ;
        RECT 231.400 48.615 232.860 49.135 ;
        RECT 226.890 41.725 227.060 48.595 ;
        RECT 229.150 41.725 229.320 48.595 ;
        RECT 232.690 48.385 232.860 48.615 ;
        RECT 232.225 48.135 232.860 48.385 ;
        RECT 232.690 47.465 232.860 48.135 ;
        RECT 232.230 47.295 232.860 47.465 ;
        RECT 232.690 46.625 232.860 47.295 ;
        RECT 232.230 46.360 232.860 46.625 ;
        RECT 232.690 46.085 232.860 46.360 ;
        RECT 232.225 45.835 232.860 46.085 ;
        RECT 232.690 45.165 232.860 45.835 ;
        RECT 232.230 44.995 232.860 45.165 ;
        RECT 232.690 44.325 232.860 44.995 ;
        RECT 232.230 44.060 232.860 44.325 ;
        RECT 232.690 43.845 232.860 44.060 ;
        RECT 231.920 41.985 232.860 43.845 ;
        RECT 226.890 41.555 229.320 41.725 ;
        RECT 231.400 40.335 232.860 41.985 ;
        RECT 232.690 40.165 232.860 40.335 ;
        RECT 231.965 39.415 232.860 40.165 ;
        RECT 232.690 39.245 232.860 39.415 ;
        RECT 231.940 38.555 232.860 39.245 ;
        RECT 226.890 38.015 229.320 38.185 ;
        RECT 231.400 38.035 232.860 38.555 ;
        RECT 226.890 31.145 227.060 38.015 ;
        RECT 229.150 31.145 229.320 38.015 ;
        RECT 232.690 37.805 232.860 38.035 ;
        RECT 232.225 37.555 232.860 37.805 ;
        RECT 232.690 36.885 232.860 37.555 ;
        RECT 232.230 36.715 232.860 36.885 ;
        RECT 232.690 36.045 232.860 36.715 ;
        RECT 232.230 35.780 232.860 36.045 ;
        RECT 232.690 35.505 232.860 35.780 ;
        RECT 232.225 35.255 232.860 35.505 ;
        RECT 232.690 34.585 232.860 35.255 ;
        RECT 232.230 34.415 232.860 34.585 ;
        RECT 232.690 33.745 232.860 34.415 ;
        RECT 232.230 33.480 232.860 33.745 ;
        RECT 232.690 33.265 232.860 33.480 ;
        RECT 231.920 31.405 232.860 33.265 ;
        RECT 226.890 30.975 229.320 31.145 ;
        RECT 231.400 29.755 232.860 31.405 ;
        RECT 232.690 29.585 232.860 29.755 ;
        RECT 231.965 28.835 232.860 29.585 ;
        RECT 232.690 28.665 232.860 28.835 ;
        RECT 231.940 27.975 232.860 28.665 ;
        RECT 226.890 27.435 229.320 27.605 ;
        RECT 231.400 27.455 232.860 27.975 ;
        RECT 226.890 20.565 227.060 27.435 ;
        RECT 229.150 20.565 229.320 27.435 ;
        RECT 232.690 27.225 232.860 27.455 ;
        RECT 232.225 26.975 232.860 27.225 ;
        RECT 232.690 26.305 232.860 26.975 ;
        RECT 232.230 26.135 232.860 26.305 ;
        RECT 232.690 25.465 232.860 26.135 ;
        RECT 232.230 25.200 232.860 25.465 ;
        RECT 232.690 24.925 232.860 25.200 ;
        RECT 232.225 24.675 232.860 24.925 ;
        RECT 232.690 24.005 232.860 24.675 ;
        RECT 232.230 23.835 232.860 24.005 ;
        RECT 232.690 23.165 232.860 23.835 ;
        RECT 232.230 22.900 232.860 23.165 ;
        RECT 232.690 22.685 232.860 22.900 ;
        RECT 231.920 20.825 232.860 22.685 ;
        RECT 226.890 20.395 229.320 20.565 ;
        RECT 231.400 19.175 232.860 20.825 ;
        RECT 232.690 19.005 232.860 19.175 ;
        RECT 231.965 18.255 232.860 19.005 ;
        RECT 232.690 18.085 232.860 18.255 ;
        RECT 231.940 17.395 232.860 18.085 ;
        RECT 226.890 16.855 229.320 17.025 ;
        RECT 231.400 16.875 232.860 17.395 ;
        RECT 226.890 9.985 227.060 16.855 ;
        RECT 229.150 9.985 229.320 16.855 ;
        RECT 232.690 16.645 232.860 16.875 ;
        RECT 232.225 16.395 232.860 16.645 ;
        RECT 232.690 15.725 232.860 16.395 ;
        RECT 232.230 15.555 232.860 15.725 ;
        RECT 232.690 14.885 232.860 15.555 ;
        RECT 232.230 14.620 232.860 14.885 ;
        RECT 232.690 14.345 232.860 14.620 ;
        RECT 232.225 14.095 232.860 14.345 ;
        RECT 232.690 13.425 232.860 14.095 ;
        RECT 232.230 13.255 232.860 13.425 ;
        RECT 232.690 12.585 232.860 13.255 ;
        RECT 232.230 12.320 232.860 12.585 ;
        RECT 232.690 12.105 232.860 12.320 ;
        RECT 231.920 10.245 232.860 12.105 ;
        RECT 226.890 9.815 229.320 9.985 ;
        RECT 231.400 8.595 232.860 10.245 ;
        RECT 232.690 8.510 232.860 8.595 ;
      LAYER mcon ;
        RECT 232.690 49.595 232.860 49.765 ;
        RECT 232.690 49.135 232.860 49.305 ;
        RECT 232.690 48.675 232.860 48.845 ;
        RECT 232.690 48.215 232.860 48.385 ;
        RECT 232.690 47.755 232.860 47.925 ;
        RECT 232.690 47.295 232.860 47.465 ;
        RECT 232.690 46.835 232.860 47.005 ;
        RECT 232.690 46.375 232.860 46.545 ;
        RECT 232.690 45.915 232.860 46.085 ;
        RECT 232.690 45.455 232.860 45.625 ;
        RECT 232.690 44.995 232.860 45.165 ;
        RECT 232.690 44.535 232.860 44.705 ;
        RECT 232.690 44.075 232.860 44.245 ;
        RECT 232.690 43.615 232.860 43.785 ;
        RECT 232.690 43.155 232.860 43.325 ;
        RECT 232.690 42.695 232.860 42.865 ;
        RECT 232.690 42.235 232.860 42.405 ;
        RECT 227.530 41.555 227.700 41.725 ;
        RECT 227.890 41.555 228.060 41.725 ;
        RECT 228.250 41.555 228.420 41.725 ;
        RECT 228.610 41.555 228.780 41.725 ;
        RECT 232.690 41.775 232.860 41.945 ;
        RECT 232.690 41.315 232.860 41.485 ;
        RECT 232.690 40.855 232.860 41.025 ;
        RECT 232.690 40.395 232.860 40.565 ;
        RECT 232.690 39.935 232.860 40.105 ;
        RECT 232.690 39.475 232.860 39.645 ;
        RECT 232.690 39.015 232.860 39.185 ;
        RECT 232.690 38.555 232.860 38.725 ;
        RECT 232.690 38.095 232.860 38.265 ;
        RECT 232.690 37.635 232.860 37.805 ;
        RECT 232.690 37.175 232.860 37.345 ;
        RECT 232.690 36.715 232.860 36.885 ;
        RECT 232.690 36.255 232.860 36.425 ;
        RECT 232.690 35.795 232.860 35.965 ;
        RECT 232.690 35.335 232.860 35.505 ;
        RECT 232.690 34.875 232.860 35.045 ;
        RECT 232.690 34.415 232.860 34.585 ;
        RECT 232.690 33.955 232.860 34.125 ;
        RECT 232.690 33.495 232.860 33.665 ;
        RECT 232.690 33.035 232.860 33.205 ;
        RECT 232.690 32.575 232.860 32.745 ;
        RECT 232.690 32.115 232.860 32.285 ;
        RECT 232.690 31.655 232.860 31.825 ;
        RECT 227.530 30.975 227.700 31.145 ;
        RECT 227.890 30.975 228.060 31.145 ;
        RECT 228.250 30.975 228.420 31.145 ;
        RECT 228.610 30.975 228.780 31.145 ;
        RECT 232.690 31.195 232.860 31.365 ;
        RECT 232.690 30.735 232.860 30.905 ;
        RECT 232.690 30.275 232.860 30.445 ;
        RECT 232.690 29.815 232.860 29.985 ;
        RECT 232.690 29.355 232.860 29.525 ;
        RECT 232.690 28.895 232.860 29.065 ;
        RECT 232.690 28.435 232.860 28.605 ;
        RECT 232.690 27.975 232.860 28.145 ;
        RECT 232.690 27.515 232.860 27.685 ;
        RECT 232.690 27.055 232.860 27.225 ;
        RECT 232.690 26.595 232.860 26.765 ;
        RECT 232.690 26.135 232.860 26.305 ;
        RECT 232.690 25.675 232.860 25.845 ;
        RECT 232.690 25.215 232.860 25.385 ;
        RECT 232.690 24.755 232.860 24.925 ;
        RECT 232.690 24.295 232.860 24.465 ;
        RECT 232.690 23.835 232.860 24.005 ;
        RECT 232.690 23.375 232.860 23.545 ;
        RECT 232.690 22.915 232.860 23.085 ;
        RECT 232.690 22.455 232.860 22.625 ;
        RECT 232.690 21.995 232.860 22.165 ;
        RECT 232.690 21.535 232.860 21.705 ;
        RECT 232.690 21.075 232.860 21.245 ;
        RECT 227.530 20.395 227.700 20.565 ;
        RECT 227.890 20.395 228.060 20.565 ;
        RECT 228.250 20.395 228.420 20.565 ;
        RECT 228.610 20.395 228.780 20.565 ;
        RECT 232.690 20.615 232.860 20.785 ;
        RECT 232.690 20.155 232.860 20.325 ;
        RECT 232.690 19.695 232.860 19.865 ;
        RECT 232.690 19.235 232.860 19.405 ;
        RECT 232.690 18.775 232.860 18.945 ;
        RECT 232.690 18.315 232.860 18.485 ;
        RECT 232.690 17.855 232.860 18.025 ;
        RECT 232.690 17.395 232.860 17.565 ;
        RECT 232.690 16.935 232.860 17.105 ;
        RECT 232.690 16.475 232.860 16.645 ;
        RECT 232.690 16.015 232.860 16.185 ;
        RECT 232.690 15.555 232.860 15.725 ;
        RECT 232.690 15.095 232.860 15.265 ;
        RECT 232.690 14.635 232.860 14.805 ;
        RECT 232.690 14.175 232.860 14.345 ;
        RECT 232.690 13.715 232.860 13.885 ;
        RECT 232.690 13.255 232.860 13.425 ;
        RECT 232.690 12.795 232.860 12.965 ;
        RECT 232.690 12.335 232.860 12.505 ;
        RECT 232.690 11.875 232.860 12.045 ;
        RECT 232.690 11.415 232.860 11.585 ;
        RECT 232.690 10.955 232.860 11.125 ;
        RECT 232.690 10.495 232.860 10.665 ;
        RECT 227.530 9.815 227.700 9.985 ;
        RECT 227.890 9.815 228.060 9.985 ;
        RECT 228.250 9.815 228.420 9.985 ;
        RECT 228.610 9.815 228.780 9.985 ;
        RECT 232.690 10.035 232.860 10.205 ;
        RECT 232.690 9.575 232.860 9.745 ;
        RECT 232.690 9.115 232.860 9.285 ;
        RECT 232.690 8.655 232.860 8.825 ;
      LAYER met1 ;
        RECT 228.740 41.755 229.440 41.790 ;
        RECT 227.295 41.525 229.440 41.755 ;
        RECT 228.740 41.490 229.440 41.525 ;
        RECT 228.740 31.175 229.440 31.210 ;
        RECT 227.295 30.945 229.440 31.175 ;
        RECT 228.740 30.910 229.440 30.945 ;
        RECT 228.740 20.595 229.440 20.630 ;
        RECT 227.295 20.365 229.440 20.595 ;
        RECT 228.740 20.330 229.440 20.365 ;
        RECT 228.740 10.015 229.440 10.050 ;
        RECT 227.295 9.785 229.440 10.015 ;
        RECT 228.740 9.750 229.440 9.785 ;
        RECT 232.535 -1.475 233.015 49.910 ;
        RECT 232.135 -2.175 233.395 -1.475 ;
      LAYER via ;
        RECT 228.800 41.510 229.060 41.770 ;
        RECT 229.120 41.510 229.380 41.770 ;
        RECT 232.660 41.670 232.920 41.930 ;
        RECT 232.660 41.350 232.920 41.610 ;
        RECT 228.800 30.930 229.060 31.190 ;
        RECT 229.120 30.930 229.380 31.190 ;
        RECT 232.660 31.090 232.920 31.350 ;
        RECT 232.660 30.770 232.920 31.030 ;
        RECT 228.800 20.350 229.060 20.610 ;
        RECT 229.120 20.350 229.380 20.610 ;
        RECT 232.660 20.510 232.920 20.770 ;
        RECT 232.660 20.190 232.920 20.450 ;
        RECT 228.800 9.770 229.060 10.030 ;
        RECT 229.120 9.770 229.380 10.030 ;
        RECT 232.660 9.930 232.920 10.190 ;
        RECT 232.660 9.610 232.920 9.870 ;
        RECT 232.155 -1.795 232.415 -1.535 ;
        RECT 232.475 -1.795 232.735 -1.535 ;
        RECT 232.795 -1.795 233.055 -1.535 ;
        RECT 233.115 -1.795 233.375 -1.535 ;
        RECT 232.155 -2.115 232.415 -1.855 ;
        RECT 232.475 -2.115 232.735 -1.855 ;
        RECT 232.795 -2.115 233.055 -1.855 ;
        RECT 233.115 -2.115 233.375 -1.855 ;
      LAYER met2 ;
        RECT 232.590 41.840 232.990 41.940 ;
        RECT 228.790 41.440 232.990 41.840 ;
        RECT 232.590 41.340 232.990 41.440 ;
        RECT 232.590 31.260 232.990 31.360 ;
        RECT 228.790 30.860 232.990 31.260 ;
        RECT 232.590 30.760 232.990 30.860 ;
        RECT 232.590 20.680 232.990 20.780 ;
        RECT 228.790 20.280 232.990 20.680 ;
        RECT 232.590 20.180 232.990 20.280 ;
        RECT 232.590 10.100 232.990 10.200 ;
        RECT 228.790 9.700 232.990 10.100 ;
        RECT 232.590 9.600 232.990 9.700 ;
        RECT 231.945 -2.325 233.545 -1.325 ;
      LAYER via2 ;
        RECT 232.005 -2.165 233.485 -1.485 ;
      LAYER met3 ;
        RECT 231.970 -2.375 235.475 -1.275 ;
    END
    PORT
      LAYER pwell ;
        RECT -11.320 14.520 -10.535 15.410 ;
        RECT -11.320 1.180 -10.535 2.070 ;
      LAYER li1 ;
        RECT -11.595 15.340 -11.425 15.425 ;
        RECT -11.595 14.590 -10.700 15.340 ;
        RECT -11.595 14.380 -11.425 14.590 ;
        RECT -11.595 14.150 -10.605 14.380 ;
        RECT -11.595 13.480 -11.425 14.150 ;
        RECT -11.595 13.270 -10.605 13.480 ;
        RECT -11.595 13.000 -11.425 13.270 ;
        RECT -11.595 12.770 -10.605 13.000 ;
        RECT -11.595 12.100 -11.425 12.770 ;
        RECT -11.595 11.890 -10.605 12.100 ;
        RECT -11.595 11.620 -11.425 11.890 ;
        RECT -11.595 11.390 -10.605 11.620 ;
        RECT -11.595 10.720 -11.425 11.390 ;
        RECT -11.595 10.510 -10.605 10.720 ;
        RECT -11.595 10.240 -11.425 10.510 ;
        RECT -11.595 10.010 -10.605 10.240 ;
        RECT -11.595 9.340 -11.425 10.010 ;
        RECT -11.595 9.130 -10.605 9.340 ;
        RECT -11.595 8.860 -11.425 9.130 ;
        RECT -11.595 8.630 -10.605 8.860 ;
        RECT -11.595 7.960 -11.425 8.630 ;
        RECT -11.595 7.750 -10.605 7.960 ;
        RECT -11.595 7.480 -11.425 7.750 ;
        RECT -11.595 7.250 -10.605 7.480 ;
        RECT -11.595 6.580 -11.425 7.250 ;
        RECT -11.595 6.370 -10.605 6.580 ;
        RECT -11.595 6.100 -11.425 6.370 ;
        RECT -11.595 5.870 -10.605 6.100 ;
        RECT -11.595 5.200 -11.425 5.870 ;
        RECT -11.595 4.990 -10.605 5.200 ;
        RECT -11.595 4.720 -11.425 4.990 ;
        RECT -11.595 4.490 -10.605 4.720 ;
        RECT -11.595 3.820 -11.425 4.490 ;
        RECT -11.595 3.610 -10.605 3.820 ;
        RECT -11.595 3.340 -11.425 3.610 ;
        RECT -11.595 3.110 -10.605 3.340 ;
        RECT -11.595 2.440 -11.425 3.110 ;
        RECT -11.595 2.230 -10.605 2.440 ;
        RECT -11.595 2.000 -11.425 2.230 ;
        RECT -11.595 1.250 -10.700 2.000 ;
        RECT -11.595 1.165 -11.425 1.250 ;
      LAYER mcon ;
        RECT -11.595 15.110 -11.425 15.280 ;
        RECT -11.595 14.650 -11.425 14.820 ;
        RECT -11.595 14.190 -11.425 14.360 ;
        RECT -11.595 13.730 -11.425 13.900 ;
        RECT -11.595 12.810 -11.425 12.980 ;
        RECT -11.595 12.350 -11.425 12.520 ;
        RECT -11.595 11.430 -11.425 11.600 ;
        RECT -11.595 10.970 -11.425 11.140 ;
        RECT -11.595 10.050 -11.425 10.220 ;
        RECT -11.595 9.590 -11.425 9.760 ;
        RECT -11.595 8.670 -11.425 8.840 ;
        RECT -11.595 8.210 -11.425 8.380 ;
        RECT -11.595 7.290 -11.425 7.460 ;
        RECT -11.595 6.830 -11.425 7.000 ;
        RECT -11.595 5.910 -11.425 6.080 ;
        RECT -11.595 5.450 -11.425 5.620 ;
        RECT -11.595 4.530 -11.425 4.700 ;
        RECT -11.595 4.070 -11.425 4.240 ;
        RECT -11.595 3.150 -11.425 3.320 ;
        RECT -11.595 2.690 -11.425 2.860 ;
        RECT -11.595 1.770 -11.425 1.940 ;
        RECT -11.595 1.310 -11.425 1.480 ;
      LAYER met1 ;
        RECT -11.750 -1.475 -11.270 15.425 ;
        RECT -12.150 -2.175 -10.890 -1.475 ;
      LAYER via ;
        RECT -12.130 -1.795 -11.870 -1.535 ;
        RECT -11.810 -1.795 -11.550 -1.535 ;
        RECT -11.490 -1.795 -11.230 -1.535 ;
        RECT -11.170 -1.795 -10.910 -1.535 ;
        RECT -12.130 -2.115 -11.870 -1.855 ;
        RECT -11.810 -2.115 -11.550 -1.855 ;
        RECT -11.490 -2.115 -11.230 -1.855 ;
        RECT -11.170 -2.115 -10.910 -1.855 ;
      LAYER met2 ;
        RECT -12.340 -2.325 -10.740 -1.325 ;
      LAYER via2 ;
        RECT -12.280 -2.165 -10.800 -1.485 ;
      LAYER met3 ;
        RECT -14.155 -2.375 -7.190 -1.275 ;
    END
  END vss
  PIN sample
    ANTENNAGATEAREA 3.960000 ;
    PORT
      LAYER li1 ;
        RECT 231.450 44.035 231.700 45.665 ;
        RECT 231.450 33.455 231.700 35.085 ;
        RECT 231.450 22.875 231.700 24.505 ;
        RECT 231.450 12.295 231.700 13.925 ;
      LAYER mcon ;
        RECT 231.500 44.075 231.670 44.245 ;
        RECT 231.500 33.495 231.670 33.665 ;
        RECT 231.500 22.915 231.670 23.085 ;
        RECT 231.500 12.335 231.670 12.505 ;
      LAYER met1 ;
        RECT 231.425 44.030 231.745 44.290 ;
        RECT 231.425 33.450 231.745 33.710 ;
        RECT 231.425 22.870 231.745 23.130 ;
        RECT 231.425 12.290 231.745 12.550 ;
      LAYER via ;
        RECT 231.455 44.030 231.715 44.290 ;
        RECT 231.455 33.450 231.715 33.710 ;
        RECT 231.455 22.870 231.715 23.130 ;
        RECT 231.455 12.290 231.715 12.550 ;
      LAYER met2 ;
        RECT 231.425 44.000 233.815 44.320 ;
        RECT 233.415 33.740 233.815 44.000 ;
        RECT 231.425 33.420 233.815 33.740 ;
        RECT 233.415 23.160 233.815 33.420 ;
        RECT 231.425 22.840 233.815 23.160 ;
        RECT 233.415 12.580 233.815 22.840 ;
        RECT 231.425 12.260 233.815 12.580 ;
        RECT 233.415 1.195 233.815 12.260 ;
        RECT 233.015 0.795 233.815 1.195 ;
      LAYER via2 ;
        RECT 233.075 0.855 233.355 1.135 ;
        RECT 233.475 0.855 233.755 1.135 ;
      LAYER met3 ;
        RECT 115.255 0.795 233.815 1.195 ;
        RECT 115.255 -0.510 115.655 0.795 ;
        RECT -14.155 -0.910 115.655 -0.510 ;
    END
  END sample
  PIN out
    ANTENNADIFFAREA 11.599999 ;
    PORT
      LAYER li1 ;
        RECT 223.570 47.435 224.610 47.605 ;
        RECT 227.430 47.435 228.470 47.605 ;
        RECT 223.570 46.255 224.610 46.425 ;
        RECT 227.430 46.255 228.470 46.425 ;
        RECT 223.570 45.075 224.610 45.245 ;
        RECT 227.430 45.075 228.470 45.245 ;
        RECT 223.570 43.895 224.610 44.065 ;
        RECT 227.430 43.895 228.470 44.065 ;
        RECT 223.570 42.715 224.610 42.885 ;
        RECT 227.430 42.715 228.470 42.885 ;
        RECT 223.570 36.855 224.610 37.025 ;
        RECT 227.430 36.855 228.470 37.025 ;
        RECT 223.570 35.675 224.610 35.845 ;
        RECT 227.430 35.675 228.470 35.845 ;
        RECT 223.570 34.495 224.610 34.665 ;
        RECT 227.430 34.495 228.470 34.665 ;
        RECT 223.570 33.315 224.610 33.485 ;
        RECT 227.430 33.315 228.470 33.485 ;
        RECT 223.570 32.135 224.610 32.305 ;
        RECT 227.430 32.135 228.470 32.305 ;
        RECT 223.570 26.275 224.610 26.445 ;
        RECT 227.430 26.275 228.470 26.445 ;
        RECT 223.570 25.095 224.610 25.265 ;
        RECT 227.430 25.095 228.470 25.265 ;
        RECT 223.570 23.915 224.610 24.085 ;
        RECT 227.430 23.915 228.470 24.085 ;
        RECT 223.570 22.735 224.610 22.905 ;
        RECT 227.430 22.735 228.470 22.905 ;
        RECT 223.570 21.555 224.610 21.725 ;
        RECT 227.430 21.555 228.470 21.725 ;
        RECT 223.570 15.695 224.610 15.865 ;
        RECT 227.430 15.695 228.470 15.865 ;
        RECT 223.570 14.515 224.610 14.685 ;
        RECT 227.430 14.515 228.470 14.685 ;
        RECT 223.570 13.335 224.610 13.505 ;
        RECT 227.430 13.335 228.470 13.505 ;
        RECT 223.570 12.155 224.610 12.325 ;
        RECT 227.430 12.155 228.470 12.325 ;
        RECT 223.570 10.975 224.610 11.145 ;
        RECT 227.430 10.975 228.470 11.145 ;
      LAYER mcon ;
        RECT 223.825 47.435 223.995 47.605 ;
        RECT 224.185 47.435 224.355 47.605 ;
        RECT 227.685 47.435 227.855 47.605 ;
        RECT 228.045 47.435 228.215 47.605 ;
        RECT 223.825 46.255 223.995 46.425 ;
        RECT 224.185 46.255 224.355 46.425 ;
        RECT 227.685 46.255 227.855 46.425 ;
        RECT 228.045 46.255 228.215 46.425 ;
        RECT 223.825 45.075 223.995 45.245 ;
        RECT 224.185 45.075 224.355 45.245 ;
        RECT 227.685 45.075 227.855 45.245 ;
        RECT 228.045 45.075 228.215 45.245 ;
        RECT 223.825 43.895 223.995 44.065 ;
        RECT 224.185 43.895 224.355 44.065 ;
        RECT 227.685 43.895 227.855 44.065 ;
        RECT 228.045 43.895 228.215 44.065 ;
        RECT 223.825 42.715 223.995 42.885 ;
        RECT 224.185 42.715 224.355 42.885 ;
        RECT 227.685 42.715 227.855 42.885 ;
        RECT 228.045 42.715 228.215 42.885 ;
        RECT 223.825 36.855 223.995 37.025 ;
        RECT 224.185 36.855 224.355 37.025 ;
        RECT 227.685 36.855 227.855 37.025 ;
        RECT 228.045 36.855 228.215 37.025 ;
        RECT 223.825 35.675 223.995 35.845 ;
        RECT 224.185 35.675 224.355 35.845 ;
        RECT 227.685 35.675 227.855 35.845 ;
        RECT 228.045 35.675 228.215 35.845 ;
        RECT 223.825 34.495 223.995 34.665 ;
        RECT 224.185 34.495 224.355 34.665 ;
        RECT 227.685 34.495 227.855 34.665 ;
        RECT 228.045 34.495 228.215 34.665 ;
        RECT 223.825 33.315 223.995 33.485 ;
        RECT 224.185 33.315 224.355 33.485 ;
        RECT 227.685 33.315 227.855 33.485 ;
        RECT 228.045 33.315 228.215 33.485 ;
        RECT 223.825 32.135 223.995 32.305 ;
        RECT 224.185 32.135 224.355 32.305 ;
        RECT 227.685 32.135 227.855 32.305 ;
        RECT 228.045 32.135 228.215 32.305 ;
        RECT 223.825 26.275 223.995 26.445 ;
        RECT 224.185 26.275 224.355 26.445 ;
        RECT 227.685 26.275 227.855 26.445 ;
        RECT 228.045 26.275 228.215 26.445 ;
        RECT 223.825 25.095 223.995 25.265 ;
        RECT 224.185 25.095 224.355 25.265 ;
        RECT 227.685 25.095 227.855 25.265 ;
        RECT 228.045 25.095 228.215 25.265 ;
        RECT 223.825 23.915 223.995 24.085 ;
        RECT 224.185 23.915 224.355 24.085 ;
        RECT 227.685 23.915 227.855 24.085 ;
        RECT 228.045 23.915 228.215 24.085 ;
        RECT 223.825 22.735 223.995 22.905 ;
        RECT 224.185 22.735 224.355 22.905 ;
        RECT 227.685 22.735 227.855 22.905 ;
        RECT 228.045 22.735 228.215 22.905 ;
        RECT 223.825 21.555 223.995 21.725 ;
        RECT 224.185 21.555 224.355 21.725 ;
        RECT 227.685 21.555 227.855 21.725 ;
        RECT 228.045 21.555 228.215 21.725 ;
        RECT 223.825 15.695 223.995 15.865 ;
        RECT 224.185 15.695 224.355 15.865 ;
        RECT 227.685 15.695 227.855 15.865 ;
        RECT 228.045 15.695 228.215 15.865 ;
        RECT 223.825 14.515 223.995 14.685 ;
        RECT 224.185 14.515 224.355 14.685 ;
        RECT 227.685 14.515 227.855 14.685 ;
        RECT 228.045 14.515 228.215 14.685 ;
        RECT 223.825 13.335 223.995 13.505 ;
        RECT 224.185 13.335 224.355 13.505 ;
        RECT 227.685 13.335 227.855 13.505 ;
        RECT 228.045 13.335 228.215 13.505 ;
        RECT 223.825 12.155 223.995 12.325 ;
        RECT 224.185 12.155 224.355 12.325 ;
        RECT 227.685 12.155 227.855 12.325 ;
        RECT 228.045 12.155 228.215 12.325 ;
        RECT 223.825 10.975 223.995 11.145 ;
        RECT 224.185 10.975 224.355 11.145 ;
        RECT 227.685 10.975 227.855 11.145 ;
        RECT 228.045 10.975 228.215 11.145 ;
      LAYER met1 ;
        RECT 225.100 47.635 225.800 47.670 ;
        RECT 223.590 47.405 228.450 47.635 ;
        RECT 225.100 47.370 225.800 47.405 ;
        RECT 225.100 46.455 225.800 46.490 ;
        RECT 223.590 46.225 228.450 46.455 ;
        RECT 225.100 46.190 225.800 46.225 ;
        RECT 225.100 45.275 225.800 45.310 ;
        RECT 223.590 45.045 228.450 45.275 ;
        RECT 225.100 45.010 225.800 45.045 ;
        RECT 225.100 44.095 225.800 44.130 ;
        RECT 223.590 43.865 228.450 44.095 ;
        RECT 225.100 43.830 225.800 43.865 ;
        RECT 225.100 42.915 225.800 42.950 ;
        RECT 223.590 42.685 228.450 42.915 ;
        RECT 225.100 42.650 225.800 42.685 ;
        RECT 225.100 37.055 225.800 37.090 ;
        RECT 223.590 36.825 228.450 37.055 ;
        RECT 225.100 36.790 225.800 36.825 ;
        RECT 225.100 35.875 225.800 35.910 ;
        RECT 223.590 35.645 228.450 35.875 ;
        RECT 225.100 35.610 225.800 35.645 ;
        RECT 225.100 34.695 225.800 34.730 ;
        RECT 223.590 34.465 228.450 34.695 ;
        RECT 225.100 34.430 225.800 34.465 ;
        RECT 225.100 33.515 225.800 33.550 ;
        RECT 223.590 33.285 228.450 33.515 ;
        RECT 225.100 33.250 225.800 33.285 ;
        RECT 225.100 32.335 225.800 32.370 ;
        RECT 223.590 32.105 228.450 32.335 ;
        RECT 225.100 32.070 225.800 32.105 ;
        RECT 225.100 26.475 225.800 26.510 ;
        RECT 223.590 26.245 228.450 26.475 ;
        RECT 225.100 26.210 225.800 26.245 ;
        RECT 225.100 25.295 225.800 25.330 ;
        RECT 223.590 25.065 228.450 25.295 ;
        RECT 225.100 25.030 225.800 25.065 ;
        RECT 225.100 24.115 225.800 24.150 ;
        RECT 223.590 23.885 228.450 24.115 ;
        RECT 225.100 23.850 225.800 23.885 ;
        RECT 225.100 22.935 225.800 22.970 ;
        RECT 223.590 22.705 228.450 22.935 ;
        RECT 225.100 22.670 225.800 22.705 ;
        RECT 225.100 21.755 225.800 21.790 ;
        RECT 223.590 21.525 228.450 21.755 ;
        RECT 225.100 21.490 225.800 21.525 ;
        RECT 225.100 15.895 225.800 15.930 ;
        RECT 223.590 15.665 228.450 15.895 ;
        RECT 225.100 15.630 225.800 15.665 ;
        RECT 225.100 14.715 225.800 14.750 ;
        RECT 223.590 14.485 228.450 14.715 ;
        RECT 225.100 14.450 225.800 14.485 ;
        RECT 225.100 13.535 225.800 13.570 ;
        RECT 223.590 13.305 228.450 13.535 ;
        RECT 225.100 13.270 225.800 13.305 ;
        RECT 225.100 12.355 225.800 12.390 ;
        RECT 223.590 12.125 228.450 12.355 ;
        RECT 225.100 12.090 225.800 12.125 ;
        RECT 225.100 11.175 225.800 11.210 ;
        RECT 223.590 10.945 228.450 11.175 ;
        RECT 225.100 10.910 225.800 10.945 ;
      LAYER via ;
        RECT 225.160 47.390 225.420 47.650 ;
        RECT 225.480 47.390 225.740 47.650 ;
        RECT 225.160 46.210 225.420 46.470 ;
        RECT 225.480 46.210 225.740 46.470 ;
        RECT 225.160 45.030 225.420 45.290 ;
        RECT 225.480 45.030 225.740 45.290 ;
        RECT 225.160 43.850 225.420 44.110 ;
        RECT 225.480 43.850 225.740 44.110 ;
        RECT 225.160 42.670 225.420 42.930 ;
        RECT 225.480 42.670 225.740 42.930 ;
        RECT 225.160 36.810 225.420 37.070 ;
        RECT 225.480 36.810 225.740 37.070 ;
        RECT 225.160 35.630 225.420 35.890 ;
        RECT 225.480 35.630 225.740 35.890 ;
        RECT 225.160 34.450 225.420 34.710 ;
        RECT 225.480 34.450 225.740 34.710 ;
        RECT 225.160 33.270 225.420 33.530 ;
        RECT 225.480 33.270 225.740 33.530 ;
        RECT 225.160 32.090 225.420 32.350 ;
        RECT 225.480 32.090 225.740 32.350 ;
        RECT 225.160 26.230 225.420 26.490 ;
        RECT 225.480 26.230 225.740 26.490 ;
        RECT 225.160 25.050 225.420 25.310 ;
        RECT 225.480 25.050 225.740 25.310 ;
        RECT 225.160 23.870 225.420 24.130 ;
        RECT 225.480 23.870 225.740 24.130 ;
        RECT 225.160 22.690 225.420 22.950 ;
        RECT 225.480 22.690 225.740 22.950 ;
        RECT 225.160 21.510 225.420 21.770 ;
        RECT 225.480 21.510 225.740 21.770 ;
        RECT 225.160 15.650 225.420 15.910 ;
        RECT 225.480 15.650 225.740 15.910 ;
        RECT 225.160 14.470 225.420 14.730 ;
        RECT 225.480 14.470 225.740 14.730 ;
        RECT 225.160 13.290 225.420 13.550 ;
        RECT 225.480 13.290 225.740 13.550 ;
        RECT 225.160 12.110 225.420 12.370 ;
        RECT 225.480 12.110 225.740 12.370 ;
        RECT 225.160 10.930 225.420 11.190 ;
        RECT 225.480 10.930 225.740 11.190 ;
      LAYER met2 ;
        RECT 225.350 47.720 225.750 48.310 ;
        RECT 225.150 47.320 225.750 47.720 ;
        RECT 225.350 46.540 225.750 47.320 ;
        RECT 221.275 45.330 221.675 46.430 ;
        RECT 225.150 46.140 225.750 46.540 ;
        RECT 225.350 45.360 225.750 46.140 ;
        RECT 225.150 45.330 225.750 45.360 ;
        RECT 221.275 44.830 225.750 45.330 ;
        RECT 225.350 44.180 225.750 44.830 ;
        RECT 225.150 43.780 225.750 44.180 ;
        RECT 225.350 43.000 225.750 43.780 ;
        RECT 225.150 42.600 225.750 43.000 ;
        RECT 225.350 37.140 225.750 37.730 ;
        RECT 225.150 36.740 225.750 37.140 ;
        RECT 225.350 35.960 225.750 36.740 ;
        RECT 221.275 34.750 221.675 35.850 ;
        RECT 225.150 35.560 225.750 35.960 ;
        RECT 225.350 34.780 225.750 35.560 ;
        RECT 225.150 34.750 225.750 34.780 ;
        RECT 221.275 34.250 225.750 34.750 ;
        RECT 225.350 33.600 225.750 34.250 ;
        RECT 225.150 33.200 225.750 33.600 ;
        RECT 225.350 32.420 225.750 33.200 ;
        RECT 225.150 32.020 225.750 32.420 ;
        RECT 225.350 26.560 225.750 27.150 ;
        RECT 225.150 26.160 225.750 26.560 ;
        RECT 225.350 25.380 225.750 26.160 ;
        RECT 221.275 24.170 221.675 25.270 ;
        RECT 225.150 24.980 225.750 25.380 ;
        RECT 225.350 24.200 225.750 24.980 ;
        RECT 225.150 24.170 225.750 24.200 ;
        RECT 221.275 23.670 225.750 24.170 ;
        RECT 225.350 23.020 225.750 23.670 ;
        RECT 225.150 22.620 225.750 23.020 ;
        RECT 225.350 21.840 225.750 22.620 ;
        RECT 225.150 21.440 225.750 21.840 ;
        RECT 225.350 15.980 225.750 16.570 ;
        RECT 225.150 15.580 225.750 15.980 ;
        RECT 225.350 14.800 225.750 15.580 ;
        RECT 221.275 13.590 221.675 14.690 ;
        RECT 225.150 14.400 225.750 14.800 ;
        RECT 225.350 13.620 225.750 14.400 ;
        RECT 225.150 13.590 225.750 13.620 ;
        RECT 221.275 13.090 225.750 13.590 ;
        RECT 225.350 12.440 225.750 13.090 ;
        RECT 225.150 12.040 225.750 12.440 ;
        RECT 225.350 11.260 225.750 12.040 ;
        RECT 225.150 10.860 225.750 11.260 ;
      LAYER via2 ;
        RECT 221.335 46.090 221.615 46.370 ;
        RECT 221.335 45.690 221.615 45.970 ;
        RECT 221.335 45.290 221.615 45.570 ;
        RECT 221.335 44.890 221.615 45.170 ;
        RECT 221.335 35.510 221.615 35.790 ;
        RECT 221.335 35.110 221.615 35.390 ;
        RECT 221.335 34.710 221.615 34.990 ;
        RECT 221.335 34.310 221.615 34.590 ;
        RECT 221.335 24.930 221.615 25.210 ;
        RECT 221.335 24.530 221.615 24.810 ;
        RECT 221.335 24.130 221.615 24.410 ;
        RECT 221.335 23.730 221.615 24.010 ;
        RECT 221.335 14.350 221.615 14.630 ;
        RECT 221.335 13.950 221.615 14.230 ;
        RECT 221.335 13.550 221.615 13.830 ;
        RECT 221.335 13.150 221.615 13.430 ;
      LAYER met3 ;
        RECT 221.275 44.830 221.675 46.430 ;
        RECT 221.275 34.250 221.675 35.850 ;
        RECT 221.275 23.670 221.675 25.270 ;
        RECT 221.275 13.090 221.675 14.690 ;
      LAYER via3 ;
        RECT 221.315 46.070 221.635 46.390 ;
        RECT 221.315 45.670 221.635 45.990 ;
        RECT 221.315 45.270 221.635 45.590 ;
        RECT 221.315 44.870 221.635 45.190 ;
        RECT 221.315 35.490 221.635 35.810 ;
        RECT 221.315 35.090 221.635 35.410 ;
        RECT 221.315 34.690 221.635 35.010 ;
        RECT 221.315 34.290 221.635 34.610 ;
        RECT 221.315 24.910 221.635 25.230 ;
        RECT 221.315 24.510 221.635 24.830 ;
        RECT 221.315 24.110 221.635 24.430 ;
        RECT 221.315 23.710 221.635 24.030 ;
        RECT 221.315 14.330 221.635 14.650 ;
        RECT 221.315 13.930 221.635 14.250 ;
        RECT 221.315 13.530 221.635 13.850 ;
        RECT 221.315 13.130 221.635 13.450 ;
      LAYER met4 ;
        RECT 221.275 49.850 221.675 50.080 ;
        RECT 3.405 49.350 221.675 49.850 ;
        RECT 3.405 48.155 3.885 49.350 ;
        RECT 9.905 48.155 10.385 49.350 ;
        RECT 16.405 48.155 16.885 49.350 ;
        RECT 22.905 48.155 23.385 49.350 ;
        RECT 29.405 48.155 29.885 49.350 ;
        RECT 35.905 48.155 36.385 49.350 ;
        RECT 42.405 48.155 42.885 49.350 ;
        RECT 48.905 48.155 49.385 49.350 ;
        RECT 55.405 48.155 55.885 49.350 ;
        RECT 61.905 48.155 62.385 49.350 ;
        RECT 68.405 48.155 68.885 49.350 ;
        RECT 74.905 48.155 75.385 49.350 ;
        RECT 81.405 48.155 81.885 49.350 ;
        RECT 87.905 48.155 88.385 49.350 ;
        RECT 94.405 48.155 94.885 49.350 ;
        RECT 100.905 48.155 101.385 49.350 ;
        RECT 107.405 48.155 107.885 49.350 ;
        RECT 113.905 48.155 114.385 49.350 ;
        RECT 120.405 48.155 120.885 49.350 ;
        RECT 126.905 48.155 127.385 49.350 ;
        RECT 133.405 48.155 133.885 49.350 ;
        RECT 139.905 48.155 140.385 49.350 ;
        RECT 146.405 48.155 146.885 49.350 ;
        RECT 152.905 48.155 153.385 49.350 ;
        RECT 159.405 48.155 159.885 49.350 ;
        RECT 165.905 48.155 166.385 49.350 ;
        RECT 172.405 48.155 172.885 49.350 ;
        RECT 178.905 48.155 179.385 49.350 ;
        RECT 185.405 48.155 185.885 49.350 ;
        RECT 191.905 48.155 192.385 49.350 ;
        RECT 198.405 48.155 198.885 49.350 ;
        RECT 204.905 48.155 205.385 49.350 ;
        RECT 211.405 48.155 211.885 49.350 ;
        RECT 217.905 48.155 218.385 49.350 ;
        RECT 2.840 46.545 4.450 48.155 ;
        RECT 9.340 46.545 10.950 48.155 ;
        RECT 15.840 46.545 17.450 48.155 ;
        RECT 22.340 46.545 23.950 48.155 ;
        RECT 28.840 46.545 30.450 48.155 ;
        RECT 35.340 46.545 36.950 48.155 ;
        RECT 41.840 46.545 43.450 48.155 ;
        RECT 48.340 46.545 49.950 48.155 ;
        RECT 54.840 46.545 56.450 48.155 ;
        RECT 61.340 46.545 62.950 48.155 ;
        RECT 67.840 46.545 69.450 48.155 ;
        RECT 74.340 46.545 75.950 48.155 ;
        RECT 80.840 46.545 82.450 48.155 ;
        RECT 87.340 46.545 88.950 48.155 ;
        RECT 93.840 46.545 95.450 48.155 ;
        RECT 100.340 46.545 101.950 48.155 ;
        RECT 106.840 46.545 108.450 48.155 ;
        RECT 113.340 46.545 114.950 48.155 ;
        RECT 119.840 46.545 121.450 48.155 ;
        RECT 126.340 46.545 127.950 48.155 ;
        RECT 132.840 46.545 134.450 48.155 ;
        RECT 139.340 46.545 140.950 48.155 ;
        RECT 145.840 46.545 147.450 48.155 ;
        RECT 152.340 46.545 153.950 48.155 ;
        RECT 158.840 46.545 160.450 48.155 ;
        RECT 165.340 46.545 166.950 48.155 ;
        RECT 171.840 46.545 173.450 48.155 ;
        RECT 178.340 46.545 179.950 48.155 ;
        RECT 184.840 46.545 186.450 48.155 ;
        RECT 191.340 46.545 192.950 48.155 ;
        RECT 197.840 46.545 199.450 48.155 ;
        RECT 204.340 46.545 205.950 48.155 ;
        RECT 210.840 46.545 212.450 48.155 ;
        RECT 217.340 46.545 218.950 48.155 ;
        RECT 3.405 43.955 3.885 46.545 ;
        RECT 9.905 43.955 10.385 46.545 ;
        RECT 16.405 43.955 16.885 46.545 ;
        RECT 22.905 43.955 23.385 46.545 ;
        RECT 29.405 43.955 29.885 46.545 ;
        RECT 35.905 43.955 36.385 46.545 ;
        RECT 42.405 43.955 42.885 46.545 ;
        RECT 48.905 43.955 49.385 46.545 ;
        RECT 55.405 43.955 55.885 46.545 ;
        RECT 61.905 43.955 62.385 46.545 ;
        RECT 68.405 43.955 68.885 46.545 ;
        RECT 74.905 43.955 75.385 46.545 ;
        RECT 81.405 43.955 81.885 46.545 ;
        RECT 87.905 43.955 88.385 46.545 ;
        RECT 94.405 43.955 94.885 46.545 ;
        RECT 100.905 43.955 101.385 46.545 ;
        RECT 107.405 43.955 107.885 46.545 ;
        RECT 113.905 43.955 114.385 46.545 ;
        RECT 120.405 43.955 120.885 46.545 ;
        RECT 126.905 43.955 127.385 46.545 ;
        RECT 133.405 43.955 133.885 46.545 ;
        RECT 139.905 43.955 140.385 46.545 ;
        RECT 146.405 43.955 146.885 46.545 ;
        RECT 152.905 43.955 153.385 46.545 ;
        RECT 159.405 43.955 159.885 46.545 ;
        RECT 165.905 43.955 166.385 46.545 ;
        RECT 172.405 43.955 172.885 46.545 ;
        RECT 178.905 43.955 179.385 46.545 ;
        RECT 185.405 43.955 185.885 46.545 ;
        RECT 191.905 43.955 192.385 46.545 ;
        RECT 198.405 43.955 198.885 46.545 ;
        RECT 204.905 43.955 205.385 46.545 ;
        RECT 211.405 43.955 211.885 46.545 ;
        RECT 217.905 43.955 218.385 46.545 ;
        RECT 2.840 42.345 4.450 43.955 ;
        RECT 9.340 42.345 10.950 43.955 ;
        RECT 15.840 42.345 17.450 43.955 ;
        RECT 22.340 42.345 23.950 43.955 ;
        RECT 28.840 42.345 30.450 43.955 ;
        RECT 35.340 42.345 36.950 43.955 ;
        RECT 41.840 42.345 43.450 43.955 ;
        RECT 48.340 42.345 49.950 43.955 ;
        RECT 54.840 42.345 56.450 43.955 ;
        RECT 61.340 42.345 62.950 43.955 ;
        RECT 67.840 42.345 69.450 43.955 ;
        RECT 74.340 42.345 75.950 43.955 ;
        RECT 80.840 42.345 82.450 43.955 ;
        RECT 87.340 42.345 88.950 43.955 ;
        RECT 93.840 42.345 95.450 43.955 ;
        RECT 100.340 42.345 101.950 43.955 ;
        RECT 106.840 42.345 108.450 43.955 ;
        RECT 113.340 42.345 114.950 43.955 ;
        RECT 119.840 42.345 121.450 43.955 ;
        RECT 126.340 42.345 127.950 43.955 ;
        RECT 132.840 42.345 134.450 43.955 ;
        RECT 139.340 42.345 140.950 43.955 ;
        RECT 145.840 42.345 147.450 43.955 ;
        RECT 152.340 42.345 153.950 43.955 ;
        RECT 158.840 42.345 160.450 43.955 ;
        RECT 165.340 42.345 166.950 43.955 ;
        RECT 171.840 42.345 173.450 43.955 ;
        RECT 178.340 42.345 179.950 43.955 ;
        RECT 184.840 42.345 186.450 43.955 ;
        RECT 191.340 42.345 192.950 43.955 ;
        RECT 197.840 42.345 199.450 43.955 ;
        RECT 204.340 42.345 205.950 43.955 ;
        RECT 210.840 42.345 212.450 43.955 ;
        RECT 217.340 42.345 218.950 43.955 ;
        RECT 3.405 39.755 3.885 42.345 ;
        RECT 9.905 39.755 10.385 42.345 ;
        RECT 16.405 39.755 16.885 42.345 ;
        RECT 22.905 39.755 23.385 42.345 ;
        RECT 29.405 39.755 29.885 42.345 ;
        RECT 35.905 39.755 36.385 42.345 ;
        RECT 42.405 39.755 42.885 42.345 ;
        RECT 48.905 39.755 49.385 42.345 ;
        RECT 55.405 39.755 55.885 42.345 ;
        RECT 61.905 39.755 62.385 42.345 ;
        RECT 68.405 39.755 68.885 42.345 ;
        RECT 74.905 39.755 75.385 42.345 ;
        RECT 81.405 39.755 81.885 42.345 ;
        RECT 87.905 39.755 88.385 42.345 ;
        RECT 94.405 39.755 94.885 42.345 ;
        RECT 100.905 39.755 101.385 42.345 ;
        RECT 107.405 39.755 107.885 42.345 ;
        RECT 113.905 39.755 114.385 42.345 ;
        RECT 120.405 39.755 120.885 42.345 ;
        RECT 126.905 39.755 127.385 42.345 ;
        RECT 133.405 39.755 133.885 42.345 ;
        RECT 139.905 39.755 140.385 42.345 ;
        RECT 146.405 39.755 146.885 42.345 ;
        RECT 152.905 39.755 153.385 42.345 ;
        RECT 159.405 39.755 159.885 42.345 ;
        RECT 165.905 39.755 166.385 42.345 ;
        RECT 172.405 39.755 172.885 42.345 ;
        RECT 178.905 39.755 179.385 42.345 ;
        RECT 185.405 39.755 185.885 42.345 ;
        RECT 191.905 39.755 192.385 42.345 ;
        RECT 198.405 39.755 198.885 42.345 ;
        RECT 204.905 39.755 205.385 42.345 ;
        RECT 211.405 39.755 211.885 42.345 ;
        RECT 217.905 39.755 218.385 42.345 ;
        RECT 2.840 38.145 4.450 39.755 ;
        RECT 9.340 38.145 10.950 39.755 ;
        RECT 15.840 38.145 17.450 39.755 ;
        RECT 22.340 38.145 23.950 39.755 ;
        RECT 28.840 38.145 30.450 39.755 ;
        RECT 35.340 38.145 36.950 39.755 ;
        RECT 41.840 38.145 43.450 39.755 ;
        RECT 48.340 38.145 49.950 39.755 ;
        RECT 54.840 38.145 56.450 39.755 ;
        RECT 61.340 38.145 62.950 39.755 ;
        RECT 67.840 38.145 69.450 39.755 ;
        RECT 74.340 38.145 75.950 39.755 ;
        RECT 80.840 38.145 82.450 39.755 ;
        RECT 87.340 38.145 88.950 39.755 ;
        RECT 93.840 38.145 95.450 39.755 ;
        RECT 100.340 38.145 101.950 39.755 ;
        RECT 106.840 38.145 108.450 39.755 ;
        RECT 113.340 38.145 114.950 39.755 ;
        RECT 119.840 38.145 121.450 39.755 ;
        RECT 126.340 38.145 127.950 39.755 ;
        RECT 132.840 38.145 134.450 39.755 ;
        RECT 139.340 38.145 140.950 39.755 ;
        RECT 145.840 38.145 147.450 39.755 ;
        RECT 152.340 38.145 153.950 39.755 ;
        RECT 158.840 38.145 160.450 39.755 ;
        RECT 165.340 38.145 166.950 39.755 ;
        RECT 171.840 38.145 173.450 39.755 ;
        RECT 178.340 38.145 179.950 39.755 ;
        RECT 184.840 38.145 186.450 39.755 ;
        RECT 191.340 38.145 192.950 39.755 ;
        RECT 197.840 38.145 199.450 39.755 ;
        RECT 204.340 38.145 205.950 39.755 ;
        RECT 210.840 38.145 212.450 39.755 ;
        RECT 217.340 38.145 218.950 39.755 ;
        RECT 3.405 35.555 3.885 38.145 ;
        RECT 9.905 35.555 10.385 38.145 ;
        RECT 16.405 35.555 16.885 38.145 ;
        RECT 22.905 35.555 23.385 38.145 ;
        RECT 29.405 35.555 29.885 38.145 ;
        RECT 35.905 35.555 36.385 38.145 ;
        RECT 42.405 35.555 42.885 38.145 ;
        RECT 48.905 35.555 49.385 38.145 ;
        RECT 55.405 35.555 55.885 38.145 ;
        RECT 61.905 35.555 62.385 38.145 ;
        RECT 68.405 35.555 68.885 38.145 ;
        RECT 74.905 35.555 75.385 38.145 ;
        RECT 81.405 35.555 81.885 38.145 ;
        RECT 87.905 35.555 88.385 38.145 ;
        RECT 94.405 35.555 94.885 38.145 ;
        RECT 100.905 35.555 101.385 38.145 ;
        RECT 107.405 35.555 107.885 38.145 ;
        RECT 113.905 35.555 114.385 38.145 ;
        RECT 120.405 35.555 120.885 38.145 ;
        RECT 126.905 35.555 127.385 38.145 ;
        RECT 133.405 35.555 133.885 38.145 ;
        RECT 139.905 35.555 140.385 38.145 ;
        RECT 146.405 35.555 146.885 38.145 ;
        RECT 152.905 35.555 153.385 38.145 ;
        RECT 159.405 35.555 159.885 38.145 ;
        RECT 165.905 35.555 166.385 38.145 ;
        RECT 172.405 35.555 172.885 38.145 ;
        RECT 178.905 35.555 179.385 38.145 ;
        RECT 185.405 35.555 185.885 38.145 ;
        RECT 191.905 35.555 192.385 38.145 ;
        RECT 198.405 35.555 198.885 38.145 ;
        RECT 204.905 35.555 205.385 38.145 ;
        RECT 211.405 35.555 211.885 38.145 ;
        RECT 217.905 35.555 218.385 38.145 ;
        RECT 2.840 33.945 4.450 35.555 ;
        RECT 9.340 33.945 10.950 35.555 ;
        RECT 15.840 33.945 17.450 35.555 ;
        RECT 22.340 33.945 23.950 35.555 ;
        RECT 28.840 33.945 30.450 35.555 ;
        RECT 35.340 33.945 36.950 35.555 ;
        RECT 41.840 33.945 43.450 35.555 ;
        RECT 48.340 33.945 49.950 35.555 ;
        RECT 54.840 33.945 56.450 35.555 ;
        RECT 61.340 33.945 62.950 35.555 ;
        RECT 67.840 33.945 69.450 35.555 ;
        RECT 74.340 33.945 75.950 35.555 ;
        RECT 80.840 33.945 82.450 35.555 ;
        RECT 87.340 33.945 88.950 35.555 ;
        RECT 93.840 33.945 95.450 35.555 ;
        RECT 100.340 33.945 101.950 35.555 ;
        RECT 106.840 33.945 108.450 35.555 ;
        RECT 113.340 33.945 114.950 35.555 ;
        RECT 119.840 33.945 121.450 35.555 ;
        RECT 126.340 33.945 127.950 35.555 ;
        RECT 132.840 33.945 134.450 35.555 ;
        RECT 139.340 33.945 140.950 35.555 ;
        RECT 145.840 33.945 147.450 35.555 ;
        RECT 152.340 33.945 153.950 35.555 ;
        RECT 158.840 33.945 160.450 35.555 ;
        RECT 165.340 33.945 166.950 35.555 ;
        RECT 171.840 33.945 173.450 35.555 ;
        RECT 178.340 33.945 179.950 35.555 ;
        RECT 184.840 33.945 186.450 35.555 ;
        RECT 191.340 33.945 192.950 35.555 ;
        RECT 197.840 33.945 199.450 35.555 ;
        RECT 204.340 33.945 205.950 35.555 ;
        RECT 210.840 33.945 212.450 35.555 ;
        RECT 217.340 33.945 218.950 35.555 ;
        RECT 3.405 31.355 3.885 33.945 ;
        RECT 9.905 31.355 10.385 33.945 ;
        RECT 16.405 31.355 16.885 33.945 ;
        RECT 22.905 31.355 23.385 33.945 ;
        RECT 29.405 31.355 29.885 33.945 ;
        RECT 35.905 31.355 36.385 33.945 ;
        RECT 42.405 31.355 42.885 33.945 ;
        RECT 48.905 31.355 49.385 33.945 ;
        RECT 55.405 31.355 55.885 33.945 ;
        RECT 61.905 31.355 62.385 33.945 ;
        RECT 68.405 31.355 68.885 33.945 ;
        RECT 74.905 31.355 75.385 33.945 ;
        RECT 81.405 31.355 81.885 33.945 ;
        RECT 87.905 31.355 88.385 33.945 ;
        RECT 94.405 31.355 94.885 33.945 ;
        RECT 100.905 31.355 101.385 33.945 ;
        RECT 107.405 31.355 107.885 33.945 ;
        RECT 113.905 31.355 114.385 33.945 ;
        RECT 120.405 31.355 120.885 33.945 ;
        RECT 126.905 31.355 127.385 33.945 ;
        RECT 133.405 31.355 133.885 33.945 ;
        RECT 139.905 31.355 140.385 33.945 ;
        RECT 146.405 31.355 146.885 33.945 ;
        RECT 152.905 31.355 153.385 33.945 ;
        RECT 159.405 31.355 159.885 33.945 ;
        RECT 165.905 31.355 166.385 33.945 ;
        RECT 172.405 31.355 172.885 33.945 ;
        RECT 178.905 31.355 179.385 33.945 ;
        RECT 185.405 31.355 185.885 33.945 ;
        RECT 191.905 31.355 192.385 33.945 ;
        RECT 198.405 31.355 198.885 33.945 ;
        RECT 204.905 31.355 205.385 33.945 ;
        RECT 211.405 31.355 211.885 33.945 ;
        RECT 217.905 31.355 218.385 33.945 ;
        RECT 2.840 29.745 4.450 31.355 ;
        RECT 9.340 29.745 10.950 31.355 ;
        RECT 15.840 29.745 17.450 31.355 ;
        RECT 22.340 29.745 23.950 31.355 ;
        RECT 28.840 29.745 30.450 31.355 ;
        RECT 35.340 29.745 36.950 31.355 ;
        RECT 41.840 29.745 43.450 31.355 ;
        RECT 48.340 29.745 49.950 31.355 ;
        RECT 54.840 29.745 56.450 31.355 ;
        RECT 61.340 29.745 62.950 31.355 ;
        RECT 67.840 29.745 69.450 31.355 ;
        RECT 74.340 29.745 75.950 31.355 ;
        RECT 80.840 29.745 82.450 31.355 ;
        RECT 87.340 29.745 88.950 31.355 ;
        RECT 93.840 29.745 95.450 31.355 ;
        RECT 100.340 29.745 101.950 31.355 ;
        RECT 106.840 29.745 108.450 31.355 ;
        RECT 113.340 29.745 114.950 31.355 ;
        RECT 119.840 29.745 121.450 31.355 ;
        RECT 126.340 29.745 127.950 31.355 ;
        RECT 132.840 29.745 134.450 31.355 ;
        RECT 139.340 29.745 140.950 31.355 ;
        RECT 145.840 29.745 147.450 31.355 ;
        RECT 152.340 29.745 153.950 31.355 ;
        RECT 158.840 29.745 160.450 31.355 ;
        RECT 165.340 29.745 166.950 31.355 ;
        RECT 171.840 29.745 173.450 31.355 ;
        RECT 178.340 29.745 179.950 31.355 ;
        RECT 184.840 29.745 186.450 31.355 ;
        RECT 191.340 29.745 192.950 31.355 ;
        RECT 197.840 29.745 199.450 31.355 ;
        RECT 204.340 29.745 205.950 31.355 ;
        RECT 210.840 29.745 212.450 31.355 ;
        RECT 217.340 29.745 218.950 31.355 ;
        RECT 3.405 27.155 3.885 29.745 ;
        RECT 9.905 27.155 10.385 29.745 ;
        RECT 16.405 27.155 16.885 29.745 ;
        RECT 22.905 27.155 23.385 29.745 ;
        RECT 29.405 27.155 29.885 29.745 ;
        RECT 35.905 27.155 36.385 29.745 ;
        RECT 42.405 27.155 42.885 29.745 ;
        RECT 48.905 27.155 49.385 29.745 ;
        RECT 55.405 27.155 55.885 29.745 ;
        RECT 61.905 27.155 62.385 29.745 ;
        RECT 68.405 27.155 68.885 29.745 ;
        RECT 74.905 27.155 75.385 29.745 ;
        RECT 81.405 27.155 81.885 29.745 ;
        RECT 87.905 27.155 88.385 29.745 ;
        RECT 94.405 27.155 94.885 29.745 ;
        RECT 100.905 27.155 101.385 29.745 ;
        RECT 107.405 27.155 107.885 29.745 ;
        RECT 113.905 27.155 114.385 29.745 ;
        RECT 120.405 27.155 120.885 29.745 ;
        RECT 126.905 27.155 127.385 29.745 ;
        RECT 133.405 27.155 133.885 29.745 ;
        RECT 139.905 27.155 140.385 29.745 ;
        RECT 146.405 27.155 146.885 29.745 ;
        RECT 152.905 27.155 153.385 29.745 ;
        RECT 159.405 27.155 159.885 29.745 ;
        RECT 165.905 27.155 166.385 29.745 ;
        RECT 172.405 27.155 172.885 29.745 ;
        RECT 178.905 27.155 179.385 29.745 ;
        RECT 185.405 27.155 185.885 29.745 ;
        RECT 191.905 27.155 192.385 29.745 ;
        RECT 198.405 27.155 198.885 29.745 ;
        RECT 204.905 27.155 205.385 29.745 ;
        RECT 211.405 27.155 211.885 29.745 ;
        RECT 217.905 27.155 218.385 29.745 ;
        RECT 2.840 25.545 4.450 27.155 ;
        RECT 9.340 25.545 10.950 27.155 ;
        RECT 15.840 25.545 17.450 27.155 ;
        RECT 22.340 25.545 23.950 27.155 ;
        RECT 28.840 25.545 30.450 27.155 ;
        RECT 35.340 25.545 36.950 27.155 ;
        RECT 41.840 25.545 43.450 27.155 ;
        RECT 48.340 25.545 49.950 27.155 ;
        RECT 54.840 25.545 56.450 27.155 ;
        RECT 61.340 25.545 62.950 27.155 ;
        RECT 67.840 25.545 69.450 27.155 ;
        RECT 74.340 25.545 75.950 27.155 ;
        RECT 80.840 25.545 82.450 27.155 ;
        RECT 87.340 25.545 88.950 27.155 ;
        RECT 93.840 25.545 95.450 27.155 ;
        RECT 100.340 25.545 101.950 27.155 ;
        RECT 106.840 25.545 108.450 27.155 ;
        RECT 113.340 25.545 114.950 27.155 ;
        RECT 119.840 25.545 121.450 27.155 ;
        RECT 126.340 25.545 127.950 27.155 ;
        RECT 132.840 25.545 134.450 27.155 ;
        RECT 139.340 25.545 140.950 27.155 ;
        RECT 145.840 25.545 147.450 27.155 ;
        RECT 152.340 25.545 153.950 27.155 ;
        RECT 158.840 25.545 160.450 27.155 ;
        RECT 165.340 25.545 166.950 27.155 ;
        RECT 171.840 25.545 173.450 27.155 ;
        RECT 178.340 25.545 179.950 27.155 ;
        RECT 184.840 25.545 186.450 27.155 ;
        RECT 191.340 25.545 192.950 27.155 ;
        RECT 197.840 25.545 199.450 27.155 ;
        RECT 204.340 25.545 205.950 27.155 ;
        RECT 210.840 25.545 212.450 27.155 ;
        RECT 217.340 25.545 218.950 27.155 ;
        RECT 3.405 22.955 3.885 25.545 ;
        RECT 9.905 22.955 10.385 25.545 ;
        RECT 16.405 22.955 16.885 25.545 ;
        RECT 22.905 22.955 23.385 25.545 ;
        RECT 29.405 22.955 29.885 25.545 ;
        RECT 35.905 22.955 36.385 25.545 ;
        RECT 42.405 22.955 42.885 25.545 ;
        RECT 48.905 22.955 49.385 25.545 ;
        RECT 55.405 22.955 55.885 25.545 ;
        RECT 61.905 22.955 62.385 25.545 ;
        RECT 68.405 22.955 68.885 25.545 ;
        RECT 74.905 22.955 75.385 25.545 ;
        RECT 81.405 22.955 81.885 25.545 ;
        RECT 87.905 22.955 88.385 25.545 ;
        RECT 94.405 22.955 94.885 25.545 ;
        RECT 100.905 22.955 101.385 25.545 ;
        RECT 107.405 22.955 107.885 25.545 ;
        RECT 113.905 22.955 114.385 25.545 ;
        RECT 120.405 22.955 120.885 25.545 ;
        RECT 126.905 22.955 127.385 25.545 ;
        RECT 133.405 22.955 133.885 25.545 ;
        RECT 139.905 22.955 140.385 25.545 ;
        RECT 146.405 22.955 146.885 25.545 ;
        RECT 152.905 22.955 153.385 25.545 ;
        RECT 159.405 22.955 159.885 25.545 ;
        RECT 165.905 22.955 166.385 25.545 ;
        RECT 172.405 22.955 172.885 25.545 ;
        RECT 178.905 22.955 179.385 25.545 ;
        RECT 185.405 22.955 185.885 25.545 ;
        RECT 191.905 22.955 192.385 25.545 ;
        RECT 198.405 22.955 198.885 25.545 ;
        RECT 204.905 22.955 205.385 25.545 ;
        RECT 211.405 22.955 211.885 25.545 ;
        RECT 217.905 22.955 218.385 25.545 ;
        RECT 2.840 21.345 4.450 22.955 ;
        RECT 9.340 21.345 10.950 22.955 ;
        RECT 15.840 21.345 17.450 22.955 ;
        RECT 22.340 21.345 23.950 22.955 ;
        RECT 28.840 21.345 30.450 22.955 ;
        RECT 35.340 21.345 36.950 22.955 ;
        RECT 41.840 21.345 43.450 22.955 ;
        RECT 48.340 21.345 49.950 22.955 ;
        RECT 54.840 21.345 56.450 22.955 ;
        RECT 61.340 21.345 62.950 22.955 ;
        RECT 67.840 21.345 69.450 22.955 ;
        RECT 74.340 21.345 75.950 22.955 ;
        RECT 80.840 21.345 82.450 22.955 ;
        RECT 87.340 21.345 88.950 22.955 ;
        RECT 93.840 21.345 95.450 22.955 ;
        RECT 100.340 21.345 101.950 22.955 ;
        RECT 106.840 21.345 108.450 22.955 ;
        RECT 113.340 21.345 114.950 22.955 ;
        RECT 119.840 21.345 121.450 22.955 ;
        RECT 126.340 21.345 127.950 22.955 ;
        RECT 132.840 21.345 134.450 22.955 ;
        RECT 139.340 21.345 140.950 22.955 ;
        RECT 145.840 21.345 147.450 22.955 ;
        RECT 152.340 21.345 153.950 22.955 ;
        RECT 158.840 21.345 160.450 22.955 ;
        RECT 165.340 21.345 166.950 22.955 ;
        RECT 171.840 21.345 173.450 22.955 ;
        RECT 178.340 21.345 179.950 22.955 ;
        RECT 184.840 21.345 186.450 22.955 ;
        RECT 191.340 21.345 192.950 22.955 ;
        RECT 197.840 21.345 199.450 22.955 ;
        RECT 204.340 21.345 205.950 22.955 ;
        RECT 210.840 21.345 212.450 22.955 ;
        RECT 217.340 21.345 218.950 22.955 ;
        RECT 3.405 18.755 3.885 21.345 ;
        RECT 9.905 18.755 10.385 21.345 ;
        RECT 16.405 18.755 16.885 21.345 ;
        RECT 22.905 18.755 23.385 21.345 ;
        RECT 29.405 18.755 29.885 21.345 ;
        RECT 35.905 18.755 36.385 21.345 ;
        RECT 42.405 18.755 42.885 21.345 ;
        RECT 48.905 18.755 49.385 21.345 ;
        RECT 55.405 18.755 55.885 21.345 ;
        RECT 61.905 18.755 62.385 21.345 ;
        RECT 68.405 18.755 68.885 21.345 ;
        RECT 74.905 18.755 75.385 21.345 ;
        RECT 81.405 18.755 81.885 21.345 ;
        RECT 87.905 18.755 88.385 21.345 ;
        RECT 94.405 18.755 94.885 21.345 ;
        RECT 100.905 18.755 101.385 21.345 ;
        RECT 107.405 18.755 107.885 21.345 ;
        RECT 113.905 18.755 114.385 21.345 ;
        RECT 120.405 18.755 120.885 21.345 ;
        RECT 126.905 18.755 127.385 21.345 ;
        RECT 133.405 18.755 133.885 21.345 ;
        RECT 139.905 18.755 140.385 21.345 ;
        RECT 146.405 18.755 146.885 21.345 ;
        RECT 152.905 18.755 153.385 21.345 ;
        RECT 159.405 18.755 159.885 21.345 ;
        RECT 165.905 18.755 166.385 21.345 ;
        RECT 172.405 18.755 172.885 21.345 ;
        RECT 178.905 18.755 179.385 21.345 ;
        RECT 185.405 18.755 185.885 21.345 ;
        RECT 191.905 18.755 192.385 21.345 ;
        RECT 198.405 18.755 198.885 21.345 ;
        RECT 204.905 18.755 205.385 21.345 ;
        RECT 211.405 18.755 211.885 21.345 ;
        RECT 217.905 18.755 218.385 21.345 ;
        RECT 2.840 17.145 4.450 18.755 ;
        RECT 9.340 17.145 10.950 18.755 ;
        RECT 15.840 17.145 17.450 18.755 ;
        RECT 22.340 17.145 23.950 18.755 ;
        RECT 28.840 17.145 30.450 18.755 ;
        RECT 35.340 17.145 36.950 18.755 ;
        RECT 41.840 17.145 43.450 18.755 ;
        RECT 48.340 17.145 49.950 18.755 ;
        RECT 54.840 17.145 56.450 18.755 ;
        RECT 61.340 17.145 62.950 18.755 ;
        RECT 67.840 17.145 69.450 18.755 ;
        RECT 74.340 17.145 75.950 18.755 ;
        RECT 80.840 17.145 82.450 18.755 ;
        RECT 87.340 17.145 88.950 18.755 ;
        RECT 93.840 17.145 95.450 18.755 ;
        RECT 100.340 17.145 101.950 18.755 ;
        RECT 106.840 17.145 108.450 18.755 ;
        RECT 113.340 17.145 114.950 18.755 ;
        RECT 119.840 17.145 121.450 18.755 ;
        RECT 126.340 17.145 127.950 18.755 ;
        RECT 132.840 17.145 134.450 18.755 ;
        RECT 139.340 17.145 140.950 18.755 ;
        RECT 145.840 17.145 147.450 18.755 ;
        RECT 152.340 17.145 153.950 18.755 ;
        RECT 158.840 17.145 160.450 18.755 ;
        RECT 165.340 17.145 166.950 18.755 ;
        RECT 171.840 17.145 173.450 18.755 ;
        RECT 178.340 17.145 179.950 18.755 ;
        RECT 184.840 17.145 186.450 18.755 ;
        RECT 191.340 17.145 192.950 18.755 ;
        RECT 197.840 17.145 199.450 18.755 ;
        RECT 204.340 17.145 205.950 18.755 ;
        RECT 210.840 17.145 212.450 18.755 ;
        RECT 217.340 17.145 218.950 18.755 ;
        RECT 3.405 14.555 3.885 17.145 ;
        RECT 9.905 14.555 10.385 17.145 ;
        RECT 16.405 14.555 16.885 17.145 ;
        RECT 22.905 14.555 23.385 17.145 ;
        RECT 29.405 14.555 29.885 17.145 ;
        RECT 35.905 14.555 36.385 17.145 ;
        RECT 42.405 14.555 42.885 17.145 ;
        RECT 48.905 14.555 49.385 17.145 ;
        RECT 55.405 14.555 55.885 17.145 ;
        RECT 61.905 14.555 62.385 17.145 ;
        RECT 68.405 14.555 68.885 17.145 ;
        RECT 74.905 14.555 75.385 17.145 ;
        RECT 81.405 14.555 81.885 17.145 ;
        RECT 87.905 14.555 88.385 17.145 ;
        RECT 94.405 14.555 94.885 17.145 ;
        RECT 100.905 14.555 101.385 17.145 ;
        RECT 107.405 14.555 107.885 17.145 ;
        RECT 113.905 14.555 114.385 17.145 ;
        RECT 120.405 14.555 120.885 17.145 ;
        RECT 126.905 14.555 127.385 17.145 ;
        RECT 133.405 14.555 133.885 17.145 ;
        RECT 139.905 14.555 140.385 17.145 ;
        RECT 146.405 14.555 146.885 17.145 ;
        RECT 152.905 14.555 153.385 17.145 ;
        RECT 159.405 14.555 159.885 17.145 ;
        RECT 165.905 14.555 166.385 17.145 ;
        RECT 172.405 14.555 172.885 17.145 ;
        RECT 178.905 14.555 179.385 17.145 ;
        RECT 185.405 14.555 185.885 17.145 ;
        RECT 191.905 14.555 192.385 17.145 ;
        RECT 198.405 14.555 198.885 17.145 ;
        RECT 204.905 14.555 205.385 17.145 ;
        RECT 211.405 14.555 211.885 17.145 ;
        RECT 217.905 14.555 218.385 17.145 ;
        RECT 2.840 12.945 4.450 14.555 ;
        RECT 9.340 12.945 10.950 14.555 ;
        RECT 15.840 12.945 17.450 14.555 ;
        RECT 22.340 12.945 23.950 14.555 ;
        RECT 28.840 12.945 30.450 14.555 ;
        RECT 35.340 12.945 36.950 14.555 ;
        RECT 41.840 12.945 43.450 14.555 ;
        RECT 48.340 12.945 49.950 14.555 ;
        RECT 54.840 12.945 56.450 14.555 ;
        RECT 61.340 12.945 62.950 14.555 ;
        RECT 67.840 12.945 69.450 14.555 ;
        RECT 74.340 12.945 75.950 14.555 ;
        RECT 80.840 12.945 82.450 14.555 ;
        RECT 87.340 12.945 88.950 14.555 ;
        RECT 93.840 12.945 95.450 14.555 ;
        RECT 100.340 12.945 101.950 14.555 ;
        RECT 106.840 12.945 108.450 14.555 ;
        RECT 113.340 12.945 114.950 14.555 ;
        RECT 119.840 12.945 121.450 14.555 ;
        RECT 126.340 12.945 127.950 14.555 ;
        RECT 132.840 12.945 134.450 14.555 ;
        RECT 139.340 12.945 140.950 14.555 ;
        RECT 145.840 12.945 147.450 14.555 ;
        RECT 152.340 12.945 153.950 14.555 ;
        RECT 158.840 12.945 160.450 14.555 ;
        RECT 165.340 12.945 166.950 14.555 ;
        RECT 171.840 12.945 173.450 14.555 ;
        RECT 178.340 12.945 179.950 14.555 ;
        RECT 184.840 12.945 186.450 14.555 ;
        RECT 191.340 12.945 192.950 14.555 ;
        RECT 197.840 12.945 199.450 14.555 ;
        RECT 204.340 12.945 205.950 14.555 ;
        RECT 210.840 12.945 212.450 14.555 ;
        RECT 217.340 12.945 218.950 14.555 ;
        RECT 221.275 13.090 221.675 49.350 ;
        RECT 3.405 10.355 3.885 12.945 ;
        RECT 9.905 10.355 10.385 12.945 ;
        RECT 16.405 10.355 16.885 12.945 ;
        RECT 22.905 10.355 23.385 12.945 ;
        RECT 29.405 10.355 29.885 12.945 ;
        RECT 35.905 10.355 36.385 12.945 ;
        RECT 42.405 10.355 42.885 12.945 ;
        RECT 48.905 10.355 49.385 12.945 ;
        RECT 55.405 10.355 55.885 12.945 ;
        RECT 61.905 10.355 62.385 12.945 ;
        RECT 68.405 10.355 68.885 12.945 ;
        RECT 74.905 10.355 75.385 12.945 ;
        RECT 81.405 10.355 81.885 12.945 ;
        RECT 87.905 10.355 88.385 12.945 ;
        RECT 94.405 10.355 94.885 12.945 ;
        RECT 100.905 10.355 101.385 12.945 ;
        RECT 107.405 10.355 107.885 12.945 ;
        RECT 113.905 10.355 114.385 12.945 ;
        RECT 120.405 10.355 120.885 12.945 ;
        RECT 126.905 10.355 127.385 12.945 ;
        RECT 133.405 10.355 133.885 12.945 ;
        RECT 139.905 10.355 140.385 12.945 ;
        RECT 146.405 10.355 146.885 12.945 ;
        RECT 152.905 10.355 153.385 12.945 ;
        RECT 159.405 10.355 159.885 12.945 ;
        RECT 165.905 10.355 166.385 12.945 ;
        RECT 172.405 10.355 172.885 12.945 ;
        RECT 178.905 10.355 179.385 12.945 ;
        RECT 185.405 10.355 185.885 12.945 ;
        RECT 191.905 10.355 192.385 12.945 ;
        RECT 198.405 10.355 198.885 12.945 ;
        RECT 204.905 10.355 205.385 12.945 ;
        RECT 211.405 10.355 211.885 12.945 ;
        RECT 217.905 10.355 218.385 12.945 ;
        RECT 2.840 8.745 4.450 10.355 ;
        RECT 9.340 8.745 10.950 10.355 ;
        RECT 15.840 8.745 17.450 10.355 ;
        RECT 22.340 8.745 23.950 10.355 ;
        RECT 28.840 8.745 30.450 10.355 ;
        RECT 35.340 8.745 36.950 10.355 ;
        RECT 41.840 8.745 43.450 10.355 ;
        RECT 48.340 8.745 49.950 10.355 ;
        RECT 54.840 8.745 56.450 10.355 ;
        RECT 61.340 8.745 62.950 10.355 ;
        RECT 67.840 8.745 69.450 10.355 ;
        RECT 74.340 8.745 75.950 10.355 ;
        RECT 80.840 8.745 82.450 10.355 ;
        RECT 87.340 8.745 88.950 10.355 ;
        RECT 93.840 8.745 95.450 10.355 ;
        RECT 100.340 8.745 101.950 10.355 ;
        RECT 106.840 8.745 108.450 10.355 ;
        RECT 113.340 8.745 114.950 10.355 ;
        RECT 119.840 8.745 121.450 10.355 ;
        RECT 126.340 8.745 127.950 10.355 ;
        RECT 132.840 8.745 134.450 10.355 ;
        RECT 139.340 8.745 140.950 10.355 ;
        RECT 145.840 8.745 147.450 10.355 ;
        RECT 152.340 8.745 153.950 10.355 ;
        RECT 158.840 8.745 160.450 10.355 ;
        RECT 165.340 8.745 166.950 10.355 ;
        RECT 171.840 8.745 173.450 10.355 ;
        RECT 178.340 8.745 179.950 10.355 ;
        RECT 184.840 8.745 186.450 10.355 ;
        RECT 191.340 8.745 192.950 10.355 ;
        RECT 197.840 8.745 199.450 10.355 ;
        RECT 204.340 8.745 205.950 10.355 ;
        RECT 210.840 8.745 212.450 10.355 ;
        RECT 217.340 8.745 218.950 10.355 ;
        RECT 3.405 8.550 3.885 8.745 ;
        RECT 9.905 8.550 10.385 8.745 ;
        RECT 16.405 8.550 16.885 8.745 ;
        RECT 22.905 8.550 23.385 8.745 ;
        RECT 29.405 8.550 29.885 8.745 ;
        RECT 35.905 8.550 36.385 8.745 ;
        RECT 42.405 8.550 42.885 8.745 ;
        RECT 48.905 8.550 49.385 8.745 ;
        RECT 55.405 8.550 55.885 8.745 ;
        RECT 61.905 8.550 62.385 8.745 ;
        RECT 68.405 8.550 68.885 8.745 ;
        RECT 74.905 8.550 75.385 8.745 ;
        RECT 81.405 8.550 81.885 8.745 ;
        RECT 87.905 8.550 88.385 8.745 ;
        RECT 94.405 8.550 94.885 8.745 ;
        RECT 100.905 8.550 101.385 8.745 ;
        RECT 107.405 8.550 107.885 8.745 ;
        RECT 113.905 8.550 114.385 8.745 ;
        RECT 120.405 8.550 120.885 8.745 ;
        RECT 126.905 8.550 127.385 8.745 ;
        RECT 133.405 8.550 133.885 8.745 ;
        RECT 139.905 8.550 140.385 8.745 ;
        RECT 146.405 8.550 146.885 8.745 ;
        RECT 152.905 8.550 153.385 8.745 ;
        RECT 159.405 8.550 159.885 8.745 ;
        RECT 165.905 8.550 166.385 8.745 ;
        RECT 172.405 8.550 172.885 8.745 ;
        RECT 178.905 8.550 179.385 8.745 ;
        RECT 185.405 8.550 185.885 8.745 ;
        RECT 191.905 8.550 192.385 8.745 ;
        RECT 198.405 8.550 198.885 8.745 ;
        RECT 204.905 8.550 205.385 8.745 ;
        RECT 211.405 8.550 211.885 8.745 ;
        RECT 217.905 8.550 218.385 8.745 ;
    END
  END out
  PIN vin
    ANTENNADIFFAREA 13.920000 ;
    PORT
      LAYER li1 ;
        RECT 223.570 48.025 224.610 48.195 ;
        RECT 227.430 48.025 228.470 48.195 ;
        RECT 223.570 46.845 224.610 47.015 ;
        RECT 227.430 46.845 228.470 47.015 ;
        RECT 223.570 45.665 224.610 45.835 ;
        RECT 227.430 45.665 228.470 45.835 ;
        RECT 223.570 44.485 224.610 44.655 ;
        RECT 227.430 44.485 228.470 44.655 ;
        RECT 223.570 43.305 224.610 43.475 ;
        RECT 227.430 43.305 228.470 43.475 ;
        RECT 223.570 42.125 224.610 42.295 ;
        RECT 227.430 42.125 228.470 42.295 ;
        RECT 223.570 37.445 224.610 37.615 ;
        RECT 227.430 37.445 228.470 37.615 ;
        RECT 223.570 36.265 224.610 36.435 ;
        RECT 227.430 36.265 228.470 36.435 ;
        RECT 223.570 35.085 224.610 35.255 ;
        RECT 227.430 35.085 228.470 35.255 ;
        RECT 223.570 33.905 224.610 34.075 ;
        RECT 227.430 33.905 228.470 34.075 ;
        RECT 223.570 32.725 224.610 32.895 ;
        RECT 227.430 32.725 228.470 32.895 ;
        RECT 223.570 31.545 224.610 31.715 ;
        RECT 227.430 31.545 228.470 31.715 ;
        RECT 223.570 26.865 224.610 27.035 ;
        RECT 227.430 26.865 228.470 27.035 ;
        RECT 223.570 25.685 224.610 25.855 ;
        RECT 227.430 25.685 228.470 25.855 ;
        RECT 223.570 24.505 224.610 24.675 ;
        RECT 227.430 24.505 228.470 24.675 ;
        RECT 223.570 23.325 224.610 23.495 ;
        RECT 227.430 23.325 228.470 23.495 ;
        RECT 223.570 22.145 224.610 22.315 ;
        RECT 227.430 22.145 228.470 22.315 ;
        RECT 223.570 20.965 224.610 21.135 ;
        RECT 227.430 20.965 228.470 21.135 ;
        RECT 223.570 16.285 224.610 16.455 ;
        RECT 227.430 16.285 228.470 16.455 ;
        RECT 223.570 15.105 224.610 15.275 ;
        RECT 227.430 15.105 228.470 15.275 ;
        RECT 223.570 13.925 224.610 14.095 ;
        RECT 227.430 13.925 228.470 14.095 ;
        RECT 223.570 12.745 224.610 12.915 ;
        RECT 227.430 12.745 228.470 12.915 ;
        RECT 223.570 11.565 224.610 11.735 ;
        RECT 227.430 11.565 228.470 11.735 ;
        RECT 223.570 10.385 224.610 10.555 ;
        RECT 227.430 10.385 228.470 10.555 ;
      LAYER mcon ;
        RECT 223.825 48.025 223.995 48.195 ;
        RECT 224.185 48.025 224.355 48.195 ;
        RECT 227.685 48.025 227.855 48.195 ;
        RECT 228.045 48.025 228.215 48.195 ;
        RECT 223.825 46.845 223.995 47.015 ;
        RECT 224.185 46.845 224.355 47.015 ;
        RECT 227.685 46.845 227.855 47.015 ;
        RECT 228.045 46.845 228.215 47.015 ;
        RECT 223.825 45.665 223.995 45.835 ;
        RECT 224.185 45.665 224.355 45.835 ;
        RECT 227.685 45.665 227.855 45.835 ;
        RECT 228.045 45.665 228.215 45.835 ;
        RECT 223.825 44.485 223.995 44.655 ;
        RECT 224.185 44.485 224.355 44.655 ;
        RECT 227.685 44.485 227.855 44.655 ;
        RECT 228.045 44.485 228.215 44.655 ;
        RECT 223.825 43.305 223.995 43.475 ;
        RECT 224.185 43.305 224.355 43.475 ;
        RECT 227.685 43.305 227.855 43.475 ;
        RECT 228.045 43.305 228.215 43.475 ;
        RECT 223.825 42.125 223.995 42.295 ;
        RECT 224.185 42.125 224.355 42.295 ;
        RECT 227.685 42.125 227.855 42.295 ;
        RECT 228.045 42.125 228.215 42.295 ;
        RECT 223.825 37.445 223.995 37.615 ;
        RECT 224.185 37.445 224.355 37.615 ;
        RECT 227.685 37.445 227.855 37.615 ;
        RECT 228.045 37.445 228.215 37.615 ;
        RECT 223.825 36.265 223.995 36.435 ;
        RECT 224.185 36.265 224.355 36.435 ;
        RECT 227.685 36.265 227.855 36.435 ;
        RECT 228.045 36.265 228.215 36.435 ;
        RECT 223.825 35.085 223.995 35.255 ;
        RECT 224.185 35.085 224.355 35.255 ;
        RECT 227.685 35.085 227.855 35.255 ;
        RECT 228.045 35.085 228.215 35.255 ;
        RECT 223.825 33.905 223.995 34.075 ;
        RECT 224.185 33.905 224.355 34.075 ;
        RECT 227.685 33.905 227.855 34.075 ;
        RECT 228.045 33.905 228.215 34.075 ;
        RECT 223.825 32.725 223.995 32.895 ;
        RECT 224.185 32.725 224.355 32.895 ;
        RECT 227.685 32.725 227.855 32.895 ;
        RECT 228.045 32.725 228.215 32.895 ;
        RECT 223.825 31.545 223.995 31.715 ;
        RECT 224.185 31.545 224.355 31.715 ;
        RECT 227.685 31.545 227.855 31.715 ;
        RECT 228.045 31.545 228.215 31.715 ;
        RECT 223.825 26.865 223.995 27.035 ;
        RECT 224.185 26.865 224.355 27.035 ;
        RECT 227.685 26.865 227.855 27.035 ;
        RECT 228.045 26.865 228.215 27.035 ;
        RECT 223.825 25.685 223.995 25.855 ;
        RECT 224.185 25.685 224.355 25.855 ;
        RECT 227.685 25.685 227.855 25.855 ;
        RECT 228.045 25.685 228.215 25.855 ;
        RECT 223.825 24.505 223.995 24.675 ;
        RECT 224.185 24.505 224.355 24.675 ;
        RECT 227.685 24.505 227.855 24.675 ;
        RECT 228.045 24.505 228.215 24.675 ;
        RECT 223.825 23.325 223.995 23.495 ;
        RECT 224.185 23.325 224.355 23.495 ;
        RECT 227.685 23.325 227.855 23.495 ;
        RECT 228.045 23.325 228.215 23.495 ;
        RECT 223.825 22.145 223.995 22.315 ;
        RECT 224.185 22.145 224.355 22.315 ;
        RECT 227.685 22.145 227.855 22.315 ;
        RECT 228.045 22.145 228.215 22.315 ;
        RECT 223.825 20.965 223.995 21.135 ;
        RECT 224.185 20.965 224.355 21.135 ;
        RECT 227.685 20.965 227.855 21.135 ;
        RECT 228.045 20.965 228.215 21.135 ;
        RECT 223.825 16.285 223.995 16.455 ;
        RECT 224.185 16.285 224.355 16.455 ;
        RECT 227.685 16.285 227.855 16.455 ;
        RECT 228.045 16.285 228.215 16.455 ;
        RECT 223.825 15.105 223.995 15.275 ;
        RECT 224.185 15.105 224.355 15.275 ;
        RECT 227.685 15.105 227.855 15.275 ;
        RECT 228.045 15.105 228.215 15.275 ;
        RECT 223.825 13.925 223.995 14.095 ;
        RECT 224.185 13.925 224.355 14.095 ;
        RECT 227.685 13.925 227.855 14.095 ;
        RECT 228.045 13.925 228.215 14.095 ;
        RECT 223.825 12.745 223.995 12.915 ;
        RECT 224.185 12.745 224.355 12.915 ;
        RECT 227.685 12.745 227.855 12.915 ;
        RECT 228.045 12.745 228.215 12.915 ;
        RECT 223.825 11.565 223.995 11.735 ;
        RECT 224.185 11.565 224.355 11.735 ;
        RECT 227.685 11.565 227.855 11.735 ;
        RECT 228.045 11.565 228.215 11.735 ;
        RECT 223.825 10.385 223.995 10.555 ;
        RECT 224.185 10.385 224.355 10.555 ;
        RECT 227.685 10.385 227.855 10.555 ;
        RECT 228.045 10.385 228.215 10.555 ;
      LAYER met1 ;
        RECT 226.240 48.225 226.940 48.260 ;
        RECT 223.590 47.995 228.450 48.225 ;
        RECT 226.240 47.960 226.940 47.995 ;
        RECT 226.240 47.045 226.940 47.080 ;
        RECT 223.590 46.815 228.450 47.045 ;
        RECT 226.240 46.780 226.940 46.815 ;
        RECT 226.240 45.865 226.940 45.900 ;
        RECT 223.590 45.635 228.450 45.865 ;
        RECT 226.240 45.600 226.940 45.635 ;
        RECT 226.240 44.685 226.940 44.720 ;
        RECT 223.590 44.455 228.450 44.685 ;
        RECT 226.240 44.420 226.940 44.455 ;
        RECT 226.240 43.505 226.940 43.540 ;
        RECT 223.590 43.275 228.450 43.505 ;
        RECT 226.240 43.240 226.940 43.275 ;
        RECT 226.240 42.325 226.940 42.360 ;
        RECT 223.590 42.095 228.450 42.325 ;
        RECT 226.240 42.060 226.940 42.095 ;
        RECT 226.240 37.645 226.940 37.680 ;
        RECT 223.590 37.415 228.450 37.645 ;
        RECT 226.240 37.380 226.940 37.415 ;
        RECT 226.240 36.465 226.940 36.500 ;
        RECT 223.590 36.235 228.450 36.465 ;
        RECT 226.240 36.200 226.940 36.235 ;
        RECT 226.240 35.285 226.940 35.320 ;
        RECT 223.590 35.055 228.450 35.285 ;
        RECT 226.240 35.020 226.940 35.055 ;
        RECT 226.240 34.105 226.940 34.140 ;
        RECT 223.590 33.875 228.450 34.105 ;
        RECT 226.240 33.840 226.940 33.875 ;
        RECT 226.240 32.925 226.940 32.960 ;
        RECT 223.590 32.695 228.450 32.925 ;
        RECT 226.240 32.660 226.940 32.695 ;
        RECT 226.240 31.745 226.940 31.780 ;
        RECT 223.590 31.515 228.450 31.745 ;
        RECT 226.240 31.480 226.940 31.515 ;
        RECT 226.240 27.065 226.940 27.100 ;
        RECT 223.590 26.835 228.450 27.065 ;
        RECT 226.240 26.800 226.940 26.835 ;
        RECT 226.240 25.885 226.940 25.920 ;
        RECT 223.590 25.655 228.450 25.885 ;
        RECT 226.240 25.620 226.940 25.655 ;
        RECT 226.240 24.705 226.940 24.740 ;
        RECT 223.590 24.475 228.450 24.705 ;
        RECT 226.240 24.440 226.940 24.475 ;
        RECT 226.240 23.525 226.940 23.560 ;
        RECT 223.590 23.295 228.450 23.525 ;
        RECT 226.240 23.260 226.940 23.295 ;
        RECT 226.240 22.345 226.940 22.380 ;
        RECT 223.590 22.115 228.450 22.345 ;
        RECT 226.240 22.080 226.940 22.115 ;
        RECT 226.240 21.165 226.940 21.200 ;
        RECT 223.590 20.935 228.450 21.165 ;
        RECT 226.240 20.900 226.940 20.935 ;
        RECT 226.240 16.485 226.940 16.520 ;
        RECT 223.590 16.255 228.450 16.485 ;
        RECT 226.240 16.220 226.940 16.255 ;
        RECT 226.240 15.305 226.940 15.340 ;
        RECT 223.590 15.075 228.450 15.305 ;
        RECT 226.240 15.040 226.940 15.075 ;
        RECT 226.240 14.125 226.940 14.160 ;
        RECT 223.590 13.895 228.450 14.125 ;
        RECT 226.240 13.860 226.940 13.895 ;
        RECT 226.240 12.945 226.940 12.980 ;
        RECT 223.590 12.715 228.450 12.945 ;
        RECT 226.240 12.680 226.940 12.715 ;
        RECT 226.240 11.765 226.940 11.800 ;
        RECT 223.590 11.535 228.450 11.765 ;
        RECT 226.240 11.500 226.940 11.535 ;
        RECT 226.240 10.585 226.940 10.620 ;
        RECT 223.590 10.355 228.450 10.585 ;
        RECT 226.240 10.320 226.940 10.355 ;
      LAYER via ;
        RECT 226.300 47.980 226.560 48.240 ;
        RECT 226.620 47.980 226.880 48.240 ;
        RECT 226.300 46.800 226.560 47.060 ;
        RECT 226.620 46.800 226.880 47.060 ;
        RECT 226.300 45.620 226.560 45.880 ;
        RECT 226.620 45.620 226.880 45.880 ;
        RECT 226.300 44.440 226.560 44.700 ;
        RECT 226.620 44.440 226.880 44.700 ;
        RECT 226.300 43.260 226.560 43.520 ;
        RECT 226.620 43.260 226.880 43.520 ;
        RECT 226.300 42.080 226.560 42.340 ;
        RECT 226.620 42.080 226.880 42.340 ;
        RECT 226.300 37.400 226.560 37.660 ;
        RECT 226.620 37.400 226.880 37.660 ;
        RECT 226.300 36.220 226.560 36.480 ;
        RECT 226.620 36.220 226.880 36.480 ;
        RECT 226.300 35.040 226.560 35.300 ;
        RECT 226.620 35.040 226.880 35.300 ;
        RECT 226.300 33.860 226.560 34.120 ;
        RECT 226.620 33.860 226.880 34.120 ;
        RECT 226.300 32.680 226.560 32.940 ;
        RECT 226.620 32.680 226.880 32.940 ;
        RECT 226.300 31.500 226.560 31.760 ;
        RECT 226.620 31.500 226.880 31.760 ;
        RECT 226.300 26.820 226.560 27.080 ;
        RECT 226.620 26.820 226.880 27.080 ;
        RECT 226.300 25.640 226.560 25.900 ;
        RECT 226.620 25.640 226.880 25.900 ;
        RECT 226.300 24.460 226.560 24.720 ;
        RECT 226.620 24.460 226.880 24.720 ;
        RECT 226.300 23.280 226.560 23.540 ;
        RECT 226.620 23.280 226.880 23.540 ;
        RECT 226.300 22.100 226.560 22.360 ;
        RECT 226.620 22.100 226.880 22.360 ;
        RECT 226.300 20.920 226.560 21.180 ;
        RECT 226.620 20.920 226.880 21.180 ;
        RECT 226.300 16.240 226.560 16.500 ;
        RECT 226.620 16.240 226.880 16.500 ;
        RECT 226.300 15.060 226.560 15.320 ;
        RECT 226.620 15.060 226.880 15.320 ;
        RECT 226.300 13.880 226.560 14.140 ;
        RECT 226.620 13.880 226.880 14.140 ;
        RECT 226.300 12.700 226.560 12.960 ;
        RECT 226.620 12.700 226.880 12.960 ;
        RECT 226.300 11.520 226.560 11.780 ;
        RECT 226.620 11.520 226.880 11.780 ;
        RECT 226.300 10.340 226.560 10.600 ;
        RECT 226.620 10.340 226.880 10.600 ;
      LAYER met2 ;
        RECT 226.190 48.310 226.990 48.710 ;
        RECT 226.290 47.910 226.890 48.310 ;
        RECT 226.290 47.130 226.690 47.910 ;
        RECT 226.290 46.730 226.890 47.130 ;
        RECT 226.290 45.950 226.690 46.730 ;
        RECT 226.290 45.550 226.890 45.950 ;
        RECT 226.290 44.770 226.690 45.550 ;
        RECT 226.290 44.370 226.890 44.770 ;
        RECT 226.290 43.590 226.690 44.370 ;
        RECT 226.290 43.190 226.890 43.590 ;
        RECT 226.290 42.410 226.690 43.190 ;
        RECT 226.290 42.010 226.890 42.410 ;
        RECT 226.190 41.610 226.990 42.010 ;
        RECT 226.190 37.730 226.990 38.130 ;
        RECT 226.290 37.330 226.890 37.730 ;
        RECT 226.290 36.550 226.690 37.330 ;
        RECT 226.290 36.150 226.890 36.550 ;
        RECT 226.290 35.370 226.690 36.150 ;
        RECT 226.290 34.970 226.890 35.370 ;
        RECT 226.290 34.190 226.690 34.970 ;
        RECT 226.290 33.790 226.890 34.190 ;
        RECT 226.290 33.010 226.690 33.790 ;
        RECT 226.290 32.610 226.890 33.010 ;
        RECT 226.290 31.830 226.690 32.610 ;
        RECT 226.290 31.430 226.890 31.830 ;
        RECT 226.190 31.030 226.990 31.430 ;
        RECT 226.190 27.150 226.990 27.550 ;
        RECT 226.290 26.750 226.890 27.150 ;
        RECT 226.290 25.970 226.690 26.750 ;
        RECT 226.290 25.570 226.890 25.970 ;
        RECT 226.290 24.790 226.690 25.570 ;
        RECT 226.290 24.390 226.890 24.790 ;
        RECT 226.290 23.610 226.690 24.390 ;
        RECT 226.290 23.210 226.890 23.610 ;
        RECT 226.290 22.430 226.690 23.210 ;
        RECT 226.290 22.030 226.890 22.430 ;
        RECT 226.290 21.250 226.690 22.030 ;
        RECT 226.290 20.850 226.890 21.250 ;
        RECT 226.190 20.450 226.990 20.850 ;
        RECT 226.190 16.570 226.990 16.970 ;
        RECT 226.290 16.170 226.890 16.570 ;
        RECT 226.290 15.390 226.690 16.170 ;
        RECT 226.290 14.990 226.890 15.390 ;
        RECT 226.290 14.210 226.690 14.990 ;
        RECT 226.290 13.810 226.890 14.210 ;
        RECT 226.290 13.030 226.690 13.810 ;
        RECT 226.290 12.630 226.890 13.030 ;
        RECT 226.290 11.850 226.690 12.630 ;
        RECT 226.290 11.450 226.890 11.850 ;
        RECT 226.290 10.670 226.690 11.450 ;
        RECT 226.290 10.270 226.890 10.670 ;
        RECT 226.190 9.870 226.990 10.270 ;
      LAYER via2 ;
        RECT 226.250 48.370 226.530 48.650 ;
        RECT 226.650 48.370 226.930 48.650 ;
        RECT 226.250 41.670 226.530 41.950 ;
        RECT 226.650 41.670 226.930 41.950 ;
        RECT 226.250 37.790 226.530 38.070 ;
        RECT 226.650 37.790 226.930 38.070 ;
        RECT 226.250 31.090 226.530 31.370 ;
        RECT 226.650 31.090 226.930 31.370 ;
        RECT 226.250 27.210 226.530 27.490 ;
        RECT 226.650 27.210 226.930 27.490 ;
        RECT 226.250 20.510 226.530 20.790 ;
        RECT 226.650 20.510 226.930 20.790 ;
        RECT 226.250 16.630 226.530 16.910 ;
        RECT 226.650 16.630 226.930 16.910 ;
        RECT 226.250 9.930 226.530 10.210 ;
        RECT 226.650 9.930 226.930 10.210 ;
      LAYER met3 ;
        RECT 226.190 9.870 226.990 48.710 ;
      LAYER via3 ;
        RECT 226.230 29.370 226.550 29.690 ;
        RECT 226.630 29.370 226.950 29.690 ;
        RECT 226.230 28.970 226.550 29.290 ;
        RECT 226.630 28.970 226.950 29.290 ;
      LAYER met4 ;
        RECT 233.915 49.050 235.475 49.850 ;
        RECT 233.915 29.730 234.715 49.050 ;
        RECT 226.190 28.930 234.715 29.730 ;
    END
  END vin
  OBS
      LAYER pwell ;
        RECT 231.860 48.535 232.670 49.905 ;
        RECT 231.760 46.285 232.670 48.475 ;
        RECT 231.760 43.985 232.670 46.175 ;
        RECT 231.860 40.255 232.670 43.925 ;
        RECT 231.860 37.955 232.670 39.325 ;
        RECT 231.760 35.705 232.670 37.895 ;
        RECT 231.760 33.405 232.670 35.595 ;
        RECT 231.860 29.675 232.670 33.345 ;
        RECT 231.860 27.375 232.670 28.745 ;
        RECT 231.760 25.125 232.670 27.315 ;
        RECT 231.760 22.825 232.670 25.015 ;
        RECT 231.860 19.095 232.670 22.765 ;
        RECT 231.860 16.795 232.670 18.165 ;
        RECT 231.760 14.545 232.670 16.735 ;
        RECT -11.405 13.140 -10.495 14.490 ;
        RECT -11.405 11.760 -10.495 13.110 ;
        RECT 231.760 12.245 232.670 14.435 ;
        RECT -11.405 10.380 -10.495 11.730 ;
        RECT -11.405 9.000 -10.495 10.350 ;
        RECT -11.405 7.620 -10.495 8.970 ;
        RECT 231.860 8.515 232.670 12.185 ;
        RECT -11.405 6.240 -10.495 7.590 ;
        RECT -11.405 4.860 -10.495 6.210 ;
        RECT -11.405 3.480 -10.495 4.830 ;
        RECT -11.405 2.100 -10.495 3.450 ;
      LAYER li1 ;
        RECT 231.090 37.555 232.050 37.820 ;
        RECT 223.185 37.070 223.355 37.400 ;
        RECT 228.640 37.070 228.810 37.400 ;
        RECT 231.090 37.385 231.280 37.555 ;
        RECT 231.870 37.385 232.050 37.555 ;
        RECT 230.310 37.055 231.280 37.385 ;
        RECT 223.185 36.480 223.355 36.810 ;
        RECT 228.640 36.480 228.810 36.810 ;
        RECT 231.110 36.545 231.280 37.055 ;
        RECT 223.185 35.890 223.355 36.220 ;
        RECT 228.640 35.890 228.810 36.220 ;
        RECT 230.310 36.215 231.280 36.545 ;
        RECT 231.450 35.755 231.700 37.385 ;
        RECT 231.870 37.055 232.520 37.385 ;
        RECT 231.870 36.545 232.050 37.055 ;
        RECT 231.870 36.215 232.520 36.545 ;
        RECT 223.185 35.300 223.355 35.630 ;
        RECT 228.640 35.300 228.810 35.630 ;
        RECT 231.090 35.255 232.050 35.520 ;
        RECT 231.090 35.085 231.280 35.255 ;
        RECT 223.185 34.710 223.355 35.040 ;
        RECT 228.640 34.710 228.810 35.040 ;
        RECT 230.310 34.755 231.280 35.085 ;
        RECT 223.185 34.120 223.355 34.450 ;
        RECT 228.640 34.120 228.810 34.450 ;
        RECT 231.110 34.245 231.280 34.755 ;
        RECT 230.310 33.915 231.280 34.245 ;
        RECT 231.870 35.085 232.050 35.255 ;
        RECT 231.870 34.755 232.520 35.085 ;
        RECT 231.870 34.245 232.050 34.755 ;
        RECT 231.870 33.915 232.520 34.245 ;
        RECT 223.185 33.530 223.355 33.860 ;
        RECT 228.640 33.530 228.810 33.860 ;
        RECT 223.185 32.940 223.355 33.270 ;
        RECT 228.640 32.940 228.810 33.270 ;
        RECT 223.185 32.350 223.355 32.680 ;
        RECT 228.640 32.350 228.810 32.680 ;
        RECT 223.185 31.760 223.355 32.090 ;
        RECT 228.640 31.760 228.810 32.090 ;
        RECT 231.090 16.395 232.050 16.660 ;
        RECT 223.185 15.910 223.355 16.240 ;
        RECT 228.640 15.910 228.810 16.240 ;
        RECT 231.090 16.225 231.280 16.395 ;
        RECT 231.870 16.225 232.050 16.395 ;
        RECT 230.310 15.895 231.280 16.225 ;
        RECT 223.185 15.320 223.355 15.650 ;
        RECT 228.640 15.320 228.810 15.650 ;
        RECT 231.110 15.385 231.280 15.895 ;
        RECT 223.185 14.730 223.355 15.060 ;
        RECT 228.640 14.730 228.810 15.060 ;
        RECT 230.310 15.055 231.280 15.385 ;
        RECT 231.450 14.595 231.700 16.225 ;
        RECT 231.870 15.895 232.520 16.225 ;
        RECT 231.870 15.385 232.050 15.895 ;
        RECT 231.870 15.055 232.520 15.385 ;
        RECT 223.185 14.140 223.355 14.470 ;
        RECT 228.640 14.140 228.810 14.470 ;
        RECT 231.090 14.095 232.050 14.360 ;
        RECT -11.255 13.900 -10.625 13.980 ;
        RECT -10.025 13.900 -9.045 13.980 ;
        RECT 231.090 13.925 231.280 14.095 ;
        RECT -11.255 13.650 -9.045 13.900 ;
        RECT 223.185 13.550 223.355 13.880 ;
        RECT 228.640 13.550 228.810 13.880 ;
        RECT 230.310 13.595 231.280 13.925 ;
        RECT 223.185 12.960 223.355 13.290 ;
        RECT 228.640 12.960 228.810 13.290 ;
        RECT 231.110 13.085 231.280 13.595 ;
        RECT 230.310 12.755 231.280 13.085 ;
        RECT 231.870 13.925 232.050 14.095 ;
        RECT 231.870 13.595 232.520 13.925 ;
        RECT 231.870 13.085 232.050 13.595 ;
        RECT 231.870 12.755 232.520 13.085 ;
        RECT -11.255 12.520 -10.625 12.600 ;
        RECT -10.025 12.520 -9.045 12.600 ;
        RECT -11.255 12.270 -9.045 12.520 ;
        RECT 223.185 12.370 223.355 12.700 ;
        RECT 228.640 12.370 228.810 12.700 ;
        RECT 223.185 11.780 223.355 12.110 ;
        RECT 228.640 11.780 228.810 12.110 ;
        RECT -11.255 11.140 -10.625 11.220 ;
        RECT -10.025 11.140 -9.045 11.220 ;
        RECT 223.185 11.190 223.355 11.520 ;
        RECT 228.640 11.190 228.810 11.520 ;
        RECT -11.255 10.890 -9.045 11.140 ;
        RECT 223.185 10.600 223.355 10.930 ;
        RECT 228.640 10.600 228.810 10.930 ;
        RECT -11.255 9.760 -10.625 9.840 ;
        RECT -10.025 9.760 -9.045 9.840 ;
        RECT -11.255 9.510 -9.045 9.760 ;
        RECT -11.255 8.380 -10.625 8.460 ;
        RECT -10.025 8.380 -9.045 8.460 ;
        RECT -11.255 8.130 -9.045 8.380 ;
        RECT -11.255 7.000 -10.625 7.080 ;
        RECT -10.025 7.000 -9.045 7.080 ;
        RECT -11.255 6.750 -9.045 7.000 ;
        RECT -11.255 5.620 -10.625 5.700 ;
        RECT -10.025 5.620 -9.045 5.700 ;
        RECT -11.255 5.370 -9.045 5.620 ;
        RECT -11.255 4.240 -10.625 4.320 ;
        RECT -10.025 4.240 -9.045 4.320 ;
        RECT -11.255 3.990 -9.045 4.240 ;
        RECT -11.255 2.860 -10.625 2.940 ;
        RECT -10.025 2.860 -9.045 2.940 ;
        RECT -11.255 2.610 -9.045 2.860 ;
      LAYER mcon ;
        RECT 231.160 37.635 231.330 37.805 ;
        RECT 223.185 37.150 223.355 37.320 ;
        RECT 228.640 37.150 228.810 37.320 ;
        RECT 223.185 36.560 223.355 36.730 ;
        RECT 228.640 36.560 228.810 36.730 ;
        RECT 223.185 35.970 223.355 36.140 ;
        RECT 228.640 35.970 228.810 36.140 ;
        RECT 231.490 35.920 231.660 36.090 ;
        RECT 223.185 35.380 223.355 35.550 ;
        RECT 228.640 35.380 228.810 35.550 ;
        RECT 231.160 35.335 231.330 35.505 ;
        RECT 223.185 34.790 223.355 34.960 ;
        RECT 228.640 34.790 228.810 34.960 ;
        RECT 223.185 34.200 223.355 34.370 ;
        RECT 228.640 34.200 228.810 34.370 ;
        RECT 223.185 33.610 223.355 33.780 ;
        RECT 228.640 33.610 228.810 33.780 ;
        RECT 223.185 33.020 223.355 33.190 ;
        RECT 228.640 33.020 228.810 33.190 ;
        RECT 223.185 32.430 223.355 32.600 ;
        RECT 228.640 32.430 228.810 32.600 ;
        RECT 223.185 31.840 223.355 32.010 ;
        RECT 228.640 31.840 228.810 32.010 ;
        RECT 231.160 16.475 231.330 16.645 ;
        RECT 223.185 15.990 223.355 16.160 ;
        RECT 228.640 15.990 228.810 16.160 ;
        RECT 223.185 15.400 223.355 15.570 ;
        RECT 228.640 15.400 228.810 15.570 ;
        RECT 223.185 14.810 223.355 14.980 ;
        RECT 228.640 14.810 228.810 14.980 ;
        RECT 231.490 14.760 231.660 14.930 ;
        RECT 223.185 14.220 223.355 14.390 ;
        RECT 228.640 14.220 228.810 14.390 ;
        RECT 231.160 14.175 231.330 14.345 ;
        RECT -9.495 13.740 -9.325 13.910 ;
        RECT 223.185 13.630 223.355 13.800 ;
        RECT 228.640 13.630 228.810 13.800 ;
        RECT 223.185 13.040 223.355 13.210 ;
        RECT 228.640 13.040 228.810 13.210 ;
        RECT -9.495 12.360 -9.325 12.530 ;
        RECT 223.185 12.450 223.355 12.620 ;
        RECT 228.640 12.450 228.810 12.620 ;
        RECT 223.185 11.860 223.355 12.030 ;
        RECT 228.640 11.860 228.810 12.030 ;
        RECT 223.185 11.270 223.355 11.440 ;
        RECT 228.640 11.270 228.810 11.440 ;
        RECT -9.495 10.980 -9.325 11.150 ;
        RECT 223.185 10.680 223.355 10.850 ;
        RECT 228.640 10.680 228.810 10.850 ;
        RECT -9.495 9.600 -9.325 9.770 ;
        RECT -9.495 8.220 -9.325 8.390 ;
        RECT -9.495 6.840 -9.325 7.010 ;
        RECT -9.495 5.460 -9.325 5.630 ;
        RECT -9.495 4.080 -9.325 4.250 ;
        RECT -9.495 2.700 -9.325 2.870 ;
      LAYER met1 ;
        RECT 223.155 38.640 223.855 38.940 ;
        RECT 104.545 34.865 104.845 35.100 ;
        RECT 106.175 34.865 106.475 35.100 ;
        RECT 104.545 34.635 106.475 34.865 ;
        RECT 104.545 34.400 104.845 34.635 ;
        RECT 106.175 34.400 106.475 34.635 ;
        RECT 115.315 34.865 115.615 35.100 ;
        RECT 116.945 34.865 117.245 35.100 ;
        RECT 115.315 34.635 117.245 34.865 ;
        RECT 115.315 34.400 115.615 34.635 ;
        RECT 116.945 34.400 117.245 34.635 ;
        RECT 223.155 31.780 223.385 38.640 ;
        RECT 231.085 37.590 231.405 37.850 ;
        RECT 228.610 34.930 228.840 37.380 ;
        RECT 231.425 35.570 231.725 36.185 ;
        RECT 231.085 35.270 231.725 35.570 ;
        RECT 228.610 34.230 228.910 34.930 ;
        RECT 228.610 31.780 228.840 34.230 ;
        RECT 108.815 30.665 109.115 30.900 ;
        RECT 110.445 30.665 110.745 30.900 ;
        RECT 108.815 30.435 110.745 30.665 ;
        RECT 108.815 30.200 109.115 30.435 ;
        RECT 110.445 30.200 110.745 30.435 ;
        RECT 111.045 26.465 111.345 26.700 ;
        RECT 112.675 26.465 112.975 26.700 ;
        RECT 111.045 26.235 112.975 26.465 ;
        RECT 111.045 26.000 111.345 26.235 ;
        RECT 112.675 26.000 112.975 26.235 ;
        RECT 104.545 22.265 104.845 22.500 ;
        RECT 106.175 22.265 106.475 22.500 ;
        RECT 104.545 22.035 106.475 22.265 ;
        RECT 104.545 21.800 104.845 22.035 ;
        RECT 106.175 21.800 106.475 22.035 ;
        RECT 115.315 22.265 115.615 22.500 ;
        RECT 116.945 22.265 117.245 22.500 ;
        RECT 115.315 22.035 117.245 22.265 ;
        RECT 115.315 21.800 115.615 22.035 ;
        RECT 116.945 21.800 117.245 22.035 ;
        RECT 223.155 17.480 223.855 17.780 ;
        RECT -9.535 13.665 -9.275 13.985 ;
        RECT -9.535 12.285 -9.275 12.605 ;
        RECT -9.535 10.905 -9.275 11.225 ;
        RECT 223.155 10.620 223.385 17.480 ;
        RECT 231.085 16.430 231.405 16.690 ;
        RECT 228.610 13.770 228.840 16.220 ;
        RECT 231.425 14.410 231.725 15.025 ;
        RECT 231.085 14.110 231.725 14.410 ;
        RECT 228.610 13.070 228.910 13.770 ;
        RECT 228.610 10.620 228.840 13.070 ;
        RECT -9.535 9.525 -9.275 9.845 ;
        RECT -9.535 8.145 -9.275 8.465 ;
        RECT -9.535 6.765 -9.275 7.085 ;
        RECT -9.535 5.385 -9.275 5.705 ;
        RECT -9.535 4.005 -9.275 4.325 ;
        RECT -9.535 2.625 -9.275 2.945 ;
      LAYER via ;
        RECT 223.215 38.660 223.475 38.920 ;
        RECT 223.535 38.660 223.795 38.920 ;
        RECT 104.565 34.780 104.825 35.040 ;
        RECT 106.195 34.780 106.455 35.040 ;
        RECT 104.565 34.460 104.825 34.720 ;
        RECT 106.195 34.460 106.455 34.720 ;
        RECT 115.335 34.780 115.595 35.040 ;
        RECT 116.965 34.780 117.225 35.040 ;
        RECT 115.335 34.460 115.595 34.720 ;
        RECT 116.965 34.460 117.225 34.720 ;
        RECT 231.115 37.590 231.375 37.850 ;
        RECT 231.115 35.290 231.375 35.550 ;
        RECT 228.630 34.610 228.890 34.870 ;
        RECT 228.630 34.290 228.890 34.550 ;
        RECT 108.835 30.580 109.095 30.840 ;
        RECT 110.465 30.580 110.725 30.840 ;
        RECT 108.835 30.260 109.095 30.520 ;
        RECT 110.465 30.260 110.725 30.520 ;
        RECT 111.065 26.380 111.325 26.640 ;
        RECT 112.695 26.380 112.955 26.640 ;
        RECT 111.065 26.060 111.325 26.320 ;
        RECT 112.695 26.060 112.955 26.320 ;
        RECT 104.565 22.180 104.825 22.440 ;
        RECT 106.195 22.180 106.455 22.440 ;
        RECT 104.565 21.860 104.825 22.120 ;
        RECT 106.195 21.860 106.455 22.120 ;
        RECT 115.335 22.180 115.595 22.440 ;
        RECT 116.965 22.180 117.225 22.440 ;
        RECT 115.335 21.860 115.595 22.120 ;
        RECT 116.965 21.860 117.225 22.120 ;
        RECT 223.215 17.500 223.475 17.760 ;
        RECT 223.535 17.500 223.795 17.760 ;
        RECT -9.535 13.695 -9.275 13.955 ;
        RECT -9.535 12.315 -9.275 12.575 ;
        RECT -9.535 10.935 -9.275 11.195 ;
        RECT 231.115 16.430 231.375 16.690 ;
        RECT 231.115 14.130 231.375 14.390 ;
        RECT 228.630 13.450 228.890 13.710 ;
        RECT 228.630 13.130 228.890 13.390 ;
        RECT -9.535 9.555 -9.275 9.815 ;
        RECT -9.535 8.175 -9.275 8.435 ;
        RECT -9.535 6.795 -9.275 7.055 ;
        RECT -9.535 5.415 -9.275 5.675 ;
        RECT -9.535 4.035 -9.275 4.295 ;
        RECT -9.535 2.655 -9.275 2.915 ;
      LAYER met2 ;
        RECT 2.125 46.950 2.525 47.750 ;
        RECT 4.765 46.950 5.165 47.750 ;
        RECT 2.125 42.750 2.525 43.550 ;
        RECT 4.765 42.750 5.165 43.550 ;
        RECT 2.125 38.550 2.525 39.350 ;
        RECT 4.765 38.550 5.165 39.350 ;
        RECT 2.125 34.350 2.525 35.150 ;
        RECT 4.765 34.350 5.165 35.150 ;
        RECT 2.125 30.150 2.525 30.950 ;
        RECT 4.765 30.150 5.165 30.950 ;
        RECT 2.125 25.950 2.525 26.750 ;
        RECT 4.765 25.950 5.165 26.750 ;
        RECT 2.125 21.750 2.525 22.550 ;
        RECT 4.765 21.750 5.165 22.550 ;
        RECT 2.125 17.550 2.525 18.350 ;
        RECT 4.765 17.550 5.165 18.350 ;
        RECT -9.620 13.620 -7.250 14.020 ;
        RECT 2.125 13.350 2.525 14.150 ;
        RECT 4.765 13.350 5.165 14.150 ;
        RECT -9.620 12.240 -7.250 12.640 ;
        RECT -9.620 10.860 -7.250 11.260 ;
        RECT -9.620 9.480 -7.250 9.880 ;
        RECT 2.125 9.150 2.525 9.950 ;
        RECT 4.765 9.150 5.165 9.950 ;
        RECT -9.620 8.100 -7.250 8.500 ;
        RECT 5.645 8.050 6.145 48.850 ;
        RECT 7.645 43.300 8.145 48.850 ;
        RECT 8.625 46.950 9.025 47.750 ;
        RECT 11.265 46.950 11.665 47.750 ;
        RECT 8.625 43.300 9.025 43.550 ;
        RECT 7.645 43.000 9.025 43.300 ;
        RECT 7.645 39.100 8.145 43.000 ;
        RECT 8.625 42.750 9.025 43.000 ;
        RECT 11.265 42.750 11.665 43.550 ;
        RECT 8.625 39.100 9.025 39.350 ;
        RECT 7.645 38.800 9.025 39.100 ;
        RECT 7.645 34.900 8.145 38.800 ;
        RECT 8.625 38.550 9.025 38.800 ;
        RECT 11.265 38.550 11.665 39.350 ;
        RECT 8.625 34.900 9.025 35.150 ;
        RECT 7.645 34.600 9.025 34.900 ;
        RECT 7.645 30.700 8.145 34.600 ;
        RECT 8.625 34.350 9.025 34.600 ;
        RECT 11.265 34.350 11.665 35.150 ;
        RECT 8.625 30.700 9.025 30.950 ;
        RECT 7.645 30.400 9.025 30.700 ;
        RECT 7.645 26.500 8.145 30.400 ;
        RECT 8.625 30.150 9.025 30.400 ;
        RECT 11.265 30.150 11.665 30.950 ;
        RECT 8.625 26.500 9.025 26.750 ;
        RECT 7.645 26.200 9.025 26.500 ;
        RECT 7.645 22.300 8.145 26.200 ;
        RECT 8.625 25.950 9.025 26.200 ;
        RECT 11.265 25.950 11.665 26.750 ;
        RECT 8.625 22.300 9.025 22.550 ;
        RECT 7.645 22.000 9.025 22.300 ;
        RECT 7.645 18.100 8.145 22.000 ;
        RECT 8.625 21.750 9.025 22.000 ;
        RECT 11.265 21.750 11.665 22.550 ;
        RECT 8.625 18.100 9.025 18.350 ;
        RECT 7.645 17.800 9.025 18.100 ;
        RECT 7.645 13.900 8.145 17.800 ;
        RECT 8.625 17.550 9.025 17.800 ;
        RECT 11.265 17.550 11.665 18.350 ;
        RECT 8.625 13.900 9.025 14.150 ;
        RECT 7.645 13.600 9.025 13.900 ;
        RECT -9.620 6.720 -7.250 7.120 ;
        RECT -9.620 5.340 -7.250 5.740 ;
        RECT -9.620 3.960 -7.250 4.360 ;
        RECT -9.620 2.580 -7.250 2.980 ;
        RECT 7.645 2.690 8.145 13.600 ;
        RECT 8.625 13.350 9.025 13.600 ;
        RECT 11.265 13.350 11.665 14.150 ;
        RECT 8.625 9.150 9.025 9.950 ;
        RECT 11.265 9.150 11.665 9.950 ;
        RECT 12.145 8.050 12.645 48.850 ;
        RECT 14.145 43.300 14.645 48.850 ;
        RECT 15.125 46.950 15.525 47.750 ;
        RECT 17.765 46.950 18.165 47.750 ;
        RECT 15.125 43.300 15.525 43.550 ;
        RECT 14.145 43.000 15.525 43.300 ;
        RECT 14.145 39.100 14.645 43.000 ;
        RECT 15.125 42.750 15.525 43.000 ;
        RECT 17.765 42.750 18.165 43.550 ;
        RECT 15.125 39.100 15.525 39.350 ;
        RECT 14.145 38.800 15.525 39.100 ;
        RECT 14.145 34.900 14.645 38.800 ;
        RECT 15.125 38.550 15.525 38.800 ;
        RECT 17.765 38.550 18.165 39.350 ;
        RECT 15.125 34.900 15.525 35.150 ;
        RECT 14.145 34.600 15.525 34.900 ;
        RECT 14.145 30.700 14.645 34.600 ;
        RECT 15.125 34.350 15.525 34.600 ;
        RECT 17.765 34.350 18.165 35.150 ;
        RECT 15.125 30.700 15.525 30.950 ;
        RECT 14.145 30.400 15.525 30.700 ;
        RECT 14.145 26.500 14.645 30.400 ;
        RECT 15.125 30.150 15.525 30.400 ;
        RECT 17.765 30.150 18.165 30.950 ;
        RECT 15.125 26.500 15.525 26.750 ;
        RECT 14.145 26.200 15.525 26.500 ;
        RECT 14.145 22.300 14.645 26.200 ;
        RECT 15.125 25.950 15.525 26.200 ;
        RECT 17.765 25.950 18.165 26.750 ;
        RECT 15.125 22.300 15.525 22.550 ;
        RECT 14.145 22.000 15.525 22.300 ;
        RECT 14.145 18.100 14.645 22.000 ;
        RECT 15.125 21.750 15.525 22.000 ;
        RECT 17.765 21.750 18.165 22.550 ;
        RECT 15.125 18.100 15.525 18.350 ;
        RECT 14.145 17.800 15.525 18.100 ;
        RECT 14.145 13.900 14.645 17.800 ;
        RECT 15.125 17.550 15.525 17.800 ;
        RECT 17.765 17.550 18.165 18.350 ;
        RECT 15.125 13.900 15.525 14.150 ;
        RECT 14.145 13.600 15.525 13.900 ;
        RECT 14.145 3.490 14.645 13.600 ;
        RECT 15.125 13.350 15.525 13.600 ;
        RECT 17.765 13.350 18.165 14.150 ;
        RECT 15.125 9.150 15.525 9.950 ;
        RECT 17.765 9.150 18.165 9.950 ;
        RECT 18.645 8.050 19.145 48.850 ;
        RECT 20.645 43.300 21.145 48.850 ;
        RECT 21.625 46.950 22.025 47.750 ;
        RECT 24.265 46.950 24.665 47.750 ;
        RECT 21.625 43.300 22.025 43.550 ;
        RECT 20.645 43.000 22.025 43.300 ;
        RECT 20.645 39.100 21.145 43.000 ;
        RECT 21.625 42.750 22.025 43.000 ;
        RECT 24.265 42.750 24.665 43.550 ;
        RECT 21.625 39.100 22.025 39.350 ;
        RECT 20.645 38.800 22.025 39.100 ;
        RECT 20.645 34.900 21.145 38.800 ;
        RECT 21.625 38.550 22.025 38.800 ;
        RECT 24.265 38.550 24.665 39.350 ;
        RECT 21.625 34.900 22.025 35.150 ;
        RECT 20.645 34.600 22.025 34.900 ;
        RECT 20.645 30.700 21.145 34.600 ;
        RECT 21.625 34.350 22.025 34.600 ;
        RECT 24.265 34.350 24.665 35.150 ;
        RECT 21.625 30.700 22.025 30.950 ;
        RECT 20.645 30.400 22.025 30.700 ;
        RECT 20.645 26.500 21.145 30.400 ;
        RECT 21.625 30.150 22.025 30.400 ;
        RECT 24.265 30.150 24.665 30.950 ;
        RECT 21.625 26.500 22.025 26.750 ;
        RECT 20.645 26.200 22.025 26.500 ;
        RECT 20.645 22.300 21.145 26.200 ;
        RECT 21.625 25.950 22.025 26.200 ;
        RECT 24.265 25.950 24.665 26.750 ;
        RECT 21.625 22.300 22.025 22.550 ;
        RECT 20.645 22.000 22.025 22.300 ;
        RECT 20.645 18.100 21.145 22.000 ;
        RECT 21.625 21.750 22.025 22.000 ;
        RECT 24.265 21.750 24.665 22.550 ;
        RECT 21.625 18.100 22.025 18.350 ;
        RECT 20.645 17.800 22.025 18.100 ;
        RECT 20.645 13.900 21.145 17.800 ;
        RECT 21.625 17.550 22.025 17.800 ;
        RECT 24.265 17.550 24.665 18.350 ;
        RECT 21.625 13.900 22.025 14.150 ;
        RECT 20.645 13.600 22.025 13.900 ;
        RECT 14.145 3.090 14.945 3.490 ;
        RECT 20.645 2.690 21.145 13.600 ;
        RECT 21.625 13.350 22.025 13.600 ;
        RECT 24.265 13.350 24.665 14.150 ;
        RECT 21.625 9.150 22.025 9.950 ;
        RECT 24.265 9.150 24.665 9.950 ;
        RECT 25.145 8.050 25.645 48.850 ;
        RECT 27.145 43.300 27.645 48.850 ;
        RECT 28.125 46.950 28.525 47.750 ;
        RECT 30.765 46.950 31.165 47.750 ;
        RECT 28.125 43.300 28.525 43.550 ;
        RECT 27.145 43.000 28.525 43.300 ;
        RECT 27.145 39.100 27.645 43.000 ;
        RECT 28.125 42.750 28.525 43.000 ;
        RECT 30.765 42.750 31.165 43.550 ;
        RECT 28.125 39.100 28.525 39.350 ;
        RECT 27.145 38.800 28.525 39.100 ;
        RECT 27.145 34.900 27.645 38.800 ;
        RECT 28.125 38.550 28.525 38.800 ;
        RECT 30.765 38.550 31.165 39.350 ;
        RECT 28.125 34.900 28.525 35.150 ;
        RECT 27.145 34.600 28.525 34.900 ;
        RECT 27.145 30.700 27.645 34.600 ;
        RECT 28.125 34.350 28.525 34.600 ;
        RECT 30.765 34.350 31.165 35.150 ;
        RECT 28.125 30.700 28.525 30.950 ;
        RECT 27.145 30.400 28.525 30.700 ;
        RECT 27.145 26.500 27.645 30.400 ;
        RECT 28.125 30.150 28.525 30.400 ;
        RECT 30.765 30.150 31.165 30.950 ;
        RECT 28.125 26.500 28.525 26.750 ;
        RECT 27.145 26.200 28.525 26.500 ;
        RECT 27.145 22.300 27.645 26.200 ;
        RECT 28.125 25.950 28.525 26.200 ;
        RECT 30.765 25.950 31.165 26.750 ;
        RECT 28.125 22.300 28.525 22.550 ;
        RECT 27.145 22.000 28.525 22.300 ;
        RECT 27.145 18.100 27.645 22.000 ;
        RECT 28.125 21.750 28.525 22.000 ;
        RECT 30.765 21.750 31.165 22.550 ;
        RECT 28.125 18.100 28.525 18.350 ;
        RECT 27.145 17.800 28.525 18.100 ;
        RECT 27.145 13.900 27.645 17.800 ;
        RECT 28.125 17.550 28.525 17.800 ;
        RECT 30.765 17.550 31.165 18.350 ;
        RECT 28.125 13.900 28.525 14.150 ;
        RECT 27.145 13.600 28.525 13.900 ;
        RECT 27.145 2.690 27.645 13.600 ;
        RECT 28.125 13.350 28.525 13.600 ;
        RECT 30.765 13.350 31.165 14.150 ;
        RECT 28.125 9.150 28.525 9.950 ;
        RECT 30.765 9.150 31.165 9.950 ;
        RECT 31.645 8.050 32.145 48.850 ;
        RECT 33.645 43.300 34.145 48.850 ;
        RECT 34.625 46.950 35.025 47.750 ;
        RECT 37.265 46.950 37.665 47.750 ;
        RECT 34.625 43.300 35.025 43.550 ;
        RECT 33.645 43.000 35.025 43.300 ;
        RECT 33.645 39.100 34.145 43.000 ;
        RECT 34.625 42.750 35.025 43.000 ;
        RECT 37.265 42.750 37.665 43.550 ;
        RECT 34.625 39.100 35.025 39.350 ;
        RECT 33.645 38.800 35.025 39.100 ;
        RECT 33.645 34.900 34.145 38.800 ;
        RECT 34.625 38.550 35.025 38.800 ;
        RECT 37.265 38.550 37.665 39.350 ;
        RECT 34.625 34.900 35.025 35.150 ;
        RECT 33.645 34.600 35.025 34.900 ;
        RECT 33.645 30.700 34.145 34.600 ;
        RECT 34.625 34.350 35.025 34.600 ;
        RECT 37.265 34.350 37.665 35.150 ;
        RECT 34.625 30.700 35.025 30.950 ;
        RECT 33.645 30.400 35.025 30.700 ;
        RECT 33.645 26.500 34.145 30.400 ;
        RECT 34.625 30.150 35.025 30.400 ;
        RECT 37.265 30.150 37.665 30.950 ;
        RECT 34.625 26.500 35.025 26.750 ;
        RECT 33.645 26.200 35.025 26.500 ;
        RECT 33.645 22.300 34.145 26.200 ;
        RECT 34.625 25.950 35.025 26.200 ;
        RECT 37.265 25.950 37.665 26.750 ;
        RECT 34.625 22.300 35.025 22.550 ;
        RECT 33.645 22.000 35.025 22.300 ;
        RECT 33.645 18.100 34.145 22.000 ;
        RECT 34.625 21.750 35.025 22.000 ;
        RECT 37.265 21.750 37.665 22.550 ;
        RECT 34.625 18.100 35.025 18.350 ;
        RECT 33.645 17.800 35.025 18.100 ;
        RECT 33.645 13.900 34.145 17.800 ;
        RECT 34.625 17.550 35.025 17.800 ;
        RECT 37.265 17.550 37.665 18.350 ;
        RECT 34.625 13.900 35.025 14.150 ;
        RECT 33.645 13.600 35.025 13.900 ;
        RECT 33.645 3.490 34.145 13.600 ;
        RECT 34.625 13.350 35.025 13.600 ;
        RECT 37.265 13.350 37.665 14.150 ;
        RECT 34.625 9.150 35.025 9.950 ;
        RECT 37.265 9.150 37.665 9.950 ;
        RECT 38.145 8.050 38.645 48.850 ;
        RECT 40.145 43.300 40.645 48.850 ;
        RECT 41.125 46.950 41.525 47.750 ;
        RECT 43.765 46.950 44.165 47.750 ;
        RECT 41.125 43.300 41.525 43.550 ;
        RECT 40.145 43.000 41.525 43.300 ;
        RECT 40.145 39.100 40.645 43.000 ;
        RECT 41.125 42.750 41.525 43.000 ;
        RECT 43.765 42.750 44.165 43.550 ;
        RECT 41.125 39.100 41.525 39.350 ;
        RECT 40.145 38.800 41.525 39.100 ;
        RECT 40.145 34.900 40.645 38.800 ;
        RECT 41.125 38.550 41.525 38.800 ;
        RECT 43.765 38.550 44.165 39.350 ;
        RECT 41.125 34.900 41.525 35.150 ;
        RECT 40.145 34.600 41.525 34.900 ;
        RECT 40.145 30.700 40.645 34.600 ;
        RECT 41.125 34.350 41.525 34.600 ;
        RECT 43.765 34.350 44.165 35.150 ;
        RECT 41.125 30.700 41.525 30.950 ;
        RECT 40.145 30.400 41.525 30.700 ;
        RECT 40.145 26.500 40.645 30.400 ;
        RECT 41.125 30.150 41.525 30.400 ;
        RECT 43.765 30.150 44.165 30.950 ;
        RECT 41.125 26.500 41.525 26.750 ;
        RECT 40.145 26.200 41.525 26.500 ;
        RECT 40.145 22.300 40.645 26.200 ;
        RECT 41.125 25.950 41.525 26.200 ;
        RECT 43.765 25.950 44.165 26.750 ;
        RECT 41.125 22.300 41.525 22.550 ;
        RECT 40.145 22.000 41.525 22.300 ;
        RECT 40.145 18.100 40.645 22.000 ;
        RECT 41.125 21.750 41.525 22.000 ;
        RECT 43.765 21.750 44.165 22.550 ;
        RECT 41.125 18.100 41.525 18.350 ;
        RECT 40.145 17.800 41.525 18.100 ;
        RECT 40.145 13.900 40.645 17.800 ;
        RECT 41.125 17.550 41.525 17.800 ;
        RECT 43.765 17.550 44.165 18.350 ;
        RECT 41.125 13.900 41.525 14.150 ;
        RECT 40.145 13.600 41.525 13.900 ;
        RECT 33.645 3.090 34.445 3.490 ;
        RECT 40.145 2.690 40.645 13.600 ;
        RECT 41.125 13.350 41.525 13.600 ;
        RECT 43.765 13.350 44.165 14.150 ;
        RECT 41.125 9.150 41.525 9.950 ;
        RECT 43.765 9.150 44.165 9.950 ;
        RECT 44.645 8.050 45.145 48.850 ;
        RECT 46.645 43.300 47.145 48.850 ;
        RECT 47.625 46.950 48.025 47.750 ;
        RECT 50.265 46.950 50.665 47.750 ;
        RECT 47.625 43.300 48.025 43.550 ;
        RECT 46.645 43.000 48.025 43.300 ;
        RECT 46.645 39.100 47.145 43.000 ;
        RECT 47.625 42.750 48.025 43.000 ;
        RECT 50.265 42.750 50.665 43.550 ;
        RECT 47.625 39.100 48.025 39.350 ;
        RECT 46.645 38.800 48.025 39.100 ;
        RECT 46.645 34.900 47.145 38.800 ;
        RECT 47.625 38.550 48.025 38.800 ;
        RECT 50.265 38.550 50.665 39.350 ;
        RECT 47.625 34.900 48.025 35.150 ;
        RECT 46.645 34.600 48.025 34.900 ;
        RECT 46.645 30.700 47.145 34.600 ;
        RECT 47.625 34.350 48.025 34.600 ;
        RECT 50.265 34.350 50.665 35.150 ;
        RECT 47.625 30.700 48.025 30.950 ;
        RECT 46.645 30.400 48.025 30.700 ;
        RECT 46.645 26.500 47.145 30.400 ;
        RECT 47.625 30.150 48.025 30.400 ;
        RECT 50.265 30.150 50.665 30.950 ;
        RECT 47.625 26.500 48.025 26.750 ;
        RECT 46.645 26.200 48.025 26.500 ;
        RECT 46.645 22.300 47.145 26.200 ;
        RECT 47.625 25.950 48.025 26.200 ;
        RECT 50.265 25.950 50.665 26.750 ;
        RECT 47.625 22.300 48.025 22.550 ;
        RECT 46.645 22.000 48.025 22.300 ;
        RECT 46.645 18.100 47.145 22.000 ;
        RECT 47.625 21.750 48.025 22.000 ;
        RECT 50.265 21.750 50.665 22.550 ;
        RECT 47.625 18.100 48.025 18.350 ;
        RECT 46.645 17.800 48.025 18.100 ;
        RECT 46.645 13.900 47.145 17.800 ;
        RECT 47.625 17.550 48.025 17.800 ;
        RECT 50.265 17.550 50.665 18.350 ;
        RECT 47.625 13.900 48.025 14.150 ;
        RECT 46.645 13.600 48.025 13.900 ;
        RECT 46.645 2.690 47.145 13.600 ;
        RECT 47.625 13.350 48.025 13.600 ;
        RECT 50.265 13.350 50.665 14.150 ;
        RECT 47.625 9.150 48.025 9.950 ;
        RECT 50.265 9.150 50.665 9.950 ;
        RECT 51.145 8.050 51.645 48.850 ;
        RECT 53.145 43.300 53.645 48.850 ;
        RECT 54.125 46.950 54.525 47.750 ;
        RECT 56.765 46.950 57.165 47.750 ;
        RECT 54.125 43.300 54.525 43.550 ;
        RECT 53.145 43.000 54.525 43.300 ;
        RECT 53.145 39.100 53.645 43.000 ;
        RECT 54.125 42.750 54.525 43.000 ;
        RECT 56.765 42.750 57.165 43.550 ;
        RECT 54.125 39.100 54.525 39.350 ;
        RECT 53.145 38.800 54.525 39.100 ;
        RECT 53.145 34.900 53.645 38.800 ;
        RECT 54.125 38.550 54.525 38.800 ;
        RECT 56.765 38.550 57.165 39.350 ;
        RECT 54.125 34.900 54.525 35.150 ;
        RECT 53.145 34.600 54.525 34.900 ;
        RECT 53.145 30.700 53.645 34.600 ;
        RECT 54.125 34.350 54.525 34.600 ;
        RECT 56.765 34.350 57.165 35.150 ;
        RECT 54.125 30.700 54.525 30.950 ;
        RECT 53.145 30.400 54.525 30.700 ;
        RECT 53.145 26.500 53.645 30.400 ;
        RECT 54.125 30.150 54.525 30.400 ;
        RECT 56.765 30.150 57.165 30.950 ;
        RECT 54.125 26.500 54.525 26.750 ;
        RECT 53.145 26.200 54.525 26.500 ;
        RECT 53.145 22.300 53.645 26.200 ;
        RECT 54.125 25.950 54.525 26.200 ;
        RECT 56.765 25.950 57.165 26.750 ;
        RECT 54.125 22.300 54.525 22.550 ;
        RECT 53.145 22.000 54.525 22.300 ;
        RECT 53.145 18.100 53.645 22.000 ;
        RECT 54.125 21.750 54.525 22.000 ;
        RECT 56.765 21.750 57.165 22.550 ;
        RECT 54.125 18.100 54.525 18.350 ;
        RECT 53.145 17.800 54.525 18.100 ;
        RECT 53.145 13.900 53.645 17.800 ;
        RECT 54.125 17.550 54.525 17.800 ;
        RECT 56.765 17.550 57.165 18.350 ;
        RECT 54.125 13.900 54.525 14.150 ;
        RECT 53.145 13.600 54.525 13.900 ;
        RECT 53.145 4.290 53.645 13.600 ;
        RECT 54.125 13.350 54.525 13.600 ;
        RECT 56.765 13.350 57.165 14.150 ;
        RECT 54.125 9.150 54.525 9.950 ;
        RECT 56.765 9.150 57.165 9.950 ;
        RECT 57.645 8.050 58.145 48.850 ;
        RECT 59.645 43.300 60.145 48.850 ;
        RECT 60.625 46.950 61.025 47.750 ;
        RECT 63.265 46.950 63.665 47.750 ;
        RECT 60.625 43.300 61.025 43.550 ;
        RECT 59.645 43.000 61.025 43.300 ;
        RECT 59.645 39.100 60.145 43.000 ;
        RECT 60.625 42.750 61.025 43.000 ;
        RECT 63.265 42.750 63.665 43.550 ;
        RECT 60.625 39.100 61.025 39.350 ;
        RECT 59.645 38.800 61.025 39.100 ;
        RECT 59.645 34.900 60.145 38.800 ;
        RECT 60.625 38.550 61.025 38.800 ;
        RECT 63.265 38.550 63.665 39.350 ;
        RECT 60.625 34.900 61.025 35.150 ;
        RECT 59.645 34.600 61.025 34.900 ;
        RECT 59.645 30.700 60.145 34.600 ;
        RECT 60.625 34.350 61.025 34.600 ;
        RECT 63.265 34.350 63.665 35.150 ;
        RECT 60.625 30.700 61.025 30.950 ;
        RECT 59.645 30.400 61.025 30.700 ;
        RECT 59.645 26.500 60.145 30.400 ;
        RECT 60.625 30.150 61.025 30.400 ;
        RECT 63.265 30.150 63.665 30.950 ;
        RECT 60.625 26.500 61.025 26.750 ;
        RECT 59.645 26.200 61.025 26.500 ;
        RECT 59.645 22.300 60.145 26.200 ;
        RECT 60.625 25.950 61.025 26.200 ;
        RECT 63.265 25.950 63.665 26.750 ;
        RECT 60.625 22.300 61.025 22.550 ;
        RECT 59.645 22.000 61.025 22.300 ;
        RECT 59.645 18.100 60.145 22.000 ;
        RECT 60.625 21.750 61.025 22.000 ;
        RECT 63.265 21.750 63.665 22.550 ;
        RECT 60.625 18.100 61.025 18.350 ;
        RECT 59.645 17.800 61.025 18.100 ;
        RECT 59.645 13.900 60.145 17.800 ;
        RECT 60.625 17.550 61.025 17.800 ;
        RECT 63.265 17.550 63.665 18.350 ;
        RECT 60.625 13.900 61.025 14.150 ;
        RECT 59.645 13.600 61.025 13.900 ;
        RECT 53.145 3.890 53.945 4.290 ;
        RECT 59.645 3.490 60.145 13.600 ;
        RECT 60.625 13.350 61.025 13.600 ;
        RECT 63.265 13.350 63.665 14.150 ;
        RECT 60.625 9.150 61.025 9.950 ;
        RECT 63.265 9.150 63.665 9.950 ;
        RECT 64.145 8.050 64.645 48.850 ;
        RECT 66.145 43.300 66.645 48.850 ;
        RECT 67.125 46.950 67.525 47.750 ;
        RECT 69.765 46.950 70.165 47.750 ;
        RECT 67.125 43.300 67.525 43.550 ;
        RECT 66.145 43.000 67.525 43.300 ;
        RECT 66.145 39.100 66.645 43.000 ;
        RECT 67.125 42.750 67.525 43.000 ;
        RECT 69.765 42.750 70.165 43.550 ;
        RECT 67.125 39.100 67.525 39.350 ;
        RECT 66.145 38.800 67.525 39.100 ;
        RECT 66.145 34.900 66.645 38.800 ;
        RECT 67.125 38.550 67.525 38.800 ;
        RECT 69.765 38.550 70.165 39.350 ;
        RECT 67.125 34.900 67.525 35.150 ;
        RECT 66.145 34.600 67.525 34.900 ;
        RECT 66.145 30.700 66.645 34.600 ;
        RECT 67.125 34.350 67.525 34.600 ;
        RECT 69.765 34.350 70.165 35.150 ;
        RECT 67.125 30.700 67.525 30.950 ;
        RECT 66.145 30.400 67.525 30.700 ;
        RECT 66.145 26.500 66.645 30.400 ;
        RECT 67.125 30.150 67.525 30.400 ;
        RECT 69.765 30.150 70.165 30.950 ;
        RECT 67.125 26.500 67.525 26.750 ;
        RECT 66.145 26.200 67.525 26.500 ;
        RECT 66.145 22.300 66.645 26.200 ;
        RECT 67.125 25.950 67.525 26.200 ;
        RECT 69.765 25.950 70.165 26.750 ;
        RECT 67.125 22.300 67.525 22.550 ;
        RECT 66.145 22.000 67.525 22.300 ;
        RECT 66.145 18.100 66.645 22.000 ;
        RECT 67.125 21.750 67.525 22.000 ;
        RECT 69.765 21.750 70.165 22.550 ;
        RECT 67.125 18.100 67.525 18.350 ;
        RECT 66.145 17.800 67.525 18.100 ;
        RECT 66.145 13.900 66.645 17.800 ;
        RECT 67.125 17.550 67.525 17.800 ;
        RECT 69.765 17.550 70.165 18.350 ;
        RECT 67.125 13.900 67.525 14.150 ;
        RECT 66.145 13.600 67.525 13.900 ;
        RECT 59.645 3.090 60.445 3.490 ;
        RECT 66.145 2.690 66.645 13.600 ;
        RECT 67.125 13.350 67.525 13.600 ;
        RECT 69.765 13.350 70.165 14.150 ;
        RECT 67.125 9.150 67.525 9.950 ;
        RECT 69.765 9.150 70.165 9.950 ;
        RECT 70.645 8.050 71.145 48.850 ;
        RECT 72.645 43.300 73.145 48.850 ;
        RECT 73.625 46.950 74.025 47.750 ;
        RECT 76.265 46.950 76.665 47.750 ;
        RECT 73.625 43.300 74.025 43.550 ;
        RECT 72.645 43.000 74.025 43.300 ;
        RECT 72.645 39.100 73.145 43.000 ;
        RECT 73.625 42.750 74.025 43.000 ;
        RECT 76.265 42.750 76.665 43.550 ;
        RECT 73.625 39.100 74.025 39.350 ;
        RECT 72.645 38.800 74.025 39.100 ;
        RECT 72.645 34.900 73.145 38.800 ;
        RECT 73.625 38.550 74.025 38.800 ;
        RECT 76.265 38.550 76.665 39.350 ;
        RECT 73.625 34.900 74.025 35.150 ;
        RECT 72.645 34.600 74.025 34.900 ;
        RECT 72.645 30.700 73.145 34.600 ;
        RECT 73.625 34.350 74.025 34.600 ;
        RECT 76.265 34.350 76.665 35.150 ;
        RECT 73.625 30.700 74.025 30.950 ;
        RECT 72.645 30.400 74.025 30.700 ;
        RECT 72.645 26.500 73.145 30.400 ;
        RECT 73.625 30.150 74.025 30.400 ;
        RECT 76.265 30.150 76.665 30.950 ;
        RECT 73.625 26.500 74.025 26.750 ;
        RECT 72.645 26.200 74.025 26.500 ;
        RECT 72.645 22.300 73.145 26.200 ;
        RECT 73.625 25.950 74.025 26.200 ;
        RECT 76.265 25.950 76.665 26.750 ;
        RECT 73.625 22.300 74.025 22.550 ;
        RECT 72.645 22.000 74.025 22.300 ;
        RECT 72.645 18.100 73.145 22.000 ;
        RECT 73.625 21.750 74.025 22.000 ;
        RECT 76.265 21.750 76.665 22.550 ;
        RECT 73.625 18.100 74.025 18.350 ;
        RECT 72.645 17.800 74.025 18.100 ;
        RECT 72.645 13.900 73.145 17.800 ;
        RECT 73.625 17.550 74.025 17.800 ;
        RECT 76.265 17.550 76.665 18.350 ;
        RECT 73.625 13.900 74.025 14.150 ;
        RECT 72.645 13.600 74.025 13.900 ;
        RECT 72.645 2.690 73.145 13.600 ;
        RECT 73.625 13.350 74.025 13.600 ;
        RECT 76.265 13.350 76.665 14.150 ;
        RECT 73.625 9.150 74.025 9.950 ;
        RECT 76.265 9.150 76.665 9.950 ;
        RECT 77.145 8.050 77.645 48.850 ;
        RECT 79.145 43.300 79.645 48.850 ;
        RECT 80.125 46.950 80.525 47.750 ;
        RECT 82.765 46.950 83.165 47.750 ;
        RECT 80.125 43.300 80.525 43.550 ;
        RECT 79.145 43.000 80.525 43.300 ;
        RECT 79.145 39.100 79.645 43.000 ;
        RECT 80.125 42.750 80.525 43.000 ;
        RECT 82.765 42.750 83.165 43.550 ;
        RECT 80.125 39.100 80.525 39.350 ;
        RECT 79.145 38.800 80.525 39.100 ;
        RECT 79.145 34.900 79.645 38.800 ;
        RECT 80.125 38.550 80.525 38.800 ;
        RECT 82.765 38.550 83.165 39.350 ;
        RECT 80.125 34.900 80.525 35.150 ;
        RECT 79.145 34.600 80.525 34.900 ;
        RECT 79.145 30.700 79.645 34.600 ;
        RECT 80.125 34.350 80.525 34.600 ;
        RECT 82.765 34.350 83.165 35.150 ;
        RECT 80.125 30.700 80.525 30.950 ;
        RECT 79.145 30.400 80.525 30.700 ;
        RECT 79.145 26.500 79.645 30.400 ;
        RECT 80.125 30.150 80.525 30.400 ;
        RECT 82.765 30.150 83.165 30.950 ;
        RECT 80.125 26.500 80.525 26.750 ;
        RECT 79.145 26.200 80.525 26.500 ;
        RECT 79.145 22.300 79.645 26.200 ;
        RECT 80.125 25.950 80.525 26.200 ;
        RECT 82.765 25.950 83.165 26.750 ;
        RECT 80.125 22.300 80.525 22.550 ;
        RECT 79.145 22.000 80.525 22.300 ;
        RECT 79.145 18.100 79.645 22.000 ;
        RECT 80.125 21.750 80.525 22.000 ;
        RECT 82.765 21.750 83.165 22.550 ;
        RECT 80.125 18.100 80.525 18.350 ;
        RECT 79.145 17.800 80.525 18.100 ;
        RECT 79.145 13.900 79.645 17.800 ;
        RECT 80.125 17.550 80.525 17.800 ;
        RECT 82.765 17.550 83.165 18.350 ;
        RECT 80.125 13.900 80.525 14.150 ;
        RECT 79.145 13.600 80.525 13.900 ;
        RECT 79.145 4.290 79.645 13.600 ;
        RECT 80.125 13.350 80.525 13.600 ;
        RECT 82.765 13.350 83.165 14.150 ;
        RECT 80.125 9.150 80.525 9.950 ;
        RECT 82.765 9.150 83.165 9.950 ;
        RECT 83.645 8.050 84.145 48.850 ;
        RECT 85.645 43.300 86.145 48.850 ;
        RECT 86.625 46.950 87.025 47.750 ;
        RECT 89.265 46.950 89.665 47.750 ;
        RECT 86.625 43.300 87.025 43.550 ;
        RECT 85.645 43.000 87.025 43.300 ;
        RECT 85.645 39.100 86.145 43.000 ;
        RECT 86.625 42.750 87.025 43.000 ;
        RECT 89.265 42.750 89.665 43.550 ;
        RECT 86.625 39.100 87.025 39.350 ;
        RECT 85.645 38.800 87.025 39.100 ;
        RECT 85.645 34.900 86.145 38.800 ;
        RECT 86.625 38.550 87.025 38.800 ;
        RECT 89.265 38.550 89.665 39.350 ;
        RECT 86.625 34.900 87.025 35.150 ;
        RECT 85.645 34.600 87.025 34.900 ;
        RECT 85.645 30.700 86.145 34.600 ;
        RECT 86.625 34.350 87.025 34.600 ;
        RECT 89.265 34.350 89.665 35.150 ;
        RECT 86.625 30.700 87.025 30.950 ;
        RECT 85.645 30.400 87.025 30.700 ;
        RECT 85.645 26.500 86.145 30.400 ;
        RECT 86.625 30.150 87.025 30.400 ;
        RECT 89.265 30.150 89.665 30.950 ;
        RECT 86.625 26.500 87.025 26.750 ;
        RECT 85.645 26.200 87.025 26.500 ;
        RECT 85.645 22.300 86.145 26.200 ;
        RECT 86.625 25.950 87.025 26.200 ;
        RECT 89.265 25.950 89.665 26.750 ;
        RECT 86.625 22.300 87.025 22.550 ;
        RECT 85.645 22.000 87.025 22.300 ;
        RECT 85.645 18.100 86.145 22.000 ;
        RECT 86.625 21.750 87.025 22.000 ;
        RECT 89.265 21.750 89.665 22.550 ;
        RECT 86.625 18.100 87.025 18.350 ;
        RECT 85.645 17.800 87.025 18.100 ;
        RECT 85.645 13.900 86.145 17.800 ;
        RECT 86.625 17.550 87.025 17.800 ;
        RECT 89.265 17.550 89.665 18.350 ;
        RECT 86.625 13.900 87.025 14.150 ;
        RECT 85.645 13.600 87.025 13.900 ;
        RECT 79.145 3.890 79.945 4.290 ;
        RECT 85.645 3.490 86.145 13.600 ;
        RECT 86.625 13.350 87.025 13.600 ;
        RECT 89.265 13.350 89.665 14.150 ;
        RECT 86.625 9.150 87.025 9.950 ;
        RECT 89.265 9.150 89.665 9.950 ;
        RECT 90.145 8.050 90.645 48.850 ;
        RECT 92.145 43.300 92.645 48.850 ;
        RECT 93.125 46.950 93.525 47.750 ;
        RECT 95.765 46.950 96.165 47.750 ;
        RECT 93.125 43.300 93.525 43.550 ;
        RECT 92.145 43.000 93.525 43.300 ;
        RECT 92.145 39.100 92.645 43.000 ;
        RECT 93.125 42.750 93.525 43.000 ;
        RECT 95.765 42.750 96.165 43.550 ;
        RECT 93.125 39.100 93.525 39.350 ;
        RECT 92.145 38.800 93.525 39.100 ;
        RECT 92.145 34.900 92.645 38.800 ;
        RECT 93.125 38.550 93.525 38.800 ;
        RECT 95.765 38.550 96.165 39.350 ;
        RECT 93.125 34.900 93.525 35.150 ;
        RECT 92.145 34.600 93.525 34.900 ;
        RECT 92.145 30.700 92.645 34.600 ;
        RECT 93.125 34.350 93.525 34.600 ;
        RECT 95.765 34.350 96.165 35.150 ;
        RECT 93.125 30.700 93.525 30.950 ;
        RECT 92.145 30.400 93.525 30.700 ;
        RECT 92.145 26.500 92.645 30.400 ;
        RECT 93.125 30.150 93.525 30.400 ;
        RECT 95.765 30.150 96.165 30.950 ;
        RECT 93.125 26.500 93.525 26.750 ;
        RECT 92.145 26.200 93.525 26.500 ;
        RECT 92.145 22.300 92.645 26.200 ;
        RECT 93.125 25.950 93.525 26.200 ;
        RECT 95.765 25.950 96.165 26.750 ;
        RECT 93.125 22.300 93.525 22.550 ;
        RECT 92.145 22.000 93.525 22.300 ;
        RECT 92.145 18.100 92.645 22.000 ;
        RECT 93.125 21.750 93.525 22.000 ;
        RECT 95.765 21.750 96.165 22.550 ;
        RECT 93.125 18.100 93.525 18.350 ;
        RECT 92.145 17.800 93.525 18.100 ;
        RECT 92.145 13.900 92.645 17.800 ;
        RECT 93.125 17.550 93.525 17.800 ;
        RECT 95.765 17.550 96.165 18.350 ;
        RECT 93.125 13.900 93.525 14.150 ;
        RECT 92.145 13.600 93.525 13.900 ;
        RECT 85.645 3.090 86.445 3.490 ;
        RECT 92.145 2.690 92.645 13.600 ;
        RECT 93.125 13.350 93.525 13.600 ;
        RECT 95.765 13.350 96.165 14.150 ;
        RECT 93.125 9.150 93.525 9.950 ;
        RECT 95.765 9.150 96.165 9.950 ;
        RECT 96.645 8.050 97.145 48.850 ;
        RECT 98.645 43.300 99.145 48.850 ;
        RECT 99.625 46.950 100.025 47.750 ;
        RECT 102.265 46.950 102.665 47.750 ;
        RECT 99.625 43.300 100.025 43.550 ;
        RECT 98.645 43.000 100.025 43.300 ;
        RECT 98.645 39.100 99.145 43.000 ;
        RECT 99.625 42.750 100.025 43.000 ;
        RECT 102.265 42.750 102.665 43.550 ;
        RECT 99.625 39.100 100.025 39.350 ;
        RECT 98.645 38.800 100.025 39.100 ;
        RECT 98.645 34.900 99.145 38.800 ;
        RECT 99.625 38.550 100.025 38.800 ;
        RECT 102.265 38.550 102.665 39.350 ;
        RECT 99.625 34.900 100.025 35.150 ;
        RECT 98.645 34.600 100.025 34.900 ;
        RECT 98.645 30.700 99.145 34.600 ;
        RECT 99.625 34.350 100.025 34.600 ;
        RECT 102.265 34.350 102.665 35.150 ;
        RECT 99.625 30.700 100.025 30.950 ;
        RECT 98.645 30.400 100.025 30.700 ;
        RECT 98.645 26.500 99.145 30.400 ;
        RECT 99.625 30.150 100.025 30.400 ;
        RECT 102.265 30.150 102.665 30.950 ;
        RECT 99.625 26.500 100.025 26.750 ;
        RECT 98.645 26.200 100.025 26.500 ;
        RECT 98.645 22.300 99.145 26.200 ;
        RECT 99.625 25.950 100.025 26.200 ;
        RECT 102.265 25.950 102.665 26.750 ;
        RECT 99.625 22.300 100.025 22.550 ;
        RECT 98.645 22.000 100.025 22.300 ;
        RECT 98.645 18.100 99.145 22.000 ;
        RECT 99.625 21.750 100.025 22.000 ;
        RECT 102.265 21.750 102.665 22.550 ;
        RECT 99.625 18.100 100.025 18.350 ;
        RECT 98.645 17.800 100.025 18.100 ;
        RECT 98.645 13.900 99.145 17.800 ;
        RECT 99.625 17.550 100.025 17.800 ;
        RECT 102.265 17.550 102.665 18.350 ;
        RECT 99.625 13.900 100.025 14.150 ;
        RECT 98.645 13.600 100.025 13.900 ;
        RECT 98.645 5.090 99.145 13.600 ;
        RECT 99.625 13.350 100.025 13.600 ;
        RECT 102.265 13.350 102.665 14.150 ;
        RECT 99.625 9.150 100.025 9.950 ;
        RECT 102.265 9.150 102.665 9.950 ;
        RECT 103.145 8.050 103.645 48.850 ;
        RECT 105.145 43.300 105.645 48.850 ;
        RECT 106.125 46.950 106.525 47.750 ;
        RECT 108.765 46.950 109.165 47.750 ;
        RECT 106.125 43.300 106.525 43.550 ;
        RECT 105.145 43.000 106.525 43.300 ;
        RECT 105.145 39.100 105.645 43.000 ;
        RECT 106.125 42.750 106.525 43.000 ;
        RECT 108.765 42.750 109.165 43.550 ;
        RECT 106.125 39.100 106.525 39.350 ;
        RECT 105.145 38.800 106.525 39.100 ;
        RECT 104.495 34.350 104.895 35.150 ;
        RECT 104.495 21.750 104.895 22.550 ;
        RECT 105.145 18.100 105.645 38.800 ;
        RECT 106.125 38.550 106.525 38.800 ;
        RECT 108.765 38.550 109.165 39.350 ;
        RECT 106.125 34.350 106.525 35.150 ;
        RECT 108.765 34.350 109.165 35.150 ;
        RECT 106.125 30.150 106.525 30.950 ;
        RECT 108.765 30.150 109.165 30.950 ;
        RECT 106.125 25.950 106.525 26.750 ;
        RECT 108.765 26.500 109.165 26.750 ;
        RECT 109.645 26.500 110.145 48.850 ;
        RECT 110.395 30.150 110.795 30.950 ;
        RECT 111.645 30.695 112.145 48.850 ;
        RECT 112.625 46.950 113.025 47.750 ;
        RECT 115.265 46.950 115.665 47.750 ;
        RECT 112.625 42.750 113.025 43.550 ;
        RECT 115.265 43.300 115.665 43.550 ;
        RECT 116.145 43.300 116.645 48.850 ;
        RECT 115.265 43.000 116.645 43.300 ;
        RECT 115.265 42.750 115.665 43.000 ;
        RECT 112.625 38.550 113.025 39.350 ;
        RECT 115.265 39.100 115.665 39.350 ;
        RECT 116.145 39.100 116.645 43.000 ;
        RECT 115.265 38.800 116.645 39.100 ;
        RECT 115.265 38.550 115.665 38.800 ;
        RECT 112.625 34.350 113.025 35.150 ;
        RECT 115.265 34.350 115.665 35.150 ;
        RECT 112.625 30.695 113.025 30.950 ;
        RECT 111.645 30.395 113.025 30.695 ;
        RECT 108.765 26.200 110.145 26.500 ;
        RECT 108.765 25.950 109.165 26.200 ;
        RECT 106.125 21.750 106.525 22.550 ;
        RECT 108.765 21.750 109.165 22.550 ;
        RECT 106.125 18.100 106.525 18.350 ;
        RECT 105.145 17.800 106.525 18.100 ;
        RECT 105.145 13.900 105.645 17.800 ;
        RECT 106.125 17.550 106.525 17.800 ;
        RECT 108.765 17.550 109.165 18.350 ;
        RECT 106.125 13.900 106.525 14.150 ;
        RECT 105.145 13.600 106.525 13.900 ;
        RECT 105.145 5.890 105.645 13.600 ;
        RECT 106.125 13.350 106.525 13.600 ;
        RECT 108.765 13.350 109.165 14.150 ;
        RECT 106.125 9.150 106.525 9.950 ;
        RECT 108.765 9.150 109.165 9.950 ;
        RECT 109.645 7.490 110.145 26.200 ;
        RECT 110.995 25.950 111.395 26.750 ;
        RECT 111.645 7.490 112.145 30.395 ;
        RECT 112.625 30.150 113.025 30.395 ;
        RECT 115.265 30.150 115.665 30.950 ;
        RECT 112.625 25.950 113.025 26.750 ;
        RECT 115.265 25.950 115.665 26.750 ;
        RECT 112.625 21.750 113.025 22.550 ;
        RECT 115.265 21.750 115.665 22.550 ;
        RECT 112.625 17.550 113.025 18.350 ;
        RECT 115.265 18.100 115.665 18.350 ;
        RECT 116.145 18.100 116.645 38.800 ;
        RECT 116.895 34.350 117.295 35.150 ;
        RECT 116.895 21.750 117.295 22.550 ;
        RECT 115.265 17.800 116.645 18.100 ;
        RECT 115.265 17.550 115.665 17.800 ;
        RECT 112.625 13.350 113.025 14.150 ;
        RECT 115.265 13.900 115.665 14.150 ;
        RECT 116.145 13.900 116.645 17.800 ;
        RECT 115.265 13.600 116.645 13.900 ;
        RECT 115.265 13.350 115.665 13.600 ;
        RECT 112.625 9.150 113.025 9.950 ;
        RECT 115.265 9.150 115.665 9.950 ;
        RECT 108.145 7.090 108.945 7.490 ;
        RECT 109.645 7.090 112.145 7.490 ;
        RECT 112.845 7.090 113.645 7.490 ;
        RECT 105.145 5.490 105.945 5.890 ;
        RECT 98.645 4.690 99.445 5.090 ;
        RECT 7.645 2.290 8.445 2.690 ;
        RECT 20.645 2.290 21.445 2.690 ;
        RECT 27.145 2.290 27.945 2.690 ;
        RECT 40.145 2.290 40.945 2.690 ;
        RECT 46.645 2.290 47.445 2.690 ;
        RECT 66.145 2.290 66.945 2.690 ;
        RECT 72.645 2.290 73.445 2.690 ;
        RECT 92.145 2.290 92.945 2.690 ;
        RECT 108.145 1.090 108.645 7.090 ;
        RECT 110.645 1.890 111.145 7.090 ;
        RECT 110.345 1.490 111.145 1.890 ;
        RECT 107.845 0.690 108.645 1.090 ;
        RECT 113.145 0.290 113.645 7.090 ;
        RECT 116.145 5.890 116.645 13.600 ;
        RECT 118.145 8.050 118.645 48.850 ;
        RECT 119.125 46.950 119.525 47.750 ;
        RECT 121.765 46.950 122.165 47.750 ;
        RECT 119.125 42.750 119.525 43.550 ;
        RECT 121.765 43.300 122.165 43.550 ;
        RECT 122.645 43.300 123.145 48.850 ;
        RECT 121.765 43.000 123.145 43.300 ;
        RECT 121.765 42.750 122.165 43.000 ;
        RECT 119.125 38.550 119.525 39.350 ;
        RECT 121.765 39.100 122.165 39.350 ;
        RECT 122.645 39.100 123.145 43.000 ;
        RECT 121.765 38.800 123.145 39.100 ;
        RECT 121.765 38.550 122.165 38.800 ;
        RECT 119.125 34.350 119.525 35.150 ;
        RECT 121.765 34.900 122.165 35.150 ;
        RECT 122.645 34.900 123.145 38.800 ;
        RECT 121.765 34.600 123.145 34.900 ;
        RECT 121.765 34.350 122.165 34.600 ;
        RECT 119.125 30.150 119.525 30.950 ;
        RECT 121.765 30.700 122.165 30.950 ;
        RECT 122.645 30.700 123.145 34.600 ;
        RECT 121.765 30.400 123.145 30.700 ;
        RECT 121.765 30.150 122.165 30.400 ;
        RECT 119.125 25.950 119.525 26.750 ;
        RECT 121.765 26.500 122.165 26.750 ;
        RECT 122.645 26.500 123.145 30.400 ;
        RECT 121.765 26.200 123.145 26.500 ;
        RECT 121.765 25.950 122.165 26.200 ;
        RECT 119.125 21.750 119.525 22.550 ;
        RECT 121.765 22.300 122.165 22.550 ;
        RECT 122.645 22.300 123.145 26.200 ;
        RECT 121.765 22.000 123.145 22.300 ;
        RECT 121.765 21.750 122.165 22.000 ;
        RECT 119.125 17.550 119.525 18.350 ;
        RECT 121.765 18.100 122.165 18.350 ;
        RECT 122.645 18.100 123.145 22.000 ;
        RECT 121.765 17.800 123.145 18.100 ;
        RECT 121.765 17.550 122.165 17.800 ;
        RECT 119.125 13.350 119.525 14.150 ;
        RECT 121.765 13.900 122.165 14.150 ;
        RECT 122.645 13.900 123.145 17.800 ;
        RECT 121.765 13.600 123.145 13.900 ;
        RECT 121.765 13.350 122.165 13.600 ;
        RECT 119.125 9.150 119.525 9.950 ;
        RECT 121.765 9.150 122.165 9.950 ;
        RECT 115.845 5.490 116.645 5.890 ;
        RECT 122.645 5.090 123.145 13.600 ;
        RECT 124.645 8.050 125.145 48.850 ;
        RECT 125.625 46.950 126.025 47.750 ;
        RECT 128.265 46.950 128.665 47.750 ;
        RECT 125.625 42.750 126.025 43.550 ;
        RECT 128.265 43.300 128.665 43.550 ;
        RECT 129.145 43.300 129.645 48.850 ;
        RECT 128.265 43.000 129.645 43.300 ;
        RECT 128.265 42.750 128.665 43.000 ;
        RECT 125.625 38.550 126.025 39.350 ;
        RECT 128.265 39.100 128.665 39.350 ;
        RECT 129.145 39.100 129.645 43.000 ;
        RECT 128.265 38.800 129.645 39.100 ;
        RECT 128.265 38.550 128.665 38.800 ;
        RECT 125.625 34.350 126.025 35.150 ;
        RECT 128.265 34.900 128.665 35.150 ;
        RECT 129.145 34.900 129.645 38.800 ;
        RECT 128.265 34.600 129.645 34.900 ;
        RECT 128.265 34.350 128.665 34.600 ;
        RECT 125.625 30.150 126.025 30.950 ;
        RECT 128.265 30.700 128.665 30.950 ;
        RECT 129.145 30.700 129.645 34.600 ;
        RECT 128.265 30.400 129.645 30.700 ;
        RECT 128.265 30.150 128.665 30.400 ;
        RECT 125.625 25.950 126.025 26.750 ;
        RECT 128.265 26.500 128.665 26.750 ;
        RECT 129.145 26.500 129.645 30.400 ;
        RECT 128.265 26.200 129.645 26.500 ;
        RECT 128.265 25.950 128.665 26.200 ;
        RECT 125.625 21.750 126.025 22.550 ;
        RECT 128.265 22.300 128.665 22.550 ;
        RECT 129.145 22.300 129.645 26.200 ;
        RECT 128.265 22.000 129.645 22.300 ;
        RECT 128.265 21.750 128.665 22.000 ;
        RECT 125.625 17.550 126.025 18.350 ;
        RECT 128.265 18.100 128.665 18.350 ;
        RECT 129.145 18.100 129.645 22.000 ;
        RECT 128.265 17.800 129.645 18.100 ;
        RECT 128.265 17.550 128.665 17.800 ;
        RECT 125.625 13.350 126.025 14.150 ;
        RECT 128.265 13.900 128.665 14.150 ;
        RECT 129.145 13.900 129.645 17.800 ;
        RECT 128.265 13.600 129.645 13.900 ;
        RECT 128.265 13.350 128.665 13.600 ;
        RECT 125.625 9.150 126.025 9.950 ;
        RECT 128.265 9.150 128.665 9.950 ;
        RECT 122.345 4.690 123.145 5.090 ;
        RECT 129.145 2.690 129.645 13.600 ;
        RECT 131.145 8.050 131.645 48.850 ;
        RECT 132.125 46.950 132.525 47.750 ;
        RECT 134.765 46.950 135.165 47.750 ;
        RECT 132.125 42.750 132.525 43.550 ;
        RECT 134.765 43.300 135.165 43.550 ;
        RECT 135.645 43.300 136.145 48.850 ;
        RECT 134.765 43.000 136.145 43.300 ;
        RECT 134.765 42.750 135.165 43.000 ;
        RECT 132.125 38.550 132.525 39.350 ;
        RECT 134.765 39.100 135.165 39.350 ;
        RECT 135.645 39.100 136.145 43.000 ;
        RECT 134.765 38.800 136.145 39.100 ;
        RECT 134.765 38.550 135.165 38.800 ;
        RECT 132.125 34.350 132.525 35.150 ;
        RECT 134.765 34.900 135.165 35.150 ;
        RECT 135.645 34.900 136.145 38.800 ;
        RECT 134.765 34.600 136.145 34.900 ;
        RECT 134.765 34.350 135.165 34.600 ;
        RECT 132.125 30.150 132.525 30.950 ;
        RECT 134.765 30.700 135.165 30.950 ;
        RECT 135.645 30.700 136.145 34.600 ;
        RECT 134.765 30.400 136.145 30.700 ;
        RECT 134.765 30.150 135.165 30.400 ;
        RECT 132.125 25.950 132.525 26.750 ;
        RECT 134.765 26.500 135.165 26.750 ;
        RECT 135.645 26.500 136.145 30.400 ;
        RECT 134.765 26.200 136.145 26.500 ;
        RECT 134.765 25.950 135.165 26.200 ;
        RECT 132.125 21.750 132.525 22.550 ;
        RECT 134.765 22.300 135.165 22.550 ;
        RECT 135.645 22.300 136.145 26.200 ;
        RECT 134.765 22.000 136.145 22.300 ;
        RECT 134.765 21.750 135.165 22.000 ;
        RECT 132.125 17.550 132.525 18.350 ;
        RECT 134.765 18.100 135.165 18.350 ;
        RECT 135.645 18.100 136.145 22.000 ;
        RECT 134.765 17.800 136.145 18.100 ;
        RECT 134.765 17.550 135.165 17.800 ;
        RECT 132.125 13.350 132.525 14.150 ;
        RECT 134.765 13.900 135.165 14.150 ;
        RECT 135.645 13.900 136.145 17.800 ;
        RECT 134.765 13.600 136.145 13.900 ;
        RECT 134.765 13.350 135.165 13.600 ;
        RECT 132.125 9.150 132.525 9.950 ;
        RECT 134.765 9.150 135.165 9.950 ;
        RECT 135.645 3.490 136.145 13.600 ;
        RECT 137.645 8.050 138.145 48.850 ;
        RECT 138.625 46.950 139.025 47.750 ;
        RECT 141.265 46.950 141.665 47.750 ;
        RECT 138.625 42.750 139.025 43.550 ;
        RECT 141.265 43.300 141.665 43.550 ;
        RECT 142.145 43.300 142.645 48.850 ;
        RECT 141.265 43.000 142.645 43.300 ;
        RECT 141.265 42.750 141.665 43.000 ;
        RECT 138.625 38.550 139.025 39.350 ;
        RECT 141.265 39.100 141.665 39.350 ;
        RECT 142.145 39.100 142.645 43.000 ;
        RECT 141.265 38.800 142.645 39.100 ;
        RECT 141.265 38.550 141.665 38.800 ;
        RECT 138.625 34.350 139.025 35.150 ;
        RECT 141.265 34.900 141.665 35.150 ;
        RECT 142.145 34.900 142.645 38.800 ;
        RECT 141.265 34.600 142.645 34.900 ;
        RECT 141.265 34.350 141.665 34.600 ;
        RECT 138.625 30.150 139.025 30.950 ;
        RECT 141.265 30.700 141.665 30.950 ;
        RECT 142.145 30.700 142.645 34.600 ;
        RECT 141.265 30.400 142.645 30.700 ;
        RECT 141.265 30.150 141.665 30.400 ;
        RECT 138.625 25.950 139.025 26.750 ;
        RECT 141.265 26.500 141.665 26.750 ;
        RECT 142.145 26.500 142.645 30.400 ;
        RECT 141.265 26.200 142.645 26.500 ;
        RECT 141.265 25.950 141.665 26.200 ;
        RECT 138.625 21.750 139.025 22.550 ;
        RECT 141.265 22.300 141.665 22.550 ;
        RECT 142.145 22.300 142.645 26.200 ;
        RECT 141.265 22.000 142.645 22.300 ;
        RECT 141.265 21.750 141.665 22.000 ;
        RECT 138.625 17.550 139.025 18.350 ;
        RECT 141.265 18.100 141.665 18.350 ;
        RECT 142.145 18.100 142.645 22.000 ;
        RECT 141.265 17.800 142.645 18.100 ;
        RECT 141.265 17.550 141.665 17.800 ;
        RECT 138.625 13.350 139.025 14.150 ;
        RECT 141.265 13.900 141.665 14.150 ;
        RECT 142.145 13.900 142.645 17.800 ;
        RECT 141.265 13.600 142.645 13.900 ;
        RECT 141.265 13.350 141.665 13.600 ;
        RECT 138.625 9.150 139.025 9.950 ;
        RECT 141.265 9.150 141.665 9.950 ;
        RECT 142.145 4.290 142.645 13.600 ;
        RECT 144.145 8.050 144.645 48.850 ;
        RECT 145.125 46.950 145.525 47.750 ;
        RECT 147.765 46.950 148.165 47.750 ;
        RECT 145.125 42.750 145.525 43.550 ;
        RECT 147.765 43.300 148.165 43.550 ;
        RECT 148.645 43.300 149.145 48.850 ;
        RECT 147.765 43.000 149.145 43.300 ;
        RECT 147.765 42.750 148.165 43.000 ;
        RECT 145.125 38.550 145.525 39.350 ;
        RECT 147.765 39.100 148.165 39.350 ;
        RECT 148.645 39.100 149.145 43.000 ;
        RECT 147.765 38.800 149.145 39.100 ;
        RECT 147.765 38.550 148.165 38.800 ;
        RECT 145.125 34.350 145.525 35.150 ;
        RECT 147.765 34.900 148.165 35.150 ;
        RECT 148.645 34.900 149.145 38.800 ;
        RECT 147.765 34.600 149.145 34.900 ;
        RECT 147.765 34.350 148.165 34.600 ;
        RECT 145.125 30.150 145.525 30.950 ;
        RECT 147.765 30.700 148.165 30.950 ;
        RECT 148.645 30.700 149.145 34.600 ;
        RECT 147.765 30.400 149.145 30.700 ;
        RECT 147.765 30.150 148.165 30.400 ;
        RECT 145.125 25.950 145.525 26.750 ;
        RECT 147.765 26.500 148.165 26.750 ;
        RECT 148.645 26.500 149.145 30.400 ;
        RECT 147.765 26.200 149.145 26.500 ;
        RECT 147.765 25.950 148.165 26.200 ;
        RECT 145.125 21.750 145.525 22.550 ;
        RECT 147.765 22.300 148.165 22.550 ;
        RECT 148.645 22.300 149.145 26.200 ;
        RECT 147.765 22.000 149.145 22.300 ;
        RECT 147.765 21.750 148.165 22.000 ;
        RECT 145.125 17.550 145.525 18.350 ;
        RECT 147.765 18.100 148.165 18.350 ;
        RECT 148.645 18.100 149.145 22.000 ;
        RECT 147.765 17.800 149.145 18.100 ;
        RECT 147.765 17.550 148.165 17.800 ;
        RECT 145.125 13.350 145.525 14.150 ;
        RECT 147.765 13.900 148.165 14.150 ;
        RECT 148.645 13.900 149.145 17.800 ;
        RECT 147.765 13.600 149.145 13.900 ;
        RECT 147.765 13.350 148.165 13.600 ;
        RECT 145.125 9.150 145.525 9.950 ;
        RECT 147.765 9.150 148.165 9.950 ;
        RECT 141.845 3.890 142.645 4.290 ;
        RECT 135.345 3.090 136.145 3.490 ;
        RECT 148.645 2.690 149.145 13.600 ;
        RECT 150.645 8.050 151.145 48.850 ;
        RECT 151.625 46.950 152.025 47.750 ;
        RECT 154.265 46.950 154.665 47.750 ;
        RECT 151.625 42.750 152.025 43.550 ;
        RECT 154.265 43.300 154.665 43.550 ;
        RECT 155.145 43.300 155.645 48.850 ;
        RECT 154.265 43.000 155.645 43.300 ;
        RECT 154.265 42.750 154.665 43.000 ;
        RECT 151.625 38.550 152.025 39.350 ;
        RECT 154.265 39.100 154.665 39.350 ;
        RECT 155.145 39.100 155.645 43.000 ;
        RECT 154.265 38.800 155.645 39.100 ;
        RECT 154.265 38.550 154.665 38.800 ;
        RECT 151.625 34.350 152.025 35.150 ;
        RECT 154.265 34.900 154.665 35.150 ;
        RECT 155.145 34.900 155.645 38.800 ;
        RECT 154.265 34.600 155.645 34.900 ;
        RECT 154.265 34.350 154.665 34.600 ;
        RECT 151.625 30.150 152.025 30.950 ;
        RECT 154.265 30.700 154.665 30.950 ;
        RECT 155.145 30.700 155.645 34.600 ;
        RECT 154.265 30.400 155.645 30.700 ;
        RECT 154.265 30.150 154.665 30.400 ;
        RECT 151.625 25.950 152.025 26.750 ;
        RECT 154.265 26.500 154.665 26.750 ;
        RECT 155.145 26.500 155.645 30.400 ;
        RECT 154.265 26.200 155.645 26.500 ;
        RECT 154.265 25.950 154.665 26.200 ;
        RECT 151.625 21.750 152.025 22.550 ;
        RECT 154.265 22.300 154.665 22.550 ;
        RECT 155.145 22.300 155.645 26.200 ;
        RECT 154.265 22.000 155.645 22.300 ;
        RECT 154.265 21.750 154.665 22.000 ;
        RECT 151.625 17.550 152.025 18.350 ;
        RECT 154.265 18.100 154.665 18.350 ;
        RECT 155.145 18.100 155.645 22.000 ;
        RECT 154.265 17.800 155.645 18.100 ;
        RECT 154.265 17.550 154.665 17.800 ;
        RECT 151.625 13.350 152.025 14.150 ;
        RECT 154.265 13.900 154.665 14.150 ;
        RECT 155.145 13.900 155.645 17.800 ;
        RECT 154.265 13.600 155.645 13.900 ;
        RECT 154.265 13.350 154.665 13.600 ;
        RECT 151.625 9.150 152.025 9.950 ;
        RECT 154.265 9.150 154.665 9.950 ;
        RECT 155.145 2.690 155.645 13.600 ;
        RECT 157.145 8.050 157.645 48.850 ;
        RECT 158.125 46.950 158.525 47.750 ;
        RECT 160.765 46.950 161.165 47.750 ;
        RECT 158.125 42.750 158.525 43.550 ;
        RECT 160.765 43.300 161.165 43.550 ;
        RECT 161.645 43.300 162.145 48.850 ;
        RECT 160.765 43.000 162.145 43.300 ;
        RECT 160.765 42.750 161.165 43.000 ;
        RECT 158.125 38.550 158.525 39.350 ;
        RECT 160.765 39.100 161.165 39.350 ;
        RECT 161.645 39.100 162.145 43.000 ;
        RECT 160.765 38.800 162.145 39.100 ;
        RECT 160.765 38.550 161.165 38.800 ;
        RECT 158.125 34.350 158.525 35.150 ;
        RECT 160.765 34.900 161.165 35.150 ;
        RECT 161.645 34.900 162.145 38.800 ;
        RECT 160.765 34.600 162.145 34.900 ;
        RECT 160.765 34.350 161.165 34.600 ;
        RECT 158.125 30.150 158.525 30.950 ;
        RECT 160.765 30.700 161.165 30.950 ;
        RECT 161.645 30.700 162.145 34.600 ;
        RECT 160.765 30.400 162.145 30.700 ;
        RECT 160.765 30.150 161.165 30.400 ;
        RECT 158.125 25.950 158.525 26.750 ;
        RECT 160.765 26.500 161.165 26.750 ;
        RECT 161.645 26.500 162.145 30.400 ;
        RECT 160.765 26.200 162.145 26.500 ;
        RECT 160.765 25.950 161.165 26.200 ;
        RECT 158.125 21.750 158.525 22.550 ;
        RECT 160.765 22.300 161.165 22.550 ;
        RECT 161.645 22.300 162.145 26.200 ;
        RECT 160.765 22.000 162.145 22.300 ;
        RECT 160.765 21.750 161.165 22.000 ;
        RECT 158.125 17.550 158.525 18.350 ;
        RECT 160.765 18.100 161.165 18.350 ;
        RECT 161.645 18.100 162.145 22.000 ;
        RECT 160.765 17.800 162.145 18.100 ;
        RECT 160.765 17.550 161.165 17.800 ;
        RECT 158.125 13.350 158.525 14.150 ;
        RECT 160.765 13.900 161.165 14.150 ;
        RECT 161.645 13.900 162.145 17.800 ;
        RECT 160.765 13.600 162.145 13.900 ;
        RECT 160.765 13.350 161.165 13.600 ;
        RECT 158.125 9.150 158.525 9.950 ;
        RECT 160.765 9.150 161.165 9.950 ;
        RECT 161.645 3.490 162.145 13.600 ;
        RECT 163.645 8.050 164.145 48.850 ;
        RECT 164.625 46.950 165.025 47.750 ;
        RECT 167.265 46.950 167.665 47.750 ;
        RECT 164.625 42.750 165.025 43.550 ;
        RECT 167.265 43.300 167.665 43.550 ;
        RECT 168.145 43.300 168.645 48.850 ;
        RECT 167.265 43.000 168.645 43.300 ;
        RECT 167.265 42.750 167.665 43.000 ;
        RECT 164.625 38.550 165.025 39.350 ;
        RECT 167.265 39.100 167.665 39.350 ;
        RECT 168.145 39.100 168.645 43.000 ;
        RECT 167.265 38.800 168.645 39.100 ;
        RECT 167.265 38.550 167.665 38.800 ;
        RECT 164.625 34.350 165.025 35.150 ;
        RECT 167.265 34.900 167.665 35.150 ;
        RECT 168.145 34.900 168.645 38.800 ;
        RECT 167.265 34.600 168.645 34.900 ;
        RECT 167.265 34.350 167.665 34.600 ;
        RECT 164.625 30.150 165.025 30.950 ;
        RECT 167.265 30.700 167.665 30.950 ;
        RECT 168.145 30.700 168.645 34.600 ;
        RECT 167.265 30.400 168.645 30.700 ;
        RECT 167.265 30.150 167.665 30.400 ;
        RECT 164.625 25.950 165.025 26.750 ;
        RECT 167.265 26.500 167.665 26.750 ;
        RECT 168.145 26.500 168.645 30.400 ;
        RECT 167.265 26.200 168.645 26.500 ;
        RECT 167.265 25.950 167.665 26.200 ;
        RECT 164.625 21.750 165.025 22.550 ;
        RECT 167.265 22.300 167.665 22.550 ;
        RECT 168.145 22.300 168.645 26.200 ;
        RECT 167.265 22.000 168.645 22.300 ;
        RECT 167.265 21.750 167.665 22.000 ;
        RECT 164.625 17.550 165.025 18.350 ;
        RECT 167.265 18.100 167.665 18.350 ;
        RECT 168.145 18.100 168.645 22.000 ;
        RECT 167.265 17.800 168.645 18.100 ;
        RECT 167.265 17.550 167.665 17.800 ;
        RECT 164.625 13.350 165.025 14.150 ;
        RECT 167.265 13.900 167.665 14.150 ;
        RECT 168.145 13.900 168.645 17.800 ;
        RECT 167.265 13.600 168.645 13.900 ;
        RECT 167.265 13.350 167.665 13.600 ;
        RECT 164.625 9.150 165.025 9.950 ;
        RECT 167.265 9.150 167.665 9.950 ;
        RECT 168.145 4.290 168.645 13.600 ;
        RECT 170.145 8.050 170.645 48.850 ;
        RECT 171.125 46.950 171.525 47.750 ;
        RECT 173.765 46.950 174.165 47.750 ;
        RECT 171.125 42.750 171.525 43.550 ;
        RECT 173.765 43.300 174.165 43.550 ;
        RECT 174.645 43.300 175.145 48.850 ;
        RECT 173.765 43.000 175.145 43.300 ;
        RECT 173.765 42.750 174.165 43.000 ;
        RECT 171.125 38.550 171.525 39.350 ;
        RECT 173.765 39.100 174.165 39.350 ;
        RECT 174.645 39.100 175.145 43.000 ;
        RECT 173.765 38.800 175.145 39.100 ;
        RECT 173.765 38.550 174.165 38.800 ;
        RECT 171.125 34.350 171.525 35.150 ;
        RECT 173.765 34.900 174.165 35.150 ;
        RECT 174.645 34.900 175.145 38.800 ;
        RECT 173.765 34.600 175.145 34.900 ;
        RECT 173.765 34.350 174.165 34.600 ;
        RECT 171.125 30.150 171.525 30.950 ;
        RECT 173.765 30.700 174.165 30.950 ;
        RECT 174.645 30.700 175.145 34.600 ;
        RECT 173.765 30.400 175.145 30.700 ;
        RECT 173.765 30.150 174.165 30.400 ;
        RECT 171.125 25.950 171.525 26.750 ;
        RECT 173.765 26.500 174.165 26.750 ;
        RECT 174.645 26.500 175.145 30.400 ;
        RECT 173.765 26.200 175.145 26.500 ;
        RECT 173.765 25.950 174.165 26.200 ;
        RECT 171.125 21.750 171.525 22.550 ;
        RECT 173.765 22.300 174.165 22.550 ;
        RECT 174.645 22.300 175.145 26.200 ;
        RECT 173.765 22.000 175.145 22.300 ;
        RECT 173.765 21.750 174.165 22.000 ;
        RECT 171.125 17.550 171.525 18.350 ;
        RECT 173.765 18.100 174.165 18.350 ;
        RECT 174.645 18.100 175.145 22.000 ;
        RECT 173.765 17.800 175.145 18.100 ;
        RECT 173.765 17.550 174.165 17.800 ;
        RECT 171.125 13.350 171.525 14.150 ;
        RECT 173.765 13.900 174.165 14.150 ;
        RECT 174.645 13.900 175.145 17.800 ;
        RECT 173.765 13.600 175.145 13.900 ;
        RECT 173.765 13.350 174.165 13.600 ;
        RECT 171.125 9.150 171.525 9.950 ;
        RECT 173.765 9.150 174.165 9.950 ;
        RECT 167.845 3.890 168.645 4.290 ;
        RECT 161.345 3.090 162.145 3.490 ;
        RECT 174.645 2.690 175.145 13.600 ;
        RECT 176.645 8.050 177.145 48.850 ;
        RECT 177.625 46.950 178.025 47.750 ;
        RECT 180.265 46.950 180.665 47.750 ;
        RECT 177.625 42.750 178.025 43.550 ;
        RECT 180.265 43.300 180.665 43.550 ;
        RECT 181.145 43.300 181.645 48.850 ;
        RECT 180.265 43.000 181.645 43.300 ;
        RECT 180.265 42.750 180.665 43.000 ;
        RECT 177.625 38.550 178.025 39.350 ;
        RECT 180.265 39.100 180.665 39.350 ;
        RECT 181.145 39.100 181.645 43.000 ;
        RECT 180.265 38.800 181.645 39.100 ;
        RECT 180.265 38.550 180.665 38.800 ;
        RECT 177.625 34.350 178.025 35.150 ;
        RECT 180.265 34.900 180.665 35.150 ;
        RECT 181.145 34.900 181.645 38.800 ;
        RECT 180.265 34.600 181.645 34.900 ;
        RECT 180.265 34.350 180.665 34.600 ;
        RECT 177.625 30.150 178.025 30.950 ;
        RECT 180.265 30.700 180.665 30.950 ;
        RECT 181.145 30.700 181.645 34.600 ;
        RECT 180.265 30.400 181.645 30.700 ;
        RECT 180.265 30.150 180.665 30.400 ;
        RECT 177.625 25.950 178.025 26.750 ;
        RECT 180.265 26.500 180.665 26.750 ;
        RECT 181.145 26.500 181.645 30.400 ;
        RECT 180.265 26.200 181.645 26.500 ;
        RECT 180.265 25.950 180.665 26.200 ;
        RECT 177.625 21.750 178.025 22.550 ;
        RECT 180.265 22.300 180.665 22.550 ;
        RECT 181.145 22.300 181.645 26.200 ;
        RECT 180.265 22.000 181.645 22.300 ;
        RECT 180.265 21.750 180.665 22.000 ;
        RECT 177.625 17.550 178.025 18.350 ;
        RECT 180.265 18.100 180.665 18.350 ;
        RECT 181.145 18.100 181.645 22.000 ;
        RECT 180.265 17.800 181.645 18.100 ;
        RECT 180.265 17.550 180.665 17.800 ;
        RECT 177.625 13.350 178.025 14.150 ;
        RECT 180.265 13.900 180.665 14.150 ;
        RECT 181.145 13.900 181.645 17.800 ;
        RECT 180.265 13.600 181.645 13.900 ;
        RECT 180.265 13.350 180.665 13.600 ;
        RECT 177.625 9.150 178.025 9.950 ;
        RECT 180.265 9.150 180.665 9.950 ;
        RECT 181.145 2.690 181.645 13.600 ;
        RECT 183.145 8.050 183.645 48.850 ;
        RECT 184.125 46.950 184.525 47.750 ;
        RECT 186.765 46.950 187.165 47.750 ;
        RECT 184.125 42.750 184.525 43.550 ;
        RECT 186.765 43.300 187.165 43.550 ;
        RECT 187.645 43.300 188.145 48.850 ;
        RECT 186.765 43.000 188.145 43.300 ;
        RECT 186.765 42.750 187.165 43.000 ;
        RECT 184.125 38.550 184.525 39.350 ;
        RECT 186.765 39.100 187.165 39.350 ;
        RECT 187.645 39.100 188.145 43.000 ;
        RECT 186.765 38.800 188.145 39.100 ;
        RECT 186.765 38.550 187.165 38.800 ;
        RECT 184.125 34.350 184.525 35.150 ;
        RECT 186.765 34.900 187.165 35.150 ;
        RECT 187.645 34.900 188.145 38.800 ;
        RECT 186.765 34.600 188.145 34.900 ;
        RECT 186.765 34.350 187.165 34.600 ;
        RECT 184.125 30.150 184.525 30.950 ;
        RECT 186.765 30.700 187.165 30.950 ;
        RECT 187.645 30.700 188.145 34.600 ;
        RECT 186.765 30.400 188.145 30.700 ;
        RECT 186.765 30.150 187.165 30.400 ;
        RECT 184.125 25.950 184.525 26.750 ;
        RECT 186.765 26.500 187.165 26.750 ;
        RECT 187.645 26.500 188.145 30.400 ;
        RECT 186.765 26.200 188.145 26.500 ;
        RECT 186.765 25.950 187.165 26.200 ;
        RECT 184.125 21.750 184.525 22.550 ;
        RECT 186.765 22.300 187.165 22.550 ;
        RECT 187.645 22.300 188.145 26.200 ;
        RECT 186.765 22.000 188.145 22.300 ;
        RECT 186.765 21.750 187.165 22.000 ;
        RECT 184.125 17.550 184.525 18.350 ;
        RECT 186.765 18.100 187.165 18.350 ;
        RECT 187.645 18.100 188.145 22.000 ;
        RECT 186.765 17.800 188.145 18.100 ;
        RECT 186.765 17.550 187.165 17.800 ;
        RECT 184.125 13.350 184.525 14.150 ;
        RECT 186.765 13.900 187.165 14.150 ;
        RECT 187.645 13.900 188.145 17.800 ;
        RECT 186.765 13.600 188.145 13.900 ;
        RECT 186.765 13.350 187.165 13.600 ;
        RECT 184.125 9.150 184.525 9.950 ;
        RECT 186.765 9.150 187.165 9.950 ;
        RECT 187.645 3.490 188.145 13.600 ;
        RECT 189.645 8.050 190.145 48.850 ;
        RECT 190.625 46.950 191.025 47.750 ;
        RECT 193.265 46.950 193.665 47.750 ;
        RECT 190.625 42.750 191.025 43.550 ;
        RECT 193.265 43.300 193.665 43.550 ;
        RECT 194.145 43.300 194.645 48.850 ;
        RECT 193.265 43.000 194.645 43.300 ;
        RECT 193.265 42.750 193.665 43.000 ;
        RECT 190.625 38.550 191.025 39.350 ;
        RECT 193.265 39.100 193.665 39.350 ;
        RECT 194.145 39.100 194.645 43.000 ;
        RECT 193.265 38.800 194.645 39.100 ;
        RECT 193.265 38.550 193.665 38.800 ;
        RECT 190.625 34.350 191.025 35.150 ;
        RECT 193.265 34.900 193.665 35.150 ;
        RECT 194.145 34.900 194.645 38.800 ;
        RECT 193.265 34.600 194.645 34.900 ;
        RECT 193.265 34.350 193.665 34.600 ;
        RECT 190.625 30.150 191.025 30.950 ;
        RECT 193.265 30.700 193.665 30.950 ;
        RECT 194.145 30.700 194.645 34.600 ;
        RECT 193.265 30.400 194.645 30.700 ;
        RECT 193.265 30.150 193.665 30.400 ;
        RECT 190.625 25.950 191.025 26.750 ;
        RECT 193.265 26.500 193.665 26.750 ;
        RECT 194.145 26.500 194.645 30.400 ;
        RECT 193.265 26.200 194.645 26.500 ;
        RECT 193.265 25.950 193.665 26.200 ;
        RECT 190.625 21.750 191.025 22.550 ;
        RECT 193.265 22.300 193.665 22.550 ;
        RECT 194.145 22.300 194.645 26.200 ;
        RECT 193.265 22.000 194.645 22.300 ;
        RECT 193.265 21.750 193.665 22.000 ;
        RECT 190.625 17.550 191.025 18.350 ;
        RECT 193.265 18.100 193.665 18.350 ;
        RECT 194.145 18.100 194.645 22.000 ;
        RECT 193.265 17.800 194.645 18.100 ;
        RECT 193.265 17.550 193.665 17.800 ;
        RECT 190.625 13.350 191.025 14.150 ;
        RECT 193.265 13.900 193.665 14.150 ;
        RECT 194.145 13.900 194.645 17.800 ;
        RECT 193.265 13.600 194.645 13.900 ;
        RECT 193.265 13.350 193.665 13.600 ;
        RECT 190.625 9.150 191.025 9.950 ;
        RECT 193.265 9.150 193.665 9.950 ;
        RECT 187.345 3.090 188.145 3.490 ;
        RECT 194.145 2.690 194.645 13.600 ;
        RECT 196.145 8.050 196.645 48.850 ;
        RECT 197.125 46.950 197.525 47.750 ;
        RECT 199.765 46.950 200.165 47.750 ;
        RECT 197.125 42.750 197.525 43.550 ;
        RECT 199.765 43.300 200.165 43.550 ;
        RECT 200.645 43.300 201.145 48.850 ;
        RECT 199.765 43.000 201.145 43.300 ;
        RECT 199.765 42.750 200.165 43.000 ;
        RECT 197.125 38.550 197.525 39.350 ;
        RECT 199.765 39.100 200.165 39.350 ;
        RECT 200.645 39.100 201.145 43.000 ;
        RECT 199.765 38.800 201.145 39.100 ;
        RECT 199.765 38.550 200.165 38.800 ;
        RECT 197.125 34.350 197.525 35.150 ;
        RECT 199.765 34.900 200.165 35.150 ;
        RECT 200.645 34.900 201.145 38.800 ;
        RECT 199.765 34.600 201.145 34.900 ;
        RECT 199.765 34.350 200.165 34.600 ;
        RECT 197.125 30.150 197.525 30.950 ;
        RECT 199.765 30.700 200.165 30.950 ;
        RECT 200.645 30.700 201.145 34.600 ;
        RECT 199.765 30.400 201.145 30.700 ;
        RECT 199.765 30.150 200.165 30.400 ;
        RECT 197.125 25.950 197.525 26.750 ;
        RECT 199.765 26.500 200.165 26.750 ;
        RECT 200.645 26.500 201.145 30.400 ;
        RECT 199.765 26.200 201.145 26.500 ;
        RECT 199.765 25.950 200.165 26.200 ;
        RECT 197.125 21.750 197.525 22.550 ;
        RECT 199.765 22.300 200.165 22.550 ;
        RECT 200.645 22.300 201.145 26.200 ;
        RECT 199.765 22.000 201.145 22.300 ;
        RECT 199.765 21.750 200.165 22.000 ;
        RECT 197.125 17.550 197.525 18.350 ;
        RECT 199.765 18.100 200.165 18.350 ;
        RECT 200.645 18.100 201.145 22.000 ;
        RECT 199.765 17.800 201.145 18.100 ;
        RECT 199.765 17.550 200.165 17.800 ;
        RECT 197.125 13.350 197.525 14.150 ;
        RECT 199.765 13.900 200.165 14.150 ;
        RECT 200.645 13.900 201.145 17.800 ;
        RECT 199.765 13.600 201.145 13.900 ;
        RECT 199.765 13.350 200.165 13.600 ;
        RECT 197.125 9.150 197.525 9.950 ;
        RECT 199.765 9.150 200.165 9.950 ;
        RECT 200.645 2.690 201.145 13.600 ;
        RECT 202.645 8.050 203.145 48.850 ;
        RECT 203.625 46.950 204.025 47.750 ;
        RECT 206.265 46.950 206.665 47.750 ;
        RECT 203.625 42.750 204.025 43.550 ;
        RECT 206.265 43.300 206.665 43.550 ;
        RECT 207.145 43.300 207.645 48.850 ;
        RECT 206.265 43.000 207.645 43.300 ;
        RECT 206.265 42.750 206.665 43.000 ;
        RECT 203.625 38.550 204.025 39.350 ;
        RECT 206.265 39.100 206.665 39.350 ;
        RECT 207.145 39.100 207.645 43.000 ;
        RECT 206.265 38.800 207.645 39.100 ;
        RECT 206.265 38.550 206.665 38.800 ;
        RECT 203.625 34.350 204.025 35.150 ;
        RECT 206.265 34.900 206.665 35.150 ;
        RECT 207.145 34.900 207.645 38.800 ;
        RECT 206.265 34.600 207.645 34.900 ;
        RECT 206.265 34.350 206.665 34.600 ;
        RECT 203.625 30.150 204.025 30.950 ;
        RECT 206.265 30.700 206.665 30.950 ;
        RECT 207.145 30.700 207.645 34.600 ;
        RECT 206.265 30.400 207.645 30.700 ;
        RECT 206.265 30.150 206.665 30.400 ;
        RECT 203.625 25.950 204.025 26.750 ;
        RECT 206.265 26.500 206.665 26.750 ;
        RECT 207.145 26.500 207.645 30.400 ;
        RECT 206.265 26.200 207.645 26.500 ;
        RECT 206.265 25.950 206.665 26.200 ;
        RECT 203.625 21.750 204.025 22.550 ;
        RECT 206.265 22.300 206.665 22.550 ;
        RECT 207.145 22.300 207.645 26.200 ;
        RECT 206.265 22.000 207.645 22.300 ;
        RECT 206.265 21.750 206.665 22.000 ;
        RECT 203.625 17.550 204.025 18.350 ;
        RECT 206.265 18.100 206.665 18.350 ;
        RECT 207.145 18.100 207.645 22.000 ;
        RECT 206.265 17.800 207.645 18.100 ;
        RECT 206.265 17.550 206.665 17.800 ;
        RECT 203.625 13.350 204.025 14.150 ;
        RECT 206.265 13.900 206.665 14.150 ;
        RECT 207.145 13.900 207.645 17.800 ;
        RECT 206.265 13.600 207.645 13.900 ;
        RECT 206.265 13.350 206.665 13.600 ;
        RECT 203.625 9.150 204.025 9.950 ;
        RECT 206.265 9.150 206.665 9.950 ;
        RECT 207.145 3.490 207.645 13.600 ;
        RECT 209.145 8.050 209.645 48.850 ;
        RECT 210.125 46.950 210.525 47.750 ;
        RECT 212.765 46.950 213.165 47.750 ;
        RECT 210.125 42.750 210.525 43.550 ;
        RECT 212.765 43.300 213.165 43.550 ;
        RECT 213.645 43.300 214.145 48.850 ;
        RECT 212.765 43.000 214.145 43.300 ;
        RECT 212.765 42.750 213.165 43.000 ;
        RECT 210.125 38.550 210.525 39.350 ;
        RECT 212.765 39.100 213.165 39.350 ;
        RECT 213.645 39.100 214.145 43.000 ;
        RECT 212.765 38.800 214.145 39.100 ;
        RECT 212.765 38.550 213.165 38.800 ;
        RECT 210.125 34.350 210.525 35.150 ;
        RECT 212.765 34.900 213.165 35.150 ;
        RECT 213.645 34.900 214.145 38.800 ;
        RECT 212.765 34.600 214.145 34.900 ;
        RECT 212.765 34.350 213.165 34.600 ;
        RECT 210.125 30.150 210.525 30.950 ;
        RECT 212.765 30.700 213.165 30.950 ;
        RECT 213.645 30.700 214.145 34.600 ;
        RECT 212.765 30.400 214.145 30.700 ;
        RECT 212.765 30.150 213.165 30.400 ;
        RECT 210.125 25.950 210.525 26.750 ;
        RECT 212.765 26.500 213.165 26.750 ;
        RECT 213.645 26.500 214.145 30.400 ;
        RECT 212.765 26.200 214.145 26.500 ;
        RECT 212.765 25.950 213.165 26.200 ;
        RECT 210.125 21.750 210.525 22.550 ;
        RECT 212.765 22.300 213.165 22.550 ;
        RECT 213.645 22.300 214.145 26.200 ;
        RECT 212.765 22.000 214.145 22.300 ;
        RECT 212.765 21.750 213.165 22.000 ;
        RECT 210.125 17.550 210.525 18.350 ;
        RECT 212.765 18.100 213.165 18.350 ;
        RECT 213.645 18.100 214.145 22.000 ;
        RECT 212.765 17.800 214.145 18.100 ;
        RECT 212.765 17.550 213.165 17.800 ;
        RECT 210.125 13.350 210.525 14.150 ;
        RECT 212.765 13.900 213.165 14.150 ;
        RECT 213.645 13.900 214.145 17.800 ;
        RECT 212.765 13.600 214.145 13.900 ;
        RECT 212.765 13.350 213.165 13.600 ;
        RECT 210.125 9.150 210.525 9.950 ;
        RECT 212.765 9.150 213.165 9.950 ;
        RECT 206.845 3.090 207.645 3.490 ;
        RECT 213.645 2.690 214.145 13.600 ;
        RECT 215.645 8.050 216.145 48.850 ;
        RECT 216.625 46.950 217.025 47.750 ;
        RECT 219.265 46.950 219.665 47.750 ;
        RECT 216.625 42.750 217.025 43.550 ;
        RECT 219.265 42.750 219.665 43.550 ;
        RECT 216.625 38.550 217.025 39.350 ;
        RECT 219.265 38.550 219.665 39.350 ;
        RECT 223.205 38.940 223.805 38.990 ;
        RECT 223.205 38.640 229.670 38.940 ;
        RECT 223.205 38.590 223.805 38.640 ;
        RECT 229.370 35.570 229.670 38.640 ;
        RECT 231.115 37.870 231.375 37.880 ;
        RECT 231.115 37.570 232.215 37.870 ;
        RECT 231.115 37.560 231.375 37.570 ;
        RECT 231.115 35.570 231.375 35.580 ;
        RECT 229.370 35.270 231.410 35.570 ;
        RECT 231.115 35.260 231.375 35.270 ;
        RECT 216.625 34.350 217.025 35.150 ;
        RECT 219.265 34.350 219.665 35.150 ;
        RECT 228.560 34.730 228.960 34.880 ;
        RECT 231.915 34.730 232.215 37.570 ;
        RECT 228.560 34.430 232.215 34.730 ;
        RECT 228.560 34.280 228.960 34.430 ;
        RECT 216.625 30.150 217.025 30.950 ;
        RECT 219.265 30.150 219.665 30.950 ;
        RECT 216.625 25.950 217.025 26.750 ;
        RECT 219.265 25.950 219.665 26.750 ;
        RECT 216.625 21.750 217.025 22.550 ;
        RECT 219.265 21.750 219.665 22.550 ;
        RECT 216.625 17.550 217.025 18.350 ;
        RECT 219.265 17.550 219.665 18.350 ;
        RECT 223.205 17.780 223.805 17.830 ;
        RECT 223.205 17.480 229.670 17.780 ;
        RECT 223.205 17.430 223.805 17.480 ;
        RECT 229.370 14.410 229.670 17.480 ;
        RECT 231.115 16.710 231.375 16.720 ;
        RECT 231.115 16.410 232.215 16.710 ;
        RECT 231.115 16.400 231.375 16.410 ;
        RECT 231.115 14.410 231.375 14.420 ;
        RECT 216.625 13.350 217.025 14.150 ;
        RECT 219.265 13.350 219.665 14.150 ;
        RECT 229.370 14.110 231.410 14.410 ;
        RECT 231.115 14.100 231.375 14.110 ;
        RECT 228.560 13.570 228.960 13.720 ;
        RECT 231.915 13.570 232.215 16.410 ;
        RECT 228.560 13.270 232.215 13.570 ;
        RECT 228.560 13.120 228.960 13.270 ;
        RECT 216.625 9.150 217.025 9.950 ;
        RECT 219.265 9.150 219.665 9.950 ;
        RECT 128.845 2.290 129.645 2.690 ;
        RECT 148.345 2.290 149.145 2.690 ;
        RECT 154.845 2.290 155.645 2.690 ;
        RECT 174.345 2.290 175.145 2.690 ;
        RECT 180.845 2.290 181.645 2.690 ;
        RECT 193.845 2.290 194.645 2.690 ;
        RECT 200.345 2.290 201.145 2.690 ;
        RECT 213.345 2.290 214.145 2.690 ;
        RECT 112.845 -0.110 113.645 0.290 ;
      LAYER via2 ;
        RECT 2.185 47.410 2.465 47.690 ;
        RECT 2.185 47.010 2.465 47.290 ;
        RECT 4.825 47.410 5.105 47.690 ;
        RECT 4.825 47.010 5.105 47.290 ;
        RECT 2.185 43.210 2.465 43.490 ;
        RECT 2.185 42.810 2.465 43.090 ;
        RECT 4.825 43.210 5.105 43.490 ;
        RECT 4.825 42.810 5.105 43.090 ;
        RECT 2.185 39.010 2.465 39.290 ;
        RECT 2.185 38.610 2.465 38.890 ;
        RECT 4.825 39.010 5.105 39.290 ;
        RECT 4.825 38.610 5.105 38.890 ;
        RECT 2.185 34.810 2.465 35.090 ;
        RECT 2.185 34.410 2.465 34.690 ;
        RECT 4.825 34.810 5.105 35.090 ;
        RECT 4.825 34.410 5.105 34.690 ;
        RECT 2.185 30.610 2.465 30.890 ;
        RECT 2.185 30.210 2.465 30.490 ;
        RECT 4.825 30.610 5.105 30.890 ;
        RECT 4.825 30.210 5.105 30.490 ;
        RECT 2.185 26.410 2.465 26.690 ;
        RECT 2.185 26.010 2.465 26.290 ;
        RECT 4.825 26.410 5.105 26.690 ;
        RECT 4.825 26.010 5.105 26.290 ;
        RECT 2.185 22.210 2.465 22.490 ;
        RECT 2.185 21.810 2.465 22.090 ;
        RECT 4.825 22.210 5.105 22.490 ;
        RECT 4.825 21.810 5.105 22.090 ;
        RECT 2.185 18.010 2.465 18.290 ;
        RECT 2.185 17.610 2.465 17.890 ;
        RECT 4.825 18.010 5.105 18.290 ;
        RECT 4.825 17.610 5.105 17.890 ;
        RECT -7.990 13.680 -7.710 13.960 ;
        RECT -7.590 13.680 -7.310 13.960 ;
        RECT 2.185 13.810 2.465 14.090 ;
        RECT 2.185 13.410 2.465 13.690 ;
        RECT 4.825 13.810 5.105 14.090 ;
        RECT 4.825 13.410 5.105 13.690 ;
        RECT -7.990 12.300 -7.710 12.580 ;
        RECT -7.590 12.300 -7.310 12.580 ;
        RECT -7.990 10.920 -7.710 11.200 ;
        RECT -7.590 10.920 -7.310 11.200 ;
        RECT -7.990 9.540 -7.710 9.820 ;
        RECT -7.590 9.540 -7.310 9.820 ;
        RECT 2.185 9.610 2.465 9.890 ;
        RECT 2.185 9.210 2.465 9.490 ;
        RECT 4.825 9.610 5.105 9.890 ;
        RECT 4.825 9.210 5.105 9.490 ;
        RECT -7.990 8.160 -7.710 8.440 ;
        RECT -7.590 8.160 -7.310 8.440 ;
        RECT 8.685 47.410 8.965 47.690 ;
        RECT 8.685 47.010 8.965 47.290 ;
        RECT 11.325 47.410 11.605 47.690 ;
        RECT 11.325 47.010 11.605 47.290 ;
        RECT 8.685 43.210 8.965 43.490 ;
        RECT 8.685 42.810 8.965 43.090 ;
        RECT 11.325 43.210 11.605 43.490 ;
        RECT 11.325 42.810 11.605 43.090 ;
        RECT 8.685 39.010 8.965 39.290 ;
        RECT 8.685 38.610 8.965 38.890 ;
        RECT 11.325 39.010 11.605 39.290 ;
        RECT 11.325 38.610 11.605 38.890 ;
        RECT 8.685 34.810 8.965 35.090 ;
        RECT 8.685 34.410 8.965 34.690 ;
        RECT 11.325 34.810 11.605 35.090 ;
        RECT 11.325 34.410 11.605 34.690 ;
        RECT 8.685 30.610 8.965 30.890 ;
        RECT 8.685 30.210 8.965 30.490 ;
        RECT 11.325 30.610 11.605 30.890 ;
        RECT 11.325 30.210 11.605 30.490 ;
        RECT 8.685 26.410 8.965 26.690 ;
        RECT 8.685 26.010 8.965 26.290 ;
        RECT 11.325 26.410 11.605 26.690 ;
        RECT 11.325 26.010 11.605 26.290 ;
        RECT 8.685 22.210 8.965 22.490 ;
        RECT 8.685 21.810 8.965 22.090 ;
        RECT 11.325 22.210 11.605 22.490 ;
        RECT 11.325 21.810 11.605 22.090 ;
        RECT 8.685 18.010 8.965 18.290 ;
        RECT 8.685 17.610 8.965 17.890 ;
        RECT 11.325 18.010 11.605 18.290 ;
        RECT 11.325 17.610 11.605 17.890 ;
        RECT 8.685 13.810 8.965 14.090 ;
        RECT -7.990 6.780 -7.710 7.060 ;
        RECT -7.590 6.780 -7.310 7.060 ;
        RECT -7.990 5.400 -7.710 5.680 ;
        RECT -7.590 5.400 -7.310 5.680 ;
        RECT -7.990 4.020 -7.710 4.300 ;
        RECT -7.590 4.020 -7.310 4.300 ;
        RECT -7.990 2.640 -7.710 2.920 ;
        RECT -7.590 2.640 -7.310 2.920 ;
        RECT 8.685 13.410 8.965 13.690 ;
        RECT 11.325 13.810 11.605 14.090 ;
        RECT 11.325 13.410 11.605 13.690 ;
        RECT 8.685 9.610 8.965 9.890 ;
        RECT 8.685 9.210 8.965 9.490 ;
        RECT 11.325 9.610 11.605 9.890 ;
        RECT 11.325 9.210 11.605 9.490 ;
        RECT 15.185 47.410 15.465 47.690 ;
        RECT 15.185 47.010 15.465 47.290 ;
        RECT 17.825 47.410 18.105 47.690 ;
        RECT 17.825 47.010 18.105 47.290 ;
        RECT 15.185 43.210 15.465 43.490 ;
        RECT 15.185 42.810 15.465 43.090 ;
        RECT 17.825 43.210 18.105 43.490 ;
        RECT 17.825 42.810 18.105 43.090 ;
        RECT 15.185 39.010 15.465 39.290 ;
        RECT 15.185 38.610 15.465 38.890 ;
        RECT 17.825 39.010 18.105 39.290 ;
        RECT 17.825 38.610 18.105 38.890 ;
        RECT 15.185 34.810 15.465 35.090 ;
        RECT 15.185 34.410 15.465 34.690 ;
        RECT 17.825 34.810 18.105 35.090 ;
        RECT 17.825 34.410 18.105 34.690 ;
        RECT 15.185 30.610 15.465 30.890 ;
        RECT 15.185 30.210 15.465 30.490 ;
        RECT 17.825 30.610 18.105 30.890 ;
        RECT 17.825 30.210 18.105 30.490 ;
        RECT 15.185 26.410 15.465 26.690 ;
        RECT 15.185 26.010 15.465 26.290 ;
        RECT 17.825 26.410 18.105 26.690 ;
        RECT 17.825 26.010 18.105 26.290 ;
        RECT 15.185 22.210 15.465 22.490 ;
        RECT 15.185 21.810 15.465 22.090 ;
        RECT 17.825 22.210 18.105 22.490 ;
        RECT 17.825 21.810 18.105 22.090 ;
        RECT 15.185 18.010 15.465 18.290 ;
        RECT 15.185 17.610 15.465 17.890 ;
        RECT 17.825 18.010 18.105 18.290 ;
        RECT 17.825 17.610 18.105 17.890 ;
        RECT 15.185 13.810 15.465 14.090 ;
        RECT 15.185 13.410 15.465 13.690 ;
        RECT 17.825 13.810 18.105 14.090 ;
        RECT 17.825 13.410 18.105 13.690 ;
        RECT 15.185 9.610 15.465 9.890 ;
        RECT 15.185 9.210 15.465 9.490 ;
        RECT 17.825 9.610 18.105 9.890 ;
        RECT 17.825 9.210 18.105 9.490 ;
        RECT 21.685 47.410 21.965 47.690 ;
        RECT 21.685 47.010 21.965 47.290 ;
        RECT 24.325 47.410 24.605 47.690 ;
        RECT 24.325 47.010 24.605 47.290 ;
        RECT 21.685 43.210 21.965 43.490 ;
        RECT 21.685 42.810 21.965 43.090 ;
        RECT 24.325 43.210 24.605 43.490 ;
        RECT 24.325 42.810 24.605 43.090 ;
        RECT 21.685 39.010 21.965 39.290 ;
        RECT 21.685 38.610 21.965 38.890 ;
        RECT 24.325 39.010 24.605 39.290 ;
        RECT 24.325 38.610 24.605 38.890 ;
        RECT 21.685 34.810 21.965 35.090 ;
        RECT 21.685 34.410 21.965 34.690 ;
        RECT 24.325 34.810 24.605 35.090 ;
        RECT 24.325 34.410 24.605 34.690 ;
        RECT 21.685 30.610 21.965 30.890 ;
        RECT 21.685 30.210 21.965 30.490 ;
        RECT 24.325 30.610 24.605 30.890 ;
        RECT 24.325 30.210 24.605 30.490 ;
        RECT 21.685 26.410 21.965 26.690 ;
        RECT 21.685 26.010 21.965 26.290 ;
        RECT 24.325 26.410 24.605 26.690 ;
        RECT 24.325 26.010 24.605 26.290 ;
        RECT 21.685 22.210 21.965 22.490 ;
        RECT 21.685 21.810 21.965 22.090 ;
        RECT 24.325 22.210 24.605 22.490 ;
        RECT 24.325 21.810 24.605 22.090 ;
        RECT 21.685 18.010 21.965 18.290 ;
        RECT 21.685 17.610 21.965 17.890 ;
        RECT 24.325 18.010 24.605 18.290 ;
        RECT 24.325 17.610 24.605 17.890 ;
        RECT 21.685 13.810 21.965 14.090 ;
        RECT 14.205 3.150 14.485 3.430 ;
        RECT 14.605 3.150 14.885 3.430 ;
        RECT 21.685 13.410 21.965 13.690 ;
        RECT 24.325 13.810 24.605 14.090 ;
        RECT 24.325 13.410 24.605 13.690 ;
        RECT 21.685 9.610 21.965 9.890 ;
        RECT 21.685 9.210 21.965 9.490 ;
        RECT 24.325 9.610 24.605 9.890 ;
        RECT 24.325 9.210 24.605 9.490 ;
        RECT 28.185 47.410 28.465 47.690 ;
        RECT 28.185 47.010 28.465 47.290 ;
        RECT 30.825 47.410 31.105 47.690 ;
        RECT 30.825 47.010 31.105 47.290 ;
        RECT 28.185 43.210 28.465 43.490 ;
        RECT 28.185 42.810 28.465 43.090 ;
        RECT 30.825 43.210 31.105 43.490 ;
        RECT 30.825 42.810 31.105 43.090 ;
        RECT 28.185 39.010 28.465 39.290 ;
        RECT 28.185 38.610 28.465 38.890 ;
        RECT 30.825 39.010 31.105 39.290 ;
        RECT 30.825 38.610 31.105 38.890 ;
        RECT 28.185 34.810 28.465 35.090 ;
        RECT 28.185 34.410 28.465 34.690 ;
        RECT 30.825 34.810 31.105 35.090 ;
        RECT 30.825 34.410 31.105 34.690 ;
        RECT 28.185 30.610 28.465 30.890 ;
        RECT 28.185 30.210 28.465 30.490 ;
        RECT 30.825 30.610 31.105 30.890 ;
        RECT 30.825 30.210 31.105 30.490 ;
        RECT 28.185 26.410 28.465 26.690 ;
        RECT 28.185 26.010 28.465 26.290 ;
        RECT 30.825 26.410 31.105 26.690 ;
        RECT 30.825 26.010 31.105 26.290 ;
        RECT 28.185 22.210 28.465 22.490 ;
        RECT 28.185 21.810 28.465 22.090 ;
        RECT 30.825 22.210 31.105 22.490 ;
        RECT 30.825 21.810 31.105 22.090 ;
        RECT 28.185 18.010 28.465 18.290 ;
        RECT 28.185 17.610 28.465 17.890 ;
        RECT 30.825 18.010 31.105 18.290 ;
        RECT 30.825 17.610 31.105 17.890 ;
        RECT 28.185 13.810 28.465 14.090 ;
        RECT 28.185 13.410 28.465 13.690 ;
        RECT 30.825 13.810 31.105 14.090 ;
        RECT 30.825 13.410 31.105 13.690 ;
        RECT 28.185 9.610 28.465 9.890 ;
        RECT 28.185 9.210 28.465 9.490 ;
        RECT 30.825 9.610 31.105 9.890 ;
        RECT 30.825 9.210 31.105 9.490 ;
        RECT 34.685 47.410 34.965 47.690 ;
        RECT 34.685 47.010 34.965 47.290 ;
        RECT 37.325 47.410 37.605 47.690 ;
        RECT 37.325 47.010 37.605 47.290 ;
        RECT 34.685 43.210 34.965 43.490 ;
        RECT 34.685 42.810 34.965 43.090 ;
        RECT 37.325 43.210 37.605 43.490 ;
        RECT 37.325 42.810 37.605 43.090 ;
        RECT 34.685 39.010 34.965 39.290 ;
        RECT 34.685 38.610 34.965 38.890 ;
        RECT 37.325 39.010 37.605 39.290 ;
        RECT 37.325 38.610 37.605 38.890 ;
        RECT 34.685 34.810 34.965 35.090 ;
        RECT 34.685 34.410 34.965 34.690 ;
        RECT 37.325 34.810 37.605 35.090 ;
        RECT 37.325 34.410 37.605 34.690 ;
        RECT 34.685 30.610 34.965 30.890 ;
        RECT 34.685 30.210 34.965 30.490 ;
        RECT 37.325 30.610 37.605 30.890 ;
        RECT 37.325 30.210 37.605 30.490 ;
        RECT 34.685 26.410 34.965 26.690 ;
        RECT 34.685 26.010 34.965 26.290 ;
        RECT 37.325 26.410 37.605 26.690 ;
        RECT 37.325 26.010 37.605 26.290 ;
        RECT 34.685 22.210 34.965 22.490 ;
        RECT 34.685 21.810 34.965 22.090 ;
        RECT 37.325 22.210 37.605 22.490 ;
        RECT 37.325 21.810 37.605 22.090 ;
        RECT 34.685 18.010 34.965 18.290 ;
        RECT 34.685 17.610 34.965 17.890 ;
        RECT 37.325 18.010 37.605 18.290 ;
        RECT 37.325 17.610 37.605 17.890 ;
        RECT 34.685 13.810 34.965 14.090 ;
        RECT 34.685 13.410 34.965 13.690 ;
        RECT 37.325 13.810 37.605 14.090 ;
        RECT 37.325 13.410 37.605 13.690 ;
        RECT 34.685 9.610 34.965 9.890 ;
        RECT 34.685 9.210 34.965 9.490 ;
        RECT 37.325 9.610 37.605 9.890 ;
        RECT 37.325 9.210 37.605 9.490 ;
        RECT 41.185 47.410 41.465 47.690 ;
        RECT 41.185 47.010 41.465 47.290 ;
        RECT 43.825 47.410 44.105 47.690 ;
        RECT 43.825 47.010 44.105 47.290 ;
        RECT 41.185 43.210 41.465 43.490 ;
        RECT 41.185 42.810 41.465 43.090 ;
        RECT 43.825 43.210 44.105 43.490 ;
        RECT 43.825 42.810 44.105 43.090 ;
        RECT 41.185 39.010 41.465 39.290 ;
        RECT 41.185 38.610 41.465 38.890 ;
        RECT 43.825 39.010 44.105 39.290 ;
        RECT 43.825 38.610 44.105 38.890 ;
        RECT 41.185 34.810 41.465 35.090 ;
        RECT 41.185 34.410 41.465 34.690 ;
        RECT 43.825 34.810 44.105 35.090 ;
        RECT 43.825 34.410 44.105 34.690 ;
        RECT 41.185 30.610 41.465 30.890 ;
        RECT 41.185 30.210 41.465 30.490 ;
        RECT 43.825 30.610 44.105 30.890 ;
        RECT 43.825 30.210 44.105 30.490 ;
        RECT 41.185 26.410 41.465 26.690 ;
        RECT 41.185 26.010 41.465 26.290 ;
        RECT 43.825 26.410 44.105 26.690 ;
        RECT 43.825 26.010 44.105 26.290 ;
        RECT 41.185 22.210 41.465 22.490 ;
        RECT 41.185 21.810 41.465 22.090 ;
        RECT 43.825 22.210 44.105 22.490 ;
        RECT 43.825 21.810 44.105 22.090 ;
        RECT 41.185 18.010 41.465 18.290 ;
        RECT 41.185 17.610 41.465 17.890 ;
        RECT 43.825 18.010 44.105 18.290 ;
        RECT 43.825 17.610 44.105 17.890 ;
        RECT 41.185 13.810 41.465 14.090 ;
        RECT 33.705 3.150 33.985 3.430 ;
        RECT 34.105 3.150 34.385 3.430 ;
        RECT 41.185 13.410 41.465 13.690 ;
        RECT 43.825 13.810 44.105 14.090 ;
        RECT 43.825 13.410 44.105 13.690 ;
        RECT 41.185 9.610 41.465 9.890 ;
        RECT 41.185 9.210 41.465 9.490 ;
        RECT 43.825 9.610 44.105 9.890 ;
        RECT 43.825 9.210 44.105 9.490 ;
        RECT 47.685 47.410 47.965 47.690 ;
        RECT 47.685 47.010 47.965 47.290 ;
        RECT 50.325 47.410 50.605 47.690 ;
        RECT 50.325 47.010 50.605 47.290 ;
        RECT 47.685 43.210 47.965 43.490 ;
        RECT 47.685 42.810 47.965 43.090 ;
        RECT 50.325 43.210 50.605 43.490 ;
        RECT 50.325 42.810 50.605 43.090 ;
        RECT 47.685 39.010 47.965 39.290 ;
        RECT 47.685 38.610 47.965 38.890 ;
        RECT 50.325 39.010 50.605 39.290 ;
        RECT 50.325 38.610 50.605 38.890 ;
        RECT 47.685 34.810 47.965 35.090 ;
        RECT 47.685 34.410 47.965 34.690 ;
        RECT 50.325 34.810 50.605 35.090 ;
        RECT 50.325 34.410 50.605 34.690 ;
        RECT 47.685 30.610 47.965 30.890 ;
        RECT 47.685 30.210 47.965 30.490 ;
        RECT 50.325 30.610 50.605 30.890 ;
        RECT 50.325 30.210 50.605 30.490 ;
        RECT 47.685 26.410 47.965 26.690 ;
        RECT 47.685 26.010 47.965 26.290 ;
        RECT 50.325 26.410 50.605 26.690 ;
        RECT 50.325 26.010 50.605 26.290 ;
        RECT 47.685 22.210 47.965 22.490 ;
        RECT 47.685 21.810 47.965 22.090 ;
        RECT 50.325 22.210 50.605 22.490 ;
        RECT 50.325 21.810 50.605 22.090 ;
        RECT 47.685 18.010 47.965 18.290 ;
        RECT 47.685 17.610 47.965 17.890 ;
        RECT 50.325 18.010 50.605 18.290 ;
        RECT 50.325 17.610 50.605 17.890 ;
        RECT 47.685 13.810 47.965 14.090 ;
        RECT 47.685 13.410 47.965 13.690 ;
        RECT 50.325 13.810 50.605 14.090 ;
        RECT 50.325 13.410 50.605 13.690 ;
        RECT 47.685 9.610 47.965 9.890 ;
        RECT 47.685 9.210 47.965 9.490 ;
        RECT 50.325 9.610 50.605 9.890 ;
        RECT 50.325 9.210 50.605 9.490 ;
        RECT 54.185 47.410 54.465 47.690 ;
        RECT 54.185 47.010 54.465 47.290 ;
        RECT 56.825 47.410 57.105 47.690 ;
        RECT 56.825 47.010 57.105 47.290 ;
        RECT 54.185 43.210 54.465 43.490 ;
        RECT 54.185 42.810 54.465 43.090 ;
        RECT 56.825 43.210 57.105 43.490 ;
        RECT 56.825 42.810 57.105 43.090 ;
        RECT 54.185 39.010 54.465 39.290 ;
        RECT 54.185 38.610 54.465 38.890 ;
        RECT 56.825 39.010 57.105 39.290 ;
        RECT 56.825 38.610 57.105 38.890 ;
        RECT 54.185 34.810 54.465 35.090 ;
        RECT 54.185 34.410 54.465 34.690 ;
        RECT 56.825 34.810 57.105 35.090 ;
        RECT 56.825 34.410 57.105 34.690 ;
        RECT 54.185 30.610 54.465 30.890 ;
        RECT 54.185 30.210 54.465 30.490 ;
        RECT 56.825 30.610 57.105 30.890 ;
        RECT 56.825 30.210 57.105 30.490 ;
        RECT 54.185 26.410 54.465 26.690 ;
        RECT 54.185 26.010 54.465 26.290 ;
        RECT 56.825 26.410 57.105 26.690 ;
        RECT 56.825 26.010 57.105 26.290 ;
        RECT 54.185 22.210 54.465 22.490 ;
        RECT 54.185 21.810 54.465 22.090 ;
        RECT 56.825 22.210 57.105 22.490 ;
        RECT 56.825 21.810 57.105 22.090 ;
        RECT 54.185 18.010 54.465 18.290 ;
        RECT 54.185 17.610 54.465 17.890 ;
        RECT 56.825 18.010 57.105 18.290 ;
        RECT 56.825 17.610 57.105 17.890 ;
        RECT 54.185 13.810 54.465 14.090 ;
        RECT 54.185 13.410 54.465 13.690 ;
        RECT 56.825 13.810 57.105 14.090 ;
        RECT 56.825 13.410 57.105 13.690 ;
        RECT 54.185 9.610 54.465 9.890 ;
        RECT 54.185 9.210 54.465 9.490 ;
        RECT 56.825 9.610 57.105 9.890 ;
        RECT 56.825 9.210 57.105 9.490 ;
        RECT 60.685 47.410 60.965 47.690 ;
        RECT 60.685 47.010 60.965 47.290 ;
        RECT 63.325 47.410 63.605 47.690 ;
        RECT 63.325 47.010 63.605 47.290 ;
        RECT 60.685 43.210 60.965 43.490 ;
        RECT 60.685 42.810 60.965 43.090 ;
        RECT 63.325 43.210 63.605 43.490 ;
        RECT 63.325 42.810 63.605 43.090 ;
        RECT 60.685 39.010 60.965 39.290 ;
        RECT 60.685 38.610 60.965 38.890 ;
        RECT 63.325 39.010 63.605 39.290 ;
        RECT 63.325 38.610 63.605 38.890 ;
        RECT 60.685 34.810 60.965 35.090 ;
        RECT 60.685 34.410 60.965 34.690 ;
        RECT 63.325 34.810 63.605 35.090 ;
        RECT 63.325 34.410 63.605 34.690 ;
        RECT 60.685 30.610 60.965 30.890 ;
        RECT 60.685 30.210 60.965 30.490 ;
        RECT 63.325 30.610 63.605 30.890 ;
        RECT 63.325 30.210 63.605 30.490 ;
        RECT 60.685 26.410 60.965 26.690 ;
        RECT 60.685 26.010 60.965 26.290 ;
        RECT 63.325 26.410 63.605 26.690 ;
        RECT 63.325 26.010 63.605 26.290 ;
        RECT 60.685 22.210 60.965 22.490 ;
        RECT 60.685 21.810 60.965 22.090 ;
        RECT 63.325 22.210 63.605 22.490 ;
        RECT 63.325 21.810 63.605 22.090 ;
        RECT 60.685 18.010 60.965 18.290 ;
        RECT 60.685 17.610 60.965 17.890 ;
        RECT 63.325 18.010 63.605 18.290 ;
        RECT 63.325 17.610 63.605 17.890 ;
        RECT 60.685 13.810 60.965 14.090 ;
        RECT 53.205 3.950 53.485 4.230 ;
        RECT 53.605 3.950 53.885 4.230 ;
        RECT 60.685 13.410 60.965 13.690 ;
        RECT 63.325 13.810 63.605 14.090 ;
        RECT 63.325 13.410 63.605 13.690 ;
        RECT 60.685 9.610 60.965 9.890 ;
        RECT 60.685 9.210 60.965 9.490 ;
        RECT 63.325 9.610 63.605 9.890 ;
        RECT 63.325 9.210 63.605 9.490 ;
        RECT 67.185 47.410 67.465 47.690 ;
        RECT 67.185 47.010 67.465 47.290 ;
        RECT 69.825 47.410 70.105 47.690 ;
        RECT 69.825 47.010 70.105 47.290 ;
        RECT 67.185 43.210 67.465 43.490 ;
        RECT 67.185 42.810 67.465 43.090 ;
        RECT 69.825 43.210 70.105 43.490 ;
        RECT 69.825 42.810 70.105 43.090 ;
        RECT 67.185 39.010 67.465 39.290 ;
        RECT 67.185 38.610 67.465 38.890 ;
        RECT 69.825 39.010 70.105 39.290 ;
        RECT 69.825 38.610 70.105 38.890 ;
        RECT 67.185 34.810 67.465 35.090 ;
        RECT 67.185 34.410 67.465 34.690 ;
        RECT 69.825 34.810 70.105 35.090 ;
        RECT 69.825 34.410 70.105 34.690 ;
        RECT 67.185 30.610 67.465 30.890 ;
        RECT 67.185 30.210 67.465 30.490 ;
        RECT 69.825 30.610 70.105 30.890 ;
        RECT 69.825 30.210 70.105 30.490 ;
        RECT 67.185 26.410 67.465 26.690 ;
        RECT 67.185 26.010 67.465 26.290 ;
        RECT 69.825 26.410 70.105 26.690 ;
        RECT 69.825 26.010 70.105 26.290 ;
        RECT 67.185 22.210 67.465 22.490 ;
        RECT 67.185 21.810 67.465 22.090 ;
        RECT 69.825 22.210 70.105 22.490 ;
        RECT 69.825 21.810 70.105 22.090 ;
        RECT 67.185 18.010 67.465 18.290 ;
        RECT 67.185 17.610 67.465 17.890 ;
        RECT 69.825 18.010 70.105 18.290 ;
        RECT 69.825 17.610 70.105 17.890 ;
        RECT 67.185 13.810 67.465 14.090 ;
        RECT 59.705 3.150 59.985 3.430 ;
        RECT 60.105 3.150 60.385 3.430 ;
        RECT 67.185 13.410 67.465 13.690 ;
        RECT 69.825 13.810 70.105 14.090 ;
        RECT 69.825 13.410 70.105 13.690 ;
        RECT 67.185 9.610 67.465 9.890 ;
        RECT 67.185 9.210 67.465 9.490 ;
        RECT 69.825 9.610 70.105 9.890 ;
        RECT 69.825 9.210 70.105 9.490 ;
        RECT 73.685 47.410 73.965 47.690 ;
        RECT 73.685 47.010 73.965 47.290 ;
        RECT 76.325 47.410 76.605 47.690 ;
        RECT 76.325 47.010 76.605 47.290 ;
        RECT 73.685 43.210 73.965 43.490 ;
        RECT 73.685 42.810 73.965 43.090 ;
        RECT 76.325 43.210 76.605 43.490 ;
        RECT 76.325 42.810 76.605 43.090 ;
        RECT 73.685 39.010 73.965 39.290 ;
        RECT 73.685 38.610 73.965 38.890 ;
        RECT 76.325 39.010 76.605 39.290 ;
        RECT 76.325 38.610 76.605 38.890 ;
        RECT 73.685 34.810 73.965 35.090 ;
        RECT 73.685 34.410 73.965 34.690 ;
        RECT 76.325 34.810 76.605 35.090 ;
        RECT 76.325 34.410 76.605 34.690 ;
        RECT 73.685 30.610 73.965 30.890 ;
        RECT 73.685 30.210 73.965 30.490 ;
        RECT 76.325 30.610 76.605 30.890 ;
        RECT 76.325 30.210 76.605 30.490 ;
        RECT 73.685 26.410 73.965 26.690 ;
        RECT 73.685 26.010 73.965 26.290 ;
        RECT 76.325 26.410 76.605 26.690 ;
        RECT 76.325 26.010 76.605 26.290 ;
        RECT 73.685 22.210 73.965 22.490 ;
        RECT 73.685 21.810 73.965 22.090 ;
        RECT 76.325 22.210 76.605 22.490 ;
        RECT 76.325 21.810 76.605 22.090 ;
        RECT 73.685 18.010 73.965 18.290 ;
        RECT 73.685 17.610 73.965 17.890 ;
        RECT 76.325 18.010 76.605 18.290 ;
        RECT 76.325 17.610 76.605 17.890 ;
        RECT 73.685 13.810 73.965 14.090 ;
        RECT 73.685 13.410 73.965 13.690 ;
        RECT 76.325 13.810 76.605 14.090 ;
        RECT 76.325 13.410 76.605 13.690 ;
        RECT 73.685 9.610 73.965 9.890 ;
        RECT 73.685 9.210 73.965 9.490 ;
        RECT 76.325 9.610 76.605 9.890 ;
        RECT 76.325 9.210 76.605 9.490 ;
        RECT 80.185 47.410 80.465 47.690 ;
        RECT 80.185 47.010 80.465 47.290 ;
        RECT 82.825 47.410 83.105 47.690 ;
        RECT 82.825 47.010 83.105 47.290 ;
        RECT 80.185 43.210 80.465 43.490 ;
        RECT 80.185 42.810 80.465 43.090 ;
        RECT 82.825 43.210 83.105 43.490 ;
        RECT 82.825 42.810 83.105 43.090 ;
        RECT 80.185 39.010 80.465 39.290 ;
        RECT 80.185 38.610 80.465 38.890 ;
        RECT 82.825 39.010 83.105 39.290 ;
        RECT 82.825 38.610 83.105 38.890 ;
        RECT 80.185 34.810 80.465 35.090 ;
        RECT 80.185 34.410 80.465 34.690 ;
        RECT 82.825 34.810 83.105 35.090 ;
        RECT 82.825 34.410 83.105 34.690 ;
        RECT 80.185 30.610 80.465 30.890 ;
        RECT 80.185 30.210 80.465 30.490 ;
        RECT 82.825 30.610 83.105 30.890 ;
        RECT 82.825 30.210 83.105 30.490 ;
        RECT 80.185 26.410 80.465 26.690 ;
        RECT 80.185 26.010 80.465 26.290 ;
        RECT 82.825 26.410 83.105 26.690 ;
        RECT 82.825 26.010 83.105 26.290 ;
        RECT 80.185 22.210 80.465 22.490 ;
        RECT 80.185 21.810 80.465 22.090 ;
        RECT 82.825 22.210 83.105 22.490 ;
        RECT 82.825 21.810 83.105 22.090 ;
        RECT 80.185 18.010 80.465 18.290 ;
        RECT 80.185 17.610 80.465 17.890 ;
        RECT 82.825 18.010 83.105 18.290 ;
        RECT 82.825 17.610 83.105 17.890 ;
        RECT 80.185 13.810 80.465 14.090 ;
        RECT 80.185 13.410 80.465 13.690 ;
        RECT 82.825 13.810 83.105 14.090 ;
        RECT 82.825 13.410 83.105 13.690 ;
        RECT 80.185 9.610 80.465 9.890 ;
        RECT 80.185 9.210 80.465 9.490 ;
        RECT 82.825 9.610 83.105 9.890 ;
        RECT 82.825 9.210 83.105 9.490 ;
        RECT 86.685 47.410 86.965 47.690 ;
        RECT 86.685 47.010 86.965 47.290 ;
        RECT 89.325 47.410 89.605 47.690 ;
        RECT 89.325 47.010 89.605 47.290 ;
        RECT 86.685 43.210 86.965 43.490 ;
        RECT 86.685 42.810 86.965 43.090 ;
        RECT 89.325 43.210 89.605 43.490 ;
        RECT 89.325 42.810 89.605 43.090 ;
        RECT 86.685 39.010 86.965 39.290 ;
        RECT 86.685 38.610 86.965 38.890 ;
        RECT 89.325 39.010 89.605 39.290 ;
        RECT 89.325 38.610 89.605 38.890 ;
        RECT 86.685 34.810 86.965 35.090 ;
        RECT 86.685 34.410 86.965 34.690 ;
        RECT 89.325 34.810 89.605 35.090 ;
        RECT 89.325 34.410 89.605 34.690 ;
        RECT 86.685 30.610 86.965 30.890 ;
        RECT 86.685 30.210 86.965 30.490 ;
        RECT 89.325 30.610 89.605 30.890 ;
        RECT 89.325 30.210 89.605 30.490 ;
        RECT 86.685 26.410 86.965 26.690 ;
        RECT 86.685 26.010 86.965 26.290 ;
        RECT 89.325 26.410 89.605 26.690 ;
        RECT 89.325 26.010 89.605 26.290 ;
        RECT 86.685 22.210 86.965 22.490 ;
        RECT 86.685 21.810 86.965 22.090 ;
        RECT 89.325 22.210 89.605 22.490 ;
        RECT 89.325 21.810 89.605 22.090 ;
        RECT 86.685 18.010 86.965 18.290 ;
        RECT 86.685 17.610 86.965 17.890 ;
        RECT 89.325 18.010 89.605 18.290 ;
        RECT 89.325 17.610 89.605 17.890 ;
        RECT 86.685 13.810 86.965 14.090 ;
        RECT 79.205 3.950 79.485 4.230 ;
        RECT 79.605 3.950 79.885 4.230 ;
        RECT 86.685 13.410 86.965 13.690 ;
        RECT 89.325 13.810 89.605 14.090 ;
        RECT 89.325 13.410 89.605 13.690 ;
        RECT 86.685 9.610 86.965 9.890 ;
        RECT 86.685 9.210 86.965 9.490 ;
        RECT 89.325 9.610 89.605 9.890 ;
        RECT 89.325 9.210 89.605 9.490 ;
        RECT 93.185 47.410 93.465 47.690 ;
        RECT 93.185 47.010 93.465 47.290 ;
        RECT 95.825 47.410 96.105 47.690 ;
        RECT 95.825 47.010 96.105 47.290 ;
        RECT 93.185 43.210 93.465 43.490 ;
        RECT 93.185 42.810 93.465 43.090 ;
        RECT 95.825 43.210 96.105 43.490 ;
        RECT 95.825 42.810 96.105 43.090 ;
        RECT 93.185 39.010 93.465 39.290 ;
        RECT 93.185 38.610 93.465 38.890 ;
        RECT 95.825 39.010 96.105 39.290 ;
        RECT 95.825 38.610 96.105 38.890 ;
        RECT 93.185 34.810 93.465 35.090 ;
        RECT 93.185 34.410 93.465 34.690 ;
        RECT 95.825 34.810 96.105 35.090 ;
        RECT 95.825 34.410 96.105 34.690 ;
        RECT 93.185 30.610 93.465 30.890 ;
        RECT 93.185 30.210 93.465 30.490 ;
        RECT 95.825 30.610 96.105 30.890 ;
        RECT 95.825 30.210 96.105 30.490 ;
        RECT 93.185 26.410 93.465 26.690 ;
        RECT 93.185 26.010 93.465 26.290 ;
        RECT 95.825 26.410 96.105 26.690 ;
        RECT 95.825 26.010 96.105 26.290 ;
        RECT 93.185 22.210 93.465 22.490 ;
        RECT 93.185 21.810 93.465 22.090 ;
        RECT 95.825 22.210 96.105 22.490 ;
        RECT 95.825 21.810 96.105 22.090 ;
        RECT 93.185 18.010 93.465 18.290 ;
        RECT 93.185 17.610 93.465 17.890 ;
        RECT 95.825 18.010 96.105 18.290 ;
        RECT 95.825 17.610 96.105 17.890 ;
        RECT 93.185 13.810 93.465 14.090 ;
        RECT 85.705 3.150 85.985 3.430 ;
        RECT 86.105 3.150 86.385 3.430 ;
        RECT 93.185 13.410 93.465 13.690 ;
        RECT 95.825 13.810 96.105 14.090 ;
        RECT 95.825 13.410 96.105 13.690 ;
        RECT 93.185 9.610 93.465 9.890 ;
        RECT 93.185 9.210 93.465 9.490 ;
        RECT 95.825 9.610 96.105 9.890 ;
        RECT 95.825 9.210 96.105 9.490 ;
        RECT 99.685 47.410 99.965 47.690 ;
        RECT 99.685 47.010 99.965 47.290 ;
        RECT 102.325 47.410 102.605 47.690 ;
        RECT 102.325 47.010 102.605 47.290 ;
        RECT 99.685 43.210 99.965 43.490 ;
        RECT 99.685 42.810 99.965 43.090 ;
        RECT 102.325 43.210 102.605 43.490 ;
        RECT 102.325 42.810 102.605 43.090 ;
        RECT 99.685 39.010 99.965 39.290 ;
        RECT 99.685 38.610 99.965 38.890 ;
        RECT 102.325 39.010 102.605 39.290 ;
        RECT 102.325 38.610 102.605 38.890 ;
        RECT 99.685 34.810 99.965 35.090 ;
        RECT 99.685 34.410 99.965 34.690 ;
        RECT 102.325 34.810 102.605 35.090 ;
        RECT 102.325 34.410 102.605 34.690 ;
        RECT 99.685 30.610 99.965 30.890 ;
        RECT 99.685 30.210 99.965 30.490 ;
        RECT 102.325 30.610 102.605 30.890 ;
        RECT 102.325 30.210 102.605 30.490 ;
        RECT 99.685 26.410 99.965 26.690 ;
        RECT 99.685 26.010 99.965 26.290 ;
        RECT 102.325 26.410 102.605 26.690 ;
        RECT 102.325 26.010 102.605 26.290 ;
        RECT 99.685 22.210 99.965 22.490 ;
        RECT 99.685 21.810 99.965 22.090 ;
        RECT 102.325 22.210 102.605 22.490 ;
        RECT 102.325 21.810 102.605 22.090 ;
        RECT 99.685 18.010 99.965 18.290 ;
        RECT 99.685 17.610 99.965 17.890 ;
        RECT 102.325 18.010 102.605 18.290 ;
        RECT 102.325 17.610 102.605 17.890 ;
        RECT 99.685 13.810 99.965 14.090 ;
        RECT 99.685 13.410 99.965 13.690 ;
        RECT 102.325 13.810 102.605 14.090 ;
        RECT 102.325 13.410 102.605 13.690 ;
        RECT 99.685 9.610 99.965 9.890 ;
        RECT 99.685 9.210 99.965 9.490 ;
        RECT 102.325 9.610 102.605 9.890 ;
        RECT 102.325 9.210 102.605 9.490 ;
        RECT 106.185 47.410 106.465 47.690 ;
        RECT 106.185 47.010 106.465 47.290 ;
        RECT 108.825 47.410 109.105 47.690 ;
        RECT 108.825 47.010 109.105 47.290 ;
        RECT 106.185 43.210 106.465 43.490 ;
        RECT 106.185 42.810 106.465 43.090 ;
        RECT 108.825 43.210 109.105 43.490 ;
        RECT 108.825 42.810 109.105 43.090 ;
        RECT 106.185 39.010 106.465 39.290 ;
        RECT 104.555 34.810 104.835 35.090 ;
        RECT 104.555 34.410 104.835 34.690 ;
        RECT 104.555 22.210 104.835 22.490 ;
        RECT 104.555 21.810 104.835 22.090 ;
        RECT 106.185 38.610 106.465 38.890 ;
        RECT 108.825 39.010 109.105 39.290 ;
        RECT 108.825 38.610 109.105 38.890 ;
        RECT 106.185 34.810 106.465 35.090 ;
        RECT 106.185 34.410 106.465 34.690 ;
        RECT 108.825 34.810 109.105 35.090 ;
        RECT 108.825 34.410 109.105 34.690 ;
        RECT 106.185 30.610 106.465 30.890 ;
        RECT 106.185 30.210 106.465 30.490 ;
        RECT 108.825 30.610 109.105 30.890 ;
        RECT 108.825 30.210 109.105 30.490 ;
        RECT 106.185 26.410 106.465 26.690 ;
        RECT 106.185 26.010 106.465 26.290 ;
        RECT 108.825 26.410 109.105 26.690 ;
        RECT 110.455 30.610 110.735 30.890 ;
        RECT 110.455 30.210 110.735 30.490 ;
        RECT 112.685 47.410 112.965 47.690 ;
        RECT 112.685 47.010 112.965 47.290 ;
        RECT 115.325 47.410 115.605 47.690 ;
        RECT 115.325 47.010 115.605 47.290 ;
        RECT 112.685 43.210 112.965 43.490 ;
        RECT 112.685 42.810 112.965 43.090 ;
        RECT 115.325 43.210 115.605 43.490 ;
        RECT 115.325 42.810 115.605 43.090 ;
        RECT 112.685 39.010 112.965 39.290 ;
        RECT 112.685 38.610 112.965 38.890 ;
        RECT 115.325 39.010 115.605 39.290 ;
        RECT 115.325 38.610 115.605 38.890 ;
        RECT 112.685 34.810 112.965 35.090 ;
        RECT 112.685 34.410 112.965 34.690 ;
        RECT 115.325 34.810 115.605 35.090 ;
        RECT 115.325 34.410 115.605 34.690 ;
        RECT 112.685 30.610 112.965 30.890 ;
        RECT 108.825 26.010 109.105 26.290 ;
        RECT 106.185 22.210 106.465 22.490 ;
        RECT 106.185 21.810 106.465 22.090 ;
        RECT 108.825 22.210 109.105 22.490 ;
        RECT 108.825 21.810 109.105 22.090 ;
        RECT 106.185 18.010 106.465 18.290 ;
        RECT 106.185 17.610 106.465 17.890 ;
        RECT 108.825 18.010 109.105 18.290 ;
        RECT 108.825 17.610 109.105 17.890 ;
        RECT 106.185 13.810 106.465 14.090 ;
        RECT 106.185 13.410 106.465 13.690 ;
        RECT 108.825 13.810 109.105 14.090 ;
        RECT 108.825 13.410 109.105 13.690 ;
        RECT 106.185 9.610 106.465 9.890 ;
        RECT 106.185 9.210 106.465 9.490 ;
        RECT 108.825 9.610 109.105 9.890 ;
        RECT 108.825 9.210 109.105 9.490 ;
        RECT 111.055 26.410 111.335 26.690 ;
        RECT 111.055 26.010 111.335 26.290 ;
        RECT 112.685 30.210 112.965 30.490 ;
        RECT 115.325 30.610 115.605 30.890 ;
        RECT 115.325 30.210 115.605 30.490 ;
        RECT 112.685 26.410 112.965 26.690 ;
        RECT 112.685 26.010 112.965 26.290 ;
        RECT 115.325 26.410 115.605 26.690 ;
        RECT 115.325 26.010 115.605 26.290 ;
        RECT 112.685 22.210 112.965 22.490 ;
        RECT 112.685 21.810 112.965 22.090 ;
        RECT 115.325 22.210 115.605 22.490 ;
        RECT 115.325 21.810 115.605 22.090 ;
        RECT 112.685 18.010 112.965 18.290 ;
        RECT 112.685 17.610 112.965 17.890 ;
        RECT 115.325 18.010 115.605 18.290 ;
        RECT 116.955 34.810 117.235 35.090 ;
        RECT 116.955 34.410 117.235 34.690 ;
        RECT 116.955 22.210 117.235 22.490 ;
        RECT 116.955 21.810 117.235 22.090 ;
        RECT 115.325 17.610 115.605 17.890 ;
        RECT 112.685 13.810 112.965 14.090 ;
        RECT 112.685 13.410 112.965 13.690 ;
        RECT 115.325 13.810 115.605 14.090 ;
        RECT 115.325 13.410 115.605 13.690 ;
        RECT 112.685 9.610 112.965 9.890 ;
        RECT 112.685 9.210 112.965 9.490 ;
        RECT 115.325 9.610 115.605 9.890 ;
        RECT 115.325 9.210 115.605 9.490 ;
        RECT 108.205 7.150 108.485 7.430 ;
        RECT 108.605 7.150 108.885 7.430 ;
        RECT 112.905 7.150 113.185 7.430 ;
        RECT 113.305 7.150 113.585 7.430 ;
        RECT 105.205 5.550 105.485 5.830 ;
        RECT 105.605 5.550 105.885 5.830 ;
        RECT 98.705 4.750 98.985 5.030 ;
        RECT 99.105 4.750 99.385 5.030 ;
        RECT 7.705 2.350 7.985 2.630 ;
        RECT 8.105 2.350 8.385 2.630 ;
        RECT 20.705 2.350 20.985 2.630 ;
        RECT 21.105 2.350 21.385 2.630 ;
        RECT 27.205 2.350 27.485 2.630 ;
        RECT 27.605 2.350 27.885 2.630 ;
        RECT 40.205 2.350 40.485 2.630 ;
        RECT 40.605 2.350 40.885 2.630 ;
        RECT 46.705 2.350 46.985 2.630 ;
        RECT 47.105 2.350 47.385 2.630 ;
        RECT 66.205 2.350 66.485 2.630 ;
        RECT 66.605 2.350 66.885 2.630 ;
        RECT 72.705 2.350 72.985 2.630 ;
        RECT 73.105 2.350 73.385 2.630 ;
        RECT 92.205 2.350 92.485 2.630 ;
        RECT 92.605 2.350 92.885 2.630 ;
        RECT 110.405 1.550 110.685 1.830 ;
        RECT 110.805 1.550 111.085 1.830 ;
        RECT 107.905 0.750 108.185 1.030 ;
        RECT 108.305 0.750 108.585 1.030 ;
        RECT 119.185 47.410 119.465 47.690 ;
        RECT 119.185 47.010 119.465 47.290 ;
        RECT 121.825 47.410 122.105 47.690 ;
        RECT 121.825 47.010 122.105 47.290 ;
        RECT 119.185 43.210 119.465 43.490 ;
        RECT 119.185 42.810 119.465 43.090 ;
        RECT 121.825 43.210 122.105 43.490 ;
        RECT 121.825 42.810 122.105 43.090 ;
        RECT 119.185 39.010 119.465 39.290 ;
        RECT 119.185 38.610 119.465 38.890 ;
        RECT 121.825 39.010 122.105 39.290 ;
        RECT 121.825 38.610 122.105 38.890 ;
        RECT 119.185 34.810 119.465 35.090 ;
        RECT 119.185 34.410 119.465 34.690 ;
        RECT 121.825 34.810 122.105 35.090 ;
        RECT 121.825 34.410 122.105 34.690 ;
        RECT 119.185 30.610 119.465 30.890 ;
        RECT 119.185 30.210 119.465 30.490 ;
        RECT 121.825 30.610 122.105 30.890 ;
        RECT 121.825 30.210 122.105 30.490 ;
        RECT 119.185 26.410 119.465 26.690 ;
        RECT 119.185 26.010 119.465 26.290 ;
        RECT 121.825 26.410 122.105 26.690 ;
        RECT 121.825 26.010 122.105 26.290 ;
        RECT 119.185 22.210 119.465 22.490 ;
        RECT 119.185 21.810 119.465 22.090 ;
        RECT 121.825 22.210 122.105 22.490 ;
        RECT 121.825 21.810 122.105 22.090 ;
        RECT 119.185 18.010 119.465 18.290 ;
        RECT 119.185 17.610 119.465 17.890 ;
        RECT 121.825 18.010 122.105 18.290 ;
        RECT 121.825 17.610 122.105 17.890 ;
        RECT 119.185 13.810 119.465 14.090 ;
        RECT 119.185 13.410 119.465 13.690 ;
        RECT 121.825 13.810 122.105 14.090 ;
        RECT 121.825 13.410 122.105 13.690 ;
        RECT 119.185 9.610 119.465 9.890 ;
        RECT 119.185 9.210 119.465 9.490 ;
        RECT 121.825 9.610 122.105 9.890 ;
        RECT 121.825 9.210 122.105 9.490 ;
        RECT 115.905 5.550 116.185 5.830 ;
        RECT 116.305 5.550 116.585 5.830 ;
        RECT 125.685 47.410 125.965 47.690 ;
        RECT 125.685 47.010 125.965 47.290 ;
        RECT 128.325 47.410 128.605 47.690 ;
        RECT 128.325 47.010 128.605 47.290 ;
        RECT 125.685 43.210 125.965 43.490 ;
        RECT 125.685 42.810 125.965 43.090 ;
        RECT 128.325 43.210 128.605 43.490 ;
        RECT 128.325 42.810 128.605 43.090 ;
        RECT 125.685 39.010 125.965 39.290 ;
        RECT 125.685 38.610 125.965 38.890 ;
        RECT 128.325 39.010 128.605 39.290 ;
        RECT 128.325 38.610 128.605 38.890 ;
        RECT 125.685 34.810 125.965 35.090 ;
        RECT 125.685 34.410 125.965 34.690 ;
        RECT 128.325 34.810 128.605 35.090 ;
        RECT 128.325 34.410 128.605 34.690 ;
        RECT 125.685 30.610 125.965 30.890 ;
        RECT 125.685 30.210 125.965 30.490 ;
        RECT 128.325 30.610 128.605 30.890 ;
        RECT 128.325 30.210 128.605 30.490 ;
        RECT 125.685 26.410 125.965 26.690 ;
        RECT 125.685 26.010 125.965 26.290 ;
        RECT 128.325 26.410 128.605 26.690 ;
        RECT 128.325 26.010 128.605 26.290 ;
        RECT 125.685 22.210 125.965 22.490 ;
        RECT 125.685 21.810 125.965 22.090 ;
        RECT 128.325 22.210 128.605 22.490 ;
        RECT 128.325 21.810 128.605 22.090 ;
        RECT 125.685 18.010 125.965 18.290 ;
        RECT 125.685 17.610 125.965 17.890 ;
        RECT 128.325 18.010 128.605 18.290 ;
        RECT 128.325 17.610 128.605 17.890 ;
        RECT 125.685 13.810 125.965 14.090 ;
        RECT 125.685 13.410 125.965 13.690 ;
        RECT 128.325 13.810 128.605 14.090 ;
        RECT 128.325 13.410 128.605 13.690 ;
        RECT 125.685 9.610 125.965 9.890 ;
        RECT 125.685 9.210 125.965 9.490 ;
        RECT 128.325 9.610 128.605 9.890 ;
        RECT 128.325 9.210 128.605 9.490 ;
        RECT 122.405 4.750 122.685 5.030 ;
        RECT 122.805 4.750 123.085 5.030 ;
        RECT 132.185 47.410 132.465 47.690 ;
        RECT 132.185 47.010 132.465 47.290 ;
        RECT 134.825 47.410 135.105 47.690 ;
        RECT 134.825 47.010 135.105 47.290 ;
        RECT 132.185 43.210 132.465 43.490 ;
        RECT 132.185 42.810 132.465 43.090 ;
        RECT 134.825 43.210 135.105 43.490 ;
        RECT 134.825 42.810 135.105 43.090 ;
        RECT 132.185 39.010 132.465 39.290 ;
        RECT 132.185 38.610 132.465 38.890 ;
        RECT 134.825 39.010 135.105 39.290 ;
        RECT 134.825 38.610 135.105 38.890 ;
        RECT 132.185 34.810 132.465 35.090 ;
        RECT 132.185 34.410 132.465 34.690 ;
        RECT 134.825 34.810 135.105 35.090 ;
        RECT 134.825 34.410 135.105 34.690 ;
        RECT 132.185 30.610 132.465 30.890 ;
        RECT 132.185 30.210 132.465 30.490 ;
        RECT 134.825 30.610 135.105 30.890 ;
        RECT 134.825 30.210 135.105 30.490 ;
        RECT 132.185 26.410 132.465 26.690 ;
        RECT 132.185 26.010 132.465 26.290 ;
        RECT 134.825 26.410 135.105 26.690 ;
        RECT 134.825 26.010 135.105 26.290 ;
        RECT 132.185 22.210 132.465 22.490 ;
        RECT 132.185 21.810 132.465 22.090 ;
        RECT 134.825 22.210 135.105 22.490 ;
        RECT 134.825 21.810 135.105 22.090 ;
        RECT 132.185 18.010 132.465 18.290 ;
        RECT 132.185 17.610 132.465 17.890 ;
        RECT 134.825 18.010 135.105 18.290 ;
        RECT 134.825 17.610 135.105 17.890 ;
        RECT 132.185 13.810 132.465 14.090 ;
        RECT 132.185 13.410 132.465 13.690 ;
        RECT 134.825 13.810 135.105 14.090 ;
        RECT 134.825 13.410 135.105 13.690 ;
        RECT 132.185 9.610 132.465 9.890 ;
        RECT 132.185 9.210 132.465 9.490 ;
        RECT 134.825 9.610 135.105 9.890 ;
        RECT 134.825 9.210 135.105 9.490 ;
        RECT 138.685 47.410 138.965 47.690 ;
        RECT 138.685 47.010 138.965 47.290 ;
        RECT 141.325 47.410 141.605 47.690 ;
        RECT 141.325 47.010 141.605 47.290 ;
        RECT 138.685 43.210 138.965 43.490 ;
        RECT 138.685 42.810 138.965 43.090 ;
        RECT 141.325 43.210 141.605 43.490 ;
        RECT 141.325 42.810 141.605 43.090 ;
        RECT 138.685 39.010 138.965 39.290 ;
        RECT 138.685 38.610 138.965 38.890 ;
        RECT 141.325 39.010 141.605 39.290 ;
        RECT 141.325 38.610 141.605 38.890 ;
        RECT 138.685 34.810 138.965 35.090 ;
        RECT 138.685 34.410 138.965 34.690 ;
        RECT 141.325 34.810 141.605 35.090 ;
        RECT 141.325 34.410 141.605 34.690 ;
        RECT 138.685 30.610 138.965 30.890 ;
        RECT 138.685 30.210 138.965 30.490 ;
        RECT 141.325 30.610 141.605 30.890 ;
        RECT 141.325 30.210 141.605 30.490 ;
        RECT 138.685 26.410 138.965 26.690 ;
        RECT 138.685 26.010 138.965 26.290 ;
        RECT 141.325 26.410 141.605 26.690 ;
        RECT 141.325 26.010 141.605 26.290 ;
        RECT 138.685 22.210 138.965 22.490 ;
        RECT 138.685 21.810 138.965 22.090 ;
        RECT 141.325 22.210 141.605 22.490 ;
        RECT 141.325 21.810 141.605 22.090 ;
        RECT 138.685 18.010 138.965 18.290 ;
        RECT 138.685 17.610 138.965 17.890 ;
        RECT 141.325 18.010 141.605 18.290 ;
        RECT 141.325 17.610 141.605 17.890 ;
        RECT 138.685 13.810 138.965 14.090 ;
        RECT 138.685 13.410 138.965 13.690 ;
        RECT 141.325 13.810 141.605 14.090 ;
        RECT 141.325 13.410 141.605 13.690 ;
        RECT 138.685 9.610 138.965 9.890 ;
        RECT 138.685 9.210 138.965 9.490 ;
        RECT 141.325 9.610 141.605 9.890 ;
        RECT 141.325 9.210 141.605 9.490 ;
        RECT 145.185 47.410 145.465 47.690 ;
        RECT 145.185 47.010 145.465 47.290 ;
        RECT 147.825 47.410 148.105 47.690 ;
        RECT 147.825 47.010 148.105 47.290 ;
        RECT 145.185 43.210 145.465 43.490 ;
        RECT 145.185 42.810 145.465 43.090 ;
        RECT 147.825 43.210 148.105 43.490 ;
        RECT 147.825 42.810 148.105 43.090 ;
        RECT 145.185 39.010 145.465 39.290 ;
        RECT 145.185 38.610 145.465 38.890 ;
        RECT 147.825 39.010 148.105 39.290 ;
        RECT 147.825 38.610 148.105 38.890 ;
        RECT 145.185 34.810 145.465 35.090 ;
        RECT 145.185 34.410 145.465 34.690 ;
        RECT 147.825 34.810 148.105 35.090 ;
        RECT 147.825 34.410 148.105 34.690 ;
        RECT 145.185 30.610 145.465 30.890 ;
        RECT 145.185 30.210 145.465 30.490 ;
        RECT 147.825 30.610 148.105 30.890 ;
        RECT 147.825 30.210 148.105 30.490 ;
        RECT 145.185 26.410 145.465 26.690 ;
        RECT 145.185 26.010 145.465 26.290 ;
        RECT 147.825 26.410 148.105 26.690 ;
        RECT 147.825 26.010 148.105 26.290 ;
        RECT 145.185 22.210 145.465 22.490 ;
        RECT 145.185 21.810 145.465 22.090 ;
        RECT 147.825 22.210 148.105 22.490 ;
        RECT 147.825 21.810 148.105 22.090 ;
        RECT 145.185 18.010 145.465 18.290 ;
        RECT 145.185 17.610 145.465 17.890 ;
        RECT 147.825 18.010 148.105 18.290 ;
        RECT 147.825 17.610 148.105 17.890 ;
        RECT 145.185 13.810 145.465 14.090 ;
        RECT 145.185 13.410 145.465 13.690 ;
        RECT 147.825 13.810 148.105 14.090 ;
        RECT 147.825 13.410 148.105 13.690 ;
        RECT 145.185 9.610 145.465 9.890 ;
        RECT 145.185 9.210 145.465 9.490 ;
        RECT 147.825 9.610 148.105 9.890 ;
        RECT 147.825 9.210 148.105 9.490 ;
        RECT 141.905 3.950 142.185 4.230 ;
        RECT 142.305 3.950 142.585 4.230 ;
        RECT 135.405 3.150 135.685 3.430 ;
        RECT 135.805 3.150 136.085 3.430 ;
        RECT 151.685 47.410 151.965 47.690 ;
        RECT 151.685 47.010 151.965 47.290 ;
        RECT 154.325 47.410 154.605 47.690 ;
        RECT 154.325 47.010 154.605 47.290 ;
        RECT 151.685 43.210 151.965 43.490 ;
        RECT 151.685 42.810 151.965 43.090 ;
        RECT 154.325 43.210 154.605 43.490 ;
        RECT 154.325 42.810 154.605 43.090 ;
        RECT 151.685 39.010 151.965 39.290 ;
        RECT 151.685 38.610 151.965 38.890 ;
        RECT 154.325 39.010 154.605 39.290 ;
        RECT 154.325 38.610 154.605 38.890 ;
        RECT 151.685 34.810 151.965 35.090 ;
        RECT 151.685 34.410 151.965 34.690 ;
        RECT 154.325 34.810 154.605 35.090 ;
        RECT 154.325 34.410 154.605 34.690 ;
        RECT 151.685 30.610 151.965 30.890 ;
        RECT 151.685 30.210 151.965 30.490 ;
        RECT 154.325 30.610 154.605 30.890 ;
        RECT 154.325 30.210 154.605 30.490 ;
        RECT 151.685 26.410 151.965 26.690 ;
        RECT 151.685 26.010 151.965 26.290 ;
        RECT 154.325 26.410 154.605 26.690 ;
        RECT 154.325 26.010 154.605 26.290 ;
        RECT 151.685 22.210 151.965 22.490 ;
        RECT 151.685 21.810 151.965 22.090 ;
        RECT 154.325 22.210 154.605 22.490 ;
        RECT 154.325 21.810 154.605 22.090 ;
        RECT 151.685 18.010 151.965 18.290 ;
        RECT 151.685 17.610 151.965 17.890 ;
        RECT 154.325 18.010 154.605 18.290 ;
        RECT 154.325 17.610 154.605 17.890 ;
        RECT 151.685 13.810 151.965 14.090 ;
        RECT 151.685 13.410 151.965 13.690 ;
        RECT 154.325 13.810 154.605 14.090 ;
        RECT 154.325 13.410 154.605 13.690 ;
        RECT 151.685 9.610 151.965 9.890 ;
        RECT 151.685 9.210 151.965 9.490 ;
        RECT 154.325 9.610 154.605 9.890 ;
        RECT 154.325 9.210 154.605 9.490 ;
        RECT 158.185 47.410 158.465 47.690 ;
        RECT 158.185 47.010 158.465 47.290 ;
        RECT 160.825 47.410 161.105 47.690 ;
        RECT 160.825 47.010 161.105 47.290 ;
        RECT 158.185 43.210 158.465 43.490 ;
        RECT 158.185 42.810 158.465 43.090 ;
        RECT 160.825 43.210 161.105 43.490 ;
        RECT 160.825 42.810 161.105 43.090 ;
        RECT 158.185 39.010 158.465 39.290 ;
        RECT 158.185 38.610 158.465 38.890 ;
        RECT 160.825 39.010 161.105 39.290 ;
        RECT 160.825 38.610 161.105 38.890 ;
        RECT 158.185 34.810 158.465 35.090 ;
        RECT 158.185 34.410 158.465 34.690 ;
        RECT 160.825 34.810 161.105 35.090 ;
        RECT 160.825 34.410 161.105 34.690 ;
        RECT 158.185 30.610 158.465 30.890 ;
        RECT 158.185 30.210 158.465 30.490 ;
        RECT 160.825 30.610 161.105 30.890 ;
        RECT 160.825 30.210 161.105 30.490 ;
        RECT 158.185 26.410 158.465 26.690 ;
        RECT 158.185 26.010 158.465 26.290 ;
        RECT 160.825 26.410 161.105 26.690 ;
        RECT 160.825 26.010 161.105 26.290 ;
        RECT 158.185 22.210 158.465 22.490 ;
        RECT 158.185 21.810 158.465 22.090 ;
        RECT 160.825 22.210 161.105 22.490 ;
        RECT 160.825 21.810 161.105 22.090 ;
        RECT 158.185 18.010 158.465 18.290 ;
        RECT 158.185 17.610 158.465 17.890 ;
        RECT 160.825 18.010 161.105 18.290 ;
        RECT 160.825 17.610 161.105 17.890 ;
        RECT 158.185 13.810 158.465 14.090 ;
        RECT 158.185 13.410 158.465 13.690 ;
        RECT 160.825 13.810 161.105 14.090 ;
        RECT 160.825 13.410 161.105 13.690 ;
        RECT 158.185 9.610 158.465 9.890 ;
        RECT 158.185 9.210 158.465 9.490 ;
        RECT 160.825 9.610 161.105 9.890 ;
        RECT 160.825 9.210 161.105 9.490 ;
        RECT 164.685 47.410 164.965 47.690 ;
        RECT 164.685 47.010 164.965 47.290 ;
        RECT 167.325 47.410 167.605 47.690 ;
        RECT 167.325 47.010 167.605 47.290 ;
        RECT 164.685 43.210 164.965 43.490 ;
        RECT 164.685 42.810 164.965 43.090 ;
        RECT 167.325 43.210 167.605 43.490 ;
        RECT 167.325 42.810 167.605 43.090 ;
        RECT 164.685 39.010 164.965 39.290 ;
        RECT 164.685 38.610 164.965 38.890 ;
        RECT 167.325 39.010 167.605 39.290 ;
        RECT 167.325 38.610 167.605 38.890 ;
        RECT 164.685 34.810 164.965 35.090 ;
        RECT 164.685 34.410 164.965 34.690 ;
        RECT 167.325 34.810 167.605 35.090 ;
        RECT 167.325 34.410 167.605 34.690 ;
        RECT 164.685 30.610 164.965 30.890 ;
        RECT 164.685 30.210 164.965 30.490 ;
        RECT 167.325 30.610 167.605 30.890 ;
        RECT 167.325 30.210 167.605 30.490 ;
        RECT 164.685 26.410 164.965 26.690 ;
        RECT 164.685 26.010 164.965 26.290 ;
        RECT 167.325 26.410 167.605 26.690 ;
        RECT 167.325 26.010 167.605 26.290 ;
        RECT 164.685 22.210 164.965 22.490 ;
        RECT 164.685 21.810 164.965 22.090 ;
        RECT 167.325 22.210 167.605 22.490 ;
        RECT 167.325 21.810 167.605 22.090 ;
        RECT 164.685 18.010 164.965 18.290 ;
        RECT 164.685 17.610 164.965 17.890 ;
        RECT 167.325 18.010 167.605 18.290 ;
        RECT 167.325 17.610 167.605 17.890 ;
        RECT 164.685 13.810 164.965 14.090 ;
        RECT 164.685 13.410 164.965 13.690 ;
        RECT 167.325 13.810 167.605 14.090 ;
        RECT 167.325 13.410 167.605 13.690 ;
        RECT 164.685 9.610 164.965 9.890 ;
        RECT 164.685 9.210 164.965 9.490 ;
        RECT 167.325 9.610 167.605 9.890 ;
        RECT 167.325 9.210 167.605 9.490 ;
        RECT 171.185 47.410 171.465 47.690 ;
        RECT 171.185 47.010 171.465 47.290 ;
        RECT 173.825 47.410 174.105 47.690 ;
        RECT 173.825 47.010 174.105 47.290 ;
        RECT 171.185 43.210 171.465 43.490 ;
        RECT 171.185 42.810 171.465 43.090 ;
        RECT 173.825 43.210 174.105 43.490 ;
        RECT 173.825 42.810 174.105 43.090 ;
        RECT 171.185 39.010 171.465 39.290 ;
        RECT 171.185 38.610 171.465 38.890 ;
        RECT 173.825 39.010 174.105 39.290 ;
        RECT 173.825 38.610 174.105 38.890 ;
        RECT 171.185 34.810 171.465 35.090 ;
        RECT 171.185 34.410 171.465 34.690 ;
        RECT 173.825 34.810 174.105 35.090 ;
        RECT 173.825 34.410 174.105 34.690 ;
        RECT 171.185 30.610 171.465 30.890 ;
        RECT 171.185 30.210 171.465 30.490 ;
        RECT 173.825 30.610 174.105 30.890 ;
        RECT 173.825 30.210 174.105 30.490 ;
        RECT 171.185 26.410 171.465 26.690 ;
        RECT 171.185 26.010 171.465 26.290 ;
        RECT 173.825 26.410 174.105 26.690 ;
        RECT 173.825 26.010 174.105 26.290 ;
        RECT 171.185 22.210 171.465 22.490 ;
        RECT 171.185 21.810 171.465 22.090 ;
        RECT 173.825 22.210 174.105 22.490 ;
        RECT 173.825 21.810 174.105 22.090 ;
        RECT 171.185 18.010 171.465 18.290 ;
        RECT 171.185 17.610 171.465 17.890 ;
        RECT 173.825 18.010 174.105 18.290 ;
        RECT 173.825 17.610 174.105 17.890 ;
        RECT 171.185 13.810 171.465 14.090 ;
        RECT 171.185 13.410 171.465 13.690 ;
        RECT 173.825 13.810 174.105 14.090 ;
        RECT 173.825 13.410 174.105 13.690 ;
        RECT 171.185 9.610 171.465 9.890 ;
        RECT 171.185 9.210 171.465 9.490 ;
        RECT 173.825 9.610 174.105 9.890 ;
        RECT 173.825 9.210 174.105 9.490 ;
        RECT 167.905 3.950 168.185 4.230 ;
        RECT 168.305 3.950 168.585 4.230 ;
        RECT 161.405 3.150 161.685 3.430 ;
        RECT 161.805 3.150 162.085 3.430 ;
        RECT 177.685 47.410 177.965 47.690 ;
        RECT 177.685 47.010 177.965 47.290 ;
        RECT 180.325 47.410 180.605 47.690 ;
        RECT 180.325 47.010 180.605 47.290 ;
        RECT 177.685 43.210 177.965 43.490 ;
        RECT 177.685 42.810 177.965 43.090 ;
        RECT 180.325 43.210 180.605 43.490 ;
        RECT 180.325 42.810 180.605 43.090 ;
        RECT 177.685 39.010 177.965 39.290 ;
        RECT 177.685 38.610 177.965 38.890 ;
        RECT 180.325 39.010 180.605 39.290 ;
        RECT 180.325 38.610 180.605 38.890 ;
        RECT 177.685 34.810 177.965 35.090 ;
        RECT 177.685 34.410 177.965 34.690 ;
        RECT 180.325 34.810 180.605 35.090 ;
        RECT 180.325 34.410 180.605 34.690 ;
        RECT 177.685 30.610 177.965 30.890 ;
        RECT 177.685 30.210 177.965 30.490 ;
        RECT 180.325 30.610 180.605 30.890 ;
        RECT 180.325 30.210 180.605 30.490 ;
        RECT 177.685 26.410 177.965 26.690 ;
        RECT 177.685 26.010 177.965 26.290 ;
        RECT 180.325 26.410 180.605 26.690 ;
        RECT 180.325 26.010 180.605 26.290 ;
        RECT 177.685 22.210 177.965 22.490 ;
        RECT 177.685 21.810 177.965 22.090 ;
        RECT 180.325 22.210 180.605 22.490 ;
        RECT 180.325 21.810 180.605 22.090 ;
        RECT 177.685 18.010 177.965 18.290 ;
        RECT 177.685 17.610 177.965 17.890 ;
        RECT 180.325 18.010 180.605 18.290 ;
        RECT 180.325 17.610 180.605 17.890 ;
        RECT 177.685 13.810 177.965 14.090 ;
        RECT 177.685 13.410 177.965 13.690 ;
        RECT 180.325 13.810 180.605 14.090 ;
        RECT 180.325 13.410 180.605 13.690 ;
        RECT 177.685 9.610 177.965 9.890 ;
        RECT 177.685 9.210 177.965 9.490 ;
        RECT 180.325 9.610 180.605 9.890 ;
        RECT 180.325 9.210 180.605 9.490 ;
        RECT 184.185 47.410 184.465 47.690 ;
        RECT 184.185 47.010 184.465 47.290 ;
        RECT 186.825 47.410 187.105 47.690 ;
        RECT 186.825 47.010 187.105 47.290 ;
        RECT 184.185 43.210 184.465 43.490 ;
        RECT 184.185 42.810 184.465 43.090 ;
        RECT 186.825 43.210 187.105 43.490 ;
        RECT 186.825 42.810 187.105 43.090 ;
        RECT 184.185 39.010 184.465 39.290 ;
        RECT 184.185 38.610 184.465 38.890 ;
        RECT 186.825 39.010 187.105 39.290 ;
        RECT 186.825 38.610 187.105 38.890 ;
        RECT 184.185 34.810 184.465 35.090 ;
        RECT 184.185 34.410 184.465 34.690 ;
        RECT 186.825 34.810 187.105 35.090 ;
        RECT 186.825 34.410 187.105 34.690 ;
        RECT 184.185 30.610 184.465 30.890 ;
        RECT 184.185 30.210 184.465 30.490 ;
        RECT 186.825 30.610 187.105 30.890 ;
        RECT 186.825 30.210 187.105 30.490 ;
        RECT 184.185 26.410 184.465 26.690 ;
        RECT 184.185 26.010 184.465 26.290 ;
        RECT 186.825 26.410 187.105 26.690 ;
        RECT 186.825 26.010 187.105 26.290 ;
        RECT 184.185 22.210 184.465 22.490 ;
        RECT 184.185 21.810 184.465 22.090 ;
        RECT 186.825 22.210 187.105 22.490 ;
        RECT 186.825 21.810 187.105 22.090 ;
        RECT 184.185 18.010 184.465 18.290 ;
        RECT 184.185 17.610 184.465 17.890 ;
        RECT 186.825 18.010 187.105 18.290 ;
        RECT 186.825 17.610 187.105 17.890 ;
        RECT 184.185 13.810 184.465 14.090 ;
        RECT 184.185 13.410 184.465 13.690 ;
        RECT 186.825 13.810 187.105 14.090 ;
        RECT 186.825 13.410 187.105 13.690 ;
        RECT 184.185 9.610 184.465 9.890 ;
        RECT 184.185 9.210 184.465 9.490 ;
        RECT 186.825 9.610 187.105 9.890 ;
        RECT 186.825 9.210 187.105 9.490 ;
        RECT 190.685 47.410 190.965 47.690 ;
        RECT 190.685 47.010 190.965 47.290 ;
        RECT 193.325 47.410 193.605 47.690 ;
        RECT 193.325 47.010 193.605 47.290 ;
        RECT 190.685 43.210 190.965 43.490 ;
        RECT 190.685 42.810 190.965 43.090 ;
        RECT 193.325 43.210 193.605 43.490 ;
        RECT 193.325 42.810 193.605 43.090 ;
        RECT 190.685 39.010 190.965 39.290 ;
        RECT 190.685 38.610 190.965 38.890 ;
        RECT 193.325 39.010 193.605 39.290 ;
        RECT 193.325 38.610 193.605 38.890 ;
        RECT 190.685 34.810 190.965 35.090 ;
        RECT 190.685 34.410 190.965 34.690 ;
        RECT 193.325 34.810 193.605 35.090 ;
        RECT 193.325 34.410 193.605 34.690 ;
        RECT 190.685 30.610 190.965 30.890 ;
        RECT 190.685 30.210 190.965 30.490 ;
        RECT 193.325 30.610 193.605 30.890 ;
        RECT 193.325 30.210 193.605 30.490 ;
        RECT 190.685 26.410 190.965 26.690 ;
        RECT 190.685 26.010 190.965 26.290 ;
        RECT 193.325 26.410 193.605 26.690 ;
        RECT 193.325 26.010 193.605 26.290 ;
        RECT 190.685 22.210 190.965 22.490 ;
        RECT 190.685 21.810 190.965 22.090 ;
        RECT 193.325 22.210 193.605 22.490 ;
        RECT 193.325 21.810 193.605 22.090 ;
        RECT 190.685 18.010 190.965 18.290 ;
        RECT 190.685 17.610 190.965 17.890 ;
        RECT 193.325 18.010 193.605 18.290 ;
        RECT 193.325 17.610 193.605 17.890 ;
        RECT 190.685 13.810 190.965 14.090 ;
        RECT 190.685 13.410 190.965 13.690 ;
        RECT 193.325 13.810 193.605 14.090 ;
        RECT 193.325 13.410 193.605 13.690 ;
        RECT 190.685 9.610 190.965 9.890 ;
        RECT 190.685 9.210 190.965 9.490 ;
        RECT 193.325 9.610 193.605 9.890 ;
        RECT 193.325 9.210 193.605 9.490 ;
        RECT 187.405 3.150 187.685 3.430 ;
        RECT 187.805 3.150 188.085 3.430 ;
        RECT 197.185 47.410 197.465 47.690 ;
        RECT 197.185 47.010 197.465 47.290 ;
        RECT 199.825 47.410 200.105 47.690 ;
        RECT 199.825 47.010 200.105 47.290 ;
        RECT 197.185 43.210 197.465 43.490 ;
        RECT 197.185 42.810 197.465 43.090 ;
        RECT 199.825 43.210 200.105 43.490 ;
        RECT 199.825 42.810 200.105 43.090 ;
        RECT 197.185 39.010 197.465 39.290 ;
        RECT 197.185 38.610 197.465 38.890 ;
        RECT 199.825 39.010 200.105 39.290 ;
        RECT 199.825 38.610 200.105 38.890 ;
        RECT 197.185 34.810 197.465 35.090 ;
        RECT 197.185 34.410 197.465 34.690 ;
        RECT 199.825 34.810 200.105 35.090 ;
        RECT 199.825 34.410 200.105 34.690 ;
        RECT 197.185 30.610 197.465 30.890 ;
        RECT 197.185 30.210 197.465 30.490 ;
        RECT 199.825 30.610 200.105 30.890 ;
        RECT 199.825 30.210 200.105 30.490 ;
        RECT 197.185 26.410 197.465 26.690 ;
        RECT 197.185 26.010 197.465 26.290 ;
        RECT 199.825 26.410 200.105 26.690 ;
        RECT 199.825 26.010 200.105 26.290 ;
        RECT 197.185 22.210 197.465 22.490 ;
        RECT 197.185 21.810 197.465 22.090 ;
        RECT 199.825 22.210 200.105 22.490 ;
        RECT 199.825 21.810 200.105 22.090 ;
        RECT 197.185 18.010 197.465 18.290 ;
        RECT 197.185 17.610 197.465 17.890 ;
        RECT 199.825 18.010 200.105 18.290 ;
        RECT 199.825 17.610 200.105 17.890 ;
        RECT 197.185 13.810 197.465 14.090 ;
        RECT 197.185 13.410 197.465 13.690 ;
        RECT 199.825 13.810 200.105 14.090 ;
        RECT 199.825 13.410 200.105 13.690 ;
        RECT 197.185 9.610 197.465 9.890 ;
        RECT 197.185 9.210 197.465 9.490 ;
        RECT 199.825 9.610 200.105 9.890 ;
        RECT 199.825 9.210 200.105 9.490 ;
        RECT 203.685 47.410 203.965 47.690 ;
        RECT 203.685 47.010 203.965 47.290 ;
        RECT 206.325 47.410 206.605 47.690 ;
        RECT 206.325 47.010 206.605 47.290 ;
        RECT 203.685 43.210 203.965 43.490 ;
        RECT 203.685 42.810 203.965 43.090 ;
        RECT 206.325 43.210 206.605 43.490 ;
        RECT 206.325 42.810 206.605 43.090 ;
        RECT 203.685 39.010 203.965 39.290 ;
        RECT 203.685 38.610 203.965 38.890 ;
        RECT 206.325 39.010 206.605 39.290 ;
        RECT 206.325 38.610 206.605 38.890 ;
        RECT 203.685 34.810 203.965 35.090 ;
        RECT 203.685 34.410 203.965 34.690 ;
        RECT 206.325 34.810 206.605 35.090 ;
        RECT 206.325 34.410 206.605 34.690 ;
        RECT 203.685 30.610 203.965 30.890 ;
        RECT 203.685 30.210 203.965 30.490 ;
        RECT 206.325 30.610 206.605 30.890 ;
        RECT 206.325 30.210 206.605 30.490 ;
        RECT 203.685 26.410 203.965 26.690 ;
        RECT 203.685 26.010 203.965 26.290 ;
        RECT 206.325 26.410 206.605 26.690 ;
        RECT 206.325 26.010 206.605 26.290 ;
        RECT 203.685 22.210 203.965 22.490 ;
        RECT 203.685 21.810 203.965 22.090 ;
        RECT 206.325 22.210 206.605 22.490 ;
        RECT 206.325 21.810 206.605 22.090 ;
        RECT 203.685 18.010 203.965 18.290 ;
        RECT 203.685 17.610 203.965 17.890 ;
        RECT 206.325 18.010 206.605 18.290 ;
        RECT 206.325 17.610 206.605 17.890 ;
        RECT 203.685 13.810 203.965 14.090 ;
        RECT 203.685 13.410 203.965 13.690 ;
        RECT 206.325 13.810 206.605 14.090 ;
        RECT 206.325 13.410 206.605 13.690 ;
        RECT 203.685 9.610 203.965 9.890 ;
        RECT 203.685 9.210 203.965 9.490 ;
        RECT 206.325 9.610 206.605 9.890 ;
        RECT 206.325 9.210 206.605 9.490 ;
        RECT 210.185 47.410 210.465 47.690 ;
        RECT 210.185 47.010 210.465 47.290 ;
        RECT 212.825 47.410 213.105 47.690 ;
        RECT 212.825 47.010 213.105 47.290 ;
        RECT 210.185 43.210 210.465 43.490 ;
        RECT 210.185 42.810 210.465 43.090 ;
        RECT 212.825 43.210 213.105 43.490 ;
        RECT 212.825 42.810 213.105 43.090 ;
        RECT 210.185 39.010 210.465 39.290 ;
        RECT 210.185 38.610 210.465 38.890 ;
        RECT 212.825 39.010 213.105 39.290 ;
        RECT 212.825 38.610 213.105 38.890 ;
        RECT 210.185 34.810 210.465 35.090 ;
        RECT 210.185 34.410 210.465 34.690 ;
        RECT 212.825 34.810 213.105 35.090 ;
        RECT 212.825 34.410 213.105 34.690 ;
        RECT 210.185 30.610 210.465 30.890 ;
        RECT 210.185 30.210 210.465 30.490 ;
        RECT 212.825 30.610 213.105 30.890 ;
        RECT 212.825 30.210 213.105 30.490 ;
        RECT 210.185 26.410 210.465 26.690 ;
        RECT 210.185 26.010 210.465 26.290 ;
        RECT 212.825 26.410 213.105 26.690 ;
        RECT 212.825 26.010 213.105 26.290 ;
        RECT 210.185 22.210 210.465 22.490 ;
        RECT 210.185 21.810 210.465 22.090 ;
        RECT 212.825 22.210 213.105 22.490 ;
        RECT 212.825 21.810 213.105 22.090 ;
        RECT 210.185 18.010 210.465 18.290 ;
        RECT 210.185 17.610 210.465 17.890 ;
        RECT 212.825 18.010 213.105 18.290 ;
        RECT 212.825 17.610 213.105 17.890 ;
        RECT 210.185 13.810 210.465 14.090 ;
        RECT 210.185 13.410 210.465 13.690 ;
        RECT 212.825 13.810 213.105 14.090 ;
        RECT 212.825 13.410 213.105 13.690 ;
        RECT 210.185 9.610 210.465 9.890 ;
        RECT 210.185 9.210 210.465 9.490 ;
        RECT 212.825 9.610 213.105 9.890 ;
        RECT 212.825 9.210 213.105 9.490 ;
        RECT 206.905 3.150 207.185 3.430 ;
        RECT 207.305 3.150 207.585 3.430 ;
        RECT 216.685 47.410 216.965 47.690 ;
        RECT 216.685 47.010 216.965 47.290 ;
        RECT 219.325 47.410 219.605 47.690 ;
        RECT 219.325 47.010 219.605 47.290 ;
        RECT 216.685 43.210 216.965 43.490 ;
        RECT 216.685 42.810 216.965 43.090 ;
        RECT 219.325 43.210 219.605 43.490 ;
        RECT 219.325 42.810 219.605 43.090 ;
        RECT 216.685 39.010 216.965 39.290 ;
        RECT 216.685 38.610 216.965 38.890 ;
        RECT 219.325 39.010 219.605 39.290 ;
        RECT 219.325 38.610 219.605 38.890 ;
        RECT 216.685 34.810 216.965 35.090 ;
        RECT 216.685 34.410 216.965 34.690 ;
        RECT 219.325 34.810 219.605 35.090 ;
        RECT 219.325 34.410 219.605 34.690 ;
        RECT 216.685 30.610 216.965 30.890 ;
        RECT 216.685 30.210 216.965 30.490 ;
        RECT 219.325 30.610 219.605 30.890 ;
        RECT 219.325 30.210 219.605 30.490 ;
        RECT 216.685 26.410 216.965 26.690 ;
        RECT 216.685 26.010 216.965 26.290 ;
        RECT 219.325 26.410 219.605 26.690 ;
        RECT 219.325 26.010 219.605 26.290 ;
        RECT 216.685 22.210 216.965 22.490 ;
        RECT 216.685 21.810 216.965 22.090 ;
        RECT 219.325 22.210 219.605 22.490 ;
        RECT 219.325 21.810 219.605 22.090 ;
        RECT 216.685 18.010 216.965 18.290 ;
        RECT 216.685 17.610 216.965 17.890 ;
        RECT 219.325 18.010 219.605 18.290 ;
        RECT 219.325 17.610 219.605 17.890 ;
        RECT 216.685 13.810 216.965 14.090 ;
        RECT 216.685 13.410 216.965 13.690 ;
        RECT 219.325 13.810 219.605 14.090 ;
        RECT 219.325 13.410 219.605 13.690 ;
        RECT 216.685 9.610 216.965 9.890 ;
        RECT 216.685 9.210 216.965 9.490 ;
        RECT 219.325 9.610 219.605 9.890 ;
        RECT 219.325 9.210 219.605 9.490 ;
        RECT 128.905 2.350 129.185 2.630 ;
        RECT 129.305 2.350 129.585 2.630 ;
        RECT 148.405 2.350 148.685 2.630 ;
        RECT 148.805 2.350 149.085 2.630 ;
        RECT 154.905 2.350 155.185 2.630 ;
        RECT 155.305 2.350 155.585 2.630 ;
        RECT 174.405 2.350 174.685 2.630 ;
        RECT 174.805 2.350 175.085 2.630 ;
        RECT 180.905 2.350 181.185 2.630 ;
        RECT 181.305 2.350 181.585 2.630 ;
        RECT 193.905 2.350 194.185 2.630 ;
        RECT 194.305 2.350 194.585 2.630 ;
        RECT 200.405 2.350 200.685 2.630 ;
        RECT 200.805 2.350 201.085 2.630 ;
        RECT 213.405 2.350 213.685 2.630 ;
        RECT 213.805 2.350 214.085 2.630 ;
        RECT 112.905 -0.050 113.185 0.230 ;
        RECT 113.305 -0.050 113.585 0.230 ;
      LAYER met3 ;
        RECT 1.645 45.850 5.645 48.850 ;
        RECT 1.645 41.650 5.645 44.650 ;
        RECT 1.645 37.450 5.645 40.450 ;
        RECT 1.645 33.250 5.645 36.250 ;
        RECT 1.645 29.050 5.645 32.050 ;
        RECT 1.645 24.850 5.645 27.850 ;
        RECT 1.645 20.650 5.645 23.650 ;
        RECT 1.645 16.450 5.645 19.450 ;
        RECT -8.050 13.620 0.670 14.020 ;
        RECT -8.050 12.240 -0.030 12.640 ;
        RECT -8.050 10.860 -0.730 11.260 ;
        RECT -8.050 9.480 -1.430 9.880 ;
        RECT -8.050 8.100 -2.130 8.500 ;
        RECT -8.050 6.720 -2.830 7.120 ;
        RECT -8.050 5.340 -3.530 5.740 ;
        RECT -8.050 3.960 -4.230 4.360 ;
        RECT -8.050 2.580 -4.930 2.980 ;
        RECT -5.330 0.290 -4.930 2.580 ;
        RECT -4.630 1.090 -4.230 3.960 ;
        RECT -3.930 1.890 -3.530 5.340 ;
        RECT -3.230 2.690 -2.830 6.720 ;
        RECT -2.530 3.490 -2.130 8.100 ;
        RECT -1.830 4.290 -1.430 9.480 ;
        RECT -1.130 5.090 -0.730 10.860 ;
        RECT -0.430 5.890 -0.030 12.240 ;
        RECT 0.270 6.690 0.670 13.620 ;
        RECT 1.645 12.250 5.645 15.250 ;
        RECT 1.645 8.050 5.645 11.050 ;
        RECT 6.145 8.050 6.645 48.850 ;
        RECT 7.145 8.050 7.645 48.850 ;
        RECT 8.145 45.850 12.145 48.850 ;
        RECT 8.145 41.650 12.145 44.650 ;
        RECT 8.145 37.450 12.145 40.450 ;
        RECT 8.145 33.250 12.145 36.250 ;
        RECT 8.145 29.050 12.145 32.050 ;
        RECT 8.145 24.850 12.145 27.850 ;
        RECT 8.145 20.650 12.145 23.650 ;
        RECT 8.145 16.450 12.145 19.450 ;
        RECT 8.145 12.250 12.145 15.250 ;
        RECT 8.145 8.050 12.145 11.050 ;
        RECT 12.645 8.050 13.145 48.850 ;
        RECT 13.645 8.050 14.145 48.850 ;
        RECT 14.645 45.850 18.645 48.850 ;
        RECT 14.645 41.650 18.645 44.650 ;
        RECT 14.645 37.450 18.645 40.450 ;
        RECT 14.645 33.250 18.645 36.250 ;
        RECT 14.645 29.050 18.645 32.050 ;
        RECT 14.645 24.850 18.645 27.850 ;
        RECT 14.645 20.650 18.645 23.650 ;
        RECT 14.645 16.450 18.645 19.450 ;
        RECT 14.645 12.250 18.645 15.250 ;
        RECT 14.645 8.050 18.645 11.050 ;
        RECT 19.145 8.050 19.645 48.850 ;
        RECT 20.145 8.050 20.645 48.850 ;
        RECT 21.145 45.850 25.145 48.850 ;
        RECT 21.145 41.650 25.145 44.650 ;
        RECT 21.145 37.450 25.145 40.450 ;
        RECT 21.145 33.250 25.145 36.250 ;
        RECT 21.145 29.050 25.145 32.050 ;
        RECT 21.145 24.850 25.145 27.850 ;
        RECT 21.145 20.650 25.145 23.650 ;
        RECT 21.145 16.450 25.145 19.450 ;
        RECT 21.145 12.250 25.145 15.250 ;
        RECT 21.145 8.050 25.145 11.050 ;
        RECT 25.645 8.050 26.145 48.850 ;
        RECT 26.645 8.050 27.145 48.850 ;
        RECT 27.645 45.850 31.645 48.850 ;
        RECT 27.645 41.650 31.645 44.650 ;
        RECT 27.645 37.450 31.645 40.450 ;
        RECT 27.645 33.250 31.645 36.250 ;
        RECT 27.645 29.050 31.645 32.050 ;
        RECT 27.645 24.850 31.645 27.850 ;
        RECT 27.645 20.650 31.645 23.650 ;
        RECT 27.645 16.450 31.645 19.450 ;
        RECT 27.645 12.250 31.645 15.250 ;
        RECT 27.645 8.050 31.645 11.050 ;
        RECT 32.145 8.050 32.645 48.850 ;
        RECT 33.145 8.050 33.645 48.850 ;
        RECT 34.145 45.850 38.145 48.850 ;
        RECT 34.145 41.650 38.145 44.650 ;
        RECT 34.145 37.450 38.145 40.450 ;
        RECT 34.145 33.250 38.145 36.250 ;
        RECT 34.145 29.050 38.145 32.050 ;
        RECT 34.145 24.850 38.145 27.850 ;
        RECT 34.145 20.650 38.145 23.650 ;
        RECT 34.145 16.450 38.145 19.450 ;
        RECT 34.145 12.250 38.145 15.250 ;
        RECT 34.145 8.050 38.145 11.050 ;
        RECT 38.645 8.050 39.145 48.850 ;
        RECT 39.645 8.050 40.145 48.850 ;
        RECT 40.645 45.850 44.645 48.850 ;
        RECT 40.645 41.650 44.645 44.650 ;
        RECT 40.645 37.450 44.645 40.450 ;
        RECT 40.645 33.250 44.645 36.250 ;
        RECT 40.645 29.050 44.645 32.050 ;
        RECT 40.645 24.850 44.645 27.850 ;
        RECT 40.645 20.650 44.645 23.650 ;
        RECT 40.645 16.450 44.645 19.450 ;
        RECT 40.645 12.250 44.645 15.250 ;
        RECT 40.645 8.050 44.645 11.050 ;
        RECT 45.145 8.050 45.645 48.850 ;
        RECT 46.145 8.050 46.645 48.850 ;
        RECT 47.145 45.850 51.145 48.850 ;
        RECT 47.145 41.650 51.145 44.650 ;
        RECT 47.145 37.450 51.145 40.450 ;
        RECT 47.145 33.250 51.145 36.250 ;
        RECT 47.145 29.050 51.145 32.050 ;
        RECT 47.145 24.850 51.145 27.850 ;
        RECT 47.145 20.650 51.145 23.650 ;
        RECT 47.145 16.450 51.145 19.450 ;
        RECT 47.145 12.250 51.145 15.250 ;
        RECT 47.145 8.050 51.145 11.050 ;
        RECT 51.645 8.050 52.145 48.850 ;
        RECT 52.645 8.050 53.145 48.850 ;
        RECT 53.645 45.850 57.645 48.850 ;
        RECT 53.645 41.650 57.645 44.650 ;
        RECT 53.645 37.450 57.645 40.450 ;
        RECT 53.645 33.250 57.645 36.250 ;
        RECT 53.645 29.050 57.645 32.050 ;
        RECT 53.645 24.850 57.645 27.850 ;
        RECT 53.645 20.650 57.645 23.650 ;
        RECT 53.645 16.450 57.645 19.450 ;
        RECT 53.645 12.250 57.645 15.250 ;
        RECT 53.645 8.050 57.645 11.050 ;
        RECT 58.145 8.050 58.645 48.850 ;
        RECT 59.145 8.050 59.645 48.850 ;
        RECT 60.145 45.850 64.145 48.850 ;
        RECT 60.145 41.650 64.145 44.650 ;
        RECT 60.145 37.450 64.145 40.450 ;
        RECT 60.145 33.250 64.145 36.250 ;
        RECT 60.145 29.050 64.145 32.050 ;
        RECT 60.145 24.850 64.145 27.850 ;
        RECT 60.145 20.650 64.145 23.650 ;
        RECT 60.145 16.450 64.145 19.450 ;
        RECT 60.145 12.250 64.145 15.250 ;
        RECT 60.145 8.050 64.145 11.050 ;
        RECT 64.645 8.050 65.145 48.850 ;
        RECT 65.645 8.050 66.145 48.850 ;
        RECT 66.645 45.850 70.645 48.850 ;
        RECT 66.645 41.650 70.645 44.650 ;
        RECT 66.645 37.450 70.645 40.450 ;
        RECT 66.645 33.250 70.645 36.250 ;
        RECT 66.645 29.050 70.645 32.050 ;
        RECT 66.645 24.850 70.645 27.850 ;
        RECT 66.645 20.650 70.645 23.650 ;
        RECT 66.645 16.450 70.645 19.450 ;
        RECT 66.645 12.250 70.645 15.250 ;
        RECT 66.645 8.050 70.645 11.050 ;
        RECT 71.145 8.050 71.645 48.850 ;
        RECT 72.145 8.050 72.645 48.850 ;
        RECT 73.145 45.850 77.145 48.850 ;
        RECT 73.145 41.650 77.145 44.650 ;
        RECT 73.145 37.450 77.145 40.450 ;
        RECT 73.145 33.250 77.145 36.250 ;
        RECT 73.145 29.050 77.145 32.050 ;
        RECT 73.145 24.850 77.145 27.850 ;
        RECT 73.145 20.650 77.145 23.650 ;
        RECT 73.145 16.450 77.145 19.450 ;
        RECT 73.145 12.250 77.145 15.250 ;
        RECT 73.145 8.050 77.145 11.050 ;
        RECT 77.645 8.050 78.145 48.850 ;
        RECT 78.645 8.050 79.145 48.850 ;
        RECT 79.645 45.850 83.645 48.850 ;
        RECT 79.645 41.650 83.645 44.650 ;
        RECT 79.645 37.450 83.645 40.450 ;
        RECT 79.645 33.250 83.645 36.250 ;
        RECT 79.645 29.050 83.645 32.050 ;
        RECT 79.645 24.850 83.645 27.850 ;
        RECT 79.645 20.650 83.645 23.650 ;
        RECT 79.645 16.450 83.645 19.450 ;
        RECT 79.645 12.250 83.645 15.250 ;
        RECT 79.645 8.050 83.645 11.050 ;
        RECT 84.145 8.050 84.645 48.850 ;
        RECT 85.145 8.050 85.645 48.850 ;
        RECT 86.145 45.850 90.145 48.850 ;
        RECT 86.145 41.650 90.145 44.650 ;
        RECT 86.145 37.450 90.145 40.450 ;
        RECT 86.145 33.250 90.145 36.250 ;
        RECT 86.145 29.050 90.145 32.050 ;
        RECT 86.145 24.850 90.145 27.850 ;
        RECT 86.145 20.650 90.145 23.650 ;
        RECT 86.145 16.450 90.145 19.450 ;
        RECT 86.145 12.250 90.145 15.250 ;
        RECT 86.145 8.050 90.145 11.050 ;
        RECT 90.645 8.050 91.145 48.850 ;
        RECT 91.645 8.050 92.145 48.850 ;
        RECT 92.645 45.850 96.645 48.850 ;
        RECT 92.645 41.650 96.645 44.650 ;
        RECT 92.645 37.450 96.645 40.450 ;
        RECT 92.645 33.250 96.645 36.250 ;
        RECT 92.645 29.050 96.645 32.050 ;
        RECT 92.645 24.850 96.645 27.850 ;
        RECT 92.645 20.650 96.645 23.650 ;
        RECT 92.645 16.450 96.645 19.450 ;
        RECT 92.645 12.250 96.645 15.250 ;
        RECT 92.645 8.050 96.645 11.050 ;
        RECT 97.145 8.050 97.645 48.850 ;
        RECT 98.145 8.050 98.645 48.850 ;
        RECT 99.145 45.850 103.145 48.850 ;
        RECT 99.145 41.650 103.145 44.650 ;
        RECT 99.145 37.450 103.145 40.450 ;
        RECT 99.145 33.250 103.145 36.250 ;
        RECT 99.145 29.050 103.145 32.050 ;
        RECT 99.145 24.850 103.145 27.850 ;
        RECT 99.145 20.650 103.145 23.650 ;
        RECT 99.145 16.450 103.145 19.450 ;
        RECT 99.145 12.250 103.145 15.250 ;
        RECT 99.145 8.050 103.145 11.050 ;
        RECT 103.645 8.050 104.145 48.850 ;
        RECT 104.645 35.150 105.145 48.850 ;
        RECT 105.645 45.850 109.645 48.850 ;
        RECT 105.645 41.650 109.645 44.650 ;
        RECT 105.645 37.450 109.645 40.450 ;
        RECT 104.495 34.350 105.145 35.150 ;
        RECT 104.645 22.550 105.145 34.350 ;
        RECT 105.645 33.250 109.645 36.250 ;
        RECT 105.645 29.050 109.645 32.050 ;
        RECT 110.145 30.950 110.645 48.850 ;
        RECT 110.145 30.150 110.795 30.950 ;
        RECT 105.645 24.850 109.645 27.850 ;
        RECT 104.495 21.750 105.145 22.550 ;
        RECT 104.645 6.690 105.145 21.750 ;
        RECT 105.645 20.650 109.645 23.650 ;
        RECT 105.645 16.450 109.645 19.450 ;
        RECT 105.645 12.250 109.645 15.250 ;
        RECT 105.645 8.050 109.645 11.050 ;
        RECT 110.145 7.490 110.645 30.150 ;
        RECT 111.145 26.750 111.645 48.850 ;
        RECT 112.145 45.850 116.145 48.850 ;
        RECT 112.145 41.650 116.145 44.650 ;
        RECT 112.145 37.450 116.145 40.450 ;
        RECT 112.145 33.250 116.145 36.250 ;
        RECT 116.645 35.150 117.145 48.850 ;
        RECT 116.645 34.350 117.295 35.150 ;
        RECT 112.145 29.050 116.145 32.050 ;
        RECT 110.995 25.950 111.645 26.750 ;
        RECT 108.145 7.090 110.645 7.490 ;
        RECT 111.145 7.490 111.645 25.950 ;
        RECT 112.145 24.850 116.145 27.850 ;
        RECT 112.145 20.650 116.145 23.650 ;
        RECT 116.645 22.550 117.145 34.350 ;
        RECT 116.645 21.750 117.295 22.550 ;
        RECT 112.145 16.450 116.145 19.450 ;
        RECT 112.145 12.250 116.145 15.250 ;
        RECT 112.145 8.050 116.145 11.050 ;
        RECT 111.145 7.090 113.645 7.490 ;
        RECT 116.645 6.690 117.145 21.750 ;
        RECT 117.645 8.050 118.145 48.850 ;
        RECT 118.645 45.850 122.645 48.850 ;
        RECT 118.645 41.650 122.645 44.650 ;
        RECT 118.645 37.450 122.645 40.450 ;
        RECT 118.645 33.250 122.645 36.250 ;
        RECT 118.645 29.050 122.645 32.050 ;
        RECT 118.645 24.850 122.645 27.850 ;
        RECT 118.645 20.650 122.645 23.650 ;
        RECT 118.645 16.450 122.645 19.450 ;
        RECT 118.645 12.250 122.645 15.250 ;
        RECT 118.645 8.050 122.645 11.050 ;
        RECT 123.145 8.050 123.645 48.850 ;
        RECT 124.145 8.050 124.645 48.850 ;
        RECT 125.145 45.850 129.145 48.850 ;
        RECT 125.145 41.650 129.145 44.650 ;
        RECT 125.145 37.450 129.145 40.450 ;
        RECT 125.145 33.250 129.145 36.250 ;
        RECT 125.145 29.050 129.145 32.050 ;
        RECT 125.145 24.850 129.145 27.850 ;
        RECT 125.145 20.650 129.145 23.650 ;
        RECT 125.145 16.450 129.145 19.450 ;
        RECT 125.145 12.250 129.145 15.250 ;
        RECT 125.145 8.050 129.145 11.050 ;
        RECT 129.645 8.050 130.145 48.850 ;
        RECT 130.645 8.050 131.145 48.850 ;
        RECT 131.645 45.850 135.645 48.850 ;
        RECT 131.645 41.650 135.645 44.650 ;
        RECT 131.645 37.450 135.645 40.450 ;
        RECT 131.645 33.250 135.645 36.250 ;
        RECT 131.645 29.050 135.645 32.050 ;
        RECT 131.645 24.850 135.645 27.850 ;
        RECT 131.645 20.650 135.645 23.650 ;
        RECT 131.645 16.450 135.645 19.450 ;
        RECT 131.645 12.250 135.645 15.250 ;
        RECT 131.645 8.050 135.645 11.050 ;
        RECT 136.145 8.050 136.645 48.850 ;
        RECT 137.145 8.050 137.645 48.850 ;
        RECT 138.145 45.850 142.145 48.850 ;
        RECT 138.145 41.650 142.145 44.650 ;
        RECT 138.145 37.450 142.145 40.450 ;
        RECT 138.145 33.250 142.145 36.250 ;
        RECT 138.145 29.050 142.145 32.050 ;
        RECT 138.145 24.850 142.145 27.850 ;
        RECT 138.145 20.650 142.145 23.650 ;
        RECT 138.145 16.450 142.145 19.450 ;
        RECT 138.145 12.250 142.145 15.250 ;
        RECT 138.145 8.050 142.145 11.050 ;
        RECT 142.645 8.050 143.145 48.850 ;
        RECT 143.645 8.050 144.145 48.850 ;
        RECT 144.645 45.850 148.645 48.850 ;
        RECT 144.645 41.650 148.645 44.650 ;
        RECT 144.645 37.450 148.645 40.450 ;
        RECT 144.645 33.250 148.645 36.250 ;
        RECT 144.645 29.050 148.645 32.050 ;
        RECT 144.645 24.850 148.645 27.850 ;
        RECT 144.645 20.650 148.645 23.650 ;
        RECT 144.645 16.450 148.645 19.450 ;
        RECT 144.645 12.250 148.645 15.250 ;
        RECT 144.645 8.050 148.645 11.050 ;
        RECT 149.145 8.050 149.645 48.850 ;
        RECT 150.145 8.050 150.645 48.850 ;
        RECT 151.145 45.850 155.145 48.850 ;
        RECT 151.145 41.650 155.145 44.650 ;
        RECT 151.145 37.450 155.145 40.450 ;
        RECT 151.145 33.250 155.145 36.250 ;
        RECT 151.145 29.050 155.145 32.050 ;
        RECT 151.145 24.850 155.145 27.850 ;
        RECT 151.145 20.650 155.145 23.650 ;
        RECT 151.145 16.450 155.145 19.450 ;
        RECT 151.145 12.250 155.145 15.250 ;
        RECT 151.145 8.050 155.145 11.050 ;
        RECT 155.645 8.050 156.145 48.850 ;
        RECT 156.645 8.050 157.145 48.850 ;
        RECT 157.645 45.850 161.645 48.850 ;
        RECT 157.645 41.650 161.645 44.650 ;
        RECT 157.645 37.450 161.645 40.450 ;
        RECT 157.645 33.250 161.645 36.250 ;
        RECT 157.645 29.050 161.645 32.050 ;
        RECT 157.645 24.850 161.645 27.850 ;
        RECT 157.645 20.650 161.645 23.650 ;
        RECT 157.645 16.450 161.645 19.450 ;
        RECT 157.645 12.250 161.645 15.250 ;
        RECT 157.645 8.050 161.645 11.050 ;
        RECT 162.145 8.050 162.645 48.850 ;
        RECT 163.145 8.050 163.645 48.850 ;
        RECT 164.145 45.850 168.145 48.850 ;
        RECT 164.145 41.650 168.145 44.650 ;
        RECT 164.145 37.450 168.145 40.450 ;
        RECT 164.145 33.250 168.145 36.250 ;
        RECT 164.145 29.050 168.145 32.050 ;
        RECT 164.145 24.850 168.145 27.850 ;
        RECT 164.145 20.650 168.145 23.650 ;
        RECT 164.145 16.450 168.145 19.450 ;
        RECT 164.145 12.250 168.145 15.250 ;
        RECT 164.145 8.050 168.145 11.050 ;
        RECT 168.645 8.050 169.145 48.850 ;
        RECT 169.645 8.050 170.145 48.850 ;
        RECT 170.645 45.850 174.645 48.850 ;
        RECT 170.645 41.650 174.645 44.650 ;
        RECT 170.645 37.450 174.645 40.450 ;
        RECT 170.645 33.250 174.645 36.250 ;
        RECT 170.645 29.050 174.645 32.050 ;
        RECT 170.645 24.850 174.645 27.850 ;
        RECT 170.645 20.650 174.645 23.650 ;
        RECT 170.645 16.450 174.645 19.450 ;
        RECT 170.645 12.250 174.645 15.250 ;
        RECT 170.645 8.050 174.645 11.050 ;
        RECT 175.145 8.050 175.645 48.850 ;
        RECT 176.145 8.050 176.645 48.850 ;
        RECT 177.145 45.850 181.145 48.850 ;
        RECT 177.145 41.650 181.145 44.650 ;
        RECT 177.145 37.450 181.145 40.450 ;
        RECT 177.145 33.250 181.145 36.250 ;
        RECT 177.145 29.050 181.145 32.050 ;
        RECT 177.145 24.850 181.145 27.850 ;
        RECT 177.145 20.650 181.145 23.650 ;
        RECT 177.145 16.450 181.145 19.450 ;
        RECT 177.145 12.250 181.145 15.250 ;
        RECT 177.145 8.050 181.145 11.050 ;
        RECT 181.645 8.050 182.145 48.850 ;
        RECT 182.645 8.050 183.145 48.850 ;
        RECT 183.645 45.850 187.645 48.850 ;
        RECT 183.645 41.650 187.645 44.650 ;
        RECT 183.645 37.450 187.645 40.450 ;
        RECT 183.645 33.250 187.645 36.250 ;
        RECT 183.645 29.050 187.645 32.050 ;
        RECT 183.645 24.850 187.645 27.850 ;
        RECT 183.645 20.650 187.645 23.650 ;
        RECT 183.645 16.450 187.645 19.450 ;
        RECT 183.645 12.250 187.645 15.250 ;
        RECT 183.645 8.050 187.645 11.050 ;
        RECT 188.145 8.050 188.645 48.850 ;
        RECT 189.145 8.050 189.645 48.850 ;
        RECT 190.145 45.850 194.145 48.850 ;
        RECT 190.145 41.650 194.145 44.650 ;
        RECT 190.145 37.450 194.145 40.450 ;
        RECT 190.145 33.250 194.145 36.250 ;
        RECT 190.145 29.050 194.145 32.050 ;
        RECT 190.145 24.850 194.145 27.850 ;
        RECT 190.145 20.650 194.145 23.650 ;
        RECT 190.145 16.450 194.145 19.450 ;
        RECT 190.145 12.250 194.145 15.250 ;
        RECT 190.145 8.050 194.145 11.050 ;
        RECT 194.645 8.050 195.145 48.850 ;
        RECT 195.645 8.050 196.145 48.850 ;
        RECT 196.645 45.850 200.645 48.850 ;
        RECT 196.645 41.650 200.645 44.650 ;
        RECT 196.645 37.450 200.645 40.450 ;
        RECT 196.645 33.250 200.645 36.250 ;
        RECT 196.645 29.050 200.645 32.050 ;
        RECT 196.645 24.850 200.645 27.850 ;
        RECT 196.645 20.650 200.645 23.650 ;
        RECT 196.645 16.450 200.645 19.450 ;
        RECT 196.645 12.250 200.645 15.250 ;
        RECT 196.645 8.050 200.645 11.050 ;
        RECT 201.145 8.050 201.645 48.850 ;
        RECT 202.145 8.050 202.645 48.850 ;
        RECT 203.145 45.850 207.145 48.850 ;
        RECT 203.145 41.650 207.145 44.650 ;
        RECT 203.145 37.450 207.145 40.450 ;
        RECT 203.145 33.250 207.145 36.250 ;
        RECT 203.145 29.050 207.145 32.050 ;
        RECT 203.145 24.850 207.145 27.850 ;
        RECT 203.145 20.650 207.145 23.650 ;
        RECT 203.145 16.450 207.145 19.450 ;
        RECT 203.145 12.250 207.145 15.250 ;
        RECT 203.145 8.050 207.145 11.050 ;
        RECT 207.645 8.050 208.145 48.850 ;
        RECT 208.645 8.050 209.145 48.850 ;
        RECT 209.645 45.850 213.645 48.850 ;
        RECT 209.645 41.650 213.645 44.650 ;
        RECT 209.645 37.450 213.645 40.450 ;
        RECT 209.645 33.250 213.645 36.250 ;
        RECT 209.645 29.050 213.645 32.050 ;
        RECT 209.645 24.850 213.645 27.850 ;
        RECT 209.645 20.650 213.645 23.650 ;
        RECT 209.645 16.450 213.645 19.450 ;
        RECT 209.645 12.250 213.645 15.250 ;
        RECT 209.645 8.050 213.645 11.050 ;
        RECT 214.145 8.050 214.645 48.850 ;
        RECT 215.145 8.050 215.645 48.850 ;
        RECT 216.145 45.850 220.145 48.850 ;
        RECT 216.145 41.650 220.145 44.650 ;
        RECT 216.145 37.450 220.145 40.450 ;
        RECT 216.145 33.250 220.145 36.250 ;
        RECT 216.145 29.050 220.145 32.050 ;
        RECT 216.145 24.850 220.145 27.850 ;
        RECT 216.145 20.650 220.145 23.650 ;
        RECT 216.145 16.450 220.145 19.450 ;
        RECT 216.145 12.250 220.145 15.250 ;
        RECT 216.145 8.050 220.145 11.050 ;
        RECT 0.270 6.290 117.145 6.690 ;
        RECT -0.430 5.490 116.645 5.890 ;
        RECT -1.130 4.690 123.145 5.090 ;
        RECT -1.830 3.890 168.645 4.290 ;
        RECT -2.530 3.090 207.645 3.490 ;
        RECT -3.230 2.290 214.145 2.690 ;
        RECT -3.930 1.490 111.145 1.890 ;
        RECT -4.630 0.690 108.645 1.090 ;
        RECT -5.330 -0.110 113.645 0.290 ;
  END
END DAC
END LIBRARY

