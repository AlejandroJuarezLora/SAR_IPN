* SPICE3 file created from sw_top_flat.ext - technology: sky130B

.subckt sw_top out en in vss vdd
X0 out.t19 en_buf in.t17 vdd.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 out.t9 net1 in.t2 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 out.t8 net1 in.t6 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 vdd.t20 vss.t32 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4 vdd.t27 en.t0 en_buf vdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 net1 en_buf vss.t17 vss.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 in.t11 en_buf out.t18 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 vdd.t23 vss.t33 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8 in.t5 net1 out.t7 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 vdd.t29 en.t1 en_buf vdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 out.t17 en_buf in.t13 vdd.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X11 en_buf en.t2 vss.t31 vss.t30 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 net1 en_buf vss.t15 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 out.t16 en_buf in.t18 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X14 net1 en_buf vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 in.t19 en_buf out.t15 vdd.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X16 en_buf en.t3 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 net1 en_buf vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 in.t3 net1 out.t6 vss.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X19 in.t7 net1 out.t5 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X20 vss.t23 vdd.t32 vss.t22 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X21 in.t4 net1 out.t4 vss.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X22 vss.t13 en_buf net1 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 out.t14 en_buf in.t14 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X24 en_buf en.t4 vss.t25 vss.t24 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 vss.t20 vdd.t33 vss.t19 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X26 out.t3 net1 in.t9 vss.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X27 out.t2 net1 in.t0 vss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X28 out.t1 net1 in.t1 vss.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X29 vss.t11 en_buf net1 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 in.t10 en_buf out.t13 vdd.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X31 in.t8 net1 out.t0 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X32 in.t12 en_buf out.t12 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X33 en_buf en.t5 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 vdd.t5 en_buf net1 vdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X35 vss.t29 en.t6 en_buf vss.t28 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 in.t15 en_buf out.t11 vdd.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X37 vss.t27 en.t7 en_buf vss.t26 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X38 out.t10 en_buf in.t16 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X39 vdd.t1 en_buf net1 vdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 in.n8 in.t12 29.3118
R1 in.n13 in.t13 29.3084
R2 in.n6 in.t16 28.5655
R3 in.n6 in.t10 28.5655
R4 in.n4 in.t17 28.5655
R5 in.n4 in.t11 28.5655
R6 in.n2 in.t18 28.5655
R7 in.n2 in.t19 28.5655
R8 in.n0 in.t14 28.5655
R9 in.n0 in.t15 28.5655
R10 in.n8 in.t7 18.1397
R11 in.n13 in.t9 18.1397
R12 in.n7 in.t0 17.4005
R13 in.n7 in.t3 17.4005
R14 in.n5 in.t1 17.4005
R15 in.n5 in.t8 17.4005
R16 in.n3 in.t2 17.4005
R17 in.n3 in.t5 17.4005
R18 in.n1 in.t6 17.4005
R19 in.n1 in.t4 17.4005
R20 in.n10 in.n9 0.811311
R21 in.n12 in.n11 0.799575
R22 in.n11 in.n10 0.794419
R23 in.n9 in.n8 0.787662
R24 in.n13 in.n12 0.773526
R25 in.n9 in.n6 0.746823
R26 in.n10 in.n4 0.746823
R27 in.n11 in.n2 0.746823
R28 in.n12 in.n0 0.743351
R29 in.n9 in.n7 0.739748
R30 in.n10 in.n5 0.739748
R31 in.n11 in.n3 0.739748
R32 in.n12 in.n1 0.739748
R33 in in.n13 0.636099
R34 out out.n14 105.326
R35 out.n11 out.n10 86.3387
R36 out.n14 out.n13 85.9532
R37 out.n10 out.n8 84.93
R38 out.n12 out.n4 83.8601
R39 out.n14 out.n0 83.6607
R40 out.n13 out.n2 83.2397
R41 out.n11 out.n6 83.0069
R42 out.n14 out.n1 81.7128
R43 out.n13 out.n3 81.5763
R44 out.n12 out.n5 81.3057
R45 out.n13 out.n12 81.2978
R46 out.n12 out.n11 80.9519
R47 out.n11 out.n7 80.2068
R48 out.n10 out.n9 80.0412
R49 out.n8 out.t11 28.5655
R50 out.n8 out.t17 28.5655
R51 out.n2 out.t13 28.5655
R52 out.n2 out.t19 28.5655
R53 out.n4 out.t18 28.5655
R54 out.n4 out.t16 28.5655
R55 out.n6 out.t15 28.5655
R56 out.n6 out.t14 28.5655
R57 out.n0 out.t12 28.5655
R58 out.n0 out.t10 28.5655
R59 out.n9 out.t4 17.4005
R60 out.n9 out.t3 17.4005
R61 out.n3 out.t6 17.4005
R62 out.n3 out.t1 17.4005
R63 out.n5 out.t0 17.4005
R64 out.n5 out.t9 17.4005
R65 out.n7 out.t7 17.4005
R66 out.n7 out.t8 17.4005
R67 out.n1 out.t5 17.4005
R68 out.n1 out.t2 17.4005
R69 vdd.n41 vdd.n36 6225.88
R70 vdd.n38 vdd.n36 3240
R71 vdd.n39 vdd.n38 3007.06
R72 vdd.t18 vdd 895.586
R73 vdd.n7 vdd.t5 584.644
R74 vdd.n18 vdd.t27 584.644
R75 vdd.n29 vdd.t19 459.192
R76 vdd.n47 vdd 420.262
R77 vdd.t4 vdd 301.551
R78 vdd.t6 vdd.n36 289.37
R79 vdd.n40 vdd.t15 289.349
R80 vdd.t26 vdd 285.68
R81 vdd vdd.t21 247.137
R82 vdd.n48 vdd.t20 243.03
R83 vdd.n49 vdd.n47 237.554
R84 vdd.n0 vdd.t22 234.554
R85 vdd.n3 vdd.t23 234.554
R86 vdd.t2 vdd.t6 197.359
R87 vdd.t7 vdd.t2 197.359
R88 vdd.t17 vdd.t7 197.359
R89 vdd.t16 vdd.t17 197.359
R90 vdd.t14 vdd.t11 197.359
R91 vdd.t11 vdd.t8 197.359
R92 vdd.t8 vdd.t3 197.359
R93 vdd.t3 vdd.t15 197.359
R94 vdd.n47 vdd.t18 192.569
R95 vdd.t9 vdd.t4 190.453
R96 vdd.t0 vdd.t9 190.453
R97 vdd.t12 vdd.t0 190.453
R98 vdd.t30 vdd.t26 190.453
R99 vdd.t28 vdd.t30 190.453
R100 vdd.t24 vdd.t28 190.453
R101 vdd.n12 vdd.n11 174.595
R102 vdd.n23 vdd.n22 174.595
R103 vdd vdd.t12 170.048
R104 vdd vdd.t24 170.048
R105 vdd.n1 vdd.t33 166.282
R106 vdd.n17 vdd.t13 151.123
R107 vdd.n28 vdd.t25 151.123
R108 vdd.n37 vdd.t16 98.6801
R109 vdd.n37 vdd.t14 98.6801
R110 vdd.n29 vdd.t32 92.9047
R111 vdd.n11 vdd.t10 26.5955
R112 vdd.n11 vdd.t1 26.5955
R113 vdd.n22 vdd.t31 26.5955
R114 vdd.n22 vdd.t29 26.5955
R115 vdd.n39 vdd.n34 22.4361
R116 vdd.n7 vdd.n6 21.8029
R117 vdd.n42 vdd.n41 21.2145
R118 vdd.n18 vdd.n17 21.0829
R119 vdd.n33 vdd.n28 15.4358
R120 vdd.n42 vdd.n35 14.5834
R121 vdd.n44 vdd.n43 4.74226
R122 vdd.n28 vdd.n27 4.6505
R123 vdd.n19 vdd.n18 4.6505
R124 vdd.n17 vdd.n16 4.6505
R125 vdd.n8 vdd.n7 4.6505
R126 vdd.n6 vdd.n5 4.6505
R127 vdd.n51 vdd.n50 4.6505
R128 vdd.n26 vdd.n25 4.6505
R129 vdd.n24 vdd.n23 4.6505
R130 vdd.n21 vdd.n20 4.6505
R131 vdd.n15 vdd.n14 4.6505
R132 vdd.n13 vdd.n12 4.6505
R133 vdd.n10 vdd.n9 4.6505
R134 vdd.n3 vdd.n2 4.36875
R135 vdd.n2 vdd.n1 3.50526
R136 vdd.n45 vdd.n44 3.23979
R137 vdd.n49 vdd.n48 3.08362
R138 vdd.n31 vdd.n29 2.61352
R139 vdd.n31 vdd.n30 2.29594
R140 vdd.n43 vdd.n34 2.19925
R141 vdd.n33 vdd.n32 1.84013
R142 vdd.n53 vdd.n33 1.09272
R143 vdd.n1 vdd.n0 0.863992
R144 vdd.n43 vdd.n42 0.847933
R145 vdd.n32 vdd.n31 0.79957
R146 vdd.n44 vdd 0.700957
R147 vdd.n50 vdd.n49 0.467369
R148 vdd.n6 vdd.n3 0.305262
R149 vdd.n53 vdd.n52 0.294492
R150 vdd vdd.n53 0.234
R151 vdd.n51 vdd.n46 0.179926
R152 vdd.n41 vdd.n40 0.134074
R153 vdd.n5 vdd.n4 0.120292
R154 vdd.n10 vdd.n8 0.120292
R155 vdd.n13 vdd.n10 0.120292
R156 vdd.n15 vdd.n13 0.120292
R157 vdd.n16 vdd.n15 0.120292
R158 vdd.n21 vdd.n19 0.120292
R159 vdd.n24 vdd.n21 0.120292
R160 vdd.n26 vdd.n24 0.120292
R161 vdd.n27 vdd.n26 0.120292
R162 vdd.n52 vdd.n51 0.120292
R163 vdd.n40 vdd.n39 0.11303
R164 vdd.n46 vdd 0.0822696
R165 vdd.n35 vdd.n34 0.0671871
R166 vdd.n8 vdd 0.0603958
R167 vdd.n19 vdd 0.0512812
R168 vdd.n45 vdd 0.0433571
R169 vdd.n5 vdd 0.0226354
R170 vdd.n16 vdd 0.0226354
R171 vdd vdd.n27 0.0226354
R172 vdd.n45 vdd 0.0226354
R173 vdd vdd.n45 0.016125
R174 vdd.n40 vdd.n35 0.0135311
R175 vdd.n38 vdd.n37 0.00492753
R176 vss.n0 vss.t18 59385
R177 vss.n3 vss.n1 5290.03
R178 vss.n4 vss.n3 4820.71
R179 vss vss.t21 4659.52
R180 vss.t21 vss 3998.93
R181 vss vss.t12 1568.9
R182 vss vss.t28 1486.33
R183 vss.n11 vss.t5 1345.97
R184 vss.t18 vss 1285.79
R185 vss.t12 vss.t14 990.885
R186 vss.t14 vss.t10 990.885
R187 vss.t10 vss.t16 990.885
R188 vss.t28 vss.t30 990.885
R189 vss.t30 vss.t26 990.885
R190 vss.t26 vss.t24 990.885
R191 vss.t5 vss.t2 928.802
R192 vss.t2 vss.t6 928.802
R193 vss.t6 vss.t1 928.802
R194 vss.t1 vss.t0 928.802
R195 vss.t9 vss.t7 928.802
R196 vss.t7 vss.t8 928.802
R197 vss.t8 vss.t4 928.802
R198 vss.t4 vss.t3 928.802
R199 vss.t16 vss 884.72
R200 vss.t24 vss 884.72
R201 vss.n2 vss.t9 464.401
R202 vss.n23 vss.t25 193.933
R203 vss.n54 vss.t17 193.933
R204 vss.n20 vss.t29 192.982
R205 vss.n60 vss.t13 192.982
R206 vss.n63 vss.t33 183.082
R207 vss.n33 vss.n32 124.692
R208 vss.n62 vss.t20 121.956
R209 vss.n15 vss.t19 121.956
R210 vss.n43 vss.t22 121.956
R211 vss.n31 vss.t23 121.956
R212 vss.n6 vss.n0 118.069
R213 vss.n49 vss.n22 114.713
R214 vss.n56 vss.n19 114.713
R215 vss.n36 vss.n27 114.398
R216 vss.n34 vss.n33 76.0005
R217 vss.n50 vss.n49 34.6358
R218 vss.n49 vss.n48 34.6358
R219 vss.n56 vss.n17 34.6358
R220 vss.n56 vss.n55 34.6358
R221 vss.n27 vss.t32 34.2973
R222 vss.n22 vss.t31 24.9236
R223 vss.n22 vss.t27 24.9236
R224 vss.n19 vss.t15 24.9236
R225 vss.n19 vss.t11 24.9236
R226 vss.n50 vss.n20 22.2123
R227 vss.n48 vss.n23 22.2123
R228 vss.n60 vss.n17 22.2123
R229 vss.n55 vss.n54 22.2123
R230 vss.n61 vss.n60 19.3355
R231 vss.n54 vss.n20 18.0711
R232 vss.n44 vss.n23 17.4103
R233 vss.n10 vss.n9 9.39653
R234 vss.n13 vss.n12 9.3005
R235 vss.n12 vss.n11 9.3005
R236 vss.n42 vss.n41 6.26433
R237 vss.n41 vss.n25 6.26433
R238 vss.n64 vss.n15 5.98311
R239 vss.n43 vss.n42 5.85582
R240 vss.n37 vss.n25 5.65809
R241 vss.n66 vss.n15 5.06789
R242 vss.n31 vss.n30 4.91351
R243 vss.n33 vss.n27 4.85762
R244 vss.n64 vss.n63 4.8005
R245 vss.n60 vss.n59 4.6505
R246 vss.n54 vss.n53 4.6505
R247 vss.n52 vss.n20 4.6505
R248 vss.n46 vss.n23 4.6505
R249 vss.n65 vss.n64 4.6505
R250 vss.n61 vss.n16 4.6505
R251 vss.n58 vss.n17 4.6505
R252 vss.n57 vss.n56 4.6505
R253 vss.n55 vss.n18 4.6505
R254 vss.n51 vss.n50 4.6505
R255 vss.n49 vss.n21 4.6505
R256 vss.n48 vss.n47 4.6505
R257 vss.n45 vss.n44 4.6505
R258 vss.n42 vss.n24 4.6505
R259 vss.n41 vss.n40 4.6505
R260 vss.n39 vss.n25 4.6505
R261 vss.n38 vss.n37 4.6505
R262 vss.n35 vss.n26 4.6505
R263 vss.n29 vss.n28 4.6505
R264 vss.n14 vss.n13 3.90461
R265 vss.n10 vss.n8 3.77398
R266 vss.n36 vss.n35 3.50735
R267 vss.n67 vss.n14 3.21121
R268 vss.n34 vss.n28 3.2005
R269 vss.n32 vss.n31 2.63064
R270 vss.n63 vss.n62 1.18311
R271 vss.n32 vss.n28 1.14023
R272 vss.n35 vss.n34 0.833377
R273 vss.n13 vss.n10 0.753441
R274 vss.n6 vss.n4 0.67602
R275 vss.n37 vss.n36 0.526527
R276 vss.n62 vss.n61 0.417891
R277 vss.n44 vss.n43 0.409011
R278 vss.n14 vss 0.314344
R279 vss.n6 vss.n5 0.288252
R280 vss vss.n66 0.19611
R281 vss.n7 vss.n6 0.134398
R282 vss.n8 vss.n7 0.12657
R283 vss vss.n67 0.1255
R284 vss.n66 vss.n65 0.120292
R285 vss.n65 vss.n16 0.120292
R286 vss.n59 vss.n58 0.120292
R287 vss.n58 vss.n57 0.120292
R288 vss.n57 vss.n18 0.120292
R289 vss.n53 vss.n18 0.120292
R290 vss.n52 vss.n51 0.120292
R291 vss.n51 vss.n21 0.120292
R292 vss.n47 vss.n21 0.120292
R293 vss.n47 vss.n46 0.120292
R294 vss.n45 vss.n24 0.120292
R295 vss.n40 vss.n24 0.120292
R296 vss.n40 vss.n39 0.120292
R297 vss.n39 vss.n38 0.120292
R298 vss.n38 vss.n26 0.120292
R299 vss.n29 vss.n26 0.120292
R300 vss.n30 vss.n29 0.120292
R301 vss.n67 vss 0.0612143
R302 vss.n59 vss 0.0603958
R303 vss vss.n45 0.0577917
R304 vss vss.n52 0.0512812
R305 vss vss.n16 0.0226354
R306 vss.n53 vss 0.0226354
R307 vss.n46 vss 0.0226354
R308 vss.n30 vss 0.0226354
R309 vss.n3 vss.n2 0.0145006
R310 en.n5 en.t0 212.081
R311 en.n7 en.t3 212.081
R312 en.n4 en.t1 212.081
R313 en.n12 en.t5 212.081
R314 en.n5 en.t6 139.78
R315 en.n7 en.t2 139.78
R316 en.n4 en.t7 139.78
R317 en.n12 en.t4 139.78
R318 en.n6 en 78.3045
R319 en.n9 en.n8 76.0005
R320 en.n11 en.n10 76.0005
R321 en.n13 en.n12 44.8017
R322 en.n6 en.n5 30.6732
R323 en.n7 en.n6 30.6732
R324 en.n8 en.n7 30.6732
R325 en.n8 en.n4 30.6732
R326 en.n11 en.n4 30.6732
R327 en.n12 en.n11 30.6732
R328 en.n9 en 19.2005
R329 en.n10 en 17.1525
R330 en en.n2 12.2885
R331 en.n10 en 6.4005
R332 en.n14 en.n2 4.6085
R333 en.n13 en.n3 4.6085
R334 en en.n9 4.3525
R335 en.n3 en 1.7925
R336 en.n19 en 0.973061
R337 en en.n19 0.767327
R338 en.n14 en.n13 0.2565
R339 en.n19 en.n18 0.0775814
R340 en.n17 en.n1 0.0437692
R341 en.n16 en.n15 0.0437692
R342 en.n17 en.n16 0.00290385
R343 en.n18 en.n17 0.00166462
R344 en.n17 en.n14 0.0011688
R345 en.n18 en.n0 0.00100408
C0 en en_buf 0.408f
C1 vdd in 0.471f
C2 out in 2.37f
C3 en net1 0.0114f
C4 vdd en 0.33f
C5 out en 3.88e-19
C6 en_buf net1 0.636f
C7 vdd en_buf 1.84f
C8 out en_buf 0.373f
C9 vdd net1 0.828f
C10 out net1 0.336f
C11 vdd out 0.305f
C12 in en 0.00149f
C13 in en_buf 0.412f
C14 in net1 0.377f
C15 en vss 0.639f
C16 out vss 0.475f
C17 in vss 0.581f
C18 vdd vss 9.34f
C19 net1 vss 1.92f
C20 en_buf vss 1.82f
C21 out.t12 vss 0.021f
C22 out.t10 vss 0.021f
C23 out.n0 vss 0.137f
C24 out.t5 vss 0.021f
C25 out.t2 vss 0.021f
C26 out.n1 vss 0.136f
C27 out.t13 vss 0.021f
C28 out.t19 vss 0.021f
C29 out.n2 vss 0.136f
C30 out.t6 vss 0.021f
C31 out.t1 vss 0.021f
C32 out.n3 vss 0.136f
C33 out.t18 vss 0.021f
C34 out.t16 vss 0.021f
C35 out.n4 vss 0.136f
C36 out.t0 vss 0.021f
C37 out.t9 vss 0.021f
C38 out.n5 vss 0.136f
C39 out.t15 vss 0.021f
C40 out.t14 vss 0.021f
C41 out.n6 vss 0.136f
C42 out.t7 vss 0.021f
C43 out.t8 vss 0.021f
C44 out.n7 vss 0.137f
C45 out.t11 vss 0.021f
C46 out.t17 vss 0.021f
C47 out.n8 vss 0.136f
C48 out.t4 vss 0.021f
C49 out.t3 vss 0.021f
C50 out.n9 vss 0.137f
C51 out.n10 vss 0.0919f
C52 out.n11 vss 0.119f
C53 out.n12 vss 0.12f
C54 out.n13 vss 0.119f
C55 out.n14 vss 0.124f
C56 in.t13 vss 0.0202f
C57 in.t9 vss 0.0223f
C58 in.t14 vss 0.0168f
C59 in.t15 vss 0.0168f
C60 in.n0 vss 0.118f
C61 in.t6 vss 0.0168f
C62 in.t4 vss 0.0168f
C63 in.n1 vss 0.118f
C64 in.t18 vss 0.0168f
C65 in.t19 vss 0.0168f
C66 in.n2 vss 0.118f
C67 in.t2 vss 0.0168f
C68 in.t5 vss 0.0168f
C69 in.n3 vss 0.118f
C70 in.t17 vss 0.0168f
C71 in.t11 vss 0.0168f
C72 in.n4 vss 0.118f
C73 in.t1 vss 0.0168f
C74 in.t8 vss 0.0168f
C75 in.n5 vss 0.118f
C76 in.t16 vss 0.0168f
C77 in.t10 vss 0.0168f
C78 in.n6 vss 0.118f
C79 in.t0 vss 0.0168f
C80 in.t3 vss 0.0168f
C81 in.n7 vss 0.118f
C82 in.t12 vss 0.0202f
C83 in.t7 vss 0.0223f
C84 in.n8 vss 0.337f
C85 in.n9 vss 0.0985f
C86 in.n10 vss 0.0987f
C87 in.n11 vss 0.0984f
C88 in.n12 vss 0.0991f
C89 in.n13 vss 0.353f
.ends

