* SPICE3 file created from sar_analog_flat.ext - technology: sky130B

.subckt sar_analog ctlp7 ctlp6 ctlp5 ctlp4 ctlp3 ctlp2 ctlp1 ctlp0 ctln7 ctln6 ctln5 ctln4 ctln3 ctln2 ctln1 ctln0     
+  trim4 trim3 trim2 trim1 trim0 trimb4 trimb3 trimb2 trimb1 trimb0 vinp vinn sample comp clkc avdd avss
X0 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 vinp.t9 dac_0.sw_top_0.en_buf comparator_0.vp.t9 avdd.t70 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X2 comparator_0.trim_0.n4.t15 trim4.t0 avss.t374 avss.t373 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 dac_1.out.t49 dac_1.sw_top_1.en_buf vinn.t48 avdd.t144 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln1.t0 avss.t294 avss.t293 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 dac_1.sw_top_0.en_buf sample.t0 avdd.t114 avdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 comparator_0.vp.t80 dac_0.carray_0.unitcap_288.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 avss.t286 trimb4.t0 comparator_0.trim_1.n4.t7 avss.t285 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X11 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 avss.t318 dac_0.sw_top_3.en_buf dac_0.sw_top_3.net1 avss.t317 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 dac_1.out dac_1.carray_0.unitcap_320.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 comparator_0.in.t3 comparator_0.trim_0.n4.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 avss.t201 trimb2.t0 comparator_0.trim_1.n2 avss.t200 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X21 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_5.Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 comparator_0.vp.t81 dac_0.carray_0.unitcap_322.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 comparator_0.vp.t77 dac_0.sw_top_1.net1 vinp.t79 avss.t358 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X27 comparator_0.vp dac_0.carray_0.unitcap_136.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 avdd.t116 sample.t1 dac_1.sw_top_3.en_buf avdd.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 dac_1.out dac_1.carray_0.unitcap_208.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 avss.t378 ctlp1.t0 dac_0.sky130_fd_sc_hd__inv_2_4.Y avss.t377 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 vinn.t25 dac_1.sw_top_0.en_buf dac_1.out.t29 avdd.t102 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X32 avdd.t10 ctln7.t0 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t3 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 comparator_0.in.t4 comparator_0.trim_0.n3.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 dac_0.sw_top_0.net1 dac_0.sw_top_0.en_buf avdd.t69 avdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 dac_1.out.t79 dac_1.sw_top_2.en_buf vinn.t76 avdd.t308 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X41 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 comparator_0.vp dac_0.carray_0.unitcap_199.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 comparator_0.vp dac_0.carray_0.unitcap_40.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 comparator_0.vp dac_0.carray_0.unitcap_31.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t2 ctlp7.t0 avdd.t156 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X49 comparator_0.outn comparator_0.outp comparator_0.in.t1 avss.t86 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X50 avss.t59 avdd.t311 avss.t58 avss.t57 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X51 vinp.t19 dac_0.sw_top_2.net1 comparator_0.vp.t13 avss.t148 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X52 comparator_0.vp.t37 dac_0.sw_top_1.en_buf vinp.t39 avdd.t182 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X53 avss.t168 ctlp2.t0 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t1 avss.t167 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X54 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 vinp.t29 dac_0.sw_top_0.net1 comparator_0.vp.t22 avss.t158 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X56 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 dac_1.out.t19 dac_1.sw_top_3.en_buf vinn.t12 avdd.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X58 avdd.t51 dac_1.sw_top_3.en_buf dac_1.sw_top_3.net1 avdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t2 ctln3.t0 avdd.t3 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t3 ctlp3.t0 avss.t176 avss.t175 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X64 dac_1.sw_top_1.en_buf sample.t2 avdd.t118 avdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 dac_1.out dac_1.carray_0.unitcap_248.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 avss.t138 dac_1.sw_top_0.en_buf dac_1.sw_top_0.net1 avss.t137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 dac_1.out.t9 dac_1.sw_top_2.net1 vinn.t9 avss.t83 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X74 comparator_0.vp dac_0.carray_0.unitcap_248.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t3 ctlp4.t0 avss.t284 avss.t283 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X76 vinn.t64 dac_1.sw_top_1.net1 dac_1.out.t69 avss.t274 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X77 dac_0.sw_top_1.en_buf sample.t3 avss.t215 avss.t214 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X78 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 dac_1.out.t39 dac_1.sw_top_0.net1 vinn.t39 avss.t211 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X80 comparator_0.vp dac_0.carray_0.unitcap_224.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 avss.t217 sample.t4 dac_0.sw_top_0.en_buf avss.t216 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X86 vinp.t8 dac_0.sw_top_0.en_buf comparator_0.vp.t8 avdd.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X87 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 dac_1.out dac_1.carray_0.unitcap_47.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 vinn.t4 dac_1.sw_top_2.net1 dac_1.out.t8 avss.t82 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X91 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 comparator_0.vp.t82 dac_0.carray_0.unitcap_337.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 comparator_0.in.t5 comparator_0.trim_0.n4.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 dac_1.out.t80 dac_1.carray_0.unitcap_14.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 vinp.t59 dac_0.sw_top_3.net1 comparator_0.vp.t52 avss.t332 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X99 avdd.t126 sample.t5 dac_0.sw_top_1.en_buf avdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X100 dac_1.sw_top_0.en_buf sample.t6 avdd.t104 avdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X101 comparator_0.in.t6 comparator_0.trim_0.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t3 ctlp2.t1 avss.t376 avss.t375 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X104 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 dac_1.out dac_1.carray_0.unitcap_223.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 dac_1.out dac_1.carray_0.unitcap_127.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 comparator_0.vp.t56 dac_0.sw_top_3.net1 vinp.t58 avss.t331 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X109 avss.t288 trimb4.t1 comparator_0.trim_1.n4.t6 avss.t287 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X110 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 comparator_0.trim_0.n4.t14 trim4.t1 avss.t372 avss.t371 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X114 comparator_0.vp dac_0.carray_0.unitcap_152.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 avss.t260 trim2.t0 comparator_0.trim_0.n2 avss.t259 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X117 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_7.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 dac_1.out.t59 dac_1.sw_top_3.net1 vinn.t56 avss.t256 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X120 vinp.t49 dac_0.sw_top_3.en_buf comparator_0.vp.t40 avdd.t257 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X121 comparator_0.vp dac_0.carray_0.unitcap_64.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 avdd.t207 avss.t409 avdd.t206 avdd.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X124 avdd.t18 clkc.t0 comparator_0.outn avdd.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X125 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 comp.t0 a_33300_5579# avss.t236 avss.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X128 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 comparator_0.vp dac_0.carray_0.unitcap_79.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 comparator_0.in.t7 comparator_0.trim_0.n3.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 a_33300_5579# comparator_0.outn avdd.t31 avdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X134 vinn.t29 dac_1.sw_top_0.en_buf dac_1.out.t28 avdd.t101 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X135 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 comparator_0.vp dac_0.carray_0.unitcap_338.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 comparator_0.vp.t30 dac_0.sw_top_1.en_buf vinp.t38 avdd.t181 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X141 dac_1.sw_top_0.net1 dac_1.sw_top_0.en_buf avss.t136 avss.t135 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 comparator_0.vp dac_0.carray_0.unitcap_159.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 avdd.t49 dac_1.sw_top_3.en_buf dac_1.sw_top_3.net1 avdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 comparator_0.vp dac_0.carray_0.unitcap_320.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 dac_1.out dac_1.carray_0.unitcap_328.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 dac_1.out dac_1.carray_0.unitcap_71.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 avdd.t210 avss.t410 avdd.t209 avdd.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X160 vinp.t69 dac_0.sw_top_2.en_buf comparator_0.vp.t64 avdd.t286 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X161 vinn.t11 dac_1.sw_top_3.en_buf dac_1.out.t18 avdd.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X162 avss.t63 ctln7.t1 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t4 avss.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X163 comparator_0.vp dac_0.carray_0.unitcap_200.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 avss.t316 dac_0.sw_top_3.en_buf dac_0.sw_top_3.net1 avss.t315 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X165 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 dac_1.out dac_1.carray_0.unitcap_167.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 avdd.t106 sample.t7 dac_0.sw_top_1.en_buf avdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X168 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t3 ctlp7.t1 avss.t230 avss.t229 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X173 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 vinn.t43 dac_1.sw_top_1.en_buf dac_1.out.t48 avdd.t143 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X176 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 vinp.t68 dac_0.sw_top_2.en_buf comparator_0.vp.t63 avdd.t285 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X178 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t3 ctln3.t1 avss.t7 avss.t6 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X179 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 comparator_0.vp dac_0.carray_0.unitcap_104.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 dac_0.sky130_fd_sc_hd__inv_2_7.Y avdd.t6 avdd.t7 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X182 comparator_0.trim_0.n4.t13 trim4.t2 avss.t370 avss.t369 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X183 dac_1.out.t47 dac_1.sw_top_1.en_buf vinn.t42 avdd.t142 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X184 avss.t162 sample.t8 dac_1.sw_top_1.en_buf avss.t161 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X185 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 dac_0.sw_top_2.en_buf sample.t9 avdd.t146 avdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X188 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 comparator_0.vp.t83 dac_0.carray_0.unitcap_331.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 avss.t306 trimb4.t2 comparator_0.trim_1.n4.t5 avss.t305 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X192 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 avdd.t155 ctlp3.t1 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t1 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X194 avss.t88 trim3.t0 comparator_0.trim_0.n3.t4 avss.t87 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X195 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 dac_1.out dac_1.carray_0.unitcap_24.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 dac_1.out.t81 dac_1.carray_0.unitcap_11.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 dac_0.sky130_fd_sc_hd__inv_2_6.Y ctlp0.t0 avdd.t2 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X201 vinp.t48 dac_0.sw_top_3.en_buf comparator_0.vp.t42 avdd.t256 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X202 dac_1.out.t78 dac_1.sw_top_2.en_buf vinn.t75 avdd.t307 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X203 avdd.t180 dac_0.sw_top_1.en_buf dac_0.sw_top_1.net1 avdd.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X204 dac_1.out.t58 dac_1.sw_top_3.net1 vinn.t55 avss.t255 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X205 comparator_0.trim_1.n3.t3 trimb3.t0 avss.t128 avss.t127 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X206 avss.t94 comparator_0.outp a_33300_6679# avss.t93 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X207 avdd.t213 avss.t411 avdd.t212 avdd.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X208 avdd.t158 ctlp4.t1 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t2 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X209 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 comparator_0.vp.t43 dac_0.sw_top_3.en_buf vinp.t47 avdd.t255 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X212 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 avss.t56 avdd.t312 avss.t55 avss.t54 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X214 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_6.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 comparator_0.vp dac_0.carray_0.unitcap_207.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 avdd.t148 sample.t10 dac_1.sw_top_3.en_buf avdd.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X218 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 comparator_0.vp dac_0.carray_0.unitcap_7.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 comparator_0.ip.t3 comparator_0.trim_1.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 dac_0.sw_top_2.net1 dac_0.sw_top_2.en_buf avdd.t284 avdd.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X222 comparator_0.vp.t18 dac_0.sw_top_2.net1 vinp.t18 avss.t147 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X223 vinp.t78 dac_0.sw_top_1.net1 comparator_0.vp.t73 avss.t357 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X224 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 comparator_0.ip.t0 clkc.t1 avdd.t20 avdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X226 dac_0.sw_top_3.net1 dac_0.sw_top_3.en_buf avss.t314 avss.t313 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 comparator_0.vp.t23 dac_0.sw_top_0.net1 vinp.t28 avss.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X228 vinn.t10 dac_1.sw_top_3.en_buf dac_1.out.t17 avdd.t46 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X229 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 avdd.t216 avss.t412 avdd.t215 avdd.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X232 vinn.t69 dac_1.sw_top_1.net1 dac_1.out.t68 avss.t273 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X233 dac_1.out dac_1.carray_0.unitcap_48.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 vinp.t17 dac_0.sw_top_2.net1 comparator_0.vp.t11 avss.t146 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X237 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 comparator_0.vp dac_0.carray_0.unitcap_231.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 comparator_0.vp dac_0.carray_0.unitcap_103.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 comparator_0.vp.t80 dac_0.carray_0.unitcap_10.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 dac_1.out.t67 dac_1.sw_top_1.net1 vinn.t68 avss.t272 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X247 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 dac_1.out dac_1.carray_0.unitcap_39.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 dac_0.sw_top_3.net1 dac_0.sw_top_3.en_buf avdd.t254 avdd.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X258 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 comparator_0.vp.t50 dac_0.sw_top_3.net1 vinp.t57 avss.t330 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X261 dac_1.out dac_1.carray_0.unitcap_104.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 dac_1.out dac_1.carray_0.unitcap_128.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 dac_1.sw_top_1.net1 dac_1.sw_top_1.en_buf avdd.t141 avdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X264 avss.t53 avdd.t313 avss.t52 avss.t51 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X265 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 avdd.t150 sample.t11 dac_1.sw_top_2.en_buf avdd.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X267 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 vinn.t38 dac_1.sw_top_0.net1 dac_1.out.t38 avss.t210 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X271 comparator_0.vp dac_0.carray_0.unitcap_208.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 dac_1.out dac_1.carray_0.unitcap_247.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 dac_1.out dac_1.carray_0.unitcap_119.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 dac_1.out dac_1.carray_0.unitcap_32.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 avss.t191 sample.t12 dac_1.sw_top_1.en_buf avss.t190 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X276 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 comparator_0.vp.t1 dac_0.sw_top_0.en_buf vinp.t7 avdd.t66 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X281 dac_1.out.t7 dac_1.sw_top_2.net1 vinn.t3 avss.t81 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X282 comparator_0.vp.t84 dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 avdd.t178 dac_0.sw_top_1.en_buf dac_0.sw_top_1.net1 avdd.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X286 comparator_0.vp.t41 dac_0.sw_top_3.en_buf vinp.t46 avdd.t252 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X287 avss.t193 sample.t13 dac_0.sw_top_1.en_buf avss.t192 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X288 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 dac_1.out.t57 dac_1.sw_top_3.net1 vinn.t54 avss.t254 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X292 dac_1.sw_top_2.en_buf sample.t14 avss.t195 avss.t194 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X293 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 dac_1.out dac_1.carray_0.unitcap_168.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 comparator_0.trim_1.n3.t2 trimb3.t1 avss.t130 avss.t129 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X299 comparator_0.trim_1.n0 trimb0.t0 avss.t160 avss.t159 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X300 avss.t174 trim1.t0 comparator_0.trim_0.n1 avss.t173 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X301 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 comparator_0.vp dac_0.carray_0.unitcap_87.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 dac_1.out.t77 dac_1.sw_top_2.en_buf vinn.t74 avdd.t306 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X305 dac_1.out dac_1.carray_0.unitcap_64.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 dac_1.out.t27 dac_1.sw_top_0.en_buf vinn.t28 avdd.t100 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X307 avss.t225 dac_1.sw_top_1.en_buf dac_1.sw_top_1.net1 avss.t224 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 comparator_0.vp dac_0.carray_0.unitcap_96.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 dac_1.out dac_1.carray_0.unitcap_112.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 dac_0.sw_top_2.net1 dac_0.sw_top_2.en_buf avdd.t282 avdd.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X311 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 comparator_0.vp dac_0.carray_0.unitcap_336.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 comparator_0.vp dac_0.carray_0.unitcap_151.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 avdd.t159 ctlp5.t0 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t0 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X321 comparator_0.vp dac_0.carray_0.unitcap_32.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 dac_1.out.t82 dac_1.carray_0.unitcap_12.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 dac_1.sw_top_2.net1 dac_1.sw_top_2.en_buf avss.t388 avss.t387 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X325 dac_0.sw_top_0.net1 dac_0.sw_top_0.en_buf avdd.t65 avdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X326 avdd.t110 ctln0.t0 dac_1.sky130_fd_sc_hd__inv_2_6.Y dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X327 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 vinn.t16 dac_1.sw_top_3.en_buf dac_1.out.t16 avdd.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X329 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 dac_1.out dac_1.carray_0.unitcap_95.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 avss.t50 avdd.t314 avss.t49 avss.t48 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X335 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 dac_1.out dac_1.carray_0.unitcap_160.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 comparator_0.vp.t66 dac_0.sw_top_2.en_buf vinp.t67 avdd.t280 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X341 vinp.t37 dac_0.sw_top_1.en_buf comparator_0.vp.t39 avdd.t176 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X342 avdd.t217 avss.t413 dac_1.sky130_fd_sc_hd__inv_2_7.Y dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X343 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 avss.t47 avdd.t315 avss.t46 avss.t45 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X345 comparator_0.vp.t2 dac_0.sw_top_0.en_buf vinp.t6 avdd.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X346 avss.t186 ctln0.t1 dac_1.sky130_fd_sc_hd__inv_2_6.Y avss.t185 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X347 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp1.t1 avss.t338 avss.t337 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X348 comparator_0.vp dac_0.carray_0.unitcap_216.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 dac_1.out dac_1.carray_0.unitcap_183.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 vinp.t66 dac_0.sw_top_2.en_buf comparator_0.vp.t60 avdd.t279 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X351 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 avdd.t34 comparator_0.outp a_33300_6679# avdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X353 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 avdd.t12 sample.t15 dac_1.sw_top_2.en_buf avdd.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X356 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 avss.t244 avss.t242 dac_1.sky130_fd_sc_hd__inv_2_7.Y avss.t243 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X361 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 dac_1.sw_top_3.net1 dac_1.sw_top_3.en_buf avss.t102 avss.t101 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X364 comparator_0.vp.t51 dac_0.sw_top_3.net1 vinp.t56 avss.t329 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X365 avss.t308 trimb4.t3 comparator_0.trim_1.n4.t4 avss.t307 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X366 avss.t368 trim4.t3 comparator_0.trim_0.n4.t12 avss.t367 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X367 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 comparator_0.diff clkc.t2 avss.t67 avss.t66 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X369 vinn.t41 dac_1.sw_top_1.en_buf dac_1.out.t46 avdd.t139 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X370 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 vinn.t37 dac_1.sw_top_0.net1 dac_1.out.t37 avss.t209 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X372 dac_1.sky130_fd_sc_hd__inv_2_6.Y ctln0.t2 avdd.t111 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X373 comparator_0.trim_1.n4.t3 trimb4.t4 avss.t182 avss.t181 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X374 avdd.t72 ctln6.t0 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t1 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X375 avdd.t14 sample.t16 dac_1.sw_top_0.en_buf avdd.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X376 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 comparator_0.vp dac_0.carray_0.unitcap_144.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_5.Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 comparator_0.vp.t47 dac_0.sw_top_3.en_buf vinp.t45 avdd.t251 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X383 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 dac_1.out dac_1.carray_0.unitcap_240.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 avss.t348 dac_0.sw_top_2.en_buf dac_0.sw_top_2.net1 avss.t347 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X386 comparator_0.ip.t4 comparator_0.trim_1.n1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 dac_0.sw_top_2.en_buf sample.t17 avdd.t16 avdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 comparator_0.vp dac_0.carray_0.unitcap_88.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 vinp.t77 dac_0.sw_top_1.net1 comparator_0.vp.t70 avss.t356 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X391 comparator_0.ip.t2 comparator_0.vp.t85 comparator_0.diff avss.t187 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X392 avss.t223 dac_1.sw_top_1.en_buf dac_1.sw_top_1.net1 avss.t222 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X393 dac_1.sky130_fd_sc_hd__inv_2_6.Y ctln0.t3 avss.t166 avss.t165 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X394 dac_1.out dac_1.carray_0.unitcap_322.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 dac_1.out.t76 dac_1.sw_top_2.en_buf vinn.t73 avdd.t305 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X396 avdd.t304 dac_1.sw_top_2.en_buf dac_1.sw_top_2.net1 avdd.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X397 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 dac_1.sw_top_3.en_buf sample.t18 avdd.t265 avdd.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X399 comparator_0.vp dac_0.carray_0.unitcap_48.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 dac_1.out.t26 dac_1.sw_top_0.en_buf vinn.t27 avdd.t99 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X404 comparator_0.vp dac_0.carray_0.unitcap_47.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 comparator_0.vp.t74 dac_0.sw_top_1.net1 vinp.t76 avss.t355 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X407 vinn.t72 dac_1.sw_top_2.en_buf dac_1.out.t75 avdd.t302 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X408 vinn.t53 dac_1.sw_top_3.net1 dac_1.out.t56 avss.t253 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X409 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t5 ctln7.t2 avdd.t239 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X410 comparator_0.in.t8 comparator_0.trim_0.n3.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 dac_1.sw_top_2.net1 dac_1.sw_top_2.en_buf avss.t386 avss.t385 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X412 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 avss.t44 avdd.t316 dac_0.sky130_fd_sc_hd__inv_2_7.Y avss.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X415 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 comparator_0.vp dac_0.carray_0.unitcap_223.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 comparator_0.vp dac_0.carray_0.unitcap_127.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 avdd.t220 avss.t414 avdd.t219 avdd.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X423 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t2 ctln6.t1 avdd.t73 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X424 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 avss.t42 avdd.t317 avss.t41 avss.t40 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X426 avss.t39 avdd.t318 avss.t38 avss.t37 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X427 avss.t36 avdd.t319 avss.t35 avss.t34 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X428 vinn.t67 dac_1.sw_top_1.net1 dac_1.out.t66 avss.t271 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X429 avss.t5 ctlp0.t1 dac_0.sky130_fd_sc_hd__inv_2_6.Y avss.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X430 comparator_0.vp.t86 dac_0.carray_0.unitcap_9.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 avdd.t223 avss.t415 avdd.t222 avdd.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X432 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 vinp.t27 dac_0.sw_top_0.net1 comparator_0.vp.t20 avss.t156 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X434 dac_1.sw_top_1.en_buf sample.t19 avdd.t267 avdd.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X435 dac_1.sw_top_0.net1 dac_1.sw_top_0.en_buf avss.t134 avss.t133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X436 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 dac_1.out dac_1.carray_0.unitcap_63.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 dac_1.out.t65 dac_1.sw_top_1.net1 vinn.t66 avss.t270 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X440 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 comparator_0.vp.t82 dac_0.carray_0.unitcap_330.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 comparator_0.vp.t10 dac_0.sw_top_2.net1 vinp.t16 avss.t145 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X448 comparator_0.outp comparator_0.outn avdd.t29 avdd.t28 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X449 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 dac_1.out.t83 dac_1.carray_0.unitcap_15.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 dac_0.sw_top_2.net1 dac_0.sw_top_2.en_buf avss.t346 avss.t345 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X452 dac_1.out.t6 dac_1.sw_top_2.net1 vinn.t2 avss.t80 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X453 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 dac_1.out dac_1.carray_0.unitcap_239.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 avss.t336 sample.t20 dac_0.sw_top_3.en_buf avss.t335 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X458 dac_1.out dac_1.carray_0.unitcap_143.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 avss.t197 sample.t21 dac_0.sw_top_1.en_buf avss.t196 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X460 avss.t246 ctlp5.t1 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t1 avss.t245 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X461 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_5.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 comparator_0.vp.t54 dac_0.sw_top_3.net1 vinp.t55 avss.t328 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X463 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 vinp.t5 dac_0.sw_top_0.en_buf comparator_0.vp.t0 avdd.t62 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X466 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 dac_1.sw_top_1.net1 dac_1.sw_top_1.en_buf avdd.t138 avdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X469 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 avdd.t120 sample.t22 dac_1.sw_top_0.en_buf avdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X471 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 avss.t366 trim4.t4 comparator_0.trim_0.n4.t11 avss.t365 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X473 avss.t110 dac_0.sw_top_0.en_buf dac_0.sw_top_0.net1 avss.t109 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X474 vinn.t40 dac_1.sw_top_1.en_buf dac_1.out.t45 avdd.t136 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X475 comparator_0.ip.t5 comparator_0.trim_1.n4.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 vinn.t52 dac_1.sw_top_3.net1 dac_1.out.t55 avss.t252 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X477 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 comparator_0.vp dac_0.carray_0.unitcap_71.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 comparator_0.vp.t44 dac_0.sw_top_3.en_buf vinp.t44 avdd.t250 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X487 avdd.t226 avss.t416 avdd.t225 avdd.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X488 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 comparator_0.ip.t6 comparator_0.trim_1.n4.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 avdd.t301 dac_1.sw_top_2.en_buf dac_1.sw_top_2.net1 avdd.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X491 dac_1.sw_top_3.en_buf sample.t23 avdd.t122 avdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X492 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 comparator_0.ip.t7 comparator_0.trim_1.n4.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 comparator_0.trim_1.n2 trimb2.t1 avss.t120 avss.t119 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X495 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 avdd.t98 dac_1.sw_top_0.en_buf dac_1.sw_top_0.net1 avdd.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X497 dac_1.sw_top_2.en_buf sample.t24 avss.t302 avss.t301 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X498 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 dac_0.sw_top_0.en_buf sample.t25 avdd.t238 avdd.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 comparator_0.vp dac_0.carray_0.unitcap_167.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 dac_1.out.t25 dac_1.sw_top_0.en_buf vinn.t26 avdd.t96 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X508 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 vinp.t36 dac_0.sw_top_1.en_buf comparator_0.vp.t38 avdd.t175 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X511 avss.t170 ctln6.t2 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t3 avss.t169 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X512 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 dac_0.sw_top_1.en_buf sample.t26 avss.t304 avss.t303 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X516 dac_1.sw_top_3.net1 dac_1.sw_top_3.en_buf avdd.t44 avdd.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 dac_1.out dac_1.carray_0.unitcap_326.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 avdd.t22 sample.t27 dac_0.sw_top_3.en_buf avdd.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 comparator_0.vp.t34 dac_0.sw_top_1.en_buf vinp.t35 avdd.t174 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X526 avss.t33 avdd.t320 avss.t32 avss.t31 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X527 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 comparator_0.vp dac_0.carray_0.unitcap_14.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 vinp.t26 dac_0.sw_top_0.net1 comparator_0.vp.t26 avss.t155 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X530 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 dac_1.out dac_1.carray_0.unitcap_23.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 avss.t108 dac_0.sw_top_0.en_buf dac_0.sw_top_0.net1 avss.t107 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X537 dac_1.out.t5 dac_1.sw_top_2.net1 vinn.t1 avss.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X538 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t6 ctln7.t3 avss.t310 avss.t309 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X546 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 comparator_0.ip.t8 comparator_0.trim_1.n4.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 avdd.t249 dac_0.sw_top_3.en_buf dac_0.sw_top_3.net1 avdd.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X549 dac_0.sw_top_1.en_buf sample.t28 avdd.t24 avdd.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 dac_1.out dac_1.carray_0.unitcap_324.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 vinp.t4 dac_0.sw_top_0.en_buf comparator_0.vp.t7 avdd.t61 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X552 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 avdd.t8 ctlp1.t2 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X554 avss.t344 dac_0.sw_top_2.en_buf dac_0.sw_top_2.net1 avss.t343 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X555 dac_1.out.t44 dac_1.sw_top_1.en_buf vinn.t47 avdd.t135 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X556 avdd.t229 avss.t417 avdd.t228 avdd.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X557 dac_1.out dac_1.carray_0.unitcap_191.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 dac_1.out.t36 dac_1.sw_top_0.net1 vinn.t36 avss.t208 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X559 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t4 ctln6.t3 avss.t172 avss.t171 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X560 dac_1.out.t84 dac_1.carray_0.unitcap_9.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 comparator_0.in.t9 comparator_0.trim_0.n4.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 comparator_0.vp.t61 dac_0.sw_top_2.en_buf vinp.t65 avdd.t278 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X563 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 comparator_0.vp.t83 dac_0.carray_0.unitcap_334.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 comparator_0.ip.t9 comparator_0.trim_1.n4.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 avss.t364 trim4.t5 comparator_0.trim_0.n4.t10 avss.t363 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X574 vinp.t54 dac_0.sw_top_3.net1 comparator_0.vp.t53 avss.t327 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X575 avdd.t287 ctlp2.t2 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X576 comparator_0.trim_0.n3.t5 trim3.t1 avss.t90 avss.t89 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X577 comparator_0.vp.t49 dac_0.sw_top_3.en_buf vinp.t43 avdd.t247 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X578 vinn.t71 dac_1.sw_top_2.en_buf dac_1.out.t74 avdd.t299 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X579 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 avdd.t232 avss.t418 avdd.t231 avdd.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X581 vinn.t51 dac_1.sw_top_3.net1 dac_1.out.t54 avss.t251 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X582 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t0 ctlp3.t2 avdd.t288 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X585 avss.t298 trimb3.t2 comparator_0.trim_1.n3.t1 avss.t297 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X586 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 comparator_0.vp dac_0.carray_0.unitcap_39.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 dac_0.sw_top_0.en_buf sample.t29 avdd.t26 avdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X590 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 vinp.t75 dac_0.sw_top_1.net1 comparator_0.vp.t78 avss.t354 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X592 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t0 ctlp4.t2 avdd.t157 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X595 avdd.t95 dac_1.sw_top_0.en_buf dac_1.sw_top_0.net1 avdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X596 comparator_0.vp dac_0.carray_0.unitcap_120.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 latch_0.Qn comp.t3 avss.t180 avss.t179 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X598 comparator_0.vp.t71 dac_0.sw_top_1.net1 vinp.t74 avss.t353 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X599 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 comparator_0.vp dac_0.carray_0.unitcap_247.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 comparator_0.vp dac_0.carray_0.unitcap_119.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 dac_1.sw_top_0.en_buf sample.t30 avss.t390 avss.t389 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X607 comparator_0.vp dac_0.carray_0.unitcap_56.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 dac_1.out dac_1.carray_0.unitcap_0.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 vinn.t24 dac_1.sw_top_0.en_buf dac_1.out.t24 avdd.t93 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X613 dac_1.out.t85 dac_1.carray_0.unitcap_288.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 dac_1.out.t64 dac_1.sw_top_1.net1 vinn.t63 avss.t269 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X615 comparator_0.vp.t16 dac_0.sw_top_2.net1 vinp.t15 avss.t144 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X616 comparator_0.vp dac_0.carray_0.unitcap_24.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 dac_0.sw_top_2.net1 dac_0.sw_top_2.en_buf avss.t342 avss.t341 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X618 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t0 ctlp2.t3 avdd.t74 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X621 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 avss.t258 trim0.t0 comparator_0.trim_0.n0 avss.t257 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X626 vinn.t62 dac_1.sw_top_1.net1 dac_1.out.t63 avss.t268 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X627 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 avss.t392 sample.t31 dac_1.sw_top_3.en_buf avss.t391 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X630 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 avdd.t235 avss.t419 avdd.t234 avdd.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X633 avdd.t153 clkc.t3 comparator_0.in.t2 avdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X634 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_7.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 comparator_0.trim_1.n1 trimb1.t0 avss.t396 avss.t395 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X636 comparator_0.vp dac_0.carray_0.unitcap_240.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 dac_1.out dac_1.carray_0.unitcap_72.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 dac_1.out dac_1.carray_0.unitcap_255.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 avdd.t246 dac_0.sw_top_3.en_buf dac_0.sw_top_3.net1 avdd.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X640 dac_1.out dac_1.carray_0.unitcap_96.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 vinp.t53 dac_0.sw_top_3.net1 comparator_0.vp.t59 avss.t326 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X642 dac_1.out dac_1.carray_0.unitcap_331.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 dac_1.out.t4 dac_1.sw_top_2.net1 vinn.t8 avss.t78 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X647 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 dac_1.out dac_1.carray_0.unitcap_111.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 dac_1.out.t35 dac_1.sw_top_0.net1 vinn.t35 avss.t207 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X653 dac_1.out dac_1.carray_0.unitcap_16.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 comparator_0.vp dac_0.carray_0.unitcap_13.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 comparator_0.outp comparator_0.outn comparator_0.ip.t1 avss.t86 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X656 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 vinp.t3 dac_0.sw_top_0.en_buf comparator_0.vp.t4 avdd.t60 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X658 dac_1.out.t43 dac_1.sw_top_1.en_buf vinn.t46 avdd.t134 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X659 vinn.t7 dac_1.sw_top_2.net1 dac_1.out.t3 avss.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X660 avss.t100 dac_1.sw_top_3.en_buf dac_1.sw_top_3.net1 avss.t99 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X661 dac_1.sw_top_1.en_buf sample.t32 avss.t394 avss.t393 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X662 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 comparator_0.vp dac_0.carray_0.unitcap_160.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 comparator_0.ip.t10 comparator_0.trim_1.n3.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 dac_1.out dac_1.carray_0.unitcap_175.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 comparator_0.vp dac_0.carray_0.unitcap_95.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 dac_0.sw_top_0.net1 dac_0.sw_top_0.en_buf avss.t106 avss.t105 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X672 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 comparator_0.in.t10 comparator_0.trim_0.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 dac_1.out dac_1.carray_0.unitcap_152.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 dac_1.sw_top_0.net1 dac_1.sw_top_0.en_buf avdd.t92 avdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X679 vinn.t50 dac_1.sw_top_3.net1 dac_1.out.t53 avss.t250 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X680 avss.t122 sample.t33 dac_0.sw_top_3.en_buf avss.t121 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X681 comparator_0.vp.t86 dac_0.carray_0.unitcap_256.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 comparator_0.in.t11 comparator_0.trim_0.n3.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 dac_1.out dac_1.carray_0.unitcap_56.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 comparator_0.vp dac_0.carray_0.unitcap_72.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 comparator_0.vp dac_0.carray_0.unitcap_183.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 vinn.t23 dac_1.sw_top_0.en_buf dac_1.out.t23 avdd.t90 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X691 avss.t30 avdd.t321 avss.t29 avss.t28 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X692 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 comparator_0.vp.t87 dac_0.carray_0.unitcap_328.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 vinp.t42 dac_0.sw_top_3.en_buf comparator_0.vp.t45 avdd.t244 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X697 comparator_0.ip.t11 comparator_0.trim_1.n4.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 dac_1.sw_top_0.en_buf sample.t34 avss.t124 avss.t123 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X700 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 dac_0.sw_top_1.net1 dac_0.sw_top_1.en_buf avss.t282 avss.t281 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X702 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 dac_0.sw_top_0.net1 dac_0.sw_top_0.en_buf avss.t104 avss.t103 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X704 dac_1.out dac_1.carray_0.unitcap_192.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_5.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t2 ctlp5.t2 avdd.t160 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X709 comparator_0.vp.t12 dac_0.sw_top_2.net1 vinp.t14 avss.t143 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X710 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 vinp.t34 dac_0.sw_top_1.en_buf comparator_0.vp.t36 avdd.t173 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X712 dac_1.out dac_1.carray_0.unitcap_88.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 vinn.t61 dac_1.sw_top_1.net1 dac_1.out.t62 avss.t267 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X714 dac_1.out dac_1.carray_0.unitcap_136.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 dac_1.out dac_1.carray_0.unitcap_224.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 avdd.t80 sample.t35 dac_0.sw_top_3.en_buf avdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X717 comparator_0.vp.t28 dac_0.sw_top_0.net1 vinp.t25 avss.t154 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X718 comparator_0.vp.t35 dac_0.sw_top_1.en_buf vinp.t33 avdd.t172 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X719 avss.t380 latch_0.Qn comp.t2 avss.t379 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X720 vinn.t15 dac_1.sw_top_3.en_buf dac_1.out.t15 avdd.t42 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X721 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 avdd.t82 sample.t36 dac_1.sw_top_1.en_buf avdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X726 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 dac_1.sky130_fd_sc_hd__inv_2_7.Y avss.t420 avdd.t236 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X730 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 comparator_0.vp.t67 dac_0.sw_top_2.en_buf vinp.t64 avdd.t277 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X734 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 dac_0.sw_top_3.en_buf sample.t37 avss.t126 avss.t125 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X736 avss.t27 avdd.t322 avss.t26 avss.t25 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X737 dac_1.out dac_1.carray_0.unitcap_215.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 vinp.t52 dac_0.sw_top_3.net1 comparator_0.vp.t58 avss.t325 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X740 avdd.t189 avss.t421 avdd.t188 avdd.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X741 avss.t98 dac_1.sw_top_3.en_buf dac_1.sw_top_3.net1 avss.t97 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X742 comparator_0.vp dac_0.carray_0.unitcap_168.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 comparator_0.ip.t12 comparator_0.trim_1.n4.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 dac_1.sky130_fd_sc_hd__inv_2_7.Y avss.t239 avss.t241 avss.t240 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X747 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 dac_1.out dac_1.carray_0.unitcap_176.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 comparator_0.trim_0.n4.t9 trim4.t6 avss.t362 avss.t361 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X752 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 dac_1.out dac_1.carray_0.unitcap_321.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 dac_1.out dac_1.carray_0.unitcap_55.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 latch_0.Qn comp.t4 avdd.t109 avdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X757 dac_1.out.t42 dac_1.sw_top_1.en_buf vinn.t45 avdd.t133 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X758 vinn.t6 dac_1.sw_top_2.net1 dac_1.out.t2 avss.t76 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X759 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 dac_1.out.t34 dac_1.sw_top_0.net1 vinn.t34 avss.t206 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X761 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 vinp.t41 dac_0.sw_top_3.en_buf comparator_0.vp.t46 avdd.t243 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X763 dac_1.out dac_1.carray_0.unitcap_184.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 avss.t280 dac_0.sw_top_1.en_buf dac_0.sw_top_1.net1 avss.t279 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X765 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 comparator_0.in.t12 comparator_0.trim_0.n0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 dac_1.out dac_1.carray_0.unitcap_337.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 dac_0.sw_top_1.net1 dac_0.sw_top_1.en_buf avdd.t171 avdd.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X770 comparator_0.trim_1.n4.t2 trimb4.t5 avss.t184 avss.t183 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X771 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 dac_1.out dac_1.carray_0.unitcap_135.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 comparator_0.vp dac_0.carray_0.unitcap_63.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 avdd.t123 ctln2.t0 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t2 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X777 avdd.t84 sample.t38 dac_0.sw_top_2.en_buf avdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X778 comparator_0.vp.t72 dac_0.sw_top_1.net1 vinp.t73 avss.t352 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X779 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X780 comparator_0.vp dac_0.carray_0.unitcap_15.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 vinn.t70 dac_1.sw_top_2.en_buf dac_1.out.t73 avdd.t298 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X782 avdd.t77 ctln5.t0 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t2 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X783 comparator_0.ip.t13 comparator_0.trim_1.n4.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 vinp.t72 dac_0.sw_top_1.net1 comparator_0.vp.t76 avss.t351 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X785 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 comparator_0.vp dac_0.carray_0.unitcap_239.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 avdd.t185 ctlp6.t0 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t1 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X788 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X789 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 comparator_0.vp dac_0.carray_0.unitcap_143.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X794 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X795 dac_1.out dac_1.carray_0.unitcap_232.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 avdd.t151 ctln4.t0 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t2 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X797 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X798 avdd.t192 avss.t422 avdd.t191 avdd.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X799 avdd.t71 ctlp7.t2 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t0 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X800 vinn.t79 dac_1.sw_top_2.en_buf dac_1.out.t72 avdd.t297 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X801 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X802 comparator_0.vp dac_0.carray_0.unitcap_8.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X803 dac_0.sky130_fd_sc_hd__inv_2_7.Y avdd.t323 avss.t24 avss.t23 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X804 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X805 dac_1.out.t61 dac_1.sw_top_1.net1 vinn.t60 avss.t266 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X806 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X807 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X808 avdd.t268 ctln3.t2 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t4 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X809 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X810 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X811 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X813 comparator_0.vp.t19 dac_0.sw_top_2.net1 vinp.t13 avss.t142 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X814 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 avss.t264 ctlp3.t3 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t2 avss.t263 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X816 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X817 dac_0.sky130_fd_sc_hd__inv_2_6.Y ctlp0.t2 avss.t164 avss.t163 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X818 avss.t22 avdd.t324 avss.t21 avss.t20 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X819 comparator_0.vp.t29 dac_0.sw_top_0.net1 vinp.t24 avss.t153 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X820 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 vinn.t14 dac_1.sw_top_3.en_buf dac_1.out.t14 avdd.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X822 avdd.t76 sample.t39 dac_1.sw_top_1.en_buf avdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X823 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t3 ctln2.t1 avdd.t124 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X824 comparator_0.in.t13 comparator_0.trim_0.n4.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X825 comparator_0.vp dac_0.carray_0.unitcap_16.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X826 vinp.t12 dac_0.sw_top_2.net1 comparator_0.vp.t14 avss.t141 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X827 dac_0.sw_top_0.en_buf sample.t40 avss.t114 avss.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X828 avss.t238 ctlp4.t3 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t1 avss.t237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X829 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X830 avss.t116 sample.t41 dac_1.sw_top_3.en_buf avss.t115 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X831 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X833 dac_1.out.t13 dac_1.sw_top_3.en_buf vinn.t13 avdd.t40 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X834 vinn.t5 dac_1.sw_top_2.net1 dac_1.out.t1 avss.t75 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X835 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X836 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X837 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X838 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X839 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X840 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X841 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t2 ctlp6.t1 avdd.t186 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X842 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X843 comparator_0.in.t14 comparator_0.trim_0.n4.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X844 comparator_0.vp.t65 dac_0.sw_top_2.en_buf vinp.t63 avdd.t276 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X845 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X846 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X847 dac_1.sw_top_2.en_buf sample.t42 avdd.t261 avdd.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X848 vinp.t51 dac_0.sw_top_3.net1 comparator_0.vp.t55 avss.t324 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X849 comparator_0.vp.t5 dac_0.sw_top_0.en_buf vinp.t2 avdd.t59 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X850 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X851 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t3 ctln4.t1 avdd.t152 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X852 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t4 ctlp5.t3 avss.t398 avss.t397 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X853 avdd.t132 dac_1.sw_top_1.en_buf dac_1.sw_top_1.net1 avdd.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X854 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X855 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X856 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X857 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 dac_1.out.t33 dac_1.sw_top_0.net1 vinn.t33 avss.t205 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X859 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X860 dac_1.out dac_1.carray_0.unitcap_199.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X861 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X863 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X864 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X865 comparator_0.outp clkc.t4 avdd.t154 avdd.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X866 avdd.t32 comparator_0.outp comparator_0.outn avdd.t28 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X867 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 dac_1.out dac_1.carray_0.unitcap_31.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X869 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X870 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X871 dac_1.out.t86 dac_1.carray_0.unitcap_256.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X872 dac_1.out.t52 dac_1.sw_top_3.net1 vinn.t59 avss.t249 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X873 vinn.t32 dac_1.sw_top_0.net1 dac_1.out.t32 avss.t204 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X874 avdd.t263 sample.t43 dac_0.sw_top_2.en_buf avdd.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X875 comparator_0.trim_1.n4.t1 trimb4.t6 avss.t233 avss.t232 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X876 vinp.t40 dac_0.sw_top_3.en_buf comparator_0.vp.t48 avdd.t242 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X877 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X878 avss.t231 a_33300_6679# latch_0.Qn avss.t93 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X879 comparator_0.trim_0.n2 trim2.t1 avss.t65 avss.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X880 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X881 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X882 dac_1.sw_top_2.net1 dac_1.sw_top_2.en_buf avdd.t296 avdd.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X884 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X885 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X886 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X888 comparator_0.vp dac_0.carray_0.unitcap_23.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X889 dac_1.sw_top_1.net1 dac_1.sw_top_1.en_buf avss.t221 avss.t220 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X890 avdd.t290 latch_0.Qn comp.t1 avdd.t289 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X891 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X892 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X893 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_6.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 vinp.t71 dac_0.sw_top_1.net1 comparator_0.vp.t79 avss.t350 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X895 avss.t334 sample.t44 dac_1.sw_top_2.en_buf avss.t333 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X896 comparator_0.vp dac_0.carray_0.unitcap_112.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X897 avdd.t162 sample.t45 dac_0.sw_top_0.en_buf avdd.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X898 comparator_0.ip.t14 comparator_0.trim_1.n3.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X899 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp1.t3 avdd.t9 dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X900 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X901 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X902 dac_1.out dac_1.carray_0.unitcap_334.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X903 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t3 ctln5.t1 avdd.t78 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X904 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X905 comparator_0.vp dac_0.carray_0.unitcap_191.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X906 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X907 dac_1.out.t22 dac_1.sw_top_0.en_buf vinn.t22 avdd.t89 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X908 avss.t19 avdd.t325 avss.t18 avss.t17 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X909 comparator_0.vp dac_0.carray_0.unitcap_0.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X910 comparator_0.vp dac_0.carray_0.unitcap_12.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 avss.t16 avdd.t326 avss.t15 avss.t14 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X912 avdd.t275 dac_0.sw_top_2.en_buf dac_0.sw_top_2.net1 avdd.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X913 dac_0.sw_top_3.en_buf sample.t46 avdd.t164 avdd.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 dac_0.sw_top_2.en_buf sample.t47 avss.t262 avss.t261 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X915 vinp.t32 dac_0.sw_top_1.en_buf comparator_0.vp.t31 avdd.t169 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X916 dac_1.sw_top_3.net1 dac_1.sw_top_3.en_buf avdd.t39 avdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X917 avss.t13 avdd.t327 avss.t12 avss.t11 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X918 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X919 dac_0.sw_top_3.en_buf sample.t48 avss.t320 avss.t319 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X920 dac_1.out.t12 dac_1.sw_top_3.en_buf vinn.t19 avdd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X921 avdd.t195 avss.t423 avdd.t194 avdd.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X922 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 comparator_0.ip.t15 comparator_0.trim_1.n3.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X924 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X926 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X927 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X928 avss.t213 ctln2.t2 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t4 avss.t212 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X930 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X931 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X932 vinp.t11 dac_0.sw_top_2.net1 comparator_0.vp.t17 avss.t140 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X933 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X934 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X935 avss.t118 ctln5.t2 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t4 avss.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X936 comparator_0.vp.t27 dac_0.sw_top_0.net1 vinp.t23 avss.t152 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X937 comparator_0.vp.t81 dac_0.carray_0.unitcap_324.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X938 comparator_0.ip.t16 comparator_0.trim_1.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 dac_0.sw_top_3.net1 dac_0.sw_top_3.en_buf avss.t312 avss.t311 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X940 comparator_0.vp dac_0.carray_0.unitcap_232.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X941 dac_0.sw_top_1.net1 dac_0.sw_top_1.en_buf avss.t278 avss.t277 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X942 avss.t296 ctlp6.t2 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t3 avss.t295 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X943 comparator_0.in.t0 dac_1.out.t87 comparator_0.diff avss.t187 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X944 avss.t276 dac_0.sw_top_1.en_buf dac_0.sw_top_1.net1 avss.t275 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X945 comparator_0.vp.t69 dac_0.sw_top_2.en_buf vinp.t62 avdd.t273 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X946 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X947 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X948 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X949 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X950 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X951 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X952 comparator_0.vp.t87 dac_0.carray_0.unitcap_326.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X953 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 dac_1.out dac_1.carray_0.unitcap_79.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X955 comparator_0.vp.t3 dac_0.sw_top_0.en_buf vinp.t1 avdd.t58 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X956 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X957 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X958 avss.t112 ctlp7.t3 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t1 avss.t111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X959 vinn.t31 dac_1.sw_top_0.net1 dac_1.out.t31 avss.t203 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X960 avdd.t130 dac_1.sw_top_1.en_buf dac_1.sw_top_1.net1 avdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X961 avss.t227 ctln4.t2 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t4 avss.t226 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X962 dac_0.sw_top_1.en_buf sample.t49 avdd.t259 avdd.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X963 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 vinp.t61 dac_0.sw_top_2.en_buf comparator_0.vp.t62 avdd.t272 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X965 avss.t340 ctln3.t3 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t5 avss.t339 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X966 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X967 avdd.t5 avdd.t4 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X968 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X969 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X971 dac_1.out dac_1.carray_0.unitcap_338.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 comparator_0.vp dac_0.carray_0.unitcap_176.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X973 dac_1.out dac_1.carray_0.unitcap_159.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X974 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X975 avss.t92 trim3.t2 comparator_0.trim_0.n3.t6 avss.t91 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X976 dac_1.sw_top_2.net1 dac_1.sw_top_2.en_buf avdd.t294 avdd.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X977 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t1 ctln2.t3 avss.t178 avss.t177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X978 dac_1.out.t71 dac_1.sw_top_2.en_buf vinn.t78 avdd.t292 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X979 vinn.t44 dac_1.sw_top_1.en_buf dac_1.out.t41 avdd.t128 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X980 avdd.t198 avss.t424 avdd.t197 avdd.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X981 comparator_0.vp dac_0.carray_0.unitcap_128.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X982 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X983 avdd.t107 ctlp0.t3 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X984 comparator_0.in.t15 comparator_0.trim_0.n1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X985 avss.t322 sample.t50 dac_0.sw_top_2.en_buf avss.t321 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X986 comparator_0.trim_1.n4.t0 trimb4.t7 avss.t235 avss.t234 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X987 dac_1.out.t21 dac_1.sw_top_0.en_buf vinn.t21 avdd.t88 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X988 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X989 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X990 comparator_0.trim_0.n3.t7 trim3.t3 avss.t189 avss.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X991 avss.t400 sample.t51 dac_1.sw_top_2.en_buf avss.t399 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X993 dac_0.sw_top_1.net1 dac_0.sw_top_1.en_buf avdd.t168 avdd.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X994 avdd.t310 sample.t52 dac_0.sw_top_0.en_buf avdd.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X995 comparator_0.vp.t75 dac_0.sw_top_1.net1 vinp.t70 avss.t349 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X996 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t0 ctlp6.t3 avss.t73 avss.t72 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X997 comparator_0.vp dac_0.carray_0.unitcap_80.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X998 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X999 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1000 comparator_0.vp dac_0.carray_0.unitcap_255.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1001 vinn.t77 dac_1.sw_top_2.en_buf dac_1.out.t70 avdd.t291 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1002 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1003 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1004 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1005 avss.t300 trimb3.t3 comparator_0.trim_1.n3.t0 avss.t299 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1006 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1007 dac_1.sw_top_0.net1 dac_1.sw_top_0.en_buf avdd.t87 avdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1008 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1009 dac_1.out.t88 dac_1.carray_0.unitcap_10.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1010 comparator_0.vp dac_0.carray_0.unitcap_111.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1011 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t1 ctln4.t3 avss.t199 avss.t198 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1012 avss.t402 sample.t53 dac_1.sw_top_0.en_buf avss.t401 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1013 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1014 avdd.t271 dac_0.sw_top_2.en_buf dac_0.sw_top_2.net1 avdd.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1015 dac_0.sw_top_3.en_buf sample.t54 avdd.t1 avdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1016 comparator_0.diff clkc.t5 avss.t228 avss.t66 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1017 comparator_0.ip.t17 comparator_0.trim_1.n0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1018 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1019 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1020 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1021 dac_0.sw_top_0.en_buf sample.t55 avss.t1 avss.t0 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1022 vinp.t10 dac_0.sw_top_2.net1 comparator_0.vp.t15 avss.t139 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1023 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1025 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1026 comparator_0.vp dac_0.carray_0.unitcap_175.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1027 dac_1.out.t11 dac_1.sw_top_3.en_buf vinn.t18 avdd.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1028 avdd.t57 dac_0.sw_top_0.en_buf dac_0.sw_top_0.net1 avdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1029 dac_1.out.t60 dac_1.sw_top_1.net1 vinn.t65 avss.t265 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1030 comparator_0.vp dac_0.carray_0.unitcap_321.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 dac_1.out dac_1.carray_0.unitcap_8.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1033 vinp.t31 dac_0.sw_top_1.en_buf comparator_0.vp.t32 avdd.t166 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1034 avss.t384 dac_1.sw_top_2.en_buf dac_1.sw_top_2.net1 avss.t383 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1035 dac_1.sw_top_3.en_buf sample.t56 avss.t3 avss.t2 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1036 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1037 dac_1.out dac_1.carray_0.unitcap_330.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1038 comparator_0.vp.t21 dac_0.sw_top_0.net1 vinp.t22 avss.t151 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1039 avdd.t112 ctln1.t1 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1040 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1041 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1043 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1044 dac_1.out dac_1.carray_0.unitcap_40.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1045 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1046 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1047 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1048 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 dac_0.sw_top_3.net1 dac_0.sw_top_3.en_buf avdd.t241 avdd.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1050 comparator_0.vp.t57 dac_0.sw_top_3.net1 vinp.t50 avss.t323 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1051 vinp.t21 dac_0.sw_top_0.net1 comparator_0.vp.t24 avss.t150 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X1052 comparator_0.vp dac_0.carray_0.unitcap_11.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1053 vinn.t0 dac_1.sw_top_2.net1 dac_1.out.t0 avss.t74 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1054 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t1 ctln5.t3 avss.t61 avss.t60 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1055 avdd.t201 avss.t425 avdd.t200 avdd.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1056 vinn.t30 dac_1.sw_top_0.net1 dac_1.out.t30 avss.t202 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1057 avss.t71 ctln1.t2 dac_1.sky130_fd_sc_hd__inv_2_4.Y avss.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1058 comparator_0.vp dac_0.carray_0.unitcap_192.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1060 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_8.Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1061 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1062 dac_1.out dac_1.carray_0.unitcap_207.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1063 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1064 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1065 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1066 dac_1.out dac_1.carray_0.unitcap_7.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1067 comparator_0.vp.t6 dac_0.sw_top_0.en_buf vinp.t0 avdd.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1068 avss.t360 trim4.t7 comparator_0.trim_0.n4.t8 avss.t359 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1069 dac_1.sw_top_2.en_buf sample.t57 avdd.t184 avdd.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1070 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1071 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1072 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1073 dac_1.sw_top_1.en_buf sample.t58 avss.t290 avss.t289 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1074 dac_1.out dac_1.carray_0.unitcap_80.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1075 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1076 dac_1.out dac_1.carray_0.unitcap_120.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1077 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1078 avss.t292 sample.t59 dac_0.sw_top_0.en_buf avss.t291 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1079 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1080 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1081 comparator_0.ip.t18 comparator_0.trim_1.n3.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1082 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1083 comparator_0.in.t16 comparator_0.trim_0.n4.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1084 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1085 dac_1.out dac_1.carray_0.unitcap_231.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1086 dac_1.out dac_1.carray_0.unitcap_103.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1087 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1088 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1089 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1090 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1091 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 vinn.t58 dac_1.sw_top_3.net1 dac_1.out.t51 avss.t248 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1093 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1094 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1095 comparator_0.vp dac_0.carray_0.unitcap_215.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1096 dac_1.sw_top_1.net1 dac_1.sw_top_1.en_buf avss.t219 avss.t218 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1097 avss.t404 sample.t60 dac_1.sw_top_0.en_buf avss.t403 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1098 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1099 dac_1.out.t50 dac_1.sw_top_3.net1 vinn.t57 avss.t247 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1100 comparator_0.in.t17 comparator_0.trim_0.n4.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1101 vinn.t20 dac_1.sw_top_0.en_buf dac_1.out.t20 avdd.t85 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1102 dac_1.out dac_1.carray_0.unitcap_144.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1103 comparator_0.vp dac_0.carray_0.unitcap_55.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1104 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1105 comparator_0.vp.t33 dac_0.sw_top_1.en_buf vinp.t30 avdd.t165 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1106 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1107 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1108 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1109 comparator_0.in.t18 comparator_0.trim_0.n4.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1110 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1111 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1112 avss.t382 dac_1.sw_top_2.en_buf dac_1.sw_top_2.net1 avss.t381 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1113 dac_1.sw_top_3.en_buf sample.t61 avss.t406 avss.t405 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1114 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1115 avdd.t54 dac_0.sw_top_0.en_buf dac_0.sw_top_0.net1 avdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1116 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1117 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1118 vinp.t20 dac_0.sw_top_0.net1 comparator_0.vp.t25 avss.t149 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1119 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1120 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1121 dac_1.out.t89 dac_1.carray_0.unitcap_13.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1122 comparator_0.vp dac_0.carray_0.unitcap_135.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1123 dac_1.out.t10 dac_1.sw_top_3.en_buf vinn.t17 avdd.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1124 avss.t132 dac_1.sw_top_0.en_buf dac_1.sw_top_0.net1 avss.t131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1125 vinp.t60 dac_0.sw_top_2.en_buf comparator_0.vp.t68 avdd.t269 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1126 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1127 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1128 dac_1.out dac_1.carray_0.unitcap_200.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1129 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1130 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1131 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1132 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1133 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1134 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1135 dac_1.out dac_1.carray_0.unitcap_87.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1136 a_33300_5579# comparator_0.outn avss.t85 avss.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X1137 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1138 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1139 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1140 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1141 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1142 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1143 avdd.t204 avss.t426 avdd.t203 avdd.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1144 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln1.t3 avdd.t27 dac_1.sky130_fd_sc_hd__inv_2_6.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1145 dac_1.out dac_1.carray_0.unitcap_216.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1146 dac_0.sw_top_2.en_buf sample.t62 avss.t408 avss.t407 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1147 dac_1.sw_top_3.net1 dac_1.sw_top_3.en_buf avss.t96 avss.t95 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1148 vinn.t49 dac_1.sw_top_1.en_buf dac_1.out.t40 avdd.t127 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1149 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1150 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1151 avss.t69 sample.t63 dac_0.sw_top_2.en_buf avss.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1152 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1153 dac_1.out dac_1.carray_0.unitcap_336.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1154 avss.t10 avdd.t328 avss.t9 avss.t8 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1155 comparator_0.vp dac_0.carray_0.unitcap_184.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1156 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1157 dac_1.out dac_1.carray_0.unitcap_151.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 comparator_0.vp.n10 comparator_0.vp.t85 130.87
R1 comparator_0.vp.n56 comparator_0.vp.t64 28.5655
R2 comparator_0.vp.n56 comparator_0.vp.t65 28.5655
R3 comparator_0.vp.n59 comparator_0.vp.t68 28.5655
R4 comparator_0.vp.n59 comparator_0.vp.t66 28.5655
R5 comparator_0.vp.n61 comparator_0.vp.t60 28.5655
R6 comparator_0.vp.n61 comparator_0.vp.t67 28.5655
R7 comparator_0.vp.n53 comparator_0.vp.t62 28.5655
R8 comparator_0.vp.n53 comparator_0.vp.t69 28.5655
R9 comparator_0.vp.n52 comparator_0.vp.t63 28.5655
R10 comparator_0.vp.n52 comparator_0.vp.t61 28.5655
R11 comparator_0.vp.n41 comparator_0.vp.t8 28.5655
R12 comparator_0.vp.n41 comparator_0.vp.t2 28.5655
R13 comparator_0.vp.n43 comparator_0.vp.t0 28.5655
R14 comparator_0.vp.n43 comparator_0.vp.t5 28.5655
R15 comparator_0.vp.n38 comparator_0.vp.t7 28.5655
R16 comparator_0.vp.n38 comparator_0.vp.t3 28.5655
R17 comparator_0.vp.n46 comparator_0.vp.t4 28.5655
R18 comparator_0.vp.n46 comparator_0.vp.t6 28.5655
R19 comparator_0.vp.n48 comparator_0.vp.t9 28.5655
R20 comparator_0.vp.n48 comparator_0.vp.t1 28.5655
R21 comparator_0.vp.n24 comparator_0.vp.t32 28.5655
R22 comparator_0.vp.n24 comparator_0.vp.t34 28.5655
R23 comparator_0.vp.n27 comparator_0.vp.t31 28.5655
R24 comparator_0.vp.n27 comparator_0.vp.t30 28.5655
R25 comparator_0.vp.n30 comparator_0.vp.t36 28.5655
R26 comparator_0.vp.n30 comparator_0.vp.t33 28.5655
R27 comparator_0.vp.n32 comparator_0.vp.t38 28.5655
R28 comparator_0.vp.n32 comparator_0.vp.t37 28.5655
R29 comparator_0.vp.n35 comparator_0.vp.t39 28.5655
R30 comparator_0.vp.n35 comparator_0.vp.t35 28.5655
R31 comparator_0.vp.n15 comparator_0.vp.t46 28.5655
R32 comparator_0.vp.n15 comparator_0.vp.t41 28.5655
R33 comparator_0.vp.n17 comparator_0.vp.t48 28.5655
R34 comparator_0.vp.n17 comparator_0.vp.t47 28.5655
R35 comparator_0.vp.n12 comparator_0.vp.t40 28.5655
R36 comparator_0.vp.n12 comparator_0.vp.t44 28.5655
R37 comparator_0.vp.n20 comparator_0.vp.t42 28.5655
R38 comparator_0.vp.n20 comparator_0.vp.t49 28.5655
R39 comparator_0.vp.n22 comparator_0.vp.t45 28.5655
R40 comparator_0.vp.n22 comparator_0.vp.t43 28.5655
R41 comparator_0.vp.n65 comparator_0.vp.n52 17.7565
R42 comparator_0.vp.n54 comparator_0.vp.t14 17.4005
R43 comparator_0.vp.n54 comparator_0.vp.t19 17.4005
R44 comparator_0.vp.n55 comparator_0.vp.t13 17.4005
R45 comparator_0.vp.n55 comparator_0.vp.t12 17.4005
R46 comparator_0.vp.n58 comparator_0.vp.t15 17.4005
R47 comparator_0.vp.n58 comparator_0.vp.t18 17.4005
R48 comparator_0.vp.n57 comparator_0.vp.t11 17.4005
R49 comparator_0.vp.n57 comparator_0.vp.t16 17.4005
R50 comparator_0.vp.n40 comparator_0.vp.t25 17.4005
R51 comparator_0.vp.n40 comparator_0.vp.t23 17.4005
R52 comparator_0.vp.n39 comparator_0.vp.t22 17.4005
R53 comparator_0.vp.n39 comparator_0.vp.t28 17.4005
R54 comparator_0.vp.n37 comparator_0.vp.t20 17.4005
R55 comparator_0.vp.n37 comparator_0.vp.t29 17.4005
R56 comparator_0.vp.n45 comparator_0.vp.t26 17.4005
R57 comparator_0.vp.n45 comparator_0.vp.t27 17.4005
R58 comparator_0.vp.n47 comparator_0.vp.t24 17.4005
R59 comparator_0.vp.n47 comparator_0.vp.t21 17.4005
R60 comparator_0.vp.n25 comparator_0.vp.t79 17.4005
R61 comparator_0.vp.n25 comparator_0.vp.t74 17.4005
R62 comparator_0.vp.n26 comparator_0.vp.t76 17.4005
R63 comparator_0.vp.n26 comparator_0.vp.t77 17.4005
R64 comparator_0.vp.n29 comparator_0.vp.t78 17.4005
R65 comparator_0.vp.n29 comparator_0.vp.t75 17.4005
R66 comparator_0.vp.n28 comparator_0.vp.t70 17.4005
R67 comparator_0.vp.n28 comparator_0.vp.t72 17.4005
R68 comparator_0.vp.n23 comparator_0.vp.t73 17.4005
R69 comparator_0.vp.n23 comparator_0.vp.t71 17.4005
R70 comparator_0.vp.n14 comparator_0.vp.t59 17.4005
R71 comparator_0.vp.n14 comparator_0.vp.t57 17.4005
R72 comparator_0.vp.n13 comparator_0.vp.t58 17.4005
R73 comparator_0.vp.n13 comparator_0.vp.t50 17.4005
R74 comparator_0.vp.n11 comparator_0.vp.t55 17.4005
R75 comparator_0.vp.n11 comparator_0.vp.t51 17.4005
R76 comparator_0.vp.n19 comparator_0.vp.t52 17.4005
R77 comparator_0.vp.n19 comparator_0.vp.t54 17.4005
R78 comparator_0.vp.n21 comparator_0.vp.t53 17.4005
R79 comparator_0.vp.n21 comparator_0.vp.t56 17.4005
R80 comparator_0.vp.n63 comparator_0.vp.t17 17.4005
R81 comparator_0.vp.n63 comparator_0.vp.t10 17.4005
R82 comparator_0.vp.n36 comparator_0.vp.n35 16.1315
R83 comparator_0.vp comparator_0.vp.n10 14.8566
R84 comparator_0.vp.n49 comparator_0.vp 8.6431
R85 comparator_0.vp.n49 comparator_0.vp 8.04326
R86 comparator_0.vp comparator_0.vp.n36 7.6255
R87 comparator_0.vp.n34 comparator_0.vp.n23 6.81045
R88 comparator_0.vp.n64 comparator_0.vp.n63 6.80945
R89 comparator_0.vp.n50 comparator_0.vp.n49 6.19787
R90 comparator_0.vp.n65 comparator_0.vp 6.0005
R91 comparator_0.vp.n51 comparator_0.vp.n50 4.3755
R92 comparator_0.vp.t86 comparator_0.vp 3.90072
R93 comparator_0.vp.t86 comparator_0.vp 3.43072
R94 comparator_0.vp.t80 comparator_0.vp 2.96072
R95 comparator_0.vp.n1 comparator_0.vp.n46 2.52713
R96 comparator_0.vp.n4 comparator_0.vp.n20 2.52713
R97 comparator_0.vp.n0 comparator_0.vp.n43 2.52031
R98 comparator_0.vp.n3 comparator_0.vp.n17 2.52031
R99 comparator_0.vp.t80 comparator_0.vp 2.49072
R100 comparator_0.vp.n10 comparator_0.vp 2.48939
R101 comparator_0.vp.n7 comparator_0.vp.n53 2.46792
R102 comparator_0.vp.n9 comparator_0.vp.n24 2.46792
R103 comparator_0.vp.n6 comparator_0.vp.n61 2.4611
R104 comparator_0.vp.n8 comparator_0.vp.n32 2.4611
R105 comparator_0.vp.n62 comparator_0.vp.n56 2.45716
R106 comparator_0.vp.n44 comparator_0.vp.n38 2.45716
R107 comparator_0.vp.n33 comparator_0.vp.n27 2.45716
R108 comparator_0.vp.n18 comparator_0.vp.n12 2.45716
R109 comparator_0.vp.n60 comparator_0.vp.n59 2.45239
R110 comparator_0.vp.n42 comparator_0.vp.n41 2.45239
R111 comparator_0.vp.n31 comparator_0.vp.n30 2.45239
R112 comparator_0.vp.n16 comparator_0.vp.n15 2.45239
R113 comparator_0.vp.n50 comparator_0.vp 2.42846
R114 comparator_0.vp.n65 comparator_0.vp.n64 1.19147
R115 comparator_0.vp.n36 comparator_0.vp.n34 1.10119
R116 comparator_0.vp comparator_0.vp.n5 1.05955
R117 comparator_0.vp.n7 comparator_0.vp.n62 0.783395
R118 comparator_0.vp.n9 comparator_0.vp.n33 0.783395
R119 comparator_0.vp.n62 comparator_0.vp.n6 0.776816
R120 comparator_0.vp.n33 comparator_0.vp.n8 0.776816
R121 comparator_0.vp.n1 comparator_0.vp.n45 0.750575
R122 comparator_0.vp.n4 comparator_0.vp.n19 0.750575
R123 comparator_0.vp.n2 comparator_0.vp.n47 0.747946
R124 comparator_0.vp.n5 comparator_0.vp.n21 0.747946
R125 comparator_0.vp.n62 comparator_0.vp.n55 0.729384
R126 comparator_0.vp.n44 comparator_0.vp.n37 0.729384
R127 comparator_0.vp.n33 comparator_0.vp.n26 0.729384
R128 comparator_0.vp.n18 comparator_0.vp.n11 0.729384
R129 comparator_0.vp.n0 comparator_0.vp.n39 0.72521
R130 comparator_0.vp.n3 comparator_0.vp.n13 0.72521
R131 comparator_0.vp.n1 comparator_0.vp.n44 0.720895
R132 comparator_0.vp.n4 comparator_0.vp.n18 0.720895
R133 comparator_0.vp.n44 comparator_0.vp.n0 0.714316
R134 comparator_0.vp.n18 comparator_0.vp.n3 0.714316
R135 comparator_0.vp.n6 comparator_0.vp.n60 0.704447
R136 comparator_0.vp.n8 comparator_0.vp.n31 0.704447
R137 comparator_0.vp.n7 comparator_0.vp.n54 0.688075
R138 comparator_0.vp.n9 comparator_0.vp.n25 0.688075
R139 comparator_0.vp.t86 comparator_0.vp 0.680248
R140 comparator_0.vp.n42 comparator_0.vp.n40 0.669405
R141 comparator_0.vp.n31 comparator_0.vp.n29 0.669405
R142 comparator_0.vp.n16 comparator_0.vp.n14 0.669405
R143 comparator_0.vp.n60 comparator_0.vp.n58 0.668426
R144 comparator_0.vp.t86 comparator_0.vp 0.592671
R145 comparator_0.vp.n2 comparator_0.vp.n48 2.52245
R146 comparator_0.vp.n5 comparator_0.vp.n22 2.52245
R147 comparator_0.vp comparator_0.vp.n51 1.90839
R148 comparator_0.vp comparator_0.vp.n2 1.07616
R149 comparator_0.vp.n3 comparator_0.vp.n16 0.711026
R150 comparator_0.vp.n0 comparator_0.vp.n42 0.711026
R151 comparator_0.vp.n8 comparator_0.vp.n28 0.665835
R152 comparator_0.vp.n6 comparator_0.vp.n57 0.665835
R153 comparator_0.vp.n5 comparator_0.vp.n4 0.658395
R154 comparator_0.vp.n2 comparator_0.vp.n1 0.658395
R155 comparator_0.vp comparator_0.vp.t86 0.554117
R156 comparator_0.vp.t82 comparator_0.vp.t83 0.530033
R157 comparator_0.vp.t83 comparator_0.vp.t87 0.530033
R158 comparator_0.vp.t87 comparator_0.vp.t81 0.530033
R159 comparator_0.vp.t81 comparator_0.vp 0.530033
R160 comparator_0.vp.t80 comparator_0.vp 0.530033
R161 comparator_0.vp.t86 comparator_0.vp.t80 0.530033
R162 comparator_0.vp.t80 comparator_0.vp 0.505093
R163 comparator_0.vp.t84 comparator_0.vp 0.442952
R164 comparator_0.vp.n51 comparator_0.vp.t84 0.438617
R165 comparator_0.vp.n36 comparator_0.vp 0.424111
R166 comparator_0.vp.t84 comparator_0.vp 0.421933
R167 comparator_0.vp comparator_0.vp.t82 0.418056
R168 comparator_0.vp.t80 comparator_0.vp 0.417516
R169 comparator_0.vp.t80 comparator_0.vp 0.398433
R170 comparator_0.vp.t80 comparator_0.vp 0.398433
R171 comparator_0.vp.t86 comparator_0.vp 0.398433
R172 comparator_0.vp.t86 comparator_0.vp 0.398433
R173 comparator_0.vp.n34 comparator_0.vp.n9 0.388493
R174 comparator_0.vp.n64 comparator_0.vp.n7 0.388493
R175 comparator_0.vp comparator_0.vp.n65 0.333833
R176 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n0 111.322
R177 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.n2 50.4671
R178 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t0 26.5955
R179 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t2 26.5955
R180 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t1 24.9236
R181 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t3 24.9236
R182 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_2.Y 13.5685
R183 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.n3 11.2645
R184 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.n4 9.41342
R185 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_2.Y 6.1445
R186 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_2.Y 4.65505
R187 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_2.Y 3.8405
R188 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.n1 2.0485
R189 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.55202
R190 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.t4 0.197458
R191 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n5 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.18982
R192 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.105455
R193 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y.n5 0.0316375
R194 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.00959054
R195 vinp.n22 vinp.t42 29.3118
R196 vinp.n37 vinp.t37 29.3118
R197 vinp.n52 vinp.t9 29.3118
R198 vinp.n8 vinp.t68 29.3118
R199 vinp.n27 vinp.t46 29.3084
R200 vinp.n42 vinp.t30 29.3084
R201 vinp.n57 vinp.t6 29.3084
R202 vinp.n13 vinp.t67 29.3084
R203 vinp.n21 vinp.t47 28.5655
R204 vinp.n21 vinp.t48 28.5655
R205 vinp.n19 vinp.t43 28.5655
R206 vinp.n19 vinp.t49 28.5655
R207 vinp.n17 vinp.t44 28.5655
R208 vinp.n17 vinp.t40 28.5655
R209 vinp.n15 vinp.t45 28.5655
R210 vinp.n15 vinp.t41 28.5655
R211 vinp.n36 vinp.t33 28.5655
R212 vinp.n36 vinp.t31 28.5655
R213 vinp.n34 vinp.t35 28.5655
R214 vinp.n34 vinp.t32 28.5655
R215 vinp.n32 vinp.t38 28.5655
R216 vinp.n32 vinp.t36 28.5655
R217 vinp.n30 vinp.t39 28.5655
R218 vinp.n30 vinp.t34 28.5655
R219 vinp.n51 vinp.t7 28.5655
R220 vinp.n51 vinp.t3 28.5655
R221 vinp.n49 vinp.t0 28.5655
R222 vinp.n49 vinp.t4 28.5655
R223 vinp.n47 vinp.t1 28.5655
R224 vinp.n47 vinp.t5 28.5655
R225 vinp.n45 vinp.t2 28.5655
R226 vinp.n45 vinp.t8 28.5655
R227 vinp.n7 vinp.t65 28.5655
R228 vinp.n7 vinp.t61 28.5655
R229 vinp.n5 vinp.t62 28.5655
R230 vinp.n5 vinp.t69 28.5655
R231 vinp.n3 vinp.t63 28.5655
R232 vinp.n3 vinp.t66 28.5655
R233 vinp.n1 vinp.t64 28.5655
R234 vinp.n1 vinp.t60 28.5655
R235 vinp.n22 vinp.t54 18.1397
R236 vinp.n27 vinp.t50 18.1397
R237 vinp.n37 vinp.t78 18.1397
R238 vinp.n42 vinp.t70 18.1397
R239 vinp.n52 vinp.t21 18.1397
R240 vinp.n57 vinp.t28 18.1397
R241 vinp.n8 vinp.t11 18.1397
R242 vinp.n13 vinp.t18 18.1397
R243 vinp.n20 vinp.t58 17.4005
R244 vinp.n20 vinp.t59 17.4005
R245 vinp.n18 vinp.t55 17.4005
R246 vinp.n18 vinp.t51 17.4005
R247 vinp.n16 vinp.t56 17.4005
R248 vinp.n16 vinp.t52 17.4005
R249 vinp.n14 vinp.t57 17.4005
R250 vinp.n14 vinp.t53 17.4005
R251 vinp.n35 vinp.t74 17.4005
R252 vinp.n35 vinp.t71 17.4005
R253 vinp.n33 vinp.t76 17.4005
R254 vinp.n33 vinp.t72 17.4005
R255 vinp.n31 vinp.t79 17.4005
R256 vinp.n31 vinp.t77 17.4005
R257 vinp.n29 vinp.t73 17.4005
R258 vinp.n29 vinp.t75 17.4005
R259 vinp.n50 vinp.t22 17.4005
R260 vinp.n50 vinp.t26 17.4005
R261 vinp.n48 vinp.t23 17.4005
R262 vinp.n48 vinp.t27 17.4005
R263 vinp.n46 vinp.t24 17.4005
R264 vinp.n46 vinp.t29 17.4005
R265 vinp.n44 vinp.t25 17.4005
R266 vinp.n44 vinp.t20 17.4005
R267 vinp.n6 vinp.t16 17.4005
R268 vinp.n6 vinp.t12 17.4005
R269 vinp.n4 vinp.t13 17.4005
R270 vinp.n4 vinp.t19 17.4005
R271 vinp.n2 vinp.t14 17.4005
R272 vinp.n2 vinp.t17 17.4005
R273 vinp.n0 vinp.t15 17.4005
R274 vinp.n0 vinp.t10 17.4005
R275 vinp.n59 vinp.n58 8.59648
R276 vinp.n61 vinp.n60 7.00774
R277 vinp.n60 vinp.n59 6.6802
R278 vinp vinp.n61 2.91369
R279 vinp.n61 vinp 2.19494
R280 vinp.n59 vinp.n43 1.91305
R281 vinp.n60 vinp.n28 1.9116
R282 vinp.n24 vinp.n23 0.811311
R283 vinp.n39 vinp.n38 0.811311
R284 vinp.n54 vinp.n53 0.811311
R285 vinp.n10 vinp.n9 0.811311
R286 vinp.n26 vinp.n25 0.799575
R287 vinp.n41 vinp.n40 0.799575
R288 vinp.n56 vinp.n55 0.799575
R289 vinp.n12 vinp.n11 0.799575
R290 vinp.n25 vinp.n24 0.794419
R291 vinp.n40 vinp.n39 0.794419
R292 vinp.n55 vinp.n54 0.794419
R293 vinp.n11 vinp.n10 0.794419
R294 vinp.n23 vinp.n22 0.787662
R295 vinp.n38 vinp.n37 0.787662
R296 vinp.n53 vinp.n52 0.787662
R297 vinp.n9 vinp.n8 0.787662
R298 vinp.n27 vinp.n26 0.773526
R299 vinp.n42 vinp.n41 0.773526
R300 vinp.n57 vinp.n56 0.773526
R301 vinp.n13 vinp.n12 0.773526
R302 vinp.n23 vinp.n21 0.746823
R303 vinp.n24 vinp.n19 0.746823
R304 vinp.n25 vinp.n17 0.746823
R305 vinp.n38 vinp.n36 0.746823
R306 vinp.n39 vinp.n34 0.746823
R307 vinp.n40 vinp.n32 0.746823
R308 vinp.n53 vinp.n51 0.746823
R309 vinp.n54 vinp.n49 0.746823
R310 vinp.n55 vinp.n47 0.746823
R311 vinp.n9 vinp.n7 0.746823
R312 vinp.n10 vinp.n5 0.746823
R313 vinp.n11 vinp.n3 0.746823
R314 vinp.n26 vinp.n15 0.743351
R315 vinp.n41 vinp.n30 0.743351
R316 vinp.n56 vinp.n45 0.743351
R317 vinp.n12 vinp.n1 0.743351
R318 vinp.n23 vinp.n20 0.739748
R319 vinp.n24 vinp.n18 0.739748
R320 vinp.n25 vinp.n16 0.739748
R321 vinp.n26 vinp.n14 0.739748
R322 vinp.n38 vinp.n35 0.739748
R323 vinp.n39 vinp.n33 0.739748
R324 vinp.n40 vinp.n31 0.739748
R325 vinp.n41 vinp.n29 0.739748
R326 vinp.n53 vinp.n50 0.739748
R327 vinp.n54 vinp.n48 0.739748
R328 vinp.n55 vinp.n46 0.739748
R329 vinp.n56 vinp.n44 0.739748
R330 vinp.n9 vinp.n6 0.739748
R331 vinp.n10 vinp.n4 0.739748
R332 vinp.n11 vinp.n2 0.739748
R333 vinp.n12 vinp.n0 0.739748
R334 vinp vinp.n13 0.627876
R335 vinp.n28 vinp.n27 0.580661
R336 vinp.n43 vinp.n42 0.579116
R337 vinp.n58 vinp.n57 0.573599
R338 vinp.n58 vinp 0.063
R339 vinp.n43 vinp 0.0583907
R340 vinp.n28 vinp 0.0567584
R341 avdd.n7447 avdd.n7443 6176.47
R342 avdd.n7486 avdd.n7482 6176.47
R343 avdd.n7546 avdd.n7542 6176.47
R344 avdd.n7586 avdd.n7582 6176.47
R345 avdd.n1813 avdd.n1812 6176.47
R346 avdd.n1639 avdd.n1638 6176.47
R347 avdd.n1723 avdd.n1722 6176.47
R348 avdd.n1675 avdd.n1674 6176.47
R349 avdd.n7448 avdd.n7447 3240
R350 avdd.n7487 avdd.n7486 3240
R351 avdd.n7547 avdd.n7546 3240
R352 avdd.n7587 avdd.n7586 3240
R353 avdd.n1812 avdd.n1811 3240
R354 avdd.n1638 avdd.n1637 3240
R355 avdd.n1722 avdd.n1721 3240
R356 avdd.n1674 avdd.n1673 3240
R357 avdd.n7448 avdd.n7446 3056.47
R358 avdd.n7487 avdd.n7485 3056.47
R359 avdd.n7547 avdd.n7545 3056.47
R360 avdd.n7587 avdd.n7585 3056.47
R361 avdd.n1811 avdd.n1807 3056.47
R362 avdd.n1637 avdd.n1633 3056.47
R363 avdd.n1721 avdd.n1717 3056.47
R364 avdd.n1673 avdd.n1669 3056.47
R365 avdd.n4765 avdd.n4764 1662.05
R366 avdd.n4756 avdd.n4486 1041.18
R367 avdd.n4652 avdd.n4582 984.707
R368 avdd.n4661 avdd.n4585 928.236
R369 avdd.t221 avdd 895.586
R370 avdd.t224 avdd 895.586
R371 avdd avdd.t202 895.586
R372 avdd.t187 avdd 895.586
R373 avdd.t205 avdd 895.586
R374 avdd.t208 avdd 895.586
R375 avdd avdd.t190 895.586
R376 avdd.t218 avdd 895.586
R377 avdd.n4492 avdd.n4490 744.707
R378 avdd.n4764 avdd 670.76
R379 avdd.n7596 avdd.t150 584.644
R380 avdd.n7619 avdd.t304 584.644
R381 avdd.n7563 avdd.t148 584.644
R382 avdd.n7556 avdd.t51 584.644
R383 avdd.n7496 avdd.t82 584.644
R384 avdd.n7519 avdd.t132 584.644
R385 avdd.n7464 avdd.t14 584.644
R386 avdd.n7457 avdd.t98 584.644
R387 avdd.n1667 avdd.t57 584.644
R388 avdd.n1700 avdd.t162 584.644
R389 avdd.n1757 avdd.t180 584.644
R390 avdd.n1750 avdd.t126 584.644
R391 avdd.n1631 avdd.t249 584.644
R392 avdd.n1790 avdd.t80 584.644
R393 avdd.n1847 avdd.t275 584.644
R394 avdd.n1840 avdd.t84 584.644
R395 avdd.n7502 avdd.t225 512.547
R396 avdd.t203 avdd.n7571 512.547
R397 avdd.n7602 avdd.t188 512.547
R398 avdd.n7472 avdd.t222 512.547
R399 avdd.n1708 avdd.t206 512.542
R400 avdd.n1741 avdd.t209 512.542
R401 avdd.n1798 avdd.t191 512.542
R402 avdd.n1831 avdd.t219 512.542
R403 avdd.t211 avdd.n7422 489.178
R404 avdd.t222 avdd.n7426 459.192
R405 avdd.n7500 avdd.t225 459.192
R406 avdd.n7572 avdd.t203 459.192
R407 avdd.n7600 avdd.t188 459.192
R408 avdd.t206 avdd.n1660 459.192
R409 avdd.n1739 avdd.t209 459.192
R410 avdd.t191 avdd.n1624 459.192
R411 avdd.n1829 avdd.t219 459.192
R412 avdd avdd.n7529 428.521
R413 avdd.n7530 avdd 428.521
R414 avdd avdd.n7629 428.521
R415 avdd.n7631 avdd 428.521
R416 avdd avdd.n1767 428.521
R417 avdd.n1768 avdd 428.521
R418 avdd avdd.n1857 428.521
R419 avdd.n1864 avdd 428.521
R420 avdd.t199 avdd.n1656 422.029
R421 avdd.t227 avdd 378.64
R422 avdd avdd.t193 378.64
R423 avdd.t196 avdd 378.64
R424 avdd.t214 avdd 378.64
R425 avdd avdd.t230 378.64
R426 avdd.t233 avdd 378.64
R427 avdd.n4759 avdd.t19 355.536
R428 avdd.t17 avdd.t28 344.103
R429 avdd.n7529 avdd.t221 340.096
R430 avdd.n7530 avdd.t224 340.096
R431 avdd.n7629 avdd.t202 340.096
R432 avdd.n7631 avdd.t187 340.096
R433 avdd.n1767 avdd.t205 340.096
R434 avdd.n1768 avdd.t208 340.096
R435 avdd.n1857 avdd.t190 340.096
R436 avdd.n1864 avdd.t218 340.096
R437 avdd.n1863 avdd.n1858 318.524
R438 avdd.n1656 avdd.n1651 318.524
R439 avdd.t97 avdd 301.551
R440 avdd.t131 avdd 301.551
R441 avdd avdd.t50 301.551
R442 avdd.t303 avdd 301.551
R443 avdd.t56 avdd 301.551
R444 avdd.t179 avdd 301.551
R445 avdd avdd.t248 301.551
R446 avdd.t274 avdd 301.551
R447 avdd.n7447 avdd.t88 289.37
R448 avdd.n7486 avdd.t135 289.37
R449 avdd.n7546 avdd.t37 289.37
R450 avdd.n7586 avdd.t292 289.37
R451 avdd.n1812 avdd.t280 289.37
R452 avdd.n1638 avdd.t252 289.37
R453 avdd.n1722 avdd.t165 289.37
R454 avdd.n1674 avdd.t63 289.37
R455 avdd.t285 avdd.n1809 287.747
R456 avdd.t244 avdd.n1635 287.747
R457 avdd.t176 avdd.n1719 287.747
R458 avdd.t70 avdd.n1671 287.747
R459 avdd.n7450 avdd.t93 287.676
R460 avdd.n7489 avdd.t128 287.676
R461 avdd.n7549 avdd.t47 287.676
R462 avdd.n7589 avdd.t297 287.676
R463 avdd.t13 avdd 285.68
R464 avdd.t81 avdd 285.68
R465 avdd avdd.t147 285.68
R466 avdd.t149 avdd 285.68
R467 avdd.t161 avdd 285.68
R468 avdd.t125 avdd 285.68
R469 avdd avdd.t79 285.68
R470 avdd.t83 avdd 285.68
R471 avdd avdd.t211 247.137
R472 avdd avdd.t227 247.137
R473 avdd.t193 avdd 247.137
R474 avdd avdd.t196 247.137
R475 avdd avdd.t199 247.137
R476 avdd avdd.t214 247.137
R477 avdd.t230 avdd 247.137
R478 avdd avdd.t233 247.137
R479 avdd.n7419 avdd.t226 243.03
R480 avdd.n7627 avdd.t204 243.03
R481 avdd.n7403 avdd.t189 243.03
R482 avdd.n7527 avdd.t223 243.03
R483 avdd.n1865 avdd.t220 243.03
R484 avdd.n1765 avdd.t207 243.03
R485 avdd.n1650 avdd.t210 243.03
R486 avdd.n1855 avdd.t192 243.03
R487 avdd avdd.n7630 242.905
R488 avdd.n4756 avdd.n4487 240
R489 avdd.n4748 avdd.n4487 240
R490 avdd.n4748 avdd.n4507 240
R491 avdd.n4744 avdd.n4507 240
R492 avdd.n4744 avdd.n4743 240
R493 avdd.n4743 avdd.n4510 240
R494 avdd.n4729 avdd.n4510 240
R495 avdd.n4729 avdd.n4529 240
R496 avdd.n4725 avdd.n4529 240
R497 avdd.n4725 avdd.n4532 240
R498 avdd.n4717 avdd.n4532 240
R499 avdd.n4717 avdd.n4543 240
R500 avdd.n4713 avdd.n4543 240
R501 avdd.n4713 avdd.n4545 240
R502 avdd.n4705 avdd.n4545 240
R503 avdd.n4705 avdd.n4551 240
R504 avdd.n4701 avdd.n4551 240
R505 avdd.n4701 avdd.n4553 240
R506 avdd.n4693 avdd.n4553 240
R507 avdd.n4693 avdd.n4559 240
R508 avdd.n4689 avdd.n4559 240
R509 avdd.n4689 avdd.n4688 240
R510 avdd.n4688 avdd.n4562 240
R511 avdd.n4577 avdd.n4562 240
R512 avdd.n4671 avdd.n4577 240
R513 avdd.n4671 avdd.n4578 240
R514 avdd.n4667 avdd.n4578 240
R515 avdd.n4667 avdd.n4582 240
R516 avdd.n4754 avdd.n4490 240
R517 avdd.n4754 avdd.n4491 240
R518 avdd.n4750 avdd.n4491 240
R519 avdd.n4723 avdd.n4535 240
R520 avdd.n4723 avdd.n4536 240
R521 avdd.n4719 avdd.n4536 240
R522 avdd.n4719 avdd.n4541 240
R523 avdd.n4711 avdd.n4541 240
R524 avdd.n4711 avdd.n4547 240
R525 avdd.n4707 avdd.n4547 240
R526 avdd.n4707 avdd.n4549 240
R527 avdd.n4699 avdd.n4549 240
R528 avdd.n4699 avdd.n4554 240
R529 avdd.n4695 avdd.n4554 240
R530 avdd.n4584 avdd.n4575 240
R531 avdd.n4665 avdd.n4584 240
R532 avdd.n4665 avdd.n4585 240
R533 avdd.n4500 avdd.n4492 240
R534 avdd.n4496 avdd.n4494 240
R535 avdd.n7578 avdd.t197 234.554
R536 avdd.n7621 avdd.t198 234.554
R537 avdd.n7537 avdd.t194 234.554
R538 avdd.n7417 avdd.t195 234.554
R539 avdd.n7478 avdd.t228 234.554
R540 avdd.n7521 avdd.t229 234.554
R541 avdd.n7438 avdd.t212 234.554
R542 avdd.n7435 avdd.t213 234.554
R543 avdd.n1685 avdd.t200 234.554
R544 avdd.n1688 avdd.t201 234.554
R545 avdd.n1714 avdd.t215 234.554
R546 avdd.n1759 avdd.t216 234.554
R547 avdd.n1775 avdd.t231 234.554
R548 avdd.n1778 avdd.t232 234.554
R549 avdd.n1804 avdd.t234 234.554
R550 avdd.n1849 avdd.t235 234.554
R551 avdd.n4537 avdd.n4535 229.412
R552 avdd.n4741 avdd.n4513 222.353
R553 avdd.n4764 avdd.n4758 221.774
R554 avdd.n4459 avdd.t6 212.081
R555 avdd.n4460 avdd.t4 212.081
R556 avdd.n4674 avdd.n4575 211.766
R557 avdd.n4695 avdd.n4556 208.236
R558 avdd.n4686 avdd.n4565 204.707
R559 avdd.n4686 avdd.n4566 201.177
R560 avdd.t93 avdd.t89 197.359
R561 avdd.t89 avdd.t101 197.359
R562 avdd.t101 avdd.t96 197.359
R563 avdd.t96 avdd.t102 197.359
R564 avdd.t85 avdd.t99 197.359
R565 avdd.t100 avdd.t85 197.359
R566 avdd.t90 avdd.t100 197.359
R567 avdd.t88 avdd.t90 197.359
R568 avdd.t128 avdd.t142 197.359
R569 avdd.t142 avdd.t136 197.359
R570 avdd.t136 avdd.t144 197.359
R571 avdd.t144 avdd.t139 197.359
R572 avdd.t127 avdd.t133 197.359
R573 avdd.t134 avdd.t127 197.359
R574 avdd.t143 avdd.t134 197.359
R575 avdd.t135 avdd.t143 197.359
R576 avdd.t47 avdd.t40 197.359
R577 avdd.t40 avdd.t41 197.359
R578 avdd.t41 avdd.t52 197.359
R579 avdd.t52 avdd.t42 197.359
R580 avdd.t45 avdd.t35 197.359
R581 avdd.t36 avdd.t45 197.359
R582 avdd.t46 avdd.t36 197.359
R583 avdd.t37 avdd.t46 197.359
R584 avdd.t297 avdd.t308 197.359
R585 avdd.t308 avdd.t302 197.359
R586 avdd.t302 avdd.t305 197.359
R587 avdd.t305 avdd.t298 197.359
R588 avdd.t291 avdd.t306 197.359
R589 avdd.t307 avdd.t291 197.359
R590 avdd.t299 avdd.t307 197.359
R591 avdd.t292 avdd.t299 197.359
R592 avdd.t278 avdd.t285 197.359
R593 avdd.t272 avdd.t278 197.359
R594 avdd.t273 avdd.t272 197.359
R595 avdd.t286 avdd.t273 197.359
R596 avdd.t276 avdd.t279 197.359
R597 avdd.t279 avdd.t277 197.359
R598 avdd.t277 avdd.t269 197.359
R599 avdd.t269 avdd.t280 197.359
R600 avdd.t255 avdd.t244 197.359
R601 avdd.t256 avdd.t255 197.359
R602 avdd.t247 avdd.t256 197.359
R603 avdd.t257 avdd.t247 197.359
R604 avdd.t250 avdd.t242 197.359
R605 avdd.t242 avdd.t251 197.359
R606 avdd.t251 avdd.t243 197.359
R607 avdd.t243 avdd.t252 197.359
R608 avdd.t172 avdd.t176 197.359
R609 avdd.t166 avdd.t172 197.359
R610 avdd.t174 avdd.t166 197.359
R611 avdd.t169 avdd.t174 197.359
R612 avdd.t181 avdd.t175 197.359
R613 avdd.t175 avdd.t182 197.359
R614 avdd.t182 avdd.t173 197.359
R615 avdd.t173 avdd.t165 197.359
R616 avdd.t66 avdd.t70 197.359
R617 avdd.t60 avdd.t66 197.359
R618 avdd.t55 avdd.t60 197.359
R619 avdd.t61 avdd.t55 197.359
R620 avdd.t58 avdd.t62 197.359
R621 avdd.t62 avdd.t59 197.359
R622 avdd.t59 avdd.t67 197.359
R623 avdd.t67 avdd.t63 197.359
R624 avdd.n4659 avdd.n4583 197.329
R625 avdd.n4750 avdd.n4505 190.589
R626 avdd.t86 avdd.t97 190.453
R627 avdd.t94 avdd.t86 190.453
R628 avdd.t91 avdd.t94 190.453
R629 avdd.t113 avdd.t13 190.453
R630 avdd.t119 avdd.t113 190.453
R631 avdd.t103 avdd.t119 190.453
R632 avdd.t137 avdd.t131 190.453
R633 avdd.t129 avdd.t137 190.453
R634 avdd.t140 avdd.t129 190.453
R635 avdd.t117 avdd.t81 190.453
R636 avdd.t75 avdd.t117 190.453
R637 avdd.t266 avdd.t75 190.453
R638 avdd.t50 avdd.t43 190.453
R639 avdd.t43 avdd.t48 190.453
R640 avdd.t48 avdd.t38 190.453
R641 avdd.t147 avdd.t264 190.453
R642 avdd.t264 avdd.t115 190.453
R643 avdd.t115 avdd.t121 190.453
R644 avdd.t295 avdd.t303 190.453
R645 avdd.t300 avdd.t295 190.453
R646 avdd.t293 avdd.t300 190.453
R647 avdd.t183 avdd.t149 190.453
R648 avdd.t11 avdd.t183 190.453
R649 avdd.t260 avdd.t11 190.453
R650 avdd.t64 avdd.t56 190.453
R651 avdd.t53 avdd.t64 190.453
R652 avdd.t68 avdd.t53 190.453
R653 avdd.t237 avdd.t161 190.453
R654 avdd.t309 avdd.t237 190.453
R655 avdd.t25 avdd.t309 190.453
R656 avdd.t167 avdd.t179 190.453
R657 avdd.t177 avdd.t167 190.453
R658 avdd.t170 avdd.t177 190.453
R659 avdd.t23 avdd.t125 190.453
R660 avdd.t105 avdd.t23 190.453
R661 avdd.t258 avdd.t105 190.453
R662 avdd.t248 avdd.t240 190.453
R663 avdd.t240 avdd.t245 190.453
R664 avdd.t245 avdd.t253 190.453
R665 avdd.t79 avdd.t163 190.453
R666 avdd.t163 avdd.t21 190.453
R667 avdd.t21 avdd.t0 190.453
R668 avdd.t283 avdd.t274 190.453
R669 avdd.t270 avdd.t283 190.453
R670 avdd.t281 avdd.t270 190.453
R671 avdd.t15 avdd.t83 190.453
R672 avdd.t262 avdd.t15 190.453
R673 avdd.t145 avdd.t262 190.453
R674 avdd.n4598 avdd.n4590 187.06
R675 avdd.n4732 avdd.n4522 187.06
R676 avdd.n4638 avdd.n4634 187.06
R677 avdd.n4678 avdd.n4569 187.06
R678 avdd.n7632 avdd.n7631 185
R679 avdd.n7629 avdd.n7628 185
R680 avdd.n7531 avdd.n7530 185
R681 avdd.n7529 avdd.n7528 185
R682 avdd.n1857 avdd.n1856 185
R683 avdd.n1769 avdd.n1768 185
R684 avdd.n1767 avdd.n1766 185
R685 avdd.n1866 avdd.n1864 185
R686 avdd.n4596 avdd.n4591 185
R687 avdd.n4591 avdd.n4509 185
R688 avdd.n4515 avdd.n4513 185
R689 avdd.n4513 avdd.n4511 185
R690 avdd.n4525 avdd.n4524 185
R691 avdd.n4526 avdd.n4525 185
R692 avdd.n4522 avdd.n4519 185
R693 avdd.n4527 avdd.n4522 185
R694 avdd.n4538 avdd.n4537 185
R695 avdd.n4537 avdd.n4528 185
R696 avdd.n4523 avdd.n4520 185
R697 avdd.n4730 avdd.n4523 185
R698 avdd.n4556 avdd.n4555 185
R699 avdd.n4558 avdd.n4556 185
R700 avdd.n4619 avdd.n4617 185
R701 avdd.n4635 avdd.n4619 185
R702 avdd.n4678 avdd.n4677 185
R703 avdd.n4679 avdd.n4678 185
R704 avdd.n4676 avdd.n4571 185
R705 avdd.n4571 avdd.n4570 185
R706 avdd.n4683 avdd.n4682 185
R707 avdd.n4682 avdd.n4681 185
R708 avdd.n4684 avdd.n4566 185
R709 avdd.n4566 avdd.n4564 185
R710 avdd.n4632 avdd.n4620 185
R711 avdd.n4620 avdd.n4561 185
R712 avdd.n4634 avdd.n4633 185
R713 avdd.n4636 avdd.n4634 185
R714 avdd.n4590 avdd.n4589 185
R715 avdd.n4600 avdd.n4590 185
R716 avdd.n4603 avdd.n4602 185
R717 avdd.n4602 avdd.n4601 185
R718 avdd.n4741 avdd.n4514 183.53
R719 avdd avdd.n1863 175.585
R720 avdd.n7608 avdd.n7598 174.595
R721 avdd.n7615 avdd.n7595 174.595
R722 avdd.n7411 avdd.n7410 174.595
R723 avdd.n7415 avdd.n7414 174.595
R724 avdd.n7508 avdd.n7498 174.595
R725 avdd.n7515 avdd.n7495 174.595
R726 avdd.n7429 avdd.n7428 174.595
R727 avdd.n7433 avdd.n7432 174.595
R728 avdd.n1695 avdd.n1666 174.595
R729 avdd.n1702 avdd.n1663 174.595
R730 avdd.n1733 avdd.n1732 174.595
R731 avdd.n1737 avdd.n1736 174.595
R732 avdd.n1785 avdd.n1630 174.595
R733 avdd.n1792 avdd.n1627 174.595
R734 avdd.n1823 avdd.n1822 174.595
R735 avdd.n1827 avdd.n1826 174.595
R736 avdd avdd.t91 170.048
R737 avdd avdd.t103 170.048
R738 avdd avdd.t140 170.048
R739 avdd avdd.t266 170.048
R740 avdd.t38 avdd 170.048
R741 avdd.t121 avdd 170.048
R742 avdd avdd.t293 170.048
R743 avdd avdd.t260 170.048
R744 avdd avdd.t68 170.048
R745 avdd avdd.t25 170.048
R746 avdd avdd.t170 170.048
R747 avdd avdd.t258 170.048
R748 avdd.t253 avdd 170.048
R749 avdd.t0 avdd 170.048
R750 avdd avdd.t281 170.048
R751 avdd avdd.t145 170.048
R752 avdd.n7579 avdd.t322 166.282
R753 avdd.n7538 avdd.t321 166.282
R754 avdd.n7479 avdd.t314 166.282
R755 avdd.n7439 avdd.t328 166.282
R756 avdd.n1686 avdd.t311 166.282
R757 avdd.n1715 avdd.t319 166.282
R758 avdd.n1776 avdd.t324 166.282
R759 avdd.n1805 avdd.t315 166.282
R760 avdd.n4769 avdd.t156 158.06
R761 avdd.n4481 avdd.t186 158.06
R762 avdd.n4777 avdd.t160 158.06
R763 avdd.n4477 avdd.t157 158.06
R764 avdd.n4785 avdd.t288 158.06
R765 avdd.n4473 avdd.t74 158.06
R766 avdd.n4793 avdd.t9 158.06
R767 avdd.n4469 avdd.t2 158.06
R768 avdd.n4801 avdd.t7 158.06
R769 avdd.n11 avdd.t10 158.06
R770 avdd.n16 avdd.t72 158.06
R771 avdd.n21 avdd.t77 158.06
R772 avdd.n26 avdd.t151 158.06
R773 avdd.n31 avdd.t268 158.06
R774 avdd.n36 avdd.t123 158.06
R775 avdd.n41 avdd.t112 158.06
R776 avdd.n46 avdd.t110 158.06
R777 avdd.n51 avdd.t217 158.06
R778 avdd.n4482 avdd.t71 155.161
R779 avdd.n4776 avdd.t185 155.161
R780 avdd.n4478 avdd.t159 155.161
R781 avdd.n4784 avdd.t158 155.161
R782 avdd.n4474 avdd.t155 155.161
R783 avdd.n4792 avdd.t287 155.161
R784 avdd.n4470 avdd.t8 155.161
R785 avdd.n4800 avdd.t107 155.161
R786 avdd.n4466 avdd.t5 155.161
R787 avdd.n15 avdd.t239 155.16
R788 avdd.n20 avdd.t73 155.16
R789 avdd.n25 avdd.t78 155.16
R790 avdd.n30 avdd.t152 155.16
R791 avdd.n35 avdd.t3 155.16
R792 avdd.n40 avdd.t124 155.16
R793 avdd.n45 avdd.t27 155.16
R794 avdd.n50 avdd.t111 155.16
R795 avdd.n0 avdd.t236 155.16
R796 avdd.n4462 avdd 152.776
R797 avdd.n7599 avdd.t261 151.123
R798 avdd.n7613 avdd.t294 151.123
R799 avdd.n7569 avdd.t122 151.123
R800 avdd.n7562 avdd.t39 151.123
R801 avdd.n7499 avdd.t267 151.123
R802 avdd.n7513 avdd.t141 151.123
R803 avdd.n7470 avdd.t104 151.123
R804 avdd.n7463 avdd.t92 151.123
R805 avdd.n1664 avdd.t69 151.123
R806 avdd.n1706 avdd.t26 151.123
R807 avdd.n1751 avdd.t171 151.123
R808 avdd.n1744 avdd.t259 151.123
R809 avdd.n1628 avdd.t254 151.123
R810 avdd.n1796 avdd.t1 151.123
R811 avdd.n1841 avdd.t282 151.123
R812 avdd.n1834 avdd.t146 151.123
R813 avdd.n4459 avdd.t323 139.78
R814 avdd.n4460 avdd.t316 139.78
R815 avdd.n4498 avdd.n4488 124.037
R816 avdd.n1816 avdd.n1808 120.001
R817 avdd.n1642 avdd.n1634 120.001
R818 avdd.n1726 avdd.n1718 120.001
R819 avdd.n1678 avdd.n1670 120.001
R820 avdd.n4653 avdd.n4581 105.035
R821 avdd.n4663 avdd.n4662 99.0123
R822 avdd.t102 avdd.n7449 98.6801
R823 avdd.n7449 avdd.t99 98.6801
R824 avdd.t139 avdd.n7488 98.6801
R825 avdd.n7488 avdd.t133 98.6801
R826 avdd.t42 avdd.n7548 98.6801
R827 avdd.n7548 avdd.t35 98.6801
R828 avdd.t298 avdd.n7588 98.6801
R829 avdd.n7588 avdd.t306 98.6801
R830 avdd.n1810 avdd.t286 98.6801
R831 avdd.n1810 avdd.t276 98.6801
R832 avdd.n1636 avdd.t257 98.6801
R833 avdd.n1636 avdd.t250 98.6801
R834 avdd.n1720 avdd.t169 98.6801
R835 avdd.n1720 avdd.t181 98.6801
R836 avdd.n1672 avdd.t61 98.6801
R837 avdd.n1672 avdd.t58 98.6801
R838 avdd.n4755 avdd.n4488 95.8462
R839 avdd.n4755 avdd.n4489 95.8462
R840 avdd.n4724 avdd.n4533 95.8462
R841 avdd.n4724 avdd.n4534 95.8462
R842 avdd.n4718 avdd.n4542 95.8462
R843 avdd.n4712 avdd.n4542 95.8462
R844 avdd.n4712 avdd.n4546 95.8462
R845 avdd.n4706 avdd.n4546 95.8462
R846 avdd.n4706 avdd.n4550 95.8462
R847 avdd.n4700 avdd.n4550 95.8462
R848 avdd.n4694 avdd.n4557 95.8462
R849 avdd.n4672 avdd.n4576 95.8462
R850 avdd.n4666 avdd.n4583 95.8462
R851 avdd.n1861 avdd.n1858 94.8302
R852 avdd.n1655 avdd.n1654 94.8302
R853 avdd.n7426 avdd.t312 92.9047
R854 avdd.n7500 avdd.t313 92.9047
R855 avdd.n7572 avdd.t327 92.9047
R856 avdd.n7600 avdd.t320 92.9047
R857 avdd.n1660 avdd.t325 92.904
R858 avdd.n1739 avdd.t318 92.904
R859 avdd.n1624 avdd.t317 92.904
R860 avdd.n1829 avdd.t326 92.904
R861 avdd.n4502 avdd.n4492 92.5005
R862 avdd.n4498 avdd.n4492 92.5005
R863 avdd.n4501 avdd.n4500 92.5005
R864 avdd.n4494 avdd.n4493 92.5005
R865 avdd.n4496 avdd.n4495 92.5005
R866 avdd.n4486 avdd.n4484 92.5005
R867 avdd.n4741 avdd.n4740 92.5005
R868 avdd.n4742 avdd.n4741 92.5005
R869 avdd.n4539 avdd.n4535 92.5005
R870 avdd.n4535 avdd.n4533 92.5005
R871 avdd.n4723 avdd.n4722 92.5005
R872 avdd.n4724 avdd.n4723 92.5005
R873 avdd.n4721 avdd.n4536 92.5005
R874 avdd.n4536 avdd.n4534 92.5005
R875 avdd.n4720 avdd.n4719 92.5005
R876 avdd.n4719 avdd.n4718 92.5005
R877 avdd.n4541 avdd.n4540 92.5005
R878 avdd.n4542 avdd.n4541 92.5005
R879 avdd.n4711 avdd.n4710 92.5005
R880 avdd.n4712 avdd.n4711 92.5005
R881 avdd.n4709 avdd.n4547 92.5005
R882 avdd.n4547 avdd.n4546 92.5005
R883 avdd.n4708 avdd.n4707 92.5005
R884 avdd.n4707 avdd.n4706 92.5005
R885 avdd.n4549 avdd.n4548 92.5005
R886 avdd.n4550 avdd.n4549 92.5005
R887 avdd.n4699 avdd.n4698 92.5005
R888 avdd.n4700 avdd.n4699 92.5005
R889 avdd.n4697 avdd.n4554 92.5005
R890 avdd.n4557 avdd.n4554 92.5005
R891 avdd.n4696 avdd.n4695 92.5005
R892 avdd.n4695 avdd.n4694 92.5005
R893 avdd.n4663 avdd.n4585 92.5005
R894 avdd.n4585 avdd.n4583 92.5005
R895 avdd.n4665 avdd.n4664 92.5005
R896 avdd.n4666 avdd.n4665 92.5005
R897 avdd.n4647 avdd.n4584 92.5005
R898 avdd.n4584 avdd.n4576 92.5005
R899 avdd.n4646 avdd.n4575 92.5005
R900 avdd.n4672 avdd.n4575 92.5005
R901 avdd.n4686 avdd.n4685 92.5005
R902 avdd.n4687 avdd.n4686 92.5005
R903 avdd.n4751 avdd.n4750 92.5005
R904 avdd.n4750 avdd.n4749 92.5005
R905 avdd.n4752 avdd.n4491 92.5005
R906 avdd.n4491 avdd.n4489 92.5005
R907 avdd.n4754 avdd.n4753 92.5005
R908 avdd.n4755 avdd.n4754 92.5005
R909 avdd.n4503 avdd.n4490 92.5005
R910 avdd.n4490 avdd.n4488 92.5005
R911 avdd.n4653 avdd.n4652 92.5005
R912 avdd.n4655 avdd.n4654 92.5005
R913 avdd.n4657 avdd.n4656 92.5005
R914 avdd.n4649 avdd.n4648 92.5005
R915 avdd.n4662 avdd.n4661 92.5005
R916 avdd.n4757 avdd.n4756 92.5005
R917 avdd.n4756 avdd.n4755 92.5005
R918 avdd.n4487 avdd.n4485 92.5005
R919 avdd.n4489 avdd.n4487 92.5005
R920 avdd.n4748 avdd.n4747 92.5005
R921 avdd.n4749 avdd.n4748 92.5005
R922 avdd.n4601 avdd.n4507 92.5005
R923 avdd.n4746 avdd.n4507 92.5005
R924 avdd.n4744 avdd.n4509 92.5005
R925 avdd.n4745 avdd.n4744 92.5005
R926 avdd.n4743 avdd.n4508 92.5005
R927 avdd.n4743 avdd.n4742 92.5005
R928 avdd.n4526 avdd.n4510 92.5005
R929 avdd.n4530 avdd.n4510 92.5005
R930 avdd.n4730 avdd.n4729 92.5005
R931 avdd.n4729 avdd.n4728 92.5005
R932 avdd.n4727 avdd.n4529 92.5005
R933 avdd.n4533 avdd.n4529 92.5005
R934 avdd.n4726 avdd.n4725 92.5005
R935 avdd.n4725 avdd.n4724 92.5005
R936 avdd.n4532 avdd.n4531 92.5005
R937 avdd.n4534 avdd.n4532 92.5005
R938 avdd.n4717 avdd.n4716 92.5005
R939 avdd.n4718 avdd.n4717 92.5005
R940 avdd.n4715 avdd.n4543 92.5005
R941 avdd.n4543 avdd.n4542 92.5005
R942 avdd.n4714 avdd.n4713 92.5005
R943 avdd.n4713 avdd.n4712 92.5005
R944 avdd.n4545 avdd.n4544 92.5005
R945 avdd.n4546 avdd.n4545 92.5005
R946 avdd.n4705 avdd.n4704 92.5005
R947 avdd.n4706 avdd.n4705 92.5005
R948 avdd.n4703 avdd.n4551 92.5005
R949 avdd.n4551 avdd.n4550 92.5005
R950 avdd.n4702 avdd.n4701 92.5005
R951 avdd.n4701 avdd.n4700 92.5005
R952 avdd.n4553 avdd.n4552 92.5005
R953 avdd.n4557 avdd.n4553 92.5005
R954 avdd.n4693 avdd.n4692 92.5005
R955 avdd.n4694 avdd.n4693 92.5005
R956 avdd.n4635 avdd.n4559 92.5005
R957 avdd.n4691 avdd.n4559 92.5005
R958 avdd.n4689 avdd.n4561 92.5005
R959 avdd.n4690 avdd.n4689 92.5005
R960 avdd.n4688 avdd.n4560 92.5005
R961 avdd.n4688 avdd.n4687 92.5005
R962 avdd.n4681 avdd.n4562 92.5005
R963 avdd.n4579 avdd.n4562 92.5005
R964 avdd.n4577 avdd.n4570 92.5005
R965 avdd.n4580 avdd.n4577 92.5005
R966 avdd.n4671 avdd.n4670 92.5005
R967 avdd.n4672 avdd.n4671 92.5005
R968 avdd.n4669 avdd.n4578 92.5005
R969 avdd.n4578 avdd.n4576 92.5005
R970 avdd.n4668 avdd.n4667 92.5005
R971 avdd.n4667 avdd.n4666 92.5005
R972 avdd.n4582 avdd.n4581 92.5005
R973 avdd.n4583 avdd.n4582 92.5005
R974 avdd.n4533 avdd.n4528 91.6177
R975 avdd.n4742 avdd.n4511 88.7987
R976 avdd.n4660 avdd.n4649 85.7988
R977 avdd.n4654 avdd.n4650 85.7981
R978 avdd.n4673 avdd.n4672 84.5702
R979 avdd.n4694 avdd.n4558 83.1607
R980 avdd.n4687 avdd.n4563 81.7512
R981 avdd.n4687 avdd.n4564 80.3417
R982 avdd.n4503 avdd.n4502 79.4358
R983 avdd avdd.n4763 79.3384
R984 avdd.n4749 avdd.t33 78.9322
R985 avdd.n7451 avdd.n7444 76.5867
R986 avdd.n7490 avdd.n7483 76.5867
R987 avdd.n7550 avdd.n7543 76.5867
R988 avdd.n7590 avdd.n7583 76.5867
R989 avdd.n4749 avdd.n4506 76.1133
R990 avdd.n4600 avdd.n4599 74.7038
R991 avdd.n4731 avdd.n4527 74.7038
R992 avdd.n4637 avdd.n4636 74.7038
R993 avdd.n4680 avdd.n4679 74.7038
R994 avdd.n4461 avdd.n4458 73.5281
R995 avdd.n4742 avdd.n4512 73.2943
R996 avdd.n4658 avdd.n4657 72.7879
R997 avdd.n4654 avdd.n4651 72.7879
R998 avdd.n4657 avdd.n4651 72.7879
R999 avdd.n4658 avdd.n4649 72.7879
R1000 avdd.n4763 avdd.n4762 69.9591
R1001 avdd.n4761 avdd.n4760 68.0792
R1002 avdd.n4557 avdd.t108 62.0183
R1003 avdd.n4759 avdd.t17 61.7334
R1004 avdd.n4460 avdd.n4459 61.346
R1005 avdd.n1862 avdd.n1861 60.1149
R1006 avdd.n1654 avdd.n1651 60.1149
R1007 avdd.n4758 avdd.n4757 57.0603
R1008 avdd.n4525 avdd.n4514 56.4711
R1009 avdd.n4718 avdd.t289 56.3803
R1010 avdd.t30 avdd.n4576 56.3803
R1011 avdd.n4659 avdd.n4651 56.1076
R1012 avdd.n4659 avdd.n4658 56.1076
R1013 avdd.n4499 avdd.n4494 52.2363
R1014 avdd.n4497 avdd.n4486 52.2363
R1015 avdd.n4500 avdd.n4499 52.2363
R1016 avdd.n4497 avdd.n4496 52.2363
R1017 avdd.n4760 avdd.t29 51.9559
R1018 avdd.n4763 avdd.t20 51.9559
R1019 avdd.n4761 avdd.t154 51.9559
R1020 avdd.n4760 avdd.t32 51.2175
R1021 avdd.n1860 avdd.n1859 50.2453
R1022 avdd.n1653 avdd.n1652 50.2453
R1023 avdd.n4763 avdd.t153 50.2329
R1024 avdd.n4761 avdd.t18 50.2329
R1025 avdd.n4602 avdd.n4505 49.4123
R1026 avdd.n4732 avdd.n4523 49.4123
R1027 avdd.n4758 avdd.n4484 47.8123
R1028 avdd.n1863 avdd.n1862 46.2505
R1029 avdd.n1656 avdd.n1655 46.2505
R1030 avdd.n4661 avdd.n4660 42.8997
R1031 avdd.n4652 avdd.n4650 42.8996
R1032 avdd.n4598 avdd.n4591 42.3534
R1033 avdd.t289 avdd.n4534 39.4664
R1034 avdd.n4666 avdd.t30 39.4664
R1035 avdd.n4806 avdd.n4465 39.2858
R1036 avdd.n57 avdd.n56 39.2858
R1037 avdd.n4682 avdd.n4566 38.824
R1038 avdd.n4643 avdd.t31 36.0994
R1039 avdd.n4615 avdd.t109 36.065
R1040 avdd.n4612 avdd.t290 36.065
R1041 avdd.n4587 avdd.t34 36.065
R1042 avdd.n4620 avdd.n4565 35.2946
R1043 avdd.n7609 avdd.n7608 34.6358
R1044 avdd.n7608 avdd.n7607 34.6358
R1045 avdd.n7615 avdd.n7580 34.6358
R1046 avdd.n7615 avdd.n7614 34.6358
R1047 avdd.n7564 avdd.n7411 34.6358
R1048 avdd.n7568 avdd.n7411 34.6358
R1049 avdd.n7557 avdd.n7415 34.6358
R1050 avdd.n7561 avdd.n7415 34.6358
R1051 avdd.n7509 avdd.n7508 34.6358
R1052 avdd.n7508 avdd.n7507 34.6358
R1053 avdd.n7515 avdd.n7480 34.6358
R1054 avdd.n7515 avdd.n7514 34.6358
R1055 avdd.n7465 avdd.n7429 34.6358
R1056 avdd.n7469 avdd.n7429 34.6358
R1057 avdd.n7458 avdd.n7433 34.6358
R1058 avdd.n7462 avdd.n7433 34.6358
R1059 avdd.n1695 avdd.n1694 34.6358
R1060 avdd.n1696 avdd.n1695 34.6358
R1061 avdd.n1702 avdd.n1701 34.6358
R1062 avdd.n1702 avdd.n1661 34.6358
R1063 avdd.n1756 avdd.n1733 34.6358
R1064 avdd.n1752 avdd.n1733 34.6358
R1065 avdd.n1749 avdd.n1737 34.6358
R1066 avdd.n1745 avdd.n1737 34.6358
R1067 avdd.n1785 avdd.n1784 34.6358
R1068 avdd.n1786 avdd.n1785 34.6358
R1069 avdd.n1792 avdd.n1791 34.6358
R1070 avdd.n1792 avdd.n1625 34.6358
R1071 avdd.n1846 avdd.n1823 34.6358
R1072 avdd.n1842 avdd.n1823 34.6358
R1073 avdd.n1839 avdd.n1827 34.6358
R1074 avdd.n1835 avdd.n1827 34.6358
R1075 avdd.n1862 avdd.n1859 34.268
R1076 avdd.n1652 avdd.n1651 34.268
R1077 avdd.n4700 avdd.t108 33.8284
R1078 avdd.n4660 avdd.n4659 33.0688
R1079 avdd.n4659 avdd.n4650 33.0686
R1080 avdd.n4619 avdd.n4556 31.7652
R1081 avdd.n4678 avdd.n4571 31.7652
R1082 avdd.n4768 avdd.n4765 31.624
R1083 avdd.n11 avdd.n10 31.2574
R1084 avdd.n1684 avdd 29.3839
R1085 avdd.n7437 avdd 29.3829
R1086 avdd.n4638 avdd.n4619 28.2358
R1087 avdd.n4674 avdd.n4571 28.2358
R1088 avdd.n7638 avdd.n7637 27.8654
R1089 avdd.n1871 avdd.n1618 27.8654
R1090 avdd.n4769 avdd.n4768 27.1064
R1091 avdd.n7598 avdd.t184 26.5955
R1092 avdd.n7598 avdd.t12 26.5955
R1093 avdd.n7595 avdd.t296 26.5955
R1094 avdd.n7595 avdd.t301 26.5955
R1095 avdd.n7410 avdd.t265 26.5955
R1096 avdd.n7410 avdd.t116 26.5955
R1097 avdd.n7414 avdd.t44 26.5955
R1098 avdd.n7414 avdd.t49 26.5955
R1099 avdd.n7498 avdd.t118 26.5955
R1100 avdd.n7498 avdd.t76 26.5955
R1101 avdd.n7495 avdd.t138 26.5955
R1102 avdd.n7495 avdd.t130 26.5955
R1103 avdd.n7428 avdd.t114 26.5955
R1104 avdd.n7428 avdd.t120 26.5955
R1105 avdd.n7432 avdd.t87 26.5955
R1106 avdd.n7432 avdd.t95 26.5955
R1107 avdd.n1666 avdd.t65 26.5955
R1108 avdd.n1666 avdd.t54 26.5955
R1109 avdd.n1663 avdd.t238 26.5955
R1110 avdd.n1663 avdd.t310 26.5955
R1111 avdd.n1732 avdd.t168 26.5955
R1112 avdd.n1732 avdd.t178 26.5955
R1113 avdd.n1736 avdd.t24 26.5955
R1114 avdd.n1736 avdd.t106 26.5955
R1115 avdd.n1630 avdd.t241 26.5955
R1116 avdd.n1630 avdd.t246 26.5955
R1117 avdd.n1627 avdd.t164 26.5955
R1118 avdd.n1627 avdd.t22 26.5955
R1119 avdd.n1822 avdd.t284 26.5955
R1120 avdd.n1822 avdd.t271 26.5955
R1121 avdd.n1826 avdd.t16 26.5955
R1122 avdd.n1826 avdd.t263 26.5955
R1123 avdd.n4502 avdd.n4501 25.6005
R1124 avdd.n4501 avdd.n4493 25.6005
R1125 avdd.n4495 avdd.n4493 25.6005
R1126 avdd.n4495 avdd.n4484 25.6005
R1127 avdd.n4753 avdd.n4503 25.6005
R1128 avdd.n4753 avdd.n4752 25.6005
R1129 avdd.n4752 avdd.n4751 25.6005
R1130 avdd.n4722 avdd.n4539 25.6005
R1131 avdd.n4722 avdd.n4721 25.6005
R1132 avdd.n4721 avdd.n4720 25.6005
R1133 avdd.n4720 avdd.n4540 25.6005
R1134 avdd.n4710 avdd.n4540 25.6005
R1135 avdd.n4710 avdd.n4709 25.6005
R1136 avdd.n4709 avdd.n4708 25.6005
R1137 avdd.n4708 avdd.n4548 25.6005
R1138 avdd.n4698 avdd.n4548 25.6005
R1139 avdd.n4698 avdd.n4697 25.6005
R1140 avdd.n4697 avdd.n4696 25.6005
R1141 avdd.n4647 avdd.n4646 25.6005
R1142 avdd.n4664 avdd.n4647 25.6005
R1143 avdd.n4664 avdd.n4663 25.6005
R1144 avdd.n4662 avdd.n4648 25.6005
R1145 avdd.n4656 avdd.n4648 25.6005
R1146 avdd.n4656 avdd.n4655 25.6005
R1147 avdd.n4655 avdd.n4653 25.6005
R1148 avdd.n4757 avdd.n4485 25.6005
R1149 avdd.n4747 avdd.n4485 25.6005
R1150 avdd.n4747 avdd.n4746 25.6005
R1151 avdd.n4746 avdd.n4745 25.6005
R1152 avdd.n4745 avdd.n4508 25.6005
R1153 avdd.n4530 avdd.n4508 25.6005
R1154 avdd.n4728 avdd.n4530 25.6005
R1155 avdd.n4728 avdd.n4727 25.6005
R1156 avdd.n4727 avdd.n4726 25.6005
R1157 avdd.n4726 avdd.n4531 25.6005
R1158 avdd.n4716 avdd.n4531 25.6005
R1159 avdd.n4716 avdd.n4715 25.6005
R1160 avdd.n4715 avdd.n4714 25.6005
R1161 avdd.n4714 avdd.n4544 25.6005
R1162 avdd.n4704 avdd.n4544 25.6005
R1163 avdd.n4704 avdd.n4703 25.6005
R1164 avdd.n4703 avdd.n4702 25.6005
R1165 avdd.n4702 avdd.n4552 25.6005
R1166 avdd.n4692 avdd.n4552 25.6005
R1167 avdd.n4692 avdd.n4691 25.6005
R1168 avdd.n4691 avdd.n4690 25.6005
R1169 avdd.n4690 avdd.n4560 25.6005
R1170 avdd.n4579 avdd.n4560 25.6005
R1171 avdd.n4580 avdd.n4579 25.6005
R1172 avdd.n4670 avdd.n4580 25.6005
R1173 avdd.n4670 avdd.n4669 25.6005
R1174 avdd.n4669 avdd.n4668 25.6005
R1175 avdd.n4668 avdd.n4581 25.6005
R1176 avdd.n4466 avdd.n4465 25.6005
R1177 avdd.n56 avdd.n0 25.6005
R1178 avdd.n4461 avdd.n4460 25.3953
R1179 avdd.n4770 avdd.n4482 25.224
R1180 avdd.n4770 avdd.n4769 25.224
R1181 avdd.n4776 avdd.n4480 25.224
R1182 avdd.n4481 avdd.n4480 25.224
R1183 avdd.n4778 avdd.n4478 25.224
R1184 avdd.n4778 avdd.n4777 25.224
R1185 avdd.n4784 avdd.n4476 25.224
R1186 avdd.n4477 avdd.n4476 25.224
R1187 avdd.n4786 avdd.n4474 25.224
R1188 avdd.n4786 avdd.n4785 25.224
R1189 avdd.n4792 avdd.n4472 25.224
R1190 avdd.n4473 avdd.n4472 25.224
R1191 avdd.n4794 avdd.n4470 25.224
R1192 avdd.n4794 avdd.n4793 25.224
R1193 avdd.n4800 avdd.n4468 25.224
R1194 avdd.n4469 avdd.n4468 25.224
R1195 avdd.n4802 avdd.n4466 25.224
R1196 avdd.n4802 avdd.n4801 25.224
R1197 avdd.n11 avdd.n9 25.224
R1198 avdd.n15 avdd.n9 25.224
R1199 avdd.n16 avdd.n8 25.224
R1200 avdd.n20 avdd.n8 25.224
R1201 avdd.n21 avdd.n7 25.224
R1202 avdd.n25 avdd.n7 25.224
R1203 avdd.n26 avdd.n6 25.224
R1204 avdd.n30 avdd.n6 25.224
R1205 avdd.n31 avdd.n5 25.224
R1206 avdd.n35 avdd.n5 25.224
R1207 avdd.n36 avdd.n4 25.224
R1208 avdd.n40 avdd.n4 25.224
R1209 avdd.n41 avdd.n3 25.224
R1210 avdd.n45 avdd.n3 25.224
R1211 avdd.n46 avdd.n2 25.224
R1212 avdd.n50 avdd.n2 25.224
R1213 avdd.n52 avdd.n51 25.224
R1214 avdd.n52 avdd.n0 25.224
R1215 avdd.n4634 avdd.n4620 24.7064
R1216 avdd.n4539 avdd.n4538 24.4711
R1217 avdd.n4740 avdd.n4515 23.7181
R1218 avdd.n4526 avdd.n4512 22.5524
R1219 avdd.n7609 avdd.n7596 22.2123
R1220 avdd.n7607 avdd.n7599 22.2123
R1221 avdd.n7619 avdd.n7580 22.2123
R1222 avdd.n7614 avdd.n7613 22.2123
R1223 avdd.n7564 avdd.n7563 22.2123
R1224 avdd.n7569 avdd.n7568 22.2123
R1225 avdd.n7557 avdd.n7556 22.2123
R1226 avdd.n7562 avdd.n7561 22.2123
R1227 avdd.n7509 avdd.n7496 22.2123
R1228 avdd.n7507 avdd.n7499 22.2123
R1229 avdd.n7519 avdd.n7480 22.2123
R1230 avdd.n7514 avdd.n7513 22.2123
R1231 avdd.n7465 avdd.n7464 22.2123
R1232 avdd.n7470 avdd.n7469 22.2123
R1233 avdd.n7458 avdd.n7457 22.2123
R1234 avdd.n7463 avdd.n7462 22.2123
R1235 avdd.n1694 avdd.n1667 22.2123
R1236 avdd.n1696 avdd.n1664 22.2123
R1237 avdd.n1701 avdd.n1700 22.2123
R1238 avdd.n1706 avdd.n1661 22.2123
R1239 avdd.n1757 avdd.n1756 22.2123
R1240 avdd.n1752 avdd.n1751 22.2123
R1241 avdd.n1750 avdd.n1749 22.2123
R1242 avdd.n1745 avdd.n1744 22.2123
R1243 avdd.n1784 avdd.n1631 22.2123
R1244 avdd.n1786 avdd.n1628 22.2123
R1245 avdd.n1791 avdd.n1790 22.2123
R1246 avdd.n1796 avdd.n1625 22.2123
R1247 avdd.n1847 avdd.n1846 22.2123
R1248 avdd.n1842 avdd.n1841 22.2123
R1249 avdd.n1840 avdd.n1839 22.2123
R1250 avdd.n1835 avdd.n1834 22.2123
R1251 avdd.n4696 avdd.n4555 22.2123
R1252 avdd.n7620 avdd.n7619 21.8029
R1253 avdd.n7556 avdd.n7555 21.8029
R1254 avdd.n7520 avdd.n7519 21.8029
R1255 avdd.n7457 avdd.n7456 21.8029
R1256 avdd.n1689 avdd.n1667 21.8029
R1257 avdd.n1758 avdd.n1757 21.8029
R1258 avdd.n1779 avdd.n1631 21.8029
R1259 avdd.n1848 avdd.n1847 21.8029
R1260 avdd.n4685 avdd.n4684 21.4593
R1261 avdd.n4682 avdd.n4569 21.177
R1262 avdd.n7613 avdd.n7596 21.0829
R1263 avdd.n7563 avdd.n7562 21.0829
R1264 avdd.n7513 avdd.n7496 21.0829
R1265 avdd.n7464 avdd.n7463 21.0829
R1266 avdd.n1700 avdd.n1664 21.0829
R1267 avdd.n1751 avdd.n1750 21.0829
R1268 avdd.n1790 avdd.n1628 21.0829
R1269 avdd.n1841 avdd.n1840 21.0829
R1270 avdd.n4474 avdd.n4473 20.3299
R1271 avdd.n36 avdd.n35 20.3299
R1272 avdd.n4499 avdd.n4498 20.1334
R1273 avdd.n4498 avdd.n4497 20.1334
R1274 avdd.n4482 avdd.n4481 19.9534
R1275 avdd.n4478 avdd.n4477 19.9534
R1276 avdd.n4785 avdd.n4784 19.9534
R1277 avdd.n4793 avdd.n4792 19.9534
R1278 avdd.n4801 avdd.n4800 19.9534
R1279 avdd.n16 avdd.n15 19.9534
R1280 avdd.n26 avdd.n25 19.9534
R1281 avdd.n31 avdd.n30 19.9534
R1282 avdd.n41 avdd.n40 19.9534
R1283 avdd.n51 avdd.n50 19.9534
R1284 avdd.n4601 avdd.n4506 19.7334
R1285 avdd.n4731 avdd.n4730 19.7334
R1286 avdd.n4777 avdd.n4776 19.577
R1287 avdd.n4470 avdd.n4469 19.577
R1288 avdd.n21 avdd.n20 19.577
R1289 avdd.n46 avdd.n45 19.577
R1290 avdd.n1817 avdd.n1807 19.0999
R1291 avdd.n1643 avdd.n1633 19.0999
R1292 avdd.n1727 avdd.n1717 19.0999
R1293 avdd.n1679 avdd.n1669 19.0999
R1294 avdd.n4591 avdd.n4513 17.6476
R1295 avdd.n7446 avdd.n7442 17.2966
R1296 avdd.n7485 avdd.n7481 17.2966
R1297 avdd.n7545 avdd.n7541 17.2966
R1298 avdd.n7585 avdd.n7581 17.2966
R1299 avdd.n1859 avdd.n1858 17.1345
R1300 avdd.n1655 avdd.n1652 17.1345
R1301 avdd.n7452 avdd.n7443 16.9954
R1302 avdd.n7491 avdd.n7482 16.9954
R1303 avdd.n7551 avdd.n7542 16.9954
R1304 avdd.n7591 avdd.n7582 16.9954
R1305 avdd.n1813 avdd.n1806 16.9954
R1306 avdd.n1639 avdd.n1632 16.9954
R1307 avdd.n1723 avdd.n1716 16.9954
R1308 avdd.n1675 avdd.n1668 16.9954
R1309 avdd.t33 avdd.n4489 16.9144
R1310 avdd.n4599 avdd.n4509 16.9144
R1311 avdd.n4646 avdd.n4645 16.1887
R1312 avdd.n4681 avdd.n4564 15.505
R1313 avdd.n7603 avdd.n7599 15.4358
R1314 avdd.n7570 avdd.n7569 15.4358
R1315 avdd.n7503 avdd.n7499 15.4358
R1316 avdd.n7471 avdd.n7470 15.4358
R1317 avdd.n1707 avdd.n1706 15.4358
R1318 avdd.n1744 avdd.n1743 15.4358
R1319 avdd.n1797 avdd.n1796 15.4358
R1320 avdd.n1834 avdd.n1833 15.4358
R1321 avdd.n4685 avdd.n4567 15.4358
R1322 avdd.n7626 avdd.n7407 14.2735
R1323 avdd.n7536 avdd.n7535 14.2735
R1324 avdd.n7526 avdd.n7424 14.2735
R1325 avdd.n1764 avdd.n1658 14.2735
R1326 avdd.n1774 avdd.n1647 14.2735
R1327 avdd.n1854 avdd.n1622 14.2735
R1328 avdd.n4563 avdd.n4561 14.0955
R1329 avdd.n4751 avdd.n4504 13.9299
R1330 avdd.n4592 avdd.n4589 13.5534
R1331 avdd.n4735 avdd.n4519 13.5534
R1332 avdd.n4633 avdd.n4621 13.5534
R1333 avdd.n4677 avdd.n4572 13.5534
R1334 avdd.n4740 avdd.n4739 13.177
R1335 avdd.n4635 avdd.n4558 12.686
R1336 avdd.n4679 avdd.n4570 12.686
R1337 avdd.n7453 avdd.n7442 12.4392
R1338 avdd.n7492 avdd.n7481 12.4392
R1339 avdd.n7552 avdd.n7541 12.4392
R1340 avdd.n7592 avdd.n7581 12.4392
R1341 avdd.n1818 avdd.n1817 12.4348
R1342 avdd.n1644 avdd.n1643 12.4348
R1343 avdd.n1728 avdd.n1727 12.4348
R1344 avdd.n1680 avdd.n1679 12.4348
R1345 avdd.n4637 avdd.n4635 11.2765
R1346 avdd.n4673 avdd.n4570 11.2765
R1347 avdd.n4762 avdd.n4761 11.2557
R1348 avdd.n4602 avdd.n4590 10.5887
R1349 avdd.n4537 avdd.n4523 10.5887
R1350 avdd.n4636 avdd.n4561 9.86697
R1351 avdd.n7451 avdd.n7450 9.3005
R1352 avdd.n7490 avdd.n7489 9.3005
R1353 avdd.n7550 avdd.n7549 9.3005
R1354 avdd.n7590 avdd.n7589 9.3005
R1355 avdd.n4463 avdd.n4462 9.3005
R1356 avdd.n4607 avdd.n4504 9.3005
R1357 avdd.n4604 avdd.n4588 9.3005
R1358 avdd.n4604 avdd.n4505 9.3005
R1359 avdd.n4506 avdd.n4505 9.3005
R1360 avdd.n4597 avdd.n4517 9.3005
R1361 avdd.n4598 avdd.n4597 9.3005
R1362 avdd.n4599 avdd.n4598 9.3005
R1363 avdd.n4734 avdd.n4518 9.3005
R1364 avdd.n4606 avdd.n4605 9.3005
R1365 avdd.n4586 avdd.n4573 9.3005
R1366 avdd.n4626 avdd.n4625 9.3005
R1367 avdd.n4629 avdd.n4622 9.3005
R1368 avdd.n4640 avdd.n4639 9.3005
R1369 avdd.n4639 avdd.n4638 9.3005
R1370 avdd.n4638 avdd.n4637 9.3005
R1371 avdd.n4631 avdd.n4630 9.3005
R1372 avdd.n4631 avdd.n4565 9.3005
R1373 avdd.n4565 avdd.n4563 9.3005
R1374 avdd.n4737 avdd.n4516 9.3005
R1375 avdd.n4516 avdd.n4514 9.3005
R1376 avdd.n4514 avdd.n4512 9.3005
R1377 avdd.n4736 avdd.n4735 9.3005
R1378 avdd.n4733 avdd.n4521 9.3005
R1379 avdd.n4733 avdd.n4732 9.3005
R1380 avdd.n4732 avdd.n4731 9.3005
R1381 avdd.n4628 avdd.n4567 9.3005
R1382 avdd.n4627 avdd.n4568 9.3005
R1383 avdd.n4569 avdd.n4568 9.3005
R1384 avdd.n4680 avdd.n4569 9.3005
R1385 avdd.n4624 avdd.n4572 9.3005
R1386 avdd.n4645 avdd.n4644 9.3005
R1387 avdd.n4675 avdd.n4574 9.3005
R1388 avdd.n4675 avdd.n4674 9.3005
R1389 avdd.n4674 avdd.n4673 9.3005
R1390 avdd.n4623 avdd.n4621 9.3005
R1391 avdd.n4618 avdd.n4616 9.3005
R1392 avdd.n4595 avdd.n4594 9.3005
R1393 avdd.n4593 avdd.n4592 9.3005
R1394 avdd.n1913 avdd.n1901 9.0005
R1395 avdd.n1918 avdd.n1917 9.0005
R1396 avdd.n1915 avdd.n1914 9.0005
R1397 avdd.n1916 avdd.n1900 9.0005
R1398 avdd.n2167 avdd.n2155 9.0005
R1399 avdd.n2172 avdd.n2171 9.0005
R1400 avdd.n2169 avdd.n2168 9.0005
R1401 avdd.n2170 avdd.n2154 9.0005
R1402 avdd.n2382 avdd.n2370 9.0005
R1403 avdd.n2387 avdd.n2386 9.0005
R1404 avdd.n2384 avdd.n2383 9.0005
R1405 avdd.n2385 avdd.n2369 9.0005
R1406 avdd.n2597 avdd.n2585 9.0005
R1407 avdd.n2602 avdd.n2601 9.0005
R1408 avdd.n2599 avdd.n2598 9.0005
R1409 avdd.n2600 avdd.n2584 9.0005
R1410 avdd.n2812 avdd.n2800 9.0005
R1411 avdd.n2817 avdd.n2816 9.0005
R1412 avdd.n2814 avdd.n2813 9.0005
R1413 avdd.n2815 avdd.n2799 9.0005
R1414 avdd.n3027 avdd.n3015 9.0005
R1415 avdd.n3032 avdd.n3031 9.0005
R1416 avdd.n3029 avdd.n3028 9.0005
R1417 avdd.n3030 avdd.n3014 9.0005
R1418 avdd.n3203 avdd.n3191 9.0005
R1419 avdd.n3208 avdd.n3207 9.0005
R1420 avdd.n3205 avdd.n3204 9.0005
R1421 avdd.n3206 avdd.n3190 9.0005
R1422 avdd.n3418 avdd.n3406 9.0005
R1423 avdd.n3423 avdd.n3422 9.0005
R1424 avdd.n3420 avdd.n3419 9.0005
R1425 avdd.n3421 avdd.n3405 9.0005
R1426 avdd.n3633 avdd.n3621 9.0005
R1427 avdd.n3638 avdd.n3637 9.0005
R1428 avdd.n3635 avdd.n3634 9.0005
R1429 avdd.n3636 avdd.n3620 9.0005
R1430 avdd.n3848 avdd.n3836 9.0005
R1431 avdd.n3853 avdd.n3852 9.0005
R1432 avdd.n3850 avdd.n3849 9.0005
R1433 avdd.n3851 avdd.n3835 9.0005
R1434 avdd.n4063 avdd.n4051 9.0005
R1435 avdd.n4068 avdd.n4067 9.0005
R1436 avdd.n4065 avdd.n4064 9.0005
R1437 avdd.n4066 avdd.n4050 9.0005
R1438 avdd.n4278 avdd.n4266 9.0005
R1439 avdd.n4283 avdd.n4282 9.0005
R1440 avdd.n4280 avdd.n4279 9.0005
R1441 avdd.n4281 avdd.n4265 9.0005
R1442 avdd.n4892 avdd.n4876 9.0005
R1443 avdd.n4891 avdd.n4890 9.0005
R1444 avdd.n4889 avdd.n4877 9.0005
R1445 avdd.n4894 avdd.n4893 9.0005
R1446 avdd.n5108 avdd.n5092 9.0005
R1447 avdd.n5107 avdd.n5106 9.0005
R1448 avdd.n5105 avdd.n5093 9.0005
R1449 avdd.n5110 avdd.n5109 9.0005
R1450 avdd.n5324 avdd.n5308 9.0005
R1451 avdd.n5323 avdd.n5322 9.0005
R1452 avdd.n5321 avdd.n5309 9.0005
R1453 avdd.n5326 avdd.n5325 9.0005
R1454 avdd.n5540 avdd.n5524 9.0005
R1455 avdd.n5539 avdd.n5538 9.0005
R1456 avdd.n5537 avdd.n5525 9.0005
R1457 avdd.n5542 avdd.n5541 9.0005
R1458 avdd.n5756 avdd.n5740 9.0005
R1459 avdd.n5755 avdd.n5754 9.0005
R1460 avdd.n5753 avdd.n5741 9.0005
R1461 avdd.n5758 avdd.n5757 9.0005
R1462 avdd.n5972 avdd.n5956 9.0005
R1463 avdd.n5971 avdd.n5970 9.0005
R1464 avdd.n5969 avdd.n5957 9.0005
R1465 avdd.n5974 avdd.n5973 9.0005
R1466 avdd.n6188 avdd.n6172 9.0005
R1467 avdd.n6187 avdd.n6186 9.0005
R1468 avdd.n6185 avdd.n6173 9.0005
R1469 avdd.n6190 avdd.n6189 9.0005
R1470 avdd.n6404 avdd.n6388 9.0005
R1471 avdd.n6403 avdd.n6402 9.0005
R1472 avdd.n6401 avdd.n6389 9.0005
R1473 avdd.n6406 avdd.n6405 9.0005
R1474 avdd.n6620 avdd.n6604 9.0005
R1475 avdd.n6619 avdd.n6618 9.0005
R1476 avdd.n6617 avdd.n6605 9.0005
R1477 avdd.n6622 avdd.n6621 9.0005
R1478 avdd.n6836 avdd.n6820 9.0005
R1479 avdd.n6835 avdd.n6834 9.0005
R1480 avdd.n6833 avdd.n6821 9.0005
R1481 avdd.n6838 avdd.n6837 9.0005
R1482 avdd.n7052 avdd.n7036 9.0005
R1483 avdd.n7051 avdd.n7050 9.0005
R1484 avdd.n7049 avdd.n7037 9.0005
R1485 avdd.n7054 avdd.n7053 9.0005
R1486 avdd.n7268 avdd.n7252 9.0005
R1487 avdd.n7267 avdd.n7266 9.0005
R1488 avdd.n7265 avdd.n7253 9.0005
R1489 avdd.n7270 avdd.n7269 9.0005
R1490 avdd.n1809 avdd.n1808 8.84285
R1491 avdd.n1635 avdd.n1634 8.84285
R1492 avdd.n1719 avdd.n1718 8.84285
R1493 avdd.n1671 avdd.n1670 8.84285
R1494 avdd.n4681 avdd.n4680 8.45747
R1495 avdd.n7535 avdd.n7419 7.70175
R1496 avdd.n7627 avdd.n7626 7.70175
R1497 avdd.n7637 avdd.n7403 7.70175
R1498 avdd.n7527 avdd.n7526 7.70175
R1499 avdd.n1865 avdd.n1618 7.70175
R1500 avdd.n1765 avdd.n1764 7.70175
R1501 avdd.n1650 avdd.n1647 7.70175
R1502 avdd.n1855 avdd.n1854 7.70175
R1503 avdd.n7452 avdd.n7451 7.66611
R1504 avdd.n7491 avdd.n7490 7.66611
R1505 avdd.n7551 avdd.n7550 7.66611
R1506 avdd.n7591 avdd.n7590 7.66611
R1507 avdd.n1808 avdd.n1806 7.66611
R1508 avdd.n1634 avdd.n1632 7.66611
R1509 avdd.n1718 avdd.n1716 7.66611
R1510 avdd.n1670 avdd.n1668 7.66611
R1511 avdd.n4462 avdd.n4461 7.13769
R1512 avdd.n4511 avdd.n4509 7.04798
R1513 avdd.n4807 avdd.n4464 7.00334
R1514 avdd.n4739 avdd.n4516 6.4005
R1515 avdd.n4524 avdd.n4516 6.02403
R1516 avdd.n4605 avdd.n4604 5.64756
R1517 avdd.n4734 avdd.n4733 5.64756
R1518 avdd.n4604 avdd.n4603 5.27109
R1519 avdd.n4733 avdd.n4520 5.27109
R1520 avdd.n4597 avdd.n4595 4.89462
R1521 avdd.n1861 avdd.n1860 4.65934
R1522 avdd.n1654 avdd.n1653 4.65934
R1523 avdd.n7457 avdd.n7434 4.6505
R1524 avdd.n7463 avdd.n7431 4.6505
R1525 avdd.n7464 avdd.n7430 4.6505
R1526 avdd.n7470 avdd.n7427 4.6505
R1527 avdd.n7524 avdd.n7424 4.6505
R1528 avdd.n7519 avdd.n7518 4.6505
R1529 avdd.n7513 avdd.n7512 4.6505
R1530 avdd.n7511 avdd.n7496 4.6505
R1531 avdd.n7505 avdd.n7499 4.6505
R1532 avdd.n7536 avdd.n7418 4.6505
R1533 avdd.n7556 avdd.n7416 4.6505
R1534 avdd.n7562 avdd.n7413 4.6505
R1535 avdd.n7563 avdd.n7412 4.6505
R1536 avdd.n7569 avdd.n7409 4.6505
R1537 avdd.n7624 avdd.n7407 4.6505
R1538 avdd.n7619 avdd.n7618 4.6505
R1539 avdd.n7613 avdd.n7612 4.6505
R1540 avdd.n7611 avdd.n7596 4.6505
R1541 avdd.n7605 avdd.n7599 4.6505
R1542 avdd.n7437 avdd.n7436 4.6505
R1543 avdd.n7441 avdd.n7440 4.6505
R1544 avdd.n7456 avdd.n7455 4.6505
R1545 avdd.n7459 avdd.n7458 4.6505
R1546 avdd.n7460 avdd.n7433 4.6505
R1547 avdd.n7462 avdd.n7461 4.6505
R1548 avdd.n7466 avdd.n7465 4.6505
R1549 avdd.n7467 avdd.n7429 4.6505
R1550 avdd.n7469 avdd.n7468 4.6505
R1551 avdd.n7475 avdd.n7474 4.6505
R1552 avdd.n7476 avdd.n7423 4.6505
R1553 avdd.n7523 avdd.n7522 4.6505
R1554 avdd.n7520 avdd.n7477 4.6505
R1555 avdd.n7517 avdd.n7480 4.6505
R1556 avdd.n7516 avdd.n7515 4.6505
R1557 avdd.n7514 avdd.n7494 4.6505
R1558 avdd.n7510 avdd.n7509 4.6505
R1559 avdd.n7508 avdd.n7497 4.6505
R1560 avdd.n7507 avdd.n7506 4.6505
R1561 avdd.n7421 avdd.n7420 4.6505
R1562 avdd.n7533 avdd.n7532 4.6505
R1563 avdd.n7540 avdd.n7539 4.6505
R1564 avdd.n7555 avdd.n7554 4.6505
R1565 avdd.n7558 avdd.n7557 4.6505
R1566 avdd.n7559 avdd.n7415 4.6505
R1567 avdd.n7561 avdd.n7560 4.6505
R1568 avdd.n7565 avdd.n7564 4.6505
R1569 avdd.n7566 avdd.n7411 4.6505
R1570 avdd.n7568 avdd.n7567 4.6505
R1571 avdd.n7575 avdd.n7574 4.6505
R1572 avdd.n7576 avdd.n7406 4.6505
R1573 avdd.n7623 avdd.n7622 4.6505
R1574 avdd.n7620 avdd.n7577 4.6505
R1575 avdd.n7617 avdd.n7580 4.6505
R1576 avdd.n7616 avdd.n7615 4.6505
R1577 avdd.n7614 avdd.n7594 4.6505
R1578 avdd.n7610 avdd.n7609 4.6505
R1579 avdd.n7608 avdd.n7597 4.6505
R1580 avdd.n7607 avdd.n7606 4.6505
R1581 avdd.n7405 avdd.n7404 4.6505
R1582 avdd.n7634 avdd.n7633 4.6505
R1583 avdd.n1834 avdd.n1828 4.6505
R1584 avdd.n1840 avdd.n1825 4.6505
R1585 avdd.n1841 avdd.n1824 4.6505
R1586 avdd.n1847 avdd.n1821 4.6505
R1587 avdd.n1796 avdd.n1795 4.6505
R1588 avdd.n1790 avdd.n1789 4.6505
R1589 avdd.n1788 avdd.n1628 4.6505
R1590 avdd.n1782 avdd.n1631 4.6505
R1591 avdd.n1744 avdd.n1738 4.6505
R1592 avdd.n1750 avdd.n1735 4.6505
R1593 avdd.n1751 avdd.n1734 4.6505
R1594 avdd.n1757 avdd.n1731 4.6505
R1595 avdd.n1706 avdd.n1705 4.6505
R1596 avdd.n1700 avdd.n1699 4.6505
R1597 avdd.n1698 avdd.n1664 4.6505
R1598 avdd.n1692 avdd.n1667 4.6505
R1599 avdd.n1711 avdd.n1710 4.6505
R1600 avdd.n1712 avdd.n1657 4.6505
R1601 avdd.n1649 avdd.n1648 4.6505
R1602 avdd.n1771 avdd.n1770 4.6505
R1603 avdd.n1801 avdd.n1800 4.6505
R1604 avdd.n1802 avdd.n1621 4.6505
R1605 avdd.n1620 avdd.n1619 4.6505
R1606 avdd.n1868 avdd.n1867 4.6505
R1607 avdd.n1836 avdd.n1835 4.6505
R1608 avdd.n1837 avdd.n1827 4.6505
R1609 avdd.n1839 avdd.n1838 4.6505
R1610 avdd.n1843 avdd.n1842 4.6505
R1611 avdd.n1844 avdd.n1823 4.6505
R1612 avdd.n1846 avdd.n1845 4.6505
R1613 avdd.n1848 avdd.n1803 4.6505
R1614 avdd.n1851 avdd.n1850 4.6505
R1615 avdd.n1852 avdd.n1622 4.6505
R1616 avdd.n1794 avdd.n1625 4.6505
R1617 avdd.n1793 avdd.n1792 4.6505
R1618 avdd.n1791 avdd.n1626 4.6505
R1619 avdd.n1787 avdd.n1786 4.6505
R1620 avdd.n1785 avdd.n1629 4.6505
R1621 avdd.n1784 avdd.n1783 4.6505
R1622 avdd.n1780 avdd.n1779 4.6505
R1623 avdd.n1777 avdd.n1646 4.6505
R1624 avdd.n1774 avdd.n1773 4.6505
R1625 avdd.n1746 avdd.n1745 4.6505
R1626 avdd.n1747 avdd.n1737 4.6505
R1627 avdd.n1749 avdd.n1748 4.6505
R1628 avdd.n1753 avdd.n1752 4.6505
R1629 avdd.n1754 avdd.n1733 4.6505
R1630 avdd.n1756 avdd.n1755 4.6505
R1631 avdd.n1758 avdd.n1713 4.6505
R1632 avdd.n1761 avdd.n1760 4.6505
R1633 avdd.n1762 avdd.n1658 4.6505
R1634 avdd.n1704 avdd.n1661 4.6505
R1635 avdd.n1703 avdd.n1702 4.6505
R1636 avdd.n1701 avdd.n1662 4.6505
R1637 avdd.n1697 avdd.n1696 4.6505
R1638 avdd.n1695 avdd.n1665 4.6505
R1639 avdd.n1694 avdd.n1693 4.6505
R1640 avdd.n1690 avdd.n1689 4.6505
R1641 avdd.n1687 avdd.n1682 4.6505
R1642 avdd.n1684 avdd.n1683 4.6505
R1643 avdd.n4739 avdd.n4738 4.6505
R1644 avdd.n4804 avdd.n4466 4.6505
R1645 avdd.n4801 avdd.n4467 4.6505
R1646 avdd.n4800 avdd.n4799 4.6505
R1647 avdd.n4797 avdd.n4469 4.6505
R1648 avdd.n4796 avdd.n4470 4.6505
R1649 avdd.n4793 avdd.n4471 4.6505
R1650 avdd.n4792 avdd.n4791 4.6505
R1651 avdd.n4789 avdd.n4473 4.6505
R1652 avdd.n4788 avdd.n4474 4.6505
R1653 avdd.n4785 avdd.n4475 4.6505
R1654 avdd.n4784 avdd.n4783 4.6505
R1655 avdd.n4781 avdd.n4477 4.6505
R1656 avdd.n4780 avdd.n4478 4.6505
R1657 avdd.n4777 avdd.n4479 4.6505
R1658 avdd.n4776 avdd.n4775 4.6505
R1659 avdd.n4773 avdd.n4481 4.6505
R1660 avdd.n4772 avdd.n4482 4.6505
R1661 avdd.n4769 avdd.n4483 4.6505
R1662 avdd.n4805 avdd.n4465 4.6505
R1663 avdd.n4803 avdd.n4802 4.6505
R1664 avdd.n4798 avdd.n4468 4.6505
R1665 avdd.n4795 avdd.n4794 4.6505
R1666 avdd.n4790 avdd.n4472 4.6505
R1667 avdd.n4787 avdd.n4786 4.6505
R1668 avdd.n4782 avdd.n4476 4.6505
R1669 avdd.n4779 avdd.n4778 4.6505
R1670 avdd.n4774 avdd.n4480 4.6505
R1671 avdd.n4771 avdd.n4770 4.6505
R1672 avdd.n4768 avdd.n4767 4.6505
R1673 avdd.n4766 avdd.n4765 4.6505
R1674 avdd.n54 avdd.n0 4.6505
R1675 avdd.n51 avdd.n1 4.6505
R1676 avdd.n50 avdd.n49 4.6505
R1677 avdd.n47 avdd.n46 4.6505
R1678 avdd.n45 avdd.n44 4.6505
R1679 avdd.n42 avdd.n41 4.6505
R1680 avdd.n40 avdd.n39 4.6505
R1681 avdd.n37 avdd.n36 4.6505
R1682 avdd.n35 avdd.n34 4.6505
R1683 avdd.n32 avdd.n31 4.6505
R1684 avdd.n30 avdd.n29 4.6505
R1685 avdd.n27 avdd.n26 4.6505
R1686 avdd.n25 avdd.n24 4.6505
R1687 avdd.n22 avdd.n21 4.6505
R1688 avdd.n20 avdd.n19 4.6505
R1689 avdd.n17 avdd.n16 4.6505
R1690 avdd.n15 avdd.n14 4.6505
R1691 avdd.n12 avdd.n11 4.6505
R1692 avdd.n56 avdd.n55 4.6505
R1693 avdd.n53 avdd.n52 4.6505
R1694 avdd.n48 avdd.n2 4.6505
R1695 avdd.n43 avdd.n3 4.6505
R1696 avdd.n38 avdd.n4 4.6505
R1697 avdd.n33 avdd.n5 4.6505
R1698 avdd.n28 avdd.n6 4.6505
R1699 avdd.n23 avdd.n7 4.6505
R1700 avdd.n18 avdd.n8 4.6505
R1701 avdd.n13 avdd.n9 4.6505
R1702 avdd.n4587 avdd 4.5906
R1703 avdd.n4615 avdd.n4614 4.56717
R1704 avdd.n4613 avdd.n4612 4.56717
R1705 avdd.n2049 avdd.n2048 4.52183
R1706 avdd.n2053 avdd.n1974 4.52183
R1707 avdd.n1936 avdd.n1933 4.52183
R1708 avdd.n2268 avdd.n2262 4.52183
R1709 avdd.n2247 avdd.n2243 4.52183
R1710 avdd.n2192 avdd.n2186 4.52183
R1711 avdd.n2483 avdd.n2477 4.52183
R1712 avdd.n2462 avdd.n2458 4.52183
R1713 avdd.n2407 avdd.n2401 4.52183
R1714 avdd.n2698 avdd.n2692 4.52183
R1715 avdd.n2677 avdd.n2673 4.52183
R1716 avdd.n2622 avdd.n2616 4.52183
R1717 avdd.n2913 avdd.n2907 4.52183
R1718 avdd.n2892 avdd.n2888 4.52183
R1719 avdd.n2837 avdd.n2831 4.52183
R1720 avdd.n3128 avdd.n3122 4.52183
R1721 avdd.n3107 avdd.n3103 4.52183
R1722 avdd.n3052 avdd.n3046 4.52183
R1723 avdd.n3338 avdd.n3337 4.52183
R1724 avdd.n3342 avdd.n3264 4.52183
R1725 avdd.n3226 avdd.n3223 4.52183
R1726 avdd.n3553 avdd.n3552 4.52183
R1727 avdd.n3557 avdd.n3479 4.52183
R1728 avdd.n3441 avdd.n3438 4.52183
R1729 avdd.n3768 avdd.n3767 4.52183
R1730 avdd.n3772 avdd.n3694 4.52183
R1731 avdd.n3656 avdd.n3653 4.52183
R1732 avdd.n3983 avdd.n3982 4.52183
R1733 avdd.n3987 avdd.n3909 4.52183
R1734 avdd.n3871 avdd.n3868 4.52183
R1735 avdd.n4198 avdd.n4197 4.52183
R1736 avdd.n4202 avdd.n4124 4.52183
R1737 avdd.n4086 avdd.n4083 4.52183
R1738 avdd.n4413 avdd.n4412 4.52183
R1739 avdd.n4417 avdd.n4339 4.52183
R1740 avdd.n4301 avdd.n4298 4.52183
R1741 avdd.n4915 avdd.n4909 4.52183
R1742 avdd.n4969 avdd.n4965 4.52183
R1743 avdd.n4990 avdd.n4984 4.52183
R1744 avdd.n5131 avdd.n5125 4.52183
R1745 avdd.n5185 avdd.n5181 4.52183
R1746 avdd.n5206 avdd.n5200 4.52183
R1747 avdd.n5347 avdd.n5341 4.52183
R1748 avdd.n5401 avdd.n5397 4.52183
R1749 avdd.n5422 avdd.n5416 4.52183
R1750 avdd.n5563 avdd.n5557 4.52183
R1751 avdd.n5617 avdd.n5613 4.52183
R1752 avdd.n5638 avdd.n5632 4.52183
R1753 avdd.n5779 avdd.n5773 4.52183
R1754 avdd.n5833 avdd.n5829 4.52183
R1755 avdd.n5854 avdd.n5848 4.52183
R1756 avdd.n5995 avdd.n5989 4.52183
R1757 avdd.n6049 avdd.n6045 4.52183
R1758 avdd.n6070 avdd.n6064 4.52183
R1759 avdd.n6211 avdd.n6205 4.52183
R1760 avdd.n6265 avdd.n6261 4.52183
R1761 avdd.n6286 avdd.n6280 4.52183
R1762 avdd.n6427 avdd.n6421 4.52183
R1763 avdd.n6481 avdd.n6477 4.52183
R1764 avdd.n6502 avdd.n6496 4.52183
R1765 avdd.n6643 avdd.n6637 4.52183
R1766 avdd.n6697 avdd.n6693 4.52183
R1767 avdd.n6718 avdd.n6712 4.52183
R1768 avdd.n6859 avdd.n6853 4.52183
R1769 avdd.n6913 avdd.n6909 4.52183
R1770 avdd.n6934 avdd.n6928 4.52183
R1771 avdd.n7075 avdd.n7069 4.52183
R1772 avdd.n7129 avdd.n7125 4.52183
R1773 avdd.n7150 avdd.n7144 4.52183
R1774 avdd.n7291 avdd.n7285 4.52183
R1775 avdd.n7345 avdd.n7341 4.52183
R1776 avdd.n7366 avdd.n7360 4.52183
R1777 avdd.n4597 avdd.n4596 4.51815
R1778 avdd.n4625 avdd.n4572 4.51815
R1779 avdd.n2019 avdd.n2018 4.51805
R1780 avdd.n1968 avdd.n1967 4.51805
R1781 avdd.n2077 avdd.n2076 4.51805
R1782 avdd.n2293 avdd.n2292 4.51805
R1783 avdd.n2222 avdd.n2126 4.51805
R1784 avdd.n2220 avdd.n2219 4.51805
R1785 avdd.n2508 avdd.n2507 4.51805
R1786 avdd.n2437 avdd.n2341 4.51805
R1787 avdd.n2435 avdd.n2434 4.51805
R1788 avdd.n2723 avdd.n2722 4.51805
R1789 avdd.n2652 avdd.n2556 4.51805
R1790 avdd.n2650 avdd.n2649 4.51805
R1791 avdd.n2938 avdd.n2937 4.51805
R1792 avdd.n2867 avdd.n2771 4.51805
R1793 avdd.n2865 avdd.n2864 4.51805
R1794 avdd.n3153 avdd.n3152 4.51805
R1795 avdd.n3082 avdd.n2986 4.51805
R1796 avdd.n3080 avdd.n3079 4.51805
R1797 avdd.n3312 avdd.n3311 4.51805
R1798 avdd.n3258 avdd.n3257 4.51805
R1799 avdd.n3366 avdd.n3365 4.51805
R1800 avdd.n3527 avdd.n3526 4.51805
R1801 avdd.n3473 avdd.n3472 4.51805
R1802 avdd.n3581 avdd.n3580 4.51805
R1803 avdd.n3742 avdd.n3741 4.51805
R1804 avdd.n3688 avdd.n3687 4.51805
R1805 avdd.n3796 avdd.n3795 4.51805
R1806 avdd.n3957 avdd.n3956 4.51805
R1807 avdd.n3903 avdd.n3902 4.51805
R1808 avdd.n4011 avdd.n4010 4.51805
R1809 avdd.n4172 avdd.n4171 4.51805
R1810 avdd.n4118 avdd.n4117 4.51805
R1811 avdd.n4226 avdd.n4225 4.51805
R1812 avdd.n4387 avdd.n4386 4.51805
R1813 avdd.n4333 avdd.n4332 4.51805
R1814 avdd.n4441 avdd.n4440 4.51805
R1815 avdd.n4942 avdd.n4941 4.51805
R1816 avdd.n4944 avdd.n4848 4.51805
R1817 avdd.n5010 avdd.n5009 4.51805
R1818 avdd.n5158 avdd.n5157 4.51805
R1819 avdd.n5160 avdd.n5064 4.51805
R1820 avdd.n5226 avdd.n5225 4.51805
R1821 avdd.n5374 avdd.n5373 4.51805
R1822 avdd.n5376 avdd.n5280 4.51805
R1823 avdd.n5442 avdd.n5441 4.51805
R1824 avdd.n5590 avdd.n5589 4.51805
R1825 avdd.n5592 avdd.n5496 4.51805
R1826 avdd.n5658 avdd.n5657 4.51805
R1827 avdd.n5806 avdd.n5805 4.51805
R1828 avdd.n5808 avdd.n5712 4.51805
R1829 avdd.n5874 avdd.n5873 4.51805
R1830 avdd.n6022 avdd.n6021 4.51805
R1831 avdd.n6024 avdd.n5928 4.51805
R1832 avdd.n6090 avdd.n6089 4.51805
R1833 avdd.n6238 avdd.n6237 4.51805
R1834 avdd.n6240 avdd.n6144 4.51805
R1835 avdd.n6306 avdd.n6305 4.51805
R1836 avdd.n6454 avdd.n6453 4.51805
R1837 avdd.n6456 avdd.n6360 4.51805
R1838 avdd.n6522 avdd.n6521 4.51805
R1839 avdd.n6670 avdd.n6669 4.51805
R1840 avdd.n6672 avdd.n6576 4.51805
R1841 avdd.n6738 avdd.n6737 4.51805
R1842 avdd.n6886 avdd.n6885 4.51805
R1843 avdd.n6888 avdd.n6792 4.51805
R1844 avdd.n6954 avdd.n6953 4.51805
R1845 avdd.n7102 avdd.n7101 4.51805
R1846 avdd.n7104 avdd.n7008 4.51805
R1847 avdd.n7170 avdd.n7169 4.51805
R1848 avdd.n7318 avdd.n7317 4.51805
R1849 avdd.n7320 avdd.n7224 4.51805
R1850 avdd.n7386 avdd.n7385 4.51805
R1851 avdd.n4642 avdd.n4641 4.5005
R1852 avdd.n4611 avdd.n4610 4.5005
R1853 avdd.n4609 avdd.n4608 4.5005
R1854 avdd.n4808 avdd.n4807 4.38235
R1855 avdd.n7622 avdd.n7621 4.36875
R1856 avdd.n7539 avdd.n7417 4.36875
R1857 avdd.n7522 avdd.n7521 4.36875
R1858 avdd.n7440 avdd.n7435 4.36875
R1859 avdd.n1688 avdd.n1687 4.36875
R1860 avdd.n1760 avdd.n1759 4.36875
R1861 avdd.n1778 avdd.n1777 4.36875
R1862 avdd.n1850 avdd.n1849 4.36875
R1863 avdd.n4601 avdd.n4600 4.22899
R1864 avdd.n4730 avdd.n4528 4.22899
R1865 avdd.n11266 avdd.n11265 4.22213
R1866 avdd.n4684 avdd.n4683 4.14168
R1867 avdd.n7630 avdd 3.97747
R1868 avdd.n4621 avdd.n4618 3.76521
R1869 avdd.n4632 avdd.n4631 3.76521
R1870 avdd.n4645 avdd.n4573 3.76521
R1871 avdd.n7402 avdd 3.62197
R1872 avdd.n7532 avdd.n7421 3.57983
R1873 avdd.n7574 avdd.n7406 3.57983
R1874 avdd.n7633 avdd.n7405 3.57983
R1875 avdd.n7474 avdd.n7423 3.57983
R1876 avdd.n1710 avdd.n1657 3.57983
R1877 avdd.n1770 avdd.n1649 3.57983
R1878 avdd.n1800 avdd.n1621 3.57983
R1879 avdd.n1867 avdd.n1620 3.57983
R1880 avdd.n4525 avdd.n4522 3.52991
R1881 avdd.n7622 avdd.n7579 3.50526
R1882 avdd.n7539 avdd.n7538 3.50526
R1883 avdd.n7522 avdd.n7479 3.50526
R1884 avdd.n7440 avdd.n7439 3.50526
R1885 avdd.n1687 avdd.n1686 3.50526
R1886 avdd.n1760 avdd.n1715 3.50526
R1887 avdd.n1777 avdd.n1776 3.50526
R1888 avdd.n1850 avdd.n1805 3.50526
R1889 avdd.n5020 avdd.n5019 3.41749
R1890 avdd.n5236 avdd.n5235 3.41749
R1891 avdd.n5452 avdd.n5451 3.41749
R1892 avdd.n5668 avdd.n5667 3.41749
R1893 avdd.n5884 avdd.n5883 3.41749
R1894 avdd.n6100 avdd.n6099 3.41749
R1895 avdd.n6316 avdd.n6315 3.41749
R1896 avdd.n6532 avdd.n6531 3.41749
R1897 avdd.n6748 avdd.n6747 3.41749
R1898 avdd.n6964 avdd.n6963 3.41749
R1899 avdd.n7180 avdd.n7179 3.41749
R1900 avdd.n7396 avdd.n7395 3.41749
R1901 avdd.n2021 avdd.n2004 3.41749
R1902 avdd.n2296 avdd.n2295 3.41749
R1903 avdd.n2511 avdd.n2510 3.41749
R1904 avdd.n2726 avdd.n2725 3.41749
R1905 avdd.n2941 avdd.n2940 3.41749
R1906 avdd.n3156 avdd.n3155 3.41749
R1907 avdd.n3315 avdd.n3294 3.41749
R1908 avdd.n3530 avdd.n3509 3.41749
R1909 avdd.n3745 avdd.n3724 3.41749
R1910 avdd.n3960 avdd.n3939 3.41749
R1911 avdd.n4175 avdd.n4154 3.41749
R1912 avdd.n4390 avdd.n4369 3.41749
R1913 avdd.n1910 avdd.n1909 3.41409
R1914 avdd.n2164 avdd.n2163 3.41409
R1915 avdd.n2379 avdd.n2378 3.41409
R1916 avdd.n2594 avdd.n2593 3.41409
R1917 avdd.n2809 avdd.n2808 3.41409
R1918 avdd.n3024 avdd.n3023 3.41409
R1919 avdd.n3200 avdd.n3199 3.41409
R1920 avdd.n3415 avdd.n3414 3.41409
R1921 avdd.n3630 avdd.n3629 3.41409
R1922 avdd.n3845 avdd.n3844 3.41409
R1923 avdd.n4060 avdd.n4059 3.41409
R1924 avdd.n4275 avdd.n4274 3.41409
R1925 avdd.n4886 avdd.n4885 3.41409
R1926 avdd.n5102 avdd.n5101 3.41409
R1927 avdd.n5318 avdd.n5317 3.41409
R1928 avdd.n5534 avdd.n5533 3.41409
R1929 avdd.n5750 avdd.n5749 3.41409
R1930 avdd.n5966 avdd.n5965 3.41409
R1931 avdd.n6182 avdd.n6181 3.41409
R1932 avdd.n6398 avdd.n6397 3.41409
R1933 avdd.n6614 avdd.n6613 3.41409
R1934 avdd.n6830 avdd.n6829 3.41409
R1935 avdd.n7046 avdd.n7045 3.41409
R1936 avdd.n7262 avdd.n7261 3.41409
R1937 avdd.n3379 avdd.n3170 3.41335
R1938 avdd.n3594 avdd.n3385 3.41335
R1939 avdd.n3809 avdd.n3600 3.41335
R1940 avdd.n4024 avdd.n3815 3.41335
R1941 avdd.n4239 avdd.n4030 3.41335
R1942 avdd.n4454 avdd.n4245 3.41335
R1943 avdd.n2036 avdd.n2009 3.4105
R1944 avdd.n2026 avdd.n2009 3.4105
R1945 avdd.n2011 avdd.n2010 3.4105
R1946 avdd.n2018 avdd.n2017 3.4105
R1947 avdd.n2015 avdd.n2014 3.4105
R1948 avdd.n2037 avdd.n2036 3.4105
R1949 avdd.n2037 avdd.n2001 3.4105
R1950 avdd.n2010 avdd.n2002 3.4105
R1951 avdd.n2033 avdd.n2031 3.4105
R1952 avdd.n2045 avdd.n2044 3.4105
R1953 avdd.n2044 avdd.n2043 3.4105
R1954 avdd.n1998 avdd.n1997 3.4105
R1955 avdd.n1992 avdd.n1991 3.4105
R1956 avdd.n2047 avdd.n2046 3.4105
R1957 avdd.n2048 avdd.n2047 3.4105
R1958 avdd.n1989 avdd.n1988 3.4105
R1959 avdd.n1984 avdd.n1972 3.4105
R1960 avdd.n1984 avdd.n1983 3.4105
R1961 avdd.n2054 avdd.n2053 3.4105
R1962 avdd.n2059 avdd.n2058 3.4105
R1963 avdd.n2066 avdd.n2065 3.4105
R1964 avdd.n2064 avdd.n2063 3.4105
R1965 avdd.n1967 avdd.n1958 3.4105
R1966 avdd.n1956 avdd.n1949 3.4105
R1967 avdd.n2070 avdd.n1950 3.4105
R1968 avdd.n1950 avdd.n1948 3.4105
R1969 avdd.n1953 avdd.n1952 3.4105
R1970 avdd.n2078 avdd.n1883 3.4105
R1971 avdd.n2078 avdd.n2077 3.4105
R1972 avdd.n2081 avdd.n2080 3.4105
R1973 avdd.n2088 avdd.n2087 3.4105
R1974 avdd.n2085 avdd.n2084 3.4105
R1975 avdd.n2084 avdd.n2083 3.4105
R1976 avdd.n1939 avdd.n1938 3.4105
R1977 avdd.n1927 avdd.n1896 3.4105
R1978 avdd.n1926 avdd.n1894 3.4105
R1979 avdd.n1894 avdd.n1893 3.4105
R1980 avdd.n1923 avdd.n1922 3.4105
R1981 avdd.n1905 avdd.n1904 3.4105
R1982 avdd.n1912 avdd.n1903 3.4105
R1983 avdd.n1912 avdd.n1911 3.4105
R1984 avdd.n1921 avdd.n1899 3.4105
R1985 avdd.n1921 avdd.n1892 3.4105
R1986 avdd.n1931 avdd.n1930 3.4105
R1987 avdd.n1937 avdd.n1891 3.4105
R1988 avdd.n1937 avdd.n1889 3.4105
R1989 avdd.n1943 avdd.n1880 3.4105
R1990 avdd.n1886 avdd.n1884 3.4105
R1991 avdd.n2079 avdd.n1887 3.4105
R1992 avdd.n1946 avdd.n1887 3.4105
R1993 avdd.n2074 avdd.n2073 3.4105
R1994 avdd.n1966 avdd.n1965 3.4105
R1995 avdd.n1966 avdd.n1947 3.4105
R1996 avdd.n1962 avdd.n1959 3.4105
R1997 avdd.n2061 avdd.n2060 3.4105
R1998 avdd.n2052 avdd.n1973 3.4105
R1999 avdd.n2052 avdd.n2051 3.4105
R2000 avdd.n1985 avdd.n1976 3.4105
R2001 avdd.n1980 avdd.n1978 3.4105
R2002 avdd.n1978 avdd.n1977 3.4105
R2003 avdd.n2042 avdd.n1996 3.4105
R2004 avdd.n2039 avdd.n2038 3.4105
R2005 avdd.n2016 avdd.n2012 3.4105
R2006 avdd.n2012 avdd.n2000 3.4105
R2007 avdd.n2028 avdd.n2027 3.4105
R2008 avdd.n2023 avdd.n2022 3.4105
R2009 avdd.n2030 avdd.n2002 3.4105
R2010 avdd.n2030 avdd.n2011 3.4105
R2011 avdd.n2030 avdd.n2029 3.4105
R2012 avdd.n2090 avdd.n1881 3.4105
R2013 avdd.n1941 avdd.n1878 3.4105
R2014 avdd.n1942 avdd.n1941 3.4105
R2015 avdd.n1936 avdd.n1935 3.4105
R2016 avdd.n1881 avdd.n1879 3.4105
R2017 avdd.n2091 avdd.n1879 3.4105
R2018 avdd.n2091 avdd.n2090 3.4105
R2019 avdd.n2301 avdd.n2093 3.4105
R2020 avdd.n2301 avdd.n2300 3.4105
R2021 avdd.n2302 avdd.n2094 3.4105
R2022 avdd.n2292 avdd.n2291 3.4105
R2023 avdd.n2288 avdd.n2287 3.4105
R2024 avdd.n2284 avdd.n2093 3.4105
R2025 avdd.n2285 avdd.n2284 3.4105
R2026 avdd.n2302 avdd.n2095 3.4105
R2027 avdd.n2275 avdd.n2106 3.4105
R2028 avdd.n2271 avdd.n2105 3.4105
R2029 avdd.n2105 avdd.n2104 3.4105
R2030 avdd.n2266 avdd.n2265 3.4105
R2031 avdd.n2253 avdd.n2252 3.4105
R2032 avdd.n2270 avdd.n2269 3.4105
R2033 avdd.n2269 avdd.n2268 3.4105
R2034 avdd.n2256 avdd.n2113 3.4105
R2035 avdd.n2251 avdd.n2112 3.4105
R2036 avdd.n2112 avdd.n2111 3.4105
R2037 avdd.n2248 avdd.n2247 3.4105
R2038 avdd.n2239 avdd.n2238 3.4105
R2039 avdd.n2232 avdd.n2120 3.4105
R2040 avdd.n2236 avdd.n2235 3.4105
R2041 avdd.n2127 avdd.n2126 3.4105
R2042 avdd.n2212 avdd.n2211 3.4105
R2043 avdd.n2228 avdd.n2227 3.4105
R2044 avdd.n2227 avdd.n2226 3.4105
R2045 avdd.n2215 avdd.n2214 3.4105
R2046 avdd.n2218 avdd.n2217 3.4105
R2047 avdd.n2219 avdd.n2218 3.4105
R2048 avdd.n2204 avdd.n2203 3.4105
R2049 avdd.n2142 avdd.n2141 3.4105
R2050 avdd.n2208 avdd.n2207 3.4105
R2051 avdd.n2207 avdd.n2206 3.4105
R2052 avdd.n2190 avdd.n2189 3.4105
R2053 avdd.n2150 avdd.n2143 3.4105
R2054 avdd.n2180 avdd.n2149 3.4105
R2055 avdd.n2149 avdd.n2148 3.4105
R2056 avdd.n2177 avdd.n2176 3.4105
R2057 avdd.n2159 avdd.n2158 3.4105
R2058 avdd.n2166 avdd.n2157 3.4105
R2059 avdd.n2166 avdd.n2165 3.4105
R2060 avdd.n2175 avdd.n2153 3.4105
R2061 avdd.n2175 avdd.n2147 3.4105
R2062 avdd.n2184 avdd.n2183 3.4105
R2063 avdd.n2191 avdd.n2146 3.4105
R2064 avdd.n2191 avdd.n2136 3.4105
R2065 avdd.n2199 avdd.n2198 3.4105
R2066 avdd.n2202 avdd.n2134 3.4105
R2067 avdd.n2131 avdd.n2130 3.4105
R2068 avdd.n2130 avdd.n2129 3.4105
R2069 avdd.n2210 avdd.n2125 3.4105
R2070 avdd.n2224 avdd.n2128 3.4105
R2071 avdd.n2224 avdd.n2223 3.4105
R2072 avdd.n2234 avdd.n2233 3.4105
R2073 avdd.n2241 avdd.n2240 3.4105
R2074 avdd.n2246 avdd.n2116 3.4105
R2075 avdd.n2246 avdd.n2110 3.4105
R2076 avdd.n2260 avdd.n2259 3.4105
R2077 avdd.n2267 avdd.n2109 3.4105
R2078 avdd.n2267 avdd.n2103 3.4105
R2079 avdd.n2279 avdd.n2278 3.4105
R2080 avdd.n2283 avdd.n2282 3.4105
R2081 avdd.n2289 avdd.n2101 3.4105
R2082 avdd.n2101 avdd.n2100 3.4105
R2083 avdd.n2099 avdd.n2097 3.4105
R2084 avdd.n2298 avdd.n2297 3.4105
R2085 avdd.n2305 avdd.n2095 3.4105
R2086 avdd.n2305 avdd.n2094 3.4105
R2087 avdd.n2305 avdd.n2304 3.4105
R2088 avdd.n2197 avdd.n2139 3.4105
R2089 avdd.n2195 avdd.n2138 3.4105
R2090 avdd.n2138 avdd.n2137 3.4105
R2091 avdd.n2193 avdd.n2192 3.4105
R2092 avdd.n2145 avdd.n2139 3.4105
R2093 avdd.n2145 avdd.n1877 3.4105
R2094 avdd.n2197 avdd.n1877 3.4105
R2095 avdd.n2516 avdd.n2308 3.4105
R2096 avdd.n2516 avdd.n2515 3.4105
R2097 avdd.n2517 avdd.n2309 3.4105
R2098 avdd.n2507 avdd.n2506 3.4105
R2099 avdd.n2503 avdd.n2502 3.4105
R2100 avdd.n2499 avdd.n2308 3.4105
R2101 avdd.n2500 avdd.n2499 3.4105
R2102 avdd.n2517 avdd.n2310 3.4105
R2103 avdd.n2490 avdd.n2321 3.4105
R2104 avdd.n2486 avdd.n2320 3.4105
R2105 avdd.n2320 avdd.n2319 3.4105
R2106 avdd.n2481 avdd.n2480 3.4105
R2107 avdd.n2468 avdd.n2467 3.4105
R2108 avdd.n2485 avdd.n2484 3.4105
R2109 avdd.n2484 avdd.n2483 3.4105
R2110 avdd.n2471 avdd.n2328 3.4105
R2111 avdd.n2466 avdd.n2327 3.4105
R2112 avdd.n2327 avdd.n2326 3.4105
R2113 avdd.n2463 avdd.n2462 3.4105
R2114 avdd.n2454 avdd.n2453 3.4105
R2115 avdd.n2447 avdd.n2335 3.4105
R2116 avdd.n2451 avdd.n2450 3.4105
R2117 avdd.n2342 avdd.n2341 3.4105
R2118 avdd.n2427 avdd.n2426 3.4105
R2119 avdd.n2443 avdd.n2442 3.4105
R2120 avdd.n2442 avdd.n2441 3.4105
R2121 avdd.n2430 avdd.n2429 3.4105
R2122 avdd.n2433 avdd.n2432 3.4105
R2123 avdd.n2434 avdd.n2433 3.4105
R2124 avdd.n2419 avdd.n2418 3.4105
R2125 avdd.n2357 avdd.n2356 3.4105
R2126 avdd.n2423 avdd.n2422 3.4105
R2127 avdd.n2422 avdd.n2421 3.4105
R2128 avdd.n2405 avdd.n2404 3.4105
R2129 avdd.n2365 avdd.n2358 3.4105
R2130 avdd.n2395 avdd.n2364 3.4105
R2131 avdd.n2364 avdd.n2363 3.4105
R2132 avdd.n2392 avdd.n2391 3.4105
R2133 avdd.n2374 avdd.n2373 3.4105
R2134 avdd.n2381 avdd.n2372 3.4105
R2135 avdd.n2381 avdd.n2380 3.4105
R2136 avdd.n2390 avdd.n2368 3.4105
R2137 avdd.n2390 avdd.n2362 3.4105
R2138 avdd.n2399 avdd.n2398 3.4105
R2139 avdd.n2406 avdd.n2361 3.4105
R2140 avdd.n2406 avdd.n2351 3.4105
R2141 avdd.n2414 avdd.n2413 3.4105
R2142 avdd.n2417 avdd.n2349 3.4105
R2143 avdd.n2346 avdd.n2345 3.4105
R2144 avdd.n2345 avdd.n2344 3.4105
R2145 avdd.n2425 avdd.n2340 3.4105
R2146 avdd.n2439 avdd.n2343 3.4105
R2147 avdd.n2439 avdd.n2438 3.4105
R2148 avdd.n2449 avdd.n2448 3.4105
R2149 avdd.n2456 avdd.n2455 3.4105
R2150 avdd.n2461 avdd.n2331 3.4105
R2151 avdd.n2461 avdd.n2325 3.4105
R2152 avdd.n2475 avdd.n2474 3.4105
R2153 avdd.n2482 avdd.n2324 3.4105
R2154 avdd.n2482 avdd.n2318 3.4105
R2155 avdd.n2494 avdd.n2493 3.4105
R2156 avdd.n2498 avdd.n2497 3.4105
R2157 avdd.n2504 avdd.n2316 3.4105
R2158 avdd.n2316 avdd.n2315 3.4105
R2159 avdd.n2314 avdd.n2312 3.4105
R2160 avdd.n2513 avdd.n2512 3.4105
R2161 avdd.n2520 avdd.n2310 3.4105
R2162 avdd.n2520 avdd.n2309 3.4105
R2163 avdd.n2520 avdd.n2519 3.4105
R2164 avdd.n2412 avdd.n2354 3.4105
R2165 avdd.n2410 avdd.n2353 3.4105
R2166 avdd.n2353 avdd.n2352 3.4105
R2167 avdd.n2408 avdd.n2407 3.4105
R2168 avdd.n2360 avdd.n2354 3.4105
R2169 avdd.n2360 avdd.n1876 3.4105
R2170 avdd.n2412 avdd.n1876 3.4105
R2171 avdd.n2731 avdd.n2523 3.4105
R2172 avdd.n2731 avdd.n2730 3.4105
R2173 avdd.n2732 avdd.n2524 3.4105
R2174 avdd.n2722 avdd.n2721 3.4105
R2175 avdd.n2718 avdd.n2717 3.4105
R2176 avdd.n2714 avdd.n2523 3.4105
R2177 avdd.n2715 avdd.n2714 3.4105
R2178 avdd.n2732 avdd.n2525 3.4105
R2179 avdd.n2705 avdd.n2536 3.4105
R2180 avdd.n2701 avdd.n2535 3.4105
R2181 avdd.n2535 avdd.n2534 3.4105
R2182 avdd.n2696 avdd.n2695 3.4105
R2183 avdd.n2683 avdd.n2682 3.4105
R2184 avdd.n2700 avdd.n2699 3.4105
R2185 avdd.n2699 avdd.n2698 3.4105
R2186 avdd.n2686 avdd.n2543 3.4105
R2187 avdd.n2681 avdd.n2542 3.4105
R2188 avdd.n2542 avdd.n2541 3.4105
R2189 avdd.n2678 avdd.n2677 3.4105
R2190 avdd.n2669 avdd.n2668 3.4105
R2191 avdd.n2662 avdd.n2550 3.4105
R2192 avdd.n2666 avdd.n2665 3.4105
R2193 avdd.n2557 avdd.n2556 3.4105
R2194 avdd.n2642 avdd.n2641 3.4105
R2195 avdd.n2658 avdd.n2657 3.4105
R2196 avdd.n2657 avdd.n2656 3.4105
R2197 avdd.n2645 avdd.n2644 3.4105
R2198 avdd.n2648 avdd.n2647 3.4105
R2199 avdd.n2649 avdd.n2648 3.4105
R2200 avdd.n2634 avdd.n2633 3.4105
R2201 avdd.n2572 avdd.n2571 3.4105
R2202 avdd.n2638 avdd.n2637 3.4105
R2203 avdd.n2637 avdd.n2636 3.4105
R2204 avdd.n2620 avdd.n2619 3.4105
R2205 avdd.n2580 avdd.n2573 3.4105
R2206 avdd.n2610 avdd.n2579 3.4105
R2207 avdd.n2579 avdd.n2578 3.4105
R2208 avdd.n2607 avdd.n2606 3.4105
R2209 avdd.n2589 avdd.n2588 3.4105
R2210 avdd.n2596 avdd.n2587 3.4105
R2211 avdd.n2596 avdd.n2595 3.4105
R2212 avdd.n2605 avdd.n2583 3.4105
R2213 avdd.n2605 avdd.n2577 3.4105
R2214 avdd.n2614 avdd.n2613 3.4105
R2215 avdd.n2621 avdd.n2576 3.4105
R2216 avdd.n2621 avdd.n2566 3.4105
R2217 avdd.n2629 avdd.n2628 3.4105
R2218 avdd.n2632 avdd.n2564 3.4105
R2219 avdd.n2561 avdd.n2560 3.4105
R2220 avdd.n2560 avdd.n2559 3.4105
R2221 avdd.n2640 avdd.n2555 3.4105
R2222 avdd.n2654 avdd.n2558 3.4105
R2223 avdd.n2654 avdd.n2653 3.4105
R2224 avdd.n2664 avdd.n2663 3.4105
R2225 avdd.n2671 avdd.n2670 3.4105
R2226 avdd.n2676 avdd.n2546 3.4105
R2227 avdd.n2676 avdd.n2540 3.4105
R2228 avdd.n2690 avdd.n2689 3.4105
R2229 avdd.n2697 avdd.n2539 3.4105
R2230 avdd.n2697 avdd.n2533 3.4105
R2231 avdd.n2709 avdd.n2708 3.4105
R2232 avdd.n2713 avdd.n2712 3.4105
R2233 avdd.n2719 avdd.n2531 3.4105
R2234 avdd.n2531 avdd.n2530 3.4105
R2235 avdd.n2529 avdd.n2527 3.4105
R2236 avdd.n2728 avdd.n2727 3.4105
R2237 avdd.n2735 avdd.n2525 3.4105
R2238 avdd.n2735 avdd.n2524 3.4105
R2239 avdd.n2735 avdd.n2734 3.4105
R2240 avdd.n2627 avdd.n2569 3.4105
R2241 avdd.n2625 avdd.n2568 3.4105
R2242 avdd.n2568 avdd.n2567 3.4105
R2243 avdd.n2623 avdd.n2622 3.4105
R2244 avdd.n2575 avdd.n2569 3.4105
R2245 avdd.n2575 avdd.n1875 3.4105
R2246 avdd.n2627 avdd.n1875 3.4105
R2247 avdd.n2946 avdd.n2738 3.4105
R2248 avdd.n2946 avdd.n2945 3.4105
R2249 avdd.n2947 avdd.n2739 3.4105
R2250 avdd.n2937 avdd.n2936 3.4105
R2251 avdd.n2933 avdd.n2932 3.4105
R2252 avdd.n2929 avdd.n2738 3.4105
R2253 avdd.n2930 avdd.n2929 3.4105
R2254 avdd.n2947 avdd.n2740 3.4105
R2255 avdd.n2920 avdd.n2751 3.4105
R2256 avdd.n2916 avdd.n2750 3.4105
R2257 avdd.n2750 avdd.n2749 3.4105
R2258 avdd.n2911 avdd.n2910 3.4105
R2259 avdd.n2898 avdd.n2897 3.4105
R2260 avdd.n2915 avdd.n2914 3.4105
R2261 avdd.n2914 avdd.n2913 3.4105
R2262 avdd.n2901 avdd.n2758 3.4105
R2263 avdd.n2896 avdd.n2757 3.4105
R2264 avdd.n2757 avdd.n2756 3.4105
R2265 avdd.n2893 avdd.n2892 3.4105
R2266 avdd.n2884 avdd.n2883 3.4105
R2267 avdd.n2877 avdd.n2765 3.4105
R2268 avdd.n2881 avdd.n2880 3.4105
R2269 avdd.n2772 avdd.n2771 3.4105
R2270 avdd.n2857 avdd.n2856 3.4105
R2271 avdd.n2873 avdd.n2872 3.4105
R2272 avdd.n2872 avdd.n2871 3.4105
R2273 avdd.n2860 avdd.n2859 3.4105
R2274 avdd.n2863 avdd.n2862 3.4105
R2275 avdd.n2864 avdd.n2863 3.4105
R2276 avdd.n2849 avdd.n2848 3.4105
R2277 avdd.n2787 avdd.n2786 3.4105
R2278 avdd.n2853 avdd.n2852 3.4105
R2279 avdd.n2852 avdd.n2851 3.4105
R2280 avdd.n2835 avdd.n2834 3.4105
R2281 avdd.n2795 avdd.n2788 3.4105
R2282 avdd.n2825 avdd.n2794 3.4105
R2283 avdd.n2794 avdd.n2793 3.4105
R2284 avdd.n2822 avdd.n2821 3.4105
R2285 avdd.n2804 avdd.n2803 3.4105
R2286 avdd.n2811 avdd.n2802 3.4105
R2287 avdd.n2811 avdd.n2810 3.4105
R2288 avdd.n2820 avdd.n2798 3.4105
R2289 avdd.n2820 avdd.n2792 3.4105
R2290 avdd.n2829 avdd.n2828 3.4105
R2291 avdd.n2836 avdd.n2791 3.4105
R2292 avdd.n2836 avdd.n2781 3.4105
R2293 avdd.n2844 avdd.n2843 3.4105
R2294 avdd.n2847 avdd.n2779 3.4105
R2295 avdd.n2776 avdd.n2775 3.4105
R2296 avdd.n2775 avdd.n2774 3.4105
R2297 avdd.n2855 avdd.n2770 3.4105
R2298 avdd.n2869 avdd.n2773 3.4105
R2299 avdd.n2869 avdd.n2868 3.4105
R2300 avdd.n2879 avdd.n2878 3.4105
R2301 avdd.n2886 avdd.n2885 3.4105
R2302 avdd.n2891 avdd.n2761 3.4105
R2303 avdd.n2891 avdd.n2755 3.4105
R2304 avdd.n2905 avdd.n2904 3.4105
R2305 avdd.n2912 avdd.n2754 3.4105
R2306 avdd.n2912 avdd.n2748 3.4105
R2307 avdd.n2924 avdd.n2923 3.4105
R2308 avdd.n2928 avdd.n2927 3.4105
R2309 avdd.n2934 avdd.n2746 3.4105
R2310 avdd.n2746 avdd.n2745 3.4105
R2311 avdd.n2744 avdd.n2742 3.4105
R2312 avdd.n2943 avdd.n2942 3.4105
R2313 avdd.n2950 avdd.n2740 3.4105
R2314 avdd.n2950 avdd.n2739 3.4105
R2315 avdd.n2950 avdd.n2949 3.4105
R2316 avdd.n2842 avdd.n2784 3.4105
R2317 avdd.n2840 avdd.n2783 3.4105
R2318 avdd.n2783 avdd.n2782 3.4105
R2319 avdd.n2838 avdd.n2837 3.4105
R2320 avdd.n2790 avdd.n2784 3.4105
R2321 avdd.n2790 avdd.n1874 3.4105
R2322 avdd.n2842 avdd.n1874 3.4105
R2323 avdd.n3161 avdd.n2953 3.4105
R2324 avdd.n3161 avdd.n3160 3.4105
R2325 avdd.n3162 avdd.n2954 3.4105
R2326 avdd.n3152 avdd.n3151 3.4105
R2327 avdd.n3148 avdd.n3147 3.4105
R2328 avdd.n3144 avdd.n2953 3.4105
R2329 avdd.n3145 avdd.n3144 3.4105
R2330 avdd.n3162 avdd.n2955 3.4105
R2331 avdd.n3135 avdd.n2966 3.4105
R2332 avdd.n3131 avdd.n2965 3.4105
R2333 avdd.n2965 avdd.n2964 3.4105
R2334 avdd.n3126 avdd.n3125 3.4105
R2335 avdd.n3113 avdd.n3112 3.4105
R2336 avdd.n3130 avdd.n3129 3.4105
R2337 avdd.n3129 avdd.n3128 3.4105
R2338 avdd.n3116 avdd.n2973 3.4105
R2339 avdd.n3111 avdd.n2972 3.4105
R2340 avdd.n2972 avdd.n2971 3.4105
R2341 avdd.n3108 avdd.n3107 3.4105
R2342 avdd.n3099 avdd.n3098 3.4105
R2343 avdd.n3092 avdd.n2980 3.4105
R2344 avdd.n3096 avdd.n3095 3.4105
R2345 avdd.n2987 avdd.n2986 3.4105
R2346 avdd.n3072 avdd.n3071 3.4105
R2347 avdd.n3088 avdd.n3087 3.4105
R2348 avdd.n3087 avdd.n3086 3.4105
R2349 avdd.n3075 avdd.n3074 3.4105
R2350 avdd.n3078 avdd.n3077 3.4105
R2351 avdd.n3079 avdd.n3078 3.4105
R2352 avdd.n3064 avdd.n3063 3.4105
R2353 avdd.n3002 avdd.n3001 3.4105
R2354 avdd.n3068 avdd.n3067 3.4105
R2355 avdd.n3067 avdd.n3066 3.4105
R2356 avdd.n3050 avdd.n3049 3.4105
R2357 avdd.n3010 avdd.n3003 3.4105
R2358 avdd.n3040 avdd.n3009 3.4105
R2359 avdd.n3009 avdd.n3008 3.4105
R2360 avdd.n3037 avdd.n3036 3.4105
R2361 avdd.n3019 avdd.n3018 3.4105
R2362 avdd.n3026 avdd.n3017 3.4105
R2363 avdd.n3026 avdd.n3025 3.4105
R2364 avdd.n3035 avdd.n3013 3.4105
R2365 avdd.n3035 avdd.n3007 3.4105
R2366 avdd.n3044 avdd.n3043 3.4105
R2367 avdd.n3051 avdd.n3006 3.4105
R2368 avdd.n3051 avdd.n2996 3.4105
R2369 avdd.n3059 avdd.n3058 3.4105
R2370 avdd.n3062 avdd.n2994 3.4105
R2371 avdd.n2991 avdd.n2990 3.4105
R2372 avdd.n2990 avdd.n2989 3.4105
R2373 avdd.n3070 avdd.n2985 3.4105
R2374 avdd.n3084 avdd.n2988 3.4105
R2375 avdd.n3084 avdd.n3083 3.4105
R2376 avdd.n3094 avdd.n3093 3.4105
R2377 avdd.n3101 avdd.n3100 3.4105
R2378 avdd.n3106 avdd.n2976 3.4105
R2379 avdd.n3106 avdd.n2970 3.4105
R2380 avdd.n3120 avdd.n3119 3.4105
R2381 avdd.n3127 avdd.n2969 3.4105
R2382 avdd.n3127 avdd.n2963 3.4105
R2383 avdd.n3139 avdd.n3138 3.4105
R2384 avdd.n3143 avdd.n3142 3.4105
R2385 avdd.n3149 avdd.n2961 3.4105
R2386 avdd.n2961 avdd.n2960 3.4105
R2387 avdd.n2959 avdd.n2957 3.4105
R2388 avdd.n3158 avdd.n3157 3.4105
R2389 avdd.n3165 avdd.n2955 3.4105
R2390 avdd.n3165 avdd.n2954 3.4105
R2391 avdd.n3165 avdd.n3164 3.4105
R2392 avdd.n3057 avdd.n2999 3.4105
R2393 avdd.n3055 avdd.n2998 3.4105
R2394 avdd.n2998 avdd.n2997 3.4105
R2395 avdd.n3053 avdd.n3052 3.4105
R2396 avdd.n3005 avdd.n2999 3.4105
R2397 avdd.n3005 avdd.n1873 3.4105
R2398 avdd.n3057 avdd.n1873 3.4105
R2399 avdd.n3308 avdd.n3307 3.4105
R2400 avdd.n3302 avdd.n3301 3.4105
R2401 avdd.n3334 avdd.n3333 3.4105
R2402 avdd.n3333 avdd.n3332 3.4105
R2403 avdd.n3288 avdd.n3287 3.4105
R2404 avdd.n3282 avdd.n3281 3.4105
R2405 avdd.n3336 avdd.n3335 3.4105
R2406 avdd.n3337 avdd.n3336 3.4105
R2407 avdd.n3279 avdd.n3278 3.4105
R2408 avdd.n3274 avdd.n3262 3.4105
R2409 avdd.n3274 avdd.n3273 3.4105
R2410 avdd.n3343 avdd.n3342 3.4105
R2411 avdd.n3348 avdd.n3347 3.4105
R2412 avdd.n3355 avdd.n3354 3.4105
R2413 avdd.n3353 avdd.n3352 3.4105
R2414 avdd.n3257 avdd.n3248 3.4105
R2415 avdd.n3246 avdd.n3239 3.4105
R2416 avdd.n3359 avdd.n3240 3.4105
R2417 avdd.n3240 avdd.n3238 3.4105
R2418 avdd.n3243 avdd.n3242 3.4105
R2419 avdd.n3367 avdd.n3173 3.4105
R2420 avdd.n3367 avdd.n3366 3.4105
R2421 avdd.n3370 avdd.n3369 3.4105
R2422 avdd.n3377 avdd.n3376 3.4105
R2423 avdd.n3374 avdd.n3373 3.4105
R2424 avdd.n3373 avdd.n3372 3.4105
R2425 avdd.n3231 avdd.n3169 3.4105
R2426 avdd.n3232 avdd.n3231 3.4105
R2427 avdd.n3229 avdd.n3228 3.4105
R2428 avdd.n3226 avdd.n3225 3.4105
R2429 avdd.n3217 avdd.n3186 3.4105
R2430 avdd.n3216 avdd.n3184 3.4105
R2431 avdd.n3184 avdd.n3183 3.4105
R2432 avdd.n3213 avdd.n3212 3.4105
R2433 avdd.n3195 avdd.n3194 3.4105
R2434 avdd.n3202 avdd.n3193 3.4105
R2435 avdd.n3202 avdd.n3201 3.4105
R2436 avdd.n3211 avdd.n3189 3.4105
R2437 avdd.n3211 avdd.n3182 3.4105
R2438 avdd.n3221 avdd.n3220 3.4105
R2439 avdd.n3227 avdd.n3181 3.4105
R2440 avdd.n3227 avdd.n3179 3.4105
R2441 avdd.n3233 avdd.n3171 3.4105
R2442 avdd.n3176 avdd.n3174 3.4105
R2443 avdd.n3368 avdd.n3177 3.4105
R2444 avdd.n3236 avdd.n3177 3.4105
R2445 avdd.n3363 avdd.n3362 3.4105
R2446 avdd.n3256 avdd.n3255 3.4105
R2447 avdd.n3256 avdd.n3237 3.4105
R2448 avdd.n3252 avdd.n3249 3.4105
R2449 avdd.n3350 avdd.n3349 3.4105
R2450 avdd.n3341 avdd.n3263 3.4105
R2451 avdd.n3341 avdd.n3340 3.4105
R2452 avdd.n3275 avdd.n3266 3.4105
R2453 avdd.n3270 avdd.n3268 3.4105
R2454 avdd.n3268 avdd.n3267 3.4105
R2455 avdd.n3331 avdd.n3286 3.4105
R2456 avdd.n3328 avdd.n3327 3.4105
R2457 avdd.n3310 avdd.n3309 3.4105
R2458 avdd.n3310 avdd.n3290 3.4105
R2459 avdd.n3322 avdd.n3321 3.4105
R2460 avdd.n3317 avdd.n3316 3.4105
R2461 avdd.n3381 avdd.n3170 3.4105
R2462 avdd.n3381 avdd.n3380 3.4105
R2463 avdd.n3320 avdd.n3319 3.4105
R2464 avdd.n3305 avdd.n3296 3.4105
R2465 avdd.n3323 avdd.n3296 3.4105
R2466 avdd.n3325 avdd.n3297 3.4105
R2467 avdd.n3311 avdd.n3297 3.4105
R2468 avdd.n3326 avdd.n3325 3.4105
R2469 avdd.n3326 avdd.n3291 3.4105
R2470 avdd.n3296 avdd.n3292 3.4105
R2471 avdd.n3299 avdd.n3292 3.4105
R2472 avdd.n3323 avdd.n3299 3.4105
R2473 avdd.n3305 avdd.n3299 3.4105
R2474 avdd.n3523 avdd.n3522 3.4105
R2475 avdd.n3517 avdd.n3516 3.4105
R2476 avdd.n3549 avdd.n3548 3.4105
R2477 avdd.n3548 avdd.n3547 3.4105
R2478 avdd.n3503 avdd.n3502 3.4105
R2479 avdd.n3497 avdd.n3496 3.4105
R2480 avdd.n3551 avdd.n3550 3.4105
R2481 avdd.n3552 avdd.n3551 3.4105
R2482 avdd.n3494 avdd.n3493 3.4105
R2483 avdd.n3489 avdd.n3477 3.4105
R2484 avdd.n3489 avdd.n3488 3.4105
R2485 avdd.n3558 avdd.n3557 3.4105
R2486 avdd.n3563 avdd.n3562 3.4105
R2487 avdd.n3570 avdd.n3569 3.4105
R2488 avdd.n3568 avdd.n3567 3.4105
R2489 avdd.n3472 avdd.n3463 3.4105
R2490 avdd.n3461 avdd.n3454 3.4105
R2491 avdd.n3574 avdd.n3455 3.4105
R2492 avdd.n3455 avdd.n3453 3.4105
R2493 avdd.n3458 avdd.n3457 3.4105
R2494 avdd.n3582 avdd.n3388 3.4105
R2495 avdd.n3582 avdd.n3581 3.4105
R2496 avdd.n3585 avdd.n3584 3.4105
R2497 avdd.n3592 avdd.n3591 3.4105
R2498 avdd.n3589 avdd.n3588 3.4105
R2499 avdd.n3588 avdd.n3587 3.4105
R2500 avdd.n3446 avdd.n3384 3.4105
R2501 avdd.n3447 avdd.n3446 3.4105
R2502 avdd.n3444 avdd.n3443 3.4105
R2503 avdd.n3441 avdd.n3440 3.4105
R2504 avdd.n3432 avdd.n3401 3.4105
R2505 avdd.n3431 avdd.n3399 3.4105
R2506 avdd.n3399 avdd.n3398 3.4105
R2507 avdd.n3428 avdd.n3427 3.4105
R2508 avdd.n3410 avdd.n3409 3.4105
R2509 avdd.n3417 avdd.n3408 3.4105
R2510 avdd.n3417 avdd.n3416 3.4105
R2511 avdd.n3426 avdd.n3404 3.4105
R2512 avdd.n3426 avdd.n3397 3.4105
R2513 avdd.n3436 avdd.n3435 3.4105
R2514 avdd.n3442 avdd.n3396 3.4105
R2515 avdd.n3442 avdd.n3394 3.4105
R2516 avdd.n3448 avdd.n3386 3.4105
R2517 avdd.n3391 avdd.n3389 3.4105
R2518 avdd.n3583 avdd.n3392 3.4105
R2519 avdd.n3451 avdd.n3392 3.4105
R2520 avdd.n3578 avdd.n3577 3.4105
R2521 avdd.n3471 avdd.n3470 3.4105
R2522 avdd.n3471 avdd.n3452 3.4105
R2523 avdd.n3467 avdd.n3464 3.4105
R2524 avdd.n3565 avdd.n3564 3.4105
R2525 avdd.n3556 avdd.n3478 3.4105
R2526 avdd.n3556 avdd.n3555 3.4105
R2527 avdd.n3490 avdd.n3481 3.4105
R2528 avdd.n3485 avdd.n3483 3.4105
R2529 avdd.n3483 avdd.n3482 3.4105
R2530 avdd.n3546 avdd.n3501 3.4105
R2531 avdd.n3543 avdd.n3542 3.4105
R2532 avdd.n3525 avdd.n3524 3.4105
R2533 avdd.n3525 avdd.n3505 3.4105
R2534 avdd.n3537 avdd.n3536 3.4105
R2535 avdd.n3532 avdd.n3531 3.4105
R2536 avdd.n3596 avdd.n3385 3.4105
R2537 avdd.n3596 avdd.n3595 3.4105
R2538 avdd.n3535 avdd.n3534 3.4105
R2539 avdd.n3520 avdd.n3511 3.4105
R2540 avdd.n3538 avdd.n3511 3.4105
R2541 avdd.n3540 avdd.n3512 3.4105
R2542 avdd.n3526 avdd.n3512 3.4105
R2543 avdd.n3541 avdd.n3540 3.4105
R2544 avdd.n3541 avdd.n3506 3.4105
R2545 avdd.n3511 avdd.n3507 3.4105
R2546 avdd.n3514 avdd.n3507 3.4105
R2547 avdd.n3538 avdd.n3514 3.4105
R2548 avdd.n3520 avdd.n3514 3.4105
R2549 avdd.n3738 avdd.n3737 3.4105
R2550 avdd.n3732 avdd.n3731 3.4105
R2551 avdd.n3764 avdd.n3763 3.4105
R2552 avdd.n3763 avdd.n3762 3.4105
R2553 avdd.n3718 avdd.n3717 3.4105
R2554 avdd.n3712 avdd.n3711 3.4105
R2555 avdd.n3766 avdd.n3765 3.4105
R2556 avdd.n3767 avdd.n3766 3.4105
R2557 avdd.n3709 avdd.n3708 3.4105
R2558 avdd.n3704 avdd.n3692 3.4105
R2559 avdd.n3704 avdd.n3703 3.4105
R2560 avdd.n3773 avdd.n3772 3.4105
R2561 avdd.n3778 avdd.n3777 3.4105
R2562 avdd.n3785 avdd.n3784 3.4105
R2563 avdd.n3783 avdd.n3782 3.4105
R2564 avdd.n3687 avdd.n3678 3.4105
R2565 avdd.n3676 avdd.n3669 3.4105
R2566 avdd.n3789 avdd.n3670 3.4105
R2567 avdd.n3670 avdd.n3668 3.4105
R2568 avdd.n3673 avdd.n3672 3.4105
R2569 avdd.n3797 avdd.n3603 3.4105
R2570 avdd.n3797 avdd.n3796 3.4105
R2571 avdd.n3800 avdd.n3799 3.4105
R2572 avdd.n3807 avdd.n3806 3.4105
R2573 avdd.n3804 avdd.n3803 3.4105
R2574 avdd.n3803 avdd.n3802 3.4105
R2575 avdd.n3661 avdd.n3599 3.4105
R2576 avdd.n3662 avdd.n3661 3.4105
R2577 avdd.n3659 avdd.n3658 3.4105
R2578 avdd.n3656 avdd.n3655 3.4105
R2579 avdd.n3647 avdd.n3616 3.4105
R2580 avdd.n3646 avdd.n3614 3.4105
R2581 avdd.n3614 avdd.n3613 3.4105
R2582 avdd.n3643 avdd.n3642 3.4105
R2583 avdd.n3625 avdd.n3624 3.4105
R2584 avdd.n3632 avdd.n3623 3.4105
R2585 avdd.n3632 avdd.n3631 3.4105
R2586 avdd.n3641 avdd.n3619 3.4105
R2587 avdd.n3641 avdd.n3612 3.4105
R2588 avdd.n3651 avdd.n3650 3.4105
R2589 avdd.n3657 avdd.n3611 3.4105
R2590 avdd.n3657 avdd.n3609 3.4105
R2591 avdd.n3663 avdd.n3601 3.4105
R2592 avdd.n3606 avdd.n3604 3.4105
R2593 avdd.n3798 avdd.n3607 3.4105
R2594 avdd.n3666 avdd.n3607 3.4105
R2595 avdd.n3793 avdd.n3792 3.4105
R2596 avdd.n3686 avdd.n3685 3.4105
R2597 avdd.n3686 avdd.n3667 3.4105
R2598 avdd.n3682 avdd.n3679 3.4105
R2599 avdd.n3780 avdd.n3779 3.4105
R2600 avdd.n3771 avdd.n3693 3.4105
R2601 avdd.n3771 avdd.n3770 3.4105
R2602 avdd.n3705 avdd.n3696 3.4105
R2603 avdd.n3700 avdd.n3698 3.4105
R2604 avdd.n3698 avdd.n3697 3.4105
R2605 avdd.n3761 avdd.n3716 3.4105
R2606 avdd.n3758 avdd.n3757 3.4105
R2607 avdd.n3740 avdd.n3739 3.4105
R2608 avdd.n3740 avdd.n3720 3.4105
R2609 avdd.n3752 avdd.n3751 3.4105
R2610 avdd.n3747 avdd.n3746 3.4105
R2611 avdd.n3811 avdd.n3600 3.4105
R2612 avdd.n3811 avdd.n3810 3.4105
R2613 avdd.n3750 avdd.n3749 3.4105
R2614 avdd.n3735 avdd.n3726 3.4105
R2615 avdd.n3753 avdd.n3726 3.4105
R2616 avdd.n3755 avdd.n3727 3.4105
R2617 avdd.n3741 avdd.n3727 3.4105
R2618 avdd.n3756 avdd.n3755 3.4105
R2619 avdd.n3756 avdd.n3721 3.4105
R2620 avdd.n3726 avdd.n3722 3.4105
R2621 avdd.n3729 avdd.n3722 3.4105
R2622 avdd.n3753 avdd.n3729 3.4105
R2623 avdd.n3735 avdd.n3729 3.4105
R2624 avdd.n3953 avdd.n3952 3.4105
R2625 avdd.n3947 avdd.n3946 3.4105
R2626 avdd.n3979 avdd.n3978 3.4105
R2627 avdd.n3978 avdd.n3977 3.4105
R2628 avdd.n3933 avdd.n3932 3.4105
R2629 avdd.n3927 avdd.n3926 3.4105
R2630 avdd.n3981 avdd.n3980 3.4105
R2631 avdd.n3982 avdd.n3981 3.4105
R2632 avdd.n3924 avdd.n3923 3.4105
R2633 avdd.n3919 avdd.n3907 3.4105
R2634 avdd.n3919 avdd.n3918 3.4105
R2635 avdd.n3988 avdd.n3987 3.4105
R2636 avdd.n3993 avdd.n3992 3.4105
R2637 avdd.n4000 avdd.n3999 3.4105
R2638 avdd.n3998 avdd.n3997 3.4105
R2639 avdd.n3902 avdd.n3893 3.4105
R2640 avdd.n3891 avdd.n3884 3.4105
R2641 avdd.n4004 avdd.n3885 3.4105
R2642 avdd.n3885 avdd.n3883 3.4105
R2643 avdd.n3888 avdd.n3887 3.4105
R2644 avdd.n4012 avdd.n3818 3.4105
R2645 avdd.n4012 avdd.n4011 3.4105
R2646 avdd.n4015 avdd.n4014 3.4105
R2647 avdd.n4022 avdd.n4021 3.4105
R2648 avdd.n4019 avdd.n4018 3.4105
R2649 avdd.n4018 avdd.n4017 3.4105
R2650 avdd.n3876 avdd.n3814 3.4105
R2651 avdd.n3877 avdd.n3876 3.4105
R2652 avdd.n3874 avdd.n3873 3.4105
R2653 avdd.n3871 avdd.n3870 3.4105
R2654 avdd.n3862 avdd.n3831 3.4105
R2655 avdd.n3861 avdd.n3829 3.4105
R2656 avdd.n3829 avdd.n3828 3.4105
R2657 avdd.n3858 avdd.n3857 3.4105
R2658 avdd.n3840 avdd.n3839 3.4105
R2659 avdd.n3847 avdd.n3838 3.4105
R2660 avdd.n3847 avdd.n3846 3.4105
R2661 avdd.n3856 avdd.n3834 3.4105
R2662 avdd.n3856 avdd.n3827 3.4105
R2663 avdd.n3866 avdd.n3865 3.4105
R2664 avdd.n3872 avdd.n3826 3.4105
R2665 avdd.n3872 avdd.n3824 3.4105
R2666 avdd.n3878 avdd.n3816 3.4105
R2667 avdd.n3821 avdd.n3819 3.4105
R2668 avdd.n4013 avdd.n3822 3.4105
R2669 avdd.n3881 avdd.n3822 3.4105
R2670 avdd.n4008 avdd.n4007 3.4105
R2671 avdd.n3901 avdd.n3900 3.4105
R2672 avdd.n3901 avdd.n3882 3.4105
R2673 avdd.n3897 avdd.n3894 3.4105
R2674 avdd.n3995 avdd.n3994 3.4105
R2675 avdd.n3986 avdd.n3908 3.4105
R2676 avdd.n3986 avdd.n3985 3.4105
R2677 avdd.n3920 avdd.n3911 3.4105
R2678 avdd.n3915 avdd.n3913 3.4105
R2679 avdd.n3913 avdd.n3912 3.4105
R2680 avdd.n3976 avdd.n3931 3.4105
R2681 avdd.n3973 avdd.n3972 3.4105
R2682 avdd.n3955 avdd.n3954 3.4105
R2683 avdd.n3955 avdd.n3935 3.4105
R2684 avdd.n3967 avdd.n3966 3.4105
R2685 avdd.n3962 avdd.n3961 3.4105
R2686 avdd.n4026 avdd.n3815 3.4105
R2687 avdd.n4026 avdd.n4025 3.4105
R2688 avdd.n3965 avdd.n3964 3.4105
R2689 avdd.n3950 avdd.n3941 3.4105
R2690 avdd.n3968 avdd.n3941 3.4105
R2691 avdd.n3970 avdd.n3942 3.4105
R2692 avdd.n3956 avdd.n3942 3.4105
R2693 avdd.n3971 avdd.n3970 3.4105
R2694 avdd.n3971 avdd.n3936 3.4105
R2695 avdd.n3941 avdd.n3937 3.4105
R2696 avdd.n3944 avdd.n3937 3.4105
R2697 avdd.n3968 avdd.n3944 3.4105
R2698 avdd.n3950 avdd.n3944 3.4105
R2699 avdd.n4168 avdd.n4167 3.4105
R2700 avdd.n4162 avdd.n4161 3.4105
R2701 avdd.n4194 avdd.n4193 3.4105
R2702 avdd.n4193 avdd.n4192 3.4105
R2703 avdd.n4148 avdd.n4147 3.4105
R2704 avdd.n4142 avdd.n4141 3.4105
R2705 avdd.n4196 avdd.n4195 3.4105
R2706 avdd.n4197 avdd.n4196 3.4105
R2707 avdd.n4139 avdd.n4138 3.4105
R2708 avdd.n4134 avdd.n4122 3.4105
R2709 avdd.n4134 avdd.n4133 3.4105
R2710 avdd.n4203 avdd.n4202 3.4105
R2711 avdd.n4208 avdd.n4207 3.4105
R2712 avdd.n4215 avdd.n4214 3.4105
R2713 avdd.n4213 avdd.n4212 3.4105
R2714 avdd.n4117 avdd.n4108 3.4105
R2715 avdd.n4106 avdd.n4099 3.4105
R2716 avdd.n4219 avdd.n4100 3.4105
R2717 avdd.n4100 avdd.n4098 3.4105
R2718 avdd.n4103 avdd.n4102 3.4105
R2719 avdd.n4227 avdd.n4033 3.4105
R2720 avdd.n4227 avdd.n4226 3.4105
R2721 avdd.n4230 avdd.n4229 3.4105
R2722 avdd.n4237 avdd.n4236 3.4105
R2723 avdd.n4234 avdd.n4233 3.4105
R2724 avdd.n4233 avdd.n4232 3.4105
R2725 avdd.n4091 avdd.n4029 3.4105
R2726 avdd.n4092 avdd.n4091 3.4105
R2727 avdd.n4089 avdd.n4088 3.4105
R2728 avdd.n4086 avdd.n4085 3.4105
R2729 avdd.n4077 avdd.n4046 3.4105
R2730 avdd.n4076 avdd.n4044 3.4105
R2731 avdd.n4044 avdd.n4043 3.4105
R2732 avdd.n4073 avdd.n4072 3.4105
R2733 avdd.n4055 avdd.n4054 3.4105
R2734 avdd.n4062 avdd.n4053 3.4105
R2735 avdd.n4062 avdd.n4061 3.4105
R2736 avdd.n4071 avdd.n4049 3.4105
R2737 avdd.n4071 avdd.n4042 3.4105
R2738 avdd.n4081 avdd.n4080 3.4105
R2739 avdd.n4087 avdd.n4041 3.4105
R2740 avdd.n4087 avdd.n4039 3.4105
R2741 avdd.n4093 avdd.n4031 3.4105
R2742 avdd.n4036 avdd.n4034 3.4105
R2743 avdd.n4228 avdd.n4037 3.4105
R2744 avdd.n4096 avdd.n4037 3.4105
R2745 avdd.n4223 avdd.n4222 3.4105
R2746 avdd.n4116 avdd.n4115 3.4105
R2747 avdd.n4116 avdd.n4097 3.4105
R2748 avdd.n4112 avdd.n4109 3.4105
R2749 avdd.n4210 avdd.n4209 3.4105
R2750 avdd.n4201 avdd.n4123 3.4105
R2751 avdd.n4201 avdd.n4200 3.4105
R2752 avdd.n4135 avdd.n4126 3.4105
R2753 avdd.n4130 avdd.n4128 3.4105
R2754 avdd.n4128 avdd.n4127 3.4105
R2755 avdd.n4191 avdd.n4146 3.4105
R2756 avdd.n4188 avdd.n4187 3.4105
R2757 avdd.n4170 avdd.n4169 3.4105
R2758 avdd.n4170 avdd.n4150 3.4105
R2759 avdd.n4182 avdd.n4181 3.4105
R2760 avdd.n4177 avdd.n4176 3.4105
R2761 avdd.n4241 avdd.n4030 3.4105
R2762 avdd.n4241 avdd.n4240 3.4105
R2763 avdd.n4180 avdd.n4179 3.4105
R2764 avdd.n4165 avdd.n4156 3.4105
R2765 avdd.n4183 avdd.n4156 3.4105
R2766 avdd.n4185 avdd.n4157 3.4105
R2767 avdd.n4171 avdd.n4157 3.4105
R2768 avdd.n4186 avdd.n4185 3.4105
R2769 avdd.n4186 avdd.n4151 3.4105
R2770 avdd.n4156 avdd.n4152 3.4105
R2771 avdd.n4159 avdd.n4152 3.4105
R2772 avdd.n4183 avdd.n4159 3.4105
R2773 avdd.n4165 avdd.n4159 3.4105
R2774 avdd.n4383 avdd.n4382 3.4105
R2775 avdd.n4377 avdd.n4376 3.4105
R2776 avdd.n4409 avdd.n4408 3.4105
R2777 avdd.n4408 avdd.n4407 3.4105
R2778 avdd.n4363 avdd.n4362 3.4105
R2779 avdd.n4357 avdd.n4356 3.4105
R2780 avdd.n4411 avdd.n4410 3.4105
R2781 avdd.n4412 avdd.n4411 3.4105
R2782 avdd.n4354 avdd.n4353 3.4105
R2783 avdd.n4349 avdd.n4337 3.4105
R2784 avdd.n4349 avdd.n4348 3.4105
R2785 avdd.n4418 avdd.n4417 3.4105
R2786 avdd.n4423 avdd.n4422 3.4105
R2787 avdd.n4430 avdd.n4429 3.4105
R2788 avdd.n4428 avdd.n4427 3.4105
R2789 avdd.n4332 avdd.n4323 3.4105
R2790 avdd.n4321 avdd.n4314 3.4105
R2791 avdd.n4434 avdd.n4315 3.4105
R2792 avdd.n4315 avdd.n4313 3.4105
R2793 avdd.n4318 avdd.n4317 3.4105
R2794 avdd.n4442 avdd.n4248 3.4105
R2795 avdd.n4442 avdd.n4441 3.4105
R2796 avdd.n4445 avdd.n4444 3.4105
R2797 avdd.n4452 avdd.n4451 3.4105
R2798 avdd.n4449 avdd.n4448 3.4105
R2799 avdd.n4448 avdd.n4447 3.4105
R2800 avdd.n4306 avdd.n4244 3.4105
R2801 avdd.n4307 avdd.n4306 3.4105
R2802 avdd.n4304 avdd.n4303 3.4105
R2803 avdd.n4301 avdd.n4300 3.4105
R2804 avdd.n4292 avdd.n4261 3.4105
R2805 avdd.n4291 avdd.n4259 3.4105
R2806 avdd.n4259 avdd.n4258 3.4105
R2807 avdd.n4288 avdd.n4287 3.4105
R2808 avdd.n4270 avdd.n4269 3.4105
R2809 avdd.n4277 avdd.n4268 3.4105
R2810 avdd.n4277 avdd.n4276 3.4105
R2811 avdd.n4286 avdd.n4264 3.4105
R2812 avdd.n4286 avdd.n4257 3.4105
R2813 avdd.n4296 avdd.n4295 3.4105
R2814 avdd.n4302 avdd.n4256 3.4105
R2815 avdd.n4302 avdd.n4254 3.4105
R2816 avdd.n4308 avdd.n4246 3.4105
R2817 avdd.n4251 avdd.n4249 3.4105
R2818 avdd.n4443 avdd.n4252 3.4105
R2819 avdd.n4311 avdd.n4252 3.4105
R2820 avdd.n4438 avdd.n4437 3.4105
R2821 avdd.n4331 avdd.n4330 3.4105
R2822 avdd.n4331 avdd.n4312 3.4105
R2823 avdd.n4327 avdd.n4324 3.4105
R2824 avdd.n4425 avdd.n4424 3.4105
R2825 avdd.n4416 avdd.n4338 3.4105
R2826 avdd.n4416 avdd.n4415 3.4105
R2827 avdd.n4350 avdd.n4341 3.4105
R2828 avdd.n4345 avdd.n4343 3.4105
R2829 avdd.n4343 avdd.n4342 3.4105
R2830 avdd.n4406 avdd.n4361 3.4105
R2831 avdd.n4403 avdd.n4402 3.4105
R2832 avdd.n4385 avdd.n4384 3.4105
R2833 avdd.n4385 avdd.n4365 3.4105
R2834 avdd.n4397 avdd.n4396 3.4105
R2835 avdd.n4392 avdd.n4391 3.4105
R2836 avdd.n4456 avdd.n4245 3.4105
R2837 avdd.n4456 avdd.n4455 3.4105
R2838 avdd.n4395 avdd.n4394 3.4105
R2839 avdd.n4380 avdd.n4371 3.4105
R2840 avdd.n4398 avdd.n4371 3.4105
R2841 avdd.n4400 avdd.n4372 3.4105
R2842 avdd.n4386 avdd.n4372 3.4105
R2843 avdd.n4401 avdd.n4400 3.4105
R2844 avdd.n4401 avdd.n4366 3.4105
R2845 avdd.n4371 avdd.n4367 3.4105
R2846 avdd.n4374 avdd.n4367 3.4105
R2847 avdd.n4398 avdd.n4374 3.4105
R2848 avdd.n4380 avdd.n4374 3.4105
R2849 avdd.n4819 avdd.n4812 3.4105
R2850 avdd.n4819 avdd.n4810 3.4105
R2851 avdd.n4819 avdd.n4811 3.4105
R2852 avdd.n5023 avdd.n4811 3.4105
R2853 avdd.n5015 avdd.n5014 3.4105
R2854 avdd.n5013 avdd.n5012 3.4105
R2855 avdd.n5018 avdd.n4820 3.4105
R2856 avdd.n4881 avdd.n4880 3.4105
R2857 avdd.n4888 avdd.n4879 3.4105
R2858 avdd.n4888 avdd.n4887 3.4105
R2859 avdd.n4897 avdd.n4875 3.4105
R2860 avdd.n4897 avdd.n4869 3.4105
R2861 avdd.n4903 avdd.n4872 3.4105
R2862 avdd.n4899 avdd.n4898 3.4105
R2863 avdd.n4902 avdd.n4871 3.4105
R2864 avdd.n4871 avdd.n4870 3.4105
R2865 avdd.n4907 avdd.n4906 3.4105
R2866 avdd.n4914 avdd.n4868 3.4105
R2867 avdd.n4914 avdd.n4858 3.4105
R2868 avdd.n4913 avdd.n4912 3.4105
R2869 avdd.n4921 avdd.n4920 3.4105
R2870 avdd.n4924 avdd.n4856 3.4105
R2871 avdd.n4937 avdd.n4936 3.4105
R2872 avdd.n4865 avdd.n4864 3.4105
R2873 avdd.n4930 avdd.n4929 3.4105
R2874 avdd.n4929 avdd.n4928 3.4105
R2875 avdd.n4926 avdd.n4925 3.4105
R2876 avdd.n4940 avdd.n4939 3.4105
R2877 avdd.n4941 avdd.n4940 3.4105
R2878 avdd.n4853 avdd.n4852 3.4105
R2879 avdd.n4852 avdd.n4851 3.4105
R2880 avdd.n4932 avdd.n4847 3.4105
R2881 avdd.n4934 avdd.n4933 3.4105
R2882 avdd.n4950 avdd.n4949 3.4105
R2883 avdd.n4949 avdd.n4948 3.4105
R2884 avdd.n4849 avdd.n4848 3.4105
R2885 avdd.n4946 avdd.n4850 3.4105
R2886 avdd.n4946 avdd.n4945 3.4105
R2887 avdd.n4956 avdd.n4955 3.4105
R2888 avdd.n4961 avdd.n4960 3.4105
R2889 avdd.n4954 avdd.n4842 3.4105
R2890 avdd.n4958 avdd.n4957 3.4105
R2891 avdd.n4963 avdd.n4962 3.4105
R2892 avdd.n4968 avdd.n4838 3.4105
R2893 avdd.n4968 avdd.n4832 3.4105
R2894 avdd.n4978 avdd.n4835 3.4105
R2895 avdd.n4970 avdd.n4969 3.4105
R2896 avdd.n4973 avdd.n4834 3.4105
R2897 avdd.n4834 avdd.n4833 3.4105
R2898 avdd.n4982 avdd.n4981 3.4105
R2899 avdd.n4989 avdd.n4831 3.4105
R2900 avdd.n4989 avdd.n4824 3.4105
R2901 avdd.n4994 avdd.n4828 3.4105
R2902 avdd.n4975 avdd.n4974 3.4105
R2903 avdd.n4992 avdd.n4991 3.4105
R2904 avdd.n4991 avdd.n4990 3.4105
R2905 avdd.n4988 avdd.n4987 3.4105
R2906 avdd.n4993 avdd.n4826 3.4105
R2907 avdd.n4826 avdd.n4825 3.4105
R2908 avdd.n4998 avdd.n4997 3.4105
R2909 avdd.n5002 avdd.n5001 3.4105
R2910 avdd.n5023 avdd.n4810 3.4105
R2911 avdd.n5021 avdd.n4816 3.4105
R2912 avdd.n5021 avdd.n4815 3.4105
R2913 avdd.n5003 avdd.n4815 3.4105
R2914 avdd.n5006 avdd.n5005 3.4105
R2915 avdd.n5009 avdd.n5008 3.4105
R2916 avdd.n5007 avdd.n4822 3.4105
R2917 avdd.n4822 avdd.n4821 3.4105
R2918 avdd.n4919 avdd.n4918 3.4105
R2919 avdd.n4918 avdd.n4917 3.4105
R2920 avdd.n4916 avdd.n4866 3.4105
R2921 avdd.n4916 avdd.n4915 3.4105
R2922 avdd.n4866 avdd.n4860 3.4105
R2923 avdd.n4860 avdd.n4859 3.4105
R2924 avdd.n5035 avdd.n5028 3.4105
R2925 avdd.n5035 avdd.n5026 3.4105
R2926 avdd.n5035 avdd.n5027 3.4105
R2927 avdd.n5239 avdd.n5027 3.4105
R2928 avdd.n5231 avdd.n5230 3.4105
R2929 avdd.n5229 avdd.n5228 3.4105
R2930 avdd.n5234 avdd.n5036 3.4105
R2931 avdd.n5097 avdd.n5096 3.4105
R2932 avdd.n5104 avdd.n5095 3.4105
R2933 avdd.n5104 avdd.n5103 3.4105
R2934 avdd.n5113 avdd.n5091 3.4105
R2935 avdd.n5113 avdd.n5085 3.4105
R2936 avdd.n5119 avdd.n5088 3.4105
R2937 avdd.n5115 avdd.n5114 3.4105
R2938 avdd.n5118 avdd.n5087 3.4105
R2939 avdd.n5087 avdd.n5086 3.4105
R2940 avdd.n5123 avdd.n5122 3.4105
R2941 avdd.n5130 avdd.n5084 3.4105
R2942 avdd.n5130 avdd.n5074 3.4105
R2943 avdd.n5129 avdd.n5128 3.4105
R2944 avdd.n5137 avdd.n5136 3.4105
R2945 avdd.n5140 avdd.n5072 3.4105
R2946 avdd.n5153 avdd.n5152 3.4105
R2947 avdd.n5081 avdd.n5080 3.4105
R2948 avdd.n5146 avdd.n5145 3.4105
R2949 avdd.n5145 avdd.n5144 3.4105
R2950 avdd.n5142 avdd.n5141 3.4105
R2951 avdd.n5156 avdd.n5155 3.4105
R2952 avdd.n5157 avdd.n5156 3.4105
R2953 avdd.n5069 avdd.n5068 3.4105
R2954 avdd.n5068 avdd.n5067 3.4105
R2955 avdd.n5148 avdd.n5063 3.4105
R2956 avdd.n5150 avdd.n5149 3.4105
R2957 avdd.n5166 avdd.n5165 3.4105
R2958 avdd.n5165 avdd.n5164 3.4105
R2959 avdd.n5065 avdd.n5064 3.4105
R2960 avdd.n5162 avdd.n5066 3.4105
R2961 avdd.n5162 avdd.n5161 3.4105
R2962 avdd.n5172 avdd.n5171 3.4105
R2963 avdd.n5177 avdd.n5176 3.4105
R2964 avdd.n5170 avdd.n5058 3.4105
R2965 avdd.n5174 avdd.n5173 3.4105
R2966 avdd.n5179 avdd.n5178 3.4105
R2967 avdd.n5184 avdd.n5054 3.4105
R2968 avdd.n5184 avdd.n5048 3.4105
R2969 avdd.n5194 avdd.n5051 3.4105
R2970 avdd.n5186 avdd.n5185 3.4105
R2971 avdd.n5189 avdd.n5050 3.4105
R2972 avdd.n5050 avdd.n5049 3.4105
R2973 avdd.n5198 avdd.n5197 3.4105
R2974 avdd.n5205 avdd.n5047 3.4105
R2975 avdd.n5205 avdd.n5040 3.4105
R2976 avdd.n5210 avdd.n5044 3.4105
R2977 avdd.n5191 avdd.n5190 3.4105
R2978 avdd.n5208 avdd.n5207 3.4105
R2979 avdd.n5207 avdd.n5206 3.4105
R2980 avdd.n5204 avdd.n5203 3.4105
R2981 avdd.n5209 avdd.n5042 3.4105
R2982 avdd.n5042 avdd.n5041 3.4105
R2983 avdd.n5214 avdd.n5213 3.4105
R2984 avdd.n5218 avdd.n5217 3.4105
R2985 avdd.n5239 avdd.n5026 3.4105
R2986 avdd.n5237 avdd.n5032 3.4105
R2987 avdd.n5237 avdd.n5031 3.4105
R2988 avdd.n5219 avdd.n5031 3.4105
R2989 avdd.n5222 avdd.n5221 3.4105
R2990 avdd.n5225 avdd.n5224 3.4105
R2991 avdd.n5223 avdd.n5038 3.4105
R2992 avdd.n5038 avdd.n5037 3.4105
R2993 avdd.n5135 avdd.n5134 3.4105
R2994 avdd.n5134 avdd.n5133 3.4105
R2995 avdd.n5132 avdd.n5082 3.4105
R2996 avdd.n5132 avdd.n5131 3.4105
R2997 avdd.n5082 avdd.n5076 3.4105
R2998 avdd.n5076 avdd.n5075 3.4105
R2999 avdd.n5251 avdd.n5244 3.4105
R3000 avdd.n5251 avdd.n5242 3.4105
R3001 avdd.n5251 avdd.n5243 3.4105
R3002 avdd.n5455 avdd.n5243 3.4105
R3003 avdd.n5447 avdd.n5446 3.4105
R3004 avdd.n5445 avdd.n5444 3.4105
R3005 avdd.n5450 avdd.n5252 3.4105
R3006 avdd.n5313 avdd.n5312 3.4105
R3007 avdd.n5320 avdd.n5311 3.4105
R3008 avdd.n5320 avdd.n5319 3.4105
R3009 avdd.n5329 avdd.n5307 3.4105
R3010 avdd.n5329 avdd.n5301 3.4105
R3011 avdd.n5335 avdd.n5304 3.4105
R3012 avdd.n5331 avdd.n5330 3.4105
R3013 avdd.n5334 avdd.n5303 3.4105
R3014 avdd.n5303 avdd.n5302 3.4105
R3015 avdd.n5339 avdd.n5338 3.4105
R3016 avdd.n5346 avdd.n5300 3.4105
R3017 avdd.n5346 avdd.n5290 3.4105
R3018 avdd.n5345 avdd.n5344 3.4105
R3019 avdd.n5353 avdd.n5352 3.4105
R3020 avdd.n5356 avdd.n5288 3.4105
R3021 avdd.n5369 avdd.n5368 3.4105
R3022 avdd.n5297 avdd.n5296 3.4105
R3023 avdd.n5362 avdd.n5361 3.4105
R3024 avdd.n5361 avdd.n5360 3.4105
R3025 avdd.n5358 avdd.n5357 3.4105
R3026 avdd.n5372 avdd.n5371 3.4105
R3027 avdd.n5373 avdd.n5372 3.4105
R3028 avdd.n5285 avdd.n5284 3.4105
R3029 avdd.n5284 avdd.n5283 3.4105
R3030 avdd.n5364 avdd.n5279 3.4105
R3031 avdd.n5366 avdd.n5365 3.4105
R3032 avdd.n5382 avdd.n5381 3.4105
R3033 avdd.n5381 avdd.n5380 3.4105
R3034 avdd.n5281 avdd.n5280 3.4105
R3035 avdd.n5378 avdd.n5282 3.4105
R3036 avdd.n5378 avdd.n5377 3.4105
R3037 avdd.n5388 avdd.n5387 3.4105
R3038 avdd.n5393 avdd.n5392 3.4105
R3039 avdd.n5386 avdd.n5274 3.4105
R3040 avdd.n5390 avdd.n5389 3.4105
R3041 avdd.n5395 avdd.n5394 3.4105
R3042 avdd.n5400 avdd.n5270 3.4105
R3043 avdd.n5400 avdd.n5264 3.4105
R3044 avdd.n5410 avdd.n5267 3.4105
R3045 avdd.n5402 avdd.n5401 3.4105
R3046 avdd.n5405 avdd.n5266 3.4105
R3047 avdd.n5266 avdd.n5265 3.4105
R3048 avdd.n5414 avdd.n5413 3.4105
R3049 avdd.n5421 avdd.n5263 3.4105
R3050 avdd.n5421 avdd.n5256 3.4105
R3051 avdd.n5426 avdd.n5260 3.4105
R3052 avdd.n5407 avdd.n5406 3.4105
R3053 avdd.n5424 avdd.n5423 3.4105
R3054 avdd.n5423 avdd.n5422 3.4105
R3055 avdd.n5420 avdd.n5419 3.4105
R3056 avdd.n5425 avdd.n5258 3.4105
R3057 avdd.n5258 avdd.n5257 3.4105
R3058 avdd.n5430 avdd.n5429 3.4105
R3059 avdd.n5434 avdd.n5433 3.4105
R3060 avdd.n5455 avdd.n5242 3.4105
R3061 avdd.n5453 avdd.n5248 3.4105
R3062 avdd.n5453 avdd.n5247 3.4105
R3063 avdd.n5435 avdd.n5247 3.4105
R3064 avdd.n5438 avdd.n5437 3.4105
R3065 avdd.n5441 avdd.n5440 3.4105
R3066 avdd.n5439 avdd.n5254 3.4105
R3067 avdd.n5254 avdd.n5253 3.4105
R3068 avdd.n5351 avdd.n5350 3.4105
R3069 avdd.n5350 avdd.n5349 3.4105
R3070 avdd.n5348 avdd.n5298 3.4105
R3071 avdd.n5348 avdd.n5347 3.4105
R3072 avdd.n5298 avdd.n5292 3.4105
R3073 avdd.n5292 avdd.n5291 3.4105
R3074 avdd.n5467 avdd.n5460 3.4105
R3075 avdd.n5467 avdd.n5458 3.4105
R3076 avdd.n5467 avdd.n5459 3.4105
R3077 avdd.n5671 avdd.n5459 3.4105
R3078 avdd.n5663 avdd.n5662 3.4105
R3079 avdd.n5661 avdd.n5660 3.4105
R3080 avdd.n5666 avdd.n5468 3.4105
R3081 avdd.n5529 avdd.n5528 3.4105
R3082 avdd.n5536 avdd.n5527 3.4105
R3083 avdd.n5536 avdd.n5535 3.4105
R3084 avdd.n5545 avdd.n5523 3.4105
R3085 avdd.n5545 avdd.n5517 3.4105
R3086 avdd.n5551 avdd.n5520 3.4105
R3087 avdd.n5547 avdd.n5546 3.4105
R3088 avdd.n5550 avdd.n5519 3.4105
R3089 avdd.n5519 avdd.n5518 3.4105
R3090 avdd.n5555 avdd.n5554 3.4105
R3091 avdd.n5562 avdd.n5516 3.4105
R3092 avdd.n5562 avdd.n5506 3.4105
R3093 avdd.n5561 avdd.n5560 3.4105
R3094 avdd.n5569 avdd.n5568 3.4105
R3095 avdd.n5572 avdd.n5504 3.4105
R3096 avdd.n5585 avdd.n5584 3.4105
R3097 avdd.n5513 avdd.n5512 3.4105
R3098 avdd.n5578 avdd.n5577 3.4105
R3099 avdd.n5577 avdd.n5576 3.4105
R3100 avdd.n5574 avdd.n5573 3.4105
R3101 avdd.n5588 avdd.n5587 3.4105
R3102 avdd.n5589 avdd.n5588 3.4105
R3103 avdd.n5501 avdd.n5500 3.4105
R3104 avdd.n5500 avdd.n5499 3.4105
R3105 avdd.n5580 avdd.n5495 3.4105
R3106 avdd.n5582 avdd.n5581 3.4105
R3107 avdd.n5598 avdd.n5597 3.4105
R3108 avdd.n5597 avdd.n5596 3.4105
R3109 avdd.n5497 avdd.n5496 3.4105
R3110 avdd.n5594 avdd.n5498 3.4105
R3111 avdd.n5594 avdd.n5593 3.4105
R3112 avdd.n5604 avdd.n5603 3.4105
R3113 avdd.n5609 avdd.n5608 3.4105
R3114 avdd.n5602 avdd.n5490 3.4105
R3115 avdd.n5606 avdd.n5605 3.4105
R3116 avdd.n5611 avdd.n5610 3.4105
R3117 avdd.n5616 avdd.n5486 3.4105
R3118 avdd.n5616 avdd.n5480 3.4105
R3119 avdd.n5626 avdd.n5483 3.4105
R3120 avdd.n5618 avdd.n5617 3.4105
R3121 avdd.n5621 avdd.n5482 3.4105
R3122 avdd.n5482 avdd.n5481 3.4105
R3123 avdd.n5630 avdd.n5629 3.4105
R3124 avdd.n5637 avdd.n5479 3.4105
R3125 avdd.n5637 avdd.n5472 3.4105
R3126 avdd.n5642 avdd.n5476 3.4105
R3127 avdd.n5623 avdd.n5622 3.4105
R3128 avdd.n5640 avdd.n5639 3.4105
R3129 avdd.n5639 avdd.n5638 3.4105
R3130 avdd.n5636 avdd.n5635 3.4105
R3131 avdd.n5641 avdd.n5474 3.4105
R3132 avdd.n5474 avdd.n5473 3.4105
R3133 avdd.n5646 avdd.n5645 3.4105
R3134 avdd.n5650 avdd.n5649 3.4105
R3135 avdd.n5671 avdd.n5458 3.4105
R3136 avdd.n5669 avdd.n5464 3.4105
R3137 avdd.n5669 avdd.n5463 3.4105
R3138 avdd.n5651 avdd.n5463 3.4105
R3139 avdd.n5654 avdd.n5653 3.4105
R3140 avdd.n5657 avdd.n5656 3.4105
R3141 avdd.n5655 avdd.n5470 3.4105
R3142 avdd.n5470 avdd.n5469 3.4105
R3143 avdd.n5567 avdd.n5566 3.4105
R3144 avdd.n5566 avdd.n5565 3.4105
R3145 avdd.n5564 avdd.n5514 3.4105
R3146 avdd.n5564 avdd.n5563 3.4105
R3147 avdd.n5514 avdd.n5508 3.4105
R3148 avdd.n5508 avdd.n5507 3.4105
R3149 avdd.n5683 avdd.n5676 3.4105
R3150 avdd.n5683 avdd.n5674 3.4105
R3151 avdd.n5683 avdd.n5675 3.4105
R3152 avdd.n5887 avdd.n5675 3.4105
R3153 avdd.n5879 avdd.n5878 3.4105
R3154 avdd.n5877 avdd.n5876 3.4105
R3155 avdd.n5882 avdd.n5684 3.4105
R3156 avdd.n5745 avdd.n5744 3.4105
R3157 avdd.n5752 avdd.n5743 3.4105
R3158 avdd.n5752 avdd.n5751 3.4105
R3159 avdd.n5761 avdd.n5739 3.4105
R3160 avdd.n5761 avdd.n5733 3.4105
R3161 avdd.n5767 avdd.n5736 3.4105
R3162 avdd.n5763 avdd.n5762 3.4105
R3163 avdd.n5766 avdd.n5735 3.4105
R3164 avdd.n5735 avdd.n5734 3.4105
R3165 avdd.n5771 avdd.n5770 3.4105
R3166 avdd.n5778 avdd.n5732 3.4105
R3167 avdd.n5778 avdd.n5722 3.4105
R3168 avdd.n5777 avdd.n5776 3.4105
R3169 avdd.n5785 avdd.n5784 3.4105
R3170 avdd.n5788 avdd.n5720 3.4105
R3171 avdd.n5801 avdd.n5800 3.4105
R3172 avdd.n5729 avdd.n5728 3.4105
R3173 avdd.n5794 avdd.n5793 3.4105
R3174 avdd.n5793 avdd.n5792 3.4105
R3175 avdd.n5790 avdd.n5789 3.4105
R3176 avdd.n5804 avdd.n5803 3.4105
R3177 avdd.n5805 avdd.n5804 3.4105
R3178 avdd.n5717 avdd.n5716 3.4105
R3179 avdd.n5716 avdd.n5715 3.4105
R3180 avdd.n5796 avdd.n5711 3.4105
R3181 avdd.n5798 avdd.n5797 3.4105
R3182 avdd.n5814 avdd.n5813 3.4105
R3183 avdd.n5813 avdd.n5812 3.4105
R3184 avdd.n5713 avdd.n5712 3.4105
R3185 avdd.n5810 avdd.n5714 3.4105
R3186 avdd.n5810 avdd.n5809 3.4105
R3187 avdd.n5820 avdd.n5819 3.4105
R3188 avdd.n5825 avdd.n5824 3.4105
R3189 avdd.n5818 avdd.n5706 3.4105
R3190 avdd.n5822 avdd.n5821 3.4105
R3191 avdd.n5827 avdd.n5826 3.4105
R3192 avdd.n5832 avdd.n5702 3.4105
R3193 avdd.n5832 avdd.n5696 3.4105
R3194 avdd.n5842 avdd.n5699 3.4105
R3195 avdd.n5834 avdd.n5833 3.4105
R3196 avdd.n5837 avdd.n5698 3.4105
R3197 avdd.n5698 avdd.n5697 3.4105
R3198 avdd.n5846 avdd.n5845 3.4105
R3199 avdd.n5853 avdd.n5695 3.4105
R3200 avdd.n5853 avdd.n5688 3.4105
R3201 avdd.n5858 avdd.n5692 3.4105
R3202 avdd.n5839 avdd.n5838 3.4105
R3203 avdd.n5856 avdd.n5855 3.4105
R3204 avdd.n5855 avdd.n5854 3.4105
R3205 avdd.n5852 avdd.n5851 3.4105
R3206 avdd.n5857 avdd.n5690 3.4105
R3207 avdd.n5690 avdd.n5689 3.4105
R3208 avdd.n5862 avdd.n5861 3.4105
R3209 avdd.n5866 avdd.n5865 3.4105
R3210 avdd.n5887 avdd.n5674 3.4105
R3211 avdd.n5885 avdd.n5680 3.4105
R3212 avdd.n5885 avdd.n5679 3.4105
R3213 avdd.n5867 avdd.n5679 3.4105
R3214 avdd.n5870 avdd.n5869 3.4105
R3215 avdd.n5873 avdd.n5872 3.4105
R3216 avdd.n5871 avdd.n5686 3.4105
R3217 avdd.n5686 avdd.n5685 3.4105
R3218 avdd.n5783 avdd.n5782 3.4105
R3219 avdd.n5782 avdd.n5781 3.4105
R3220 avdd.n5780 avdd.n5730 3.4105
R3221 avdd.n5780 avdd.n5779 3.4105
R3222 avdd.n5730 avdd.n5724 3.4105
R3223 avdd.n5724 avdd.n5723 3.4105
R3224 avdd.n5899 avdd.n5892 3.4105
R3225 avdd.n5899 avdd.n5890 3.4105
R3226 avdd.n5899 avdd.n5891 3.4105
R3227 avdd.n6103 avdd.n5891 3.4105
R3228 avdd.n6095 avdd.n6094 3.4105
R3229 avdd.n6093 avdd.n6092 3.4105
R3230 avdd.n6098 avdd.n5900 3.4105
R3231 avdd.n5961 avdd.n5960 3.4105
R3232 avdd.n5968 avdd.n5959 3.4105
R3233 avdd.n5968 avdd.n5967 3.4105
R3234 avdd.n5977 avdd.n5955 3.4105
R3235 avdd.n5977 avdd.n5949 3.4105
R3236 avdd.n5983 avdd.n5952 3.4105
R3237 avdd.n5979 avdd.n5978 3.4105
R3238 avdd.n5982 avdd.n5951 3.4105
R3239 avdd.n5951 avdd.n5950 3.4105
R3240 avdd.n5987 avdd.n5986 3.4105
R3241 avdd.n5994 avdd.n5948 3.4105
R3242 avdd.n5994 avdd.n5938 3.4105
R3243 avdd.n5993 avdd.n5992 3.4105
R3244 avdd.n6001 avdd.n6000 3.4105
R3245 avdd.n6004 avdd.n5936 3.4105
R3246 avdd.n6017 avdd.n6016 3.4105
R3247 avdd.n5945 avdd.n5944 3.4105
R3248 avdd.n6010 avdd.n6009 3.4105
R3249 avdd.n6009 avdd.n6008 3.4105
R3250 avdd.n6006 avdd.n6005 3.4105
R3251 avdd.n6020 avdd.n6019 3.4105
R3252 avdd.n6021 avdd.n6020 3.4105
R3253 avdd.n5933 avdd.n5932 3.4105
R3254 avdd.n5932 avdd.n5931 3.4105
R3255 avdd.n6012 avdd.n5927 3.4105
R3256 avdd.n6014 avdd.n6013 3.4105
R3257 avdd.n6030 avdd.n6029 3.4105
R3258 avdd.n6029 avdd.n6028 3.4105
R3259 avdd.n5929 avdd.n5928 3.4105
R3260 avdd.n6026 avdd.n5930 3.4105
R3261 avdd.n6026 avdd.n6025 3.4105
R3262 avdd.n6036 avdd.n6035 3.4105
R3263 avdd.n6041 avdd.n6040 3.4105
R3264 avdd.n6034 avdd.n5922 3.4105
R3265 avdd.n6038 avdd.n6037 3.4105
R3266 avdd.n6043 avdd.n6042 3.4105
R3267 avdd.n6048 avdd.n5918 3.4105
R3268 avdd.n6048 avdd.n5912 3.4105
R3269 avdd.n6058 avdd.n5915 3.4105
R3270 avdd.n6050 avdd.n6049 3.4105
R3271 avdd.n6053 avdd.n5914 3.4105
R3272 avdd.n5914 avdd.n5913 3.4105
R3273 avdd.n6062 avdd.n6061 3.4105
R3274 avdd.n6069 avdd.n5911 3.4105
R3275 avdd.n6069 avdd.n5904 3.4105
R3276 avdd.n6074 avdd.n5908 3.4105
R3277 avdd.n6055 avdd.n6054 3.4105
R3278 avdd.n6072 avdd.n6071 3.4105
R3279 avdd.n6071 avdd.n6070 3.4105
R3280 avdd.n6068 avdd.n6067 3.4105
R3281 avdd.n6073 avdd.n5906 3.4105
R3282 avdd.n5906 avdd.n5905 3.4105
R3283 avdd.n6078 avdd.n6077 3.4105
R3284 avdd.n6082 avdd.n6081 3.4105
R3285 avdd.n6103 avdd.n5890 3.4105
R3286 avdd.n6101 avdd.n5896 3.4105
R3287 avdd.n6101 avdd.n5895 3.4105
R3288 avdd.n6083 avdd.n5895 3.4105
R3289 avdd.n6086 avdd.n6085 3.4105
R3290 avdd.n6089 avdd.n6088 3.4105
R3291 avdd.n6087 avdd.n5902 3.4105
R3292 avdd.n5902 avdd.n5901 3.4105
R3293 avdd.n5999 avdd.n5998 3.4105
R3294 avdd.n5998 avdd.n5997 3.4105
R3295 avdd.n5996 avdd.n5946 3.4105
R3296 avdd.n5996 avdd.n5995 3.4105
R3297 avdd.n5946 avdd.n5940 3.4105
R3298 avdd.n5940 avdd.n5939 3.4105
R3299 avdd.n6115 avdd.n6108 3.4105
R3300 avdd.n6115 avdd.n6106 3.4105
R3301 avdd.n6115 avdd.n6107 3.4105
R3302 avdd.n6319 avdd.n6107 3.4105
R3303 avdd.n6311 avdd.n6310 3.4105
R3304 avdd.n6309 avdd.n6308 3.4105
R3305 avdd.n6314 avdd.n6116 3.4105
R3306 avdd.n6177 avdd.n6176 3.4105
R3307 avdd.n6184 avdd.n6175 3.4105
R3308 avdd.n6184 avdd.n6183 3.4105
R3309 avdd.n6193 avdd.n6171 3.4105
R3310 avdd.n6193 avdd.n6165 3.4105
R3311 avdd.n6199 avdd.n6168 3.4105
R3312 avdd.n6195 avdd.n6194 3.4105
R3313 avdd.n6198 avdd.n6167 3.4105
R3314 avdd.n6167 avdd.n6166 3.4105
R3315 avdd.n6203 avdd.n6202 3.4105
R3316 avdd.n6210 avdd.n6164 3.4105
R3317 avdd.n6210 avdd.n6154 3.4105
R3318 avdd.n6209 avdd.n6208 3.4105
R3319 avdd.n6217 avdd.n6216 3.4105
R3320 avdd.n6220 avdd.n6152 3.4105
R3321 avdd.n6233 avdd.n6232 3.4105
R3322 avdd.n6161 avdd.n6160 3.4105
R3323 avdd.n6226 avdd.n6225 3.4105
R3324 avdd.n6225 avdd.n6224 3.4105
R3325 avdd.n6222 avdd.n6221 3.4105
R3326 avdd.n6236 avdd.n6235 3.4105
R3327 avdd.n6237 avdd.n6236 3.4105
R3328 avdd.n6149 avdd.n6148 3.4105
R3329 avdd.n6148 avdd.n6147 3.4105
R3330 avdd.n6228 avdd.n6143 3.4105
R3331 avdd.n6230 avdd.n6229 3.4105
R3332 avdd.n6246 avdd.n6245 3.4105
R3333 avdd.n6245 avdd.n6244 3.4105
R3334 avdd.n6145 avdd.n6144 3.4105
R3335 avdd.n6242 avdd.n6146 3.4105
R3336 avdd.n6242 avdd.n6241 3.4105
R3337 avdd.n6252 avdd.n6251 3.4105
R3338 avdd.n6257 avdd.n6256 3.4105
R3339 avdd.n6250 avdd.n6138 3.4105
R3340 avdd.n6254 avdd.n6253 3.4105
R3341 avdd.n6259 avdd.n6258 3.4105
R3342 avdd.n6264 avdd.n6134 3.4105
R3343 avdd.n6264 avdd.n6128 3.4105
R3344 avdd.n6274 avdd.n6131 3.4105
R3345 avdd.n6266 avdd.n6265 3.4105
R3346 avdd.n6269 avdd.n6130 3.4105
R3347 avdd.n6130 avdd.n6129 3.4105
R3348 avdd.n6278 avdd.n6277 3.4105
R3349 avdd.n6285 avdd.n6127 3.4105
R3350 avdd.n6285 avdd.n6120 3.4105
R3351 avdd.n6290 avdd.n6124 3.4105
R3352 avdd.n6271 avdd.n6270 3.4105
R3353 avdd.n6288 avdd.n6287 3.4105
R3354 avdd.n6287 avdd.n6286 3.4105
R3355 avdd.n6284 avdd.n6283 3.4105
R3356 avdd.n6289 avdd.n6122 3.4105
R3357 avdd.n6122 avdd.n6121 3.4105
R3358 avdd.n6294 avdd.n6293 3.4105
R3359 avdd.n6298 avdd.n6297 3.4105
R3360 avdd.n6319 avdd.n6106 3.4105
R3361 avdd.n6317 avdd.n6112 3.4105
R3362 avdd.n6317 avdd.n6111 3.4105
R3363 avdd.n6299 avdd.n6111 3.4105
R3364 avdd.n6302 avdd.n6301 3.4105
R3365 avdd.n6305 avdd.n6304 3.4105
R3366 avdd.n6303 avdd.n6118 3.4105
R3367 avdd.n6118 avdd.n6117 3.4105
R3368 avdd.n6215 avdd.n6214 3.4105
R3369 avdd.n6214 avdd.n6213 3.4105
R3370 avdd.n6212 avdd.n6162 3.4105
R3371 avdd.n6212 avdd.n6211 3.4105
R3372 avdd.n6162 avdd.n6156 3.4105
R3373 avdd.n6156 avdd.n6155 3.4105
R3374 avdd.n6331 avdd.n6324 3.4105
R3375 avdd.n6331 avdd.n6322 3.4105
R3376 avdd.n6331 avdd.n6323 3.4105
R3377 avdd.n6535 avdd.n6323 3.4105
R3378 avdd.n6527 avdd.n6526 3.4105
R3379 avdd.n6525 avdd.n6524 3.4105
R3380 avdd.n6530 avdd.n6332 3.4105
R3381 avdd.n6393 avdd.n6392 3.4105
R3382 avdd.n6400 avdd.n6391 3.4105
R3383 avdd.n6400 avdd.n6399 3.4105
R3384 avdd.n6409 avdd.n6387 3.4105
R3385 avdd.n6409 avdd.n6381 3.4105
R3386 avdd.n6415 avdd.n6384 3.4105
R3387 avdd.n6411 avdd.n6410 3.4105
R3388 avdd.n6414 avdd.n6383 3.4105
R3389 avdd.n6383 avdd.n6382 3.4105
R3390 avdd.n6419 avdd.n6418 3.4105
R3391 avdd.n6426 avdd.n6380 3.4105
R3392 avdd.n6426 avdd.n6370 3.4105
R3393 avdd.n6425 avdd.n6424 3.4105
R3394 avdd.n6433 avdd.n6432 3.4105
R3395 avdd.n6436 avdd.n6368 3.4105
R3396 avdd.n6449 avdd.n6448 3.4105
R3397 avdd.n6377 avdd.n6376 3.4105
R3398 avdd.n6442 avdd.n6441 3.4105
R3399 avdd.n6441 avdd.n6440 3.4105
R3400 avdd.n6438 avdd.n6437 3.4105
R3401 avdd.n6452 avdd.n6451 3.4105
R3402 avdd.n6453 avdd.n6452 3.4105
R3403 avdd.n6365 avdd.n6364 3.4105
R3404 avdd.n6364 avdd.n6363 3.4105
R3405 avdd.n6444 avdd.n6359 3.4105
R3406 avdd.n6446 avdd.n6445 3.4105
R3407 avdd.n6462 avdd.n6461 3.4105
R3408 avdd.n6461 avdd.n6460 3.4105
R3409 avdd.n6361 avdd.n6360 3.4105
R3410 avdd.n6458 avdd.n6362 3.4105
R3411 avdd.n6458 avdd.n6457 3.4105
R3412 avdd.n6468 avdd.n6467 3.4105
R3413 avdd.n6473 avdd.n6472 3.4105
R3414 avdd.n6466 avdd.n6354 3.4105
R3415 avdd.n6470 avdd.n6469 3.4105
R3416 avdd.n6475 avdd.n6474 3.4105
R3417 avdd.n6480 avdd.n6350 3.4105
R3418 avdd.n6480 avdd.n6344 3.4105
R3419 avdd.n6490 avdd.n6347 3.4105
R3420 avdd.n6482 avdd.n6481 3.4105
R3421 avdd.n6485 avdd.n6346 3.4105
R3422 avdd.n6346 avdd.n6345 3.4105
R3423 avdd.n6494 avdd.n6493 3.4105
R3424 avdd.n6501 avdd.n6343 3.4105
R3425 avdd.n6501 avdd.n6336 3.4105
R3426 avdd.n6506 avdd.n6340 3.4105
R3427 avdd.n6487 avdd.n6486 3.4105
R3428 avdd.n6504 avdd.n6503 3.4105
R3429 avdd.n6503 avdd.n6502 3.4105
R3430 avdd.n6500 avdd.n6499 3.4105
R3431 avdd.n6505 avdd.n6338 3.4105
R3432 avdd.n6338 avdd.n6337 3.4105
R3433 avdd.n6510 avdd.n6509 3.4105
R3434 avdd.n6514 avdd.n6513 3.4105
R3435 avdd.n6535 avdd.n6322 3.4105
R3436 avdd.n6533 avdd.n6328 3.4105
R3437 avdd.n6533 avdd.n6327 3.4105
R3438 avdd.n6515 avdd.n6327 3.4105
R3439 avdd.n6518 avdd.n6517 3.4105
R3440 avdd.n6521 avdd.n6520 3.4105
R3441 avdd.n6519 avdd.n6334 3.4105
R3442 avdd.n6334 avdd.n6333 3.4105
R3443 avdd.n6431 avdd.n6430 3.4105
R3444 avdd.n6430 avdd.n6429 3.4105
R3445 avdd.n6428 avdd.n6378 3.4105
R3446 avdd.n6428 avdd.n6427 3.4105
R3447 avdd.n6378 avdd.n6372 3.4105
R3448 avdd.n6372 avdd.n6371 3.4105
R3449 avdd.n6547 avdd.n6540 3.4105
R3450 avdd.n6547 avdd.n6538 3.4105
R3451 avdd.n6547 avdd.n6539 3.4105
R3452 avdd.n6751 avdd.n6539 3.4105
R3453 avdd.n6743 avdd.n6742 3.4105
R3454 avdd.n6741 avdd.n6740 3.4105
R3455 avdd.n6746 avdd.n6548 3.4105
R3456 avdd.n6609 avdd.n6608 3.4105
R3457 avdd.n6616 avdd.n6607 3.4105
R3458 avdd.n6616 avdd.n6615 3.4105
R3459 avdd.n6625 avdd.n6603 3.4105
R3460 avdd.n6625 avdd.n6597 3.4105
R3461 avdd.n6631 avdd.n6600 3.4105
R3462 avdd.n6627 avdd.n6626 3.4105
R3463 avdd.n6630 avdd.n6599 3.4105
R3464 avdd.n6599 avdd.n6598 3.4105
R3465 avdd.n6635 avdd.n6634 3.4105
R3466 avdd.n6642 avdd.n6596 3.4105
R3467 avdd.n6642 avdd.n6586 3.4105
R3468 avdd.n6641 avdd.n6640 3.4105
R3469 avdd.n6649 avdd.n6648 3.4105
R3470 avdd.n6652 avdd.n6584 3.4105
R3471 avdd.n6665 avdd.n6664 3.4105
R3472 avdd.n6593 avdd.n6592 3.4105
R3473 avdd.n6658 avdd.n6657 3.4105
R3474 avdd.n6657 avdd.n6656 3.4105
R3475 avdd.n6654 avdd.n6653 3.4105
R3476 avdd.n6668 avdd.n6667 3.4105
R3477 avdd.n6669 avdd.n6668 3.4105
R3478 avdd.n6581 avdd.n6580 3.4105
R3479 avdd.n6580 avdd.n6579 3.4105
R3480 avdd.n6660 avdd.n6575 3.4105
R3481 avdd.n6662 avdd.n6661 3.4105
R3482 avdd.n6678 avdd.n6677 3.4105
R3483 avdd.n6677 avdd.n6676 3.4105
R3484 avdd.n6577 avdd.n6576 3.4105
R3485 avdd.n6674 avdd.n6578 3.4105
R3486 avdd.n6674 avdd.n6673 3.4105
R3487 avdd.n6684 avdd.n6683 3.4105
R3488 avdd.n6689 avdd.n6688 3.4105
R3489 avdd.n6682 avdd.n6570 3.4105
R3490 avdd.n6686 avdd.n6685 3.4105
R3491 avdd.n6691 avdd.n6690 3.4105
R3492 avdd.n6696 avdd.n6566 3.4105
R3493 avdd.n6696 avdd.n6560 3.4105
R3494 avdd.n6706 avdd.n6563 3.4105
R3495 avdd.n6698 avdd.n6697 3.4105
R3496 avdd.n6701 avdd.n6562 3.4105
R3497 avdd.n6562 avdd.n6561 3.4105
R3498 avdd.n6710 avdd.n6709 3.4105
R3499 avdd.n6717 avdd.n6559 3.4105
R3500 avdd.n6717 avdd.n6552 3.4105
R3501 avdd.n6722 avdd.n6556 3.4105
R3502 avdd.n6703 avdd.n6702 3.4105
R3503 avdd.n6720 avdd.n6719 3.4105
R3504 avdd.n6719 avdd.n6718 3.4105
R3505 avdd.n6716 avdd.n6715 3.4105
R3506 avdd.n6721 avdd.n6554 3.4105
R3507 avdd.n6554 avdd.n6553 3.4105
R3508 avdd.n6726 avdd.n6725 3.4105
R3509 avdd.n6730 avdd.n6729 3.4105
R3510 avdd.n6751 avdd.n6538 3.4105
R3511 avdd.n6749 avdd.n6544 3.4105
R3512 avdd.n6749 avdd.n6543 3.4105
R3513 avdd.n6731 avdd.n6543 3.4105
R3514 avdd.n6734 avdd.n6733 3.4105
R3515 avdd.n6737 avdd.n6736 3.4105
R3516 avdd.n6735 avdd.n6550 3.4105
R3517 avdd.n6550 avdd.n6549 3.4105
R3518 avdd.n6647 avdd.n6646 3.4105
R3519 avdd.n6646 avdd.n6645 3.4105
R3520 avdd.n6644 avdd.n6594 3.4105
R3521 avdd.n6644 avdd.n6643 3.4105
R3522 avdd.n6594 avdd.n6588 3.4105
R3523 avdd.n6588 avdd.n6587 3.4105
R3524 avdd.n6763 avdd.n6756 3.4105
R3525 avdd.n6763 avdd.n6754 3.4105
R3526 avdd.n6763 avdd.n6755 3.4105
R3527 avdd.n6967 avdd.n6755 3.4105
R3528 avdd.n6959 avdd.n6958 3.4105
R3529 avdd.n6957 avdd.n6956 3.4105
R3530 avdd.n6962 avdd.n6764 3.4105
R3531 avdd.n6825 avdd.n6824 3.4105
R3532 avdd.n6832 avdd.n6823 3.4105
R3533 avdd.n6832 avdd.n6831 3.4105
R3534 avdd.n6841 avdd.n6819 3.4105
R3535 avdd.n6841 avdd.n6813 3.4105
R3536 avdd.n6847 avdd.n6816 3.4105
R3537 avdd.n6843 avdd.n6842 3.4105
R3538 avdd.n6846 avdd.n6815 3.4105
R3539 avdd.n6815 avdd.n6814 3.4105
R3540 avdd.n6851 avdd.n6850 3.4105
R3541 avdd.n6858 avdd.n6812 3.4105
R3542 avdd.n6858 avdd.n6802 3.4105
R3543 avdd.n6857 avdd.n6856 3.4105
R3544 avdd.n6865 avdd.n6864 3.4105
R3545 avdd.n6868 avdd.n6800 3.4105
R3546 avdd.n6881 avdd.n6880 3.4105
R3547 avdd.n6809 avdd.n6808 3.4105
R3548 avdd.n6874 avdd.n6873 3.4105
R3549 avdd.n6873 avdd.n6872 3.4105
R3550 avdd.n6870 avdd.n6869 3.4105
R3551 avdd.n6884 avdd.n6883 3.4105
R3552 avdd.n6885 avdd.n6884 3.4105
R3553 avdd.n6797 avdd.n6796 3.4105
R3554 avdd.n6796 avdd.n6795 3.4105
R3555 avdd.n6876 avdd.n6791 3.4105
R3556 avdd.n6878 avdd.n6877 3.4105
R3557 avdd.n6894 avdd.n6893 3.4105
R3558 avdd.n6893 avdd.n6892 3.4105
R3559 avdd.n6793 avdd.n6792 3.4105
R3560 avdd.n6890 avdd.n6794 3.4105
R3561 avdd.n6890 avdd.n6889 3.4105
R3562 avdd.n6900 avdd.n6899 3.4105
R3563 avdd.n6905 avdd.n6904 3.4105
R3564 avdd.n6898 avdd.n6786 3.4105
R3565 avdd.n6902 avdd.n6901 3.4105
R3566 avdd.n6907 avdd.n6906 3.4105
R3567 avdd.n6912 avdd.n6782 3.4105
R3568 avdd.n6912 avdd.n6776 3.4105
R3569 avdd.n6922 avdd.n6779 3.4105
R3570 avdd.n6914 avdd.n6913 3.4105
R3571 avdd.n6917 avdd.n6778 3.4105
R3572 avdd.n6778 avdd.n6777 3.4105
R3573 avdd.n6926 avdd.n6925 3.4105
R3574 avdd.n6933 avdd.n6775 3.4105
R3575 avdd.n6933 avdd.n6768 3.4105
R3576 avdd.n6938 avdd.n6772 3.4105
R3577 avdd.n6919 avdd.n6918 3.4105
R3578 avdd.n6936 avdd.n6935 3.4105
R3579 avdd.n6935 avdd.n6934 3.4105
R3580 avdd.n6932 avdd.n6931 3.4105
R3581 avdd.n6937 avdd.n6770 3.4105
R3582 avdd.n6770 avdd.n6769 3.4105
R3583 avdd.n6942 avdd.n6941 3.4105
R3584 avdd.n6946 avdd.n6945 3.4105
R3585 avdd.n6967 avdd.n6754 3.4105
R3586 avdd.n6965 avdd.n6760 3.4105
R3587 avdd.n6965 avdd.n6759 3.4105
R3588 avdd.n6947 avdd.n6759 3.4105
R3589 avdd.n6950 avdd.n6949 3.4105
R3590 avdd.n6953 avdd.n6952 3.4105
R3591 avdd.n6951 avdd.n6766 3.4105
R3592 avdd.n6766 avdd.n6765 3.4105
R3593 avdd.n6863 avdd.n6862 3.4105
R3594 avdd.n6862 avdd.n6861 3.4105
R3595 avdd.n6860 avdd.n6810 3.4105
R3596 avdd.n6860 avdd.n6859 3.4105
R3597 avdd.n6810 avdd.n6804 3.4105
R3598 avdd.n6804 avdd.n6803 3.4105
R3599 avdd.n6979 avdd.n6972 3.4105
R3600 avdd.n6979 avdd.n6970 3.4105
R3601 avdd.n6979 avdd.n6971 3.4105
R3602 avdd.n7183 avdd.n6971 3.4105
R3603 avdd.n7175 avdd.n7174 3.4105
R3604 avdd.n7173 avdd.n7172 3.4105
R3605 avdd.n7178 avdd.n6980 3.4105
R3606 avdd.n7041 avdd.n7040 3.4105
R3607 avdd.n7048 avdd.n7039 3.4105
R3608 avdd.n7048 avdd.n7047 3.4105
R3609 avdd.n7057 avdd.n7035 3.4105
R3610 avdd.n7057 avdd.n7029 3.4105
R3611 avdd.n7063 avdd.n7032 3.4105
R3612 avdd.n7059 avdd.n7058 3.4105
R3613 avdd.n7062 avdd.n7031 3.4105
R3614 avdd.n7031 avdd.n7030 3.4105
R3615 avdd.n7067 avdd.n7066 3.4105
R3616 avdd.n7074 avdd.n7028 3.4105
R3617 avdd.n7074 avdd.n7018 3.4105
R3618 avdd.n7073 avdd.n7072 3.4105
R3619 avdd.n7081 avdd.n7080 3.4105
R3620 avdd.n7084 avdd.n7016 3.4105
R3621 avdd.n7097 avdd.n7096 3.4105
R3622 avdd.n7025 avdd.n7024 3.4105
R3623 avdd.n7090 avdd.n7089 3.4105
R3624 avdd.n7089 avdd.n7088 3.4105
R3625 avdd.n7086 avdd.n7085 3.4105
R3626 avdd.n7100 avdd.n7099 3.4105
R3627 avdd.n7101 avdd.n7100 3.4105
R3628 avdd.n7013 avdd.n7012 3.4105
R3629 avdd.n7012 avdd.n7011 3.4105
R3630 avdd.n7092 avdd.n7007 3.4105
R3631 avdd.n7094 avdd.n7093 3.4105
R3632 avdd.n7110 avdd.n7109 3.4105
R3633 avdd.n7109 avdd.n7108 3.4105
R3634 avdd.n7009 avdd.n7008 3.4105
R3635 avdd.n7106 avdd.n7010 3.4105
R3636 avdd.n7106 avdd.n7105 3.4105
R3637 avdd.n7116 avdd.n7115 3.4105
R3638 avdd.n7121 avdd.n7120 3.4105
R3639 avdd.n7114 avdd.n7002 3.4105
R3640 avdd.n7118 avdd.n7117 3.4105
R3641 avdd.n7123 avdd.n7122 3.4105
R3642 avdd.n7128 avdd.n6998 3.4105
R3643 avdd.n7128 avdd.n6992 3.4105
R3644 avdd.n7138 avdd.n6995 3.4105
R3645 avdd.n7130 avdd.n7129 3.4105
R3646 avdd.n7133 avdd.n6994 3.4105
R3647 avdd.n6994 avdd.n6993 3.4105
R3648 avdd.n7142 avdd.n7141 3.4105
R3649 avdd.n7149 avdd.n6991 3.4105
R3650 avdd.n7149 avdd.n6984 3.4105
R3651 avdd.n7154 avdd.n6988 3.4105
R3652 avdd.n7135 avdd.n7134 3.4105
R3653 avdd.n7152 avdd.n7151 3.4105
R3654 avdd.n7151 avdd.n7150 3.4105
R3655 avdd.n7148 avdd.n7147 3.4105
R3656 avdd.n7153 avdd.n6986 3.4105
R3657 avdd.n6986 avdd.n6985 3.4105
R3658 avdd.n7158 avdd.n7157 3.4105
R3659 avdd.n7162 avdd.n7161 3.4105
R3660 avdd.n7183 avdd.n6970 3.4105
R3661 avdd.n7181 avdd.n6976 3.4105
R3662 avdd.n7181 avdd.n6975 3.4105
R3663 avdd.n7163 avdd.n6975 3.4105
R3664 avdd.n7166 avdd.n7165 3.4105
R3665 avdd.n7169 avdd.n7168 3.4105
R3666 avdd.n7167 avdd.n6982 3.4105
R3667 avdd.n6982 avdd.n6981 3.4105
R3668 avdd.n7079 avdd.n7078 3.4105
R3669 avdd.n7078 avdd.n7077 3.4105
R3670 avdd.n7076 avdd.n7026 3.4105
R3671 avdd.n7076 avdd.n7075 3.4105
R3672 avdd.n7026 avdd.n7020 3.4105
R3673 avdd.n7020 avdd.n7019 3.4105
R3674 avdd.n7195 avdd.n7188 3.4105
R3675 avdd.n7195 avdd.n7186 3.4105
R3676 avdd.n7195 avdd.n7187 3.4105
R3677 avdd.n7399 avdd.n7187 3.4105
R3678 avdd.n7391 avdd.n7390 3.4105
R3679 avdd.n7389 avdd.n7388 3.4105
R3680 avdd.n7394 avdd.n7196 3.4105
R3681 avdd.n7257 avdd.n7256 3.4105
R3682 avdd.n7264 avdd.n7255 3.4105
R3683 avdd.n7264 avdd.n7263 3.4105
R3684 avdd.n7273 avdd.n7251 3.4105
R3685 avdd.n7273 avdd.n7245 3.4105
R3686 avdd.n7279 avdd.n7248 3.4105
R3687 avdd.n7275 avdd.n7274 3.4105
R3688 avdd.n7278 avdd.n7247 3.4105
R3689 avdd.n7247 avdd.n7246 3.4105
R3690 avdd.n7283 avdd.n7282 3.4105
R3691 avdd.n7290 avdd.n7244 3.4105
R3692 avdd.n7290 avdd.n7234 3.4105
R3693 avdd.n7289 avdd.n7288 3.4105
R3694 avdd.n7297 avdd.n7296 3.4105
R3695 avdd.n7300 avdd.n7232 3.4105
R3696 avdd.n7313 avdd.n7312 3.4105
R3697 avdd.n7241 avdd.n7240 3.4105
R3698 avdd.n7306 avdd.n7305 3.4105
R3699 avdd.n7305 avdd.n7304 3.4105
R3700 avdd.n7302 avdd.n7301 3.4105
R3701 avdd.n7316 avdd.n7315 3.4105
R3702 avdd.n7317 avdd.n7316 3.4105
R3703 avdd.n7229 avdd.n7228 3.4105
R3704 avdd.n7228 avdd.n7227 3.4105
R3705 avdd.n7308 avdd.n7223 3.4105
R3706 avdd.n7310 avdd.n7309 3.4105
R3707 avdd.n7326 avdd.n7325 3.4105
R3708 avdd.n7325 avdd.n7324 3.4105
R3709 avdd.n7225 avdd.n7224 3.4105
R3710 avdd.n7322 avdd.n7226 3.4105
R3711 avdd.n7322 avdd.n7321 3.4105
R3712 avdd.n7332 avdd.n7331 3.4105
R3713 avdd.n7337 avdd.n7336 3.4105
R3714 avdd.n7330 avdd.n7218 3.4105
R3715 avdd.n7334 avdd.n7333 3.4105
R3716 avdd.n7339 avdd.n7338 3.4105
R3717 avdd.n7344 avdd.n7214 3.4105
R3718 avdd.n7344 avdd.n7208 3.4105
R3719 avdd.n7354 avdd.n7211 3.4105
R3720 avdd.n7346 avdd.n7345 3.4105
R3721 avdd.n7349 avdd.n7210 3.4105
R3722 avdd.n7210 avdd.n7209 3.4105
R3723 avdd.n7358 avdd.n7357 3.4105
R3724 avdd.n7365 avdd.n7207 3.4105
R3725 avdd.n7365 avdd.n7200 3.4105
R3726 avdd.n7370 avdd.n7204 3.4105
R3727 avdd.n7351 avdd.n7350 3.4105
R3728 avdd.n7368 avdd.n7367 3.4105
R3729 avdd.n7367 avdd.n7366 3.4105
R3730 avdd.n7364 avdd.n7363 3.4105
R3731 avdd.n7369 avdd.n7202 3.4105
R3732 avdd.n7202 avdd.n7201 3.4105
R3733 avdd.n7374 avdd.n7373 3.4105
R3734 avdd.n7378 avdd.n7377 3.4105
R3735 avdd.n7399 avdd.n7186 3.4105
R3736 avdd.n7397 avdd.n7192 3.4105
R3737 avdd.n7397 avdd.n7191 3.4105
R3738 avdd.n7379 avdd.n7191 3.4105
R3739 avdd.n7382 avdd.n7381 3.4105
R3740 avdd.n7385 avdd.n7384 3.4105
R3741 avdd.n7383 avdd.n7198 3.4105
R3742 avdd.n7198 avdd.n7197 3.4105
R3743 avdd.n7295 avdd.n7294 3.4105
R3744 avdd.n7294 avdd.n7293 3.4105
R3745 avdd.n7292 avdd.n7242 3.4105
R3746 avdd.n7292 avdd.n7291 3.4105
R3747 avdd.n7242 avdd.n7236 3.4105
R3748 avdd.n7236 avdd.n7235 3.4105
R3749 avdd.n4617 avdd.n4555 3.38874
R3750 avdd.n4631 avdd.n4622 3.38874
R3751 avdd.n4677 avdd.n4676 3.38874
R3752 avdd avdd.n7453 3.35086
R3753 avdd avdd.n7492 3.35086
R3754 avdd avdd.n7552 3.35086
R3755 avdd avdd.n7592 3.35086
R3756 avdd avdd.n1818 3.35086
R3757 avdd avdd.n1644 3.35086
R3758 avdd avdd.n1728 3.35086
R3759 avdd avdd.n1680 3.35086
R3760 avdd.n7422 avdd 3.28549
R3761 avdd.n1820 avdd.n1819 3.23579
R3762 avdd.n1781 avdd.n1645 3.23579
R3763 avdd.n1730 avdd.n1729 3.23579
R3764 avdd.n1691 avdd.n1681 3.23579
R3765 avdd.n7454 avdd 3.20271
R3766 avdd.n7493 avdd 3.20271
R3767 avdd.n7553 avdd 3.20271
R3768 avdd.n7593 avdd 3.20271
R3769 avdd.n4643 avdd.n4642 3.15662
R3770 avdd.n7531 avdd.n7419 3.08362
R3771 avdd.n7628 avdd.n7627 3.08362
R3772 avdd.n7632 avdd.n7403 3.08362
R3773 avdd.n7528 avdd.n7527 3.08362
R3774 avdd.n1766 avdd.n1765 3.08362
R3775 avdd.n1769 avdd.n1650 3.08362
R3776 avdd.n1856 avdd.n1855 3.08362
R3777 avdd.n1866 avdd.n1865 3.08362
R3778 avdd.n7639 avdd 3.05331
R3779 avdd.n4639 avdd.n4617 3.01226
R3780 avdd.n4622 avdd.n4567 3.01226
R3781 avdd.n4676 avdd.n4675 3.01226
R3782 avdd.n4639 avdd.n4618 2.63579
R3783 avdd.n4633 avdd.n4632 2.63579
R3784 avdd.n4675 avdd.n4573 2.63579
R3785 avdd.n7501 avdd.n7500 2.61352
R3786 avdd.n7573 avdd.n7572 2.61352
R3787 avdd.n7601 avdd.n7600 2.61352
R3788 avdd.n7473 avdd.n7426 2.61352
R3789 avdd.n1709 avdd.n1660 2.61352
R3790 avdd.n1740 avdd.n1739 2.61352
R3791 avdd.n1799 avdd.n1624 2.61352
R3792 avdd.n1830 avdd.n1829 2.61352
R3793 avdd.n7422 avdd 2.57272
R3794 avdd.n7526 avdd.n7525 2.29662
R3795 avdd.n7535 avdd.n7534 2.29662
R3796 avdd.n7626 avdd.n7625 2.29662
R3797 avdd.n7637 avdd.n7636 2.29662
R3798 avdd.n1854 avdd.n1853 2.29662
R3799 avdd.n1772 avdd.n1647 2.29662
R3800 avdd.n1764 avdd.n1763 2.29662
R3801 avdd.n1869 avdd.n1618 2.29643
R3802 avdd.n7501 avdd.n7421 2.29594
R3803 avdd.n7574 avdd.n7573 2.29594
R3804 avdd.n7601 avdd.n7405 2.29594
R3805 avdd.n7474 avdd.n7473 2.29594
R3806 avdd.n1710 avdd.n1709 2.29594
R3807 avdd.n1740 avdd.n1649 2.29594
R3808 avdd.n1800 avdd.n1799 2.29594
R3809 avdd.n1830 avdd.n1620 2.29594
R3810 avdd.n4683 avdd.n4568 2.25932
R3811 avdd avdd.n7402 2.15303
R3812 avdd avdd.n4458 2.13383
R3813 avdd.n1860 avdd 2.0485
R3814 avdd.n1653 avdd 2.0485
R3815 avdd.n5019 avdd.n5011 2.03035
R3816 avdd.n5235 avdd.n5227 2.03035
R3817 avdd.n5451 avdd.n5443 2.03035
R3818 avdd.n5667 avdd.n5659 2.03035
R3819 avdd.n5883 avdd.n5875 2.03035
R3820 avdd.n6099 avdd.n6091 2.03035
R3821 avdd.n6315 avdd.n6307 2.03035
R3822 avdd.n6531 avdd.n6523 2.03035
R3823 avdd.n6747 avdd.n6739 2.03035
R3824 avdd.n6963 avdd.n6955 2.03035
R3825 avdd.n7179 avdd.n7171 2.03035
R3826 avdd.n7395 avdd.n7387 2.03035
R3827 avdd.n2021 avdd.n2020 2.03017
R3828 avdd.n2295 avdd.n2294 2.03017
R3829 avdd.n2510 avdd.n2509 2.03017
R3830 avdd.n2725 avdd.n2724 2.03017
R3831 avdd.n2940 avdd.n2939 2.03017
R3832 avdd.n3155 avdd.n3154 2.03017
R3833 avdd.n3315 avdd.n3313 2.03017
R3834 avdd.n3530 avdd.n3528 2.03017
R3835 avdd.n3745 avdd.n3743 2.03017
R3836 avdd.n3960 avdd.n3958 2.03017
R3837 avdd.n4175 avdd.n4173 2.03017
R3838 avdd.n4390 avdd.n4388 2.03017
R3839 avdd.n1911 avdd.n1910 2.01741
R3840 avdd.n2165 avdd.n2164 2.01741
R3841 avdd.n2380 avdd.n2379 2.01741
R3842 avdd.n2595 avdd.n2594 2.01741
R3843 avdd.n2810 avdd.n2809 2.01741
R3844 avdd.n3025 avdd.n3024 2.01741
R3845 avdd.n3201 avdd.n3200 2.01741
R3846 avdd.n3416 avdd.n3415 2.01741
R3847 avdd.n3631 avdd.n3630 2.01741
R3848 avdd.n3846 avdd.n3845 2.01741
R3849 avdd.n4061 avdd.n4060 2.01741
R3850 avdd.n4276 avdd.n4275 2.01741
R3851 avdd.n81 avdd.n80 2.01741
R3852 avdd.n211 avdd.n210 2.01741
R3853 avdd.n341 avdd.n340 2.01741
R3854 avdd.n471 avdd.n470 2.01741
R3855 avdd.n601 avdd.n600 2.01741
R3856 avdd.n731 avdd.n730 2.01741
R3857 avdd.n861 avdd.n860 2.01741
R3858 avdd.n991 avdd.n990 2.01741
R3859 avdd.n1121 avdd.n1120 2.01741
R3860 avdd.n1251 avdd.n1250 2.01741
R3861 avdd.n1381 avdd.n1380 2.01741
R3862 avdd.n1511 avdd.n1510 2.01741
R3863 avdd.n4887 avdd.n4886 2.01723
R3864 avdd.n5103 avdd.n5102 2.01723
R3865 avdd.n5319 avdd.n5318 2.01723
R3866 avdd.n5535 avdd.n5534 2.01723
R3867 avdd.n5751 avdd.n5750 2.01723
R3868 avdd.n5967 avdd.n5966 2.01723
R3869 avdd.n6183 avdd.n6182 2.01723
R3870 avdd.n6399 avdd.n6398 2.01723
R3871 avdd.n6615 avdd.n6614 2.01723
R3872 avdd.n6831 avdd.n6830 2.01723
R3873 avdd.n7047 avdd.n7046 2.01723
R3874 avdd.n7263 avdd.n7262 2.01723
R3875 avdd.n7748 avdd.n7747 2.01723
R3876 avdd.n10227 avdd.n10226 2.01723
R3877 avdd.n9977 avdd.n9976 2.01723
R3878 avdd.n9863 avdd.n9862 2.01723
R3879 avdd.n9749 avdd.n9748 2.01723
R3880 avdd.n9636 avdd.n9635 2.01723
R3881 avdd.n9521 avdd.n9520 2.01723
R3882 avdd.n9407 avdd.n9406 2.01723
R3883 avdd.n9293 avdd.n9292 2.01723
R3884 avdd.n9179 avdd.n9178 2.01723
R3885 avdd.n9065 avdd.n9064 2.01723
R3886 avdd.n8951 avdd.n8950 2.01723
R3887 avdd.n2040 avdd.n2039 1.93672
R3888 avdd.n2042 avdd.n2041 1.93672
R3889 avdd.n2050 avdd.n1976 1.93672
R3890 avdd.n1969 avdd.n1962 1.93672
R3891 avdd.n2061 avdd.n1970 1.93672
R3892 avdd.n2075 avdd.n2074 1.93672
R3893 avdd.n1945 avdd.n1886 1.93672
R3894 avdd.n1944 avdd.n1943 1.93672
R3895 avdd.n1932 avdd.n1931 1.93672
R3896 avdd.n2027 avdd.n2020 1.93672
R3897 avdd.n2282 avdd.n2281 1.93672
R3898 avdd.n2280 avdd.n2279 1.93672
R3899 avdd.n2261 avdd.n2260 1.93672
R3900 avdd.n2233 avdd.n2117 1.93672
R3901 avdd.n2242 avdd.n2241 1.93672
R3902 avdd.n2221 avdd.n2125 1.93672
R3903 avdd.n2202 avdd.n2201 1.93672
R3904 avdd.n2200 avdd.n2199 1.93672
R3905 avdd.n2185 avdd.n2184 1.93672
R3906 avdd.n2294 avdd.n2099 1.93672
R3907 avdd.n2497 avdd.n2496 1.93672
R3908 avdd.n2495 avdd.n2494 1.93672
R3909 avdd.n2476 avdd.n2475 1.93672
R3910 avdd.n2448 avdd.n2332 1.93672
R3911 avdd.n2457 avdd.n2456 1.93672
R3912 avdd.n2436 avdd.n2340 1.93672
R3913 avdd.n2417 avdd.n2416 1.93672
R3914 avdd.n2415 avdd.n2414 1.93672
R3915 avdd.n2400 avdd.n2399 1.93672
R3916 avdd.n2509 avdd.n2314 1.93672
R3917 avdd.n2712 avdd.n2711 1.93672
R3918 avdd.n2710 avdd.n2709 1.93672
R3919 avdd.n2691 avdd.n2690 1.93672
R3920 avdd.n2663 avdd.n2547 1.93672
R3921 avdd.n2672 avdd.n2671 1.93672
R3922 avdd.n2651 avdd.n2555 1.93672
R3923 avdd.n2632 avdd.n2631 1.93672
R3924 avdd.n2630 avdd.n2629 1.93672
R3925 avdd.n2615 avdd.n2614 1.93672
R3926 avdd.n2724 avdd.n2529 1.93672
R3927 avdd.n2927 avdd.n2926 1.93672
R3928 avdd.n2925 avdd.n2924 1.93672
R3929 avdd.n2906 avdd.n2905 1.93672
R3930 avdd.n2878 avdd.n2762 1.93672
R3931 avdd.n2887 avdd.n2886 1.93672
R3932 avdd.n2866 avdd.n2770 1.93672
R3933 avdd.n2847 avdd.n2846 1.93672
R3934 avdd.n2845 avdd.n2844 1.93672
R3935 avdd.n2830 avdd.n2829 1.93672
R3936 avdd.n2939 avdd.n2744 1.93672
R3937 avdd.n3142 avdd.n3141 1.93672
R3938 avdd.n3140 avdd.n3139 1.93672
R3939 avdd.n3121 avdd.n3120 1.93672
R3940 avdd.n3093 avdd.n2977 1.93672
R3941 avdd.n3102 avdd.n3101 1.93672
R3942 avdd.n3081 avdd.n2985 1.93672
R3943 avdd.n3062 avdd.n3061 1.93672
R3944 avdd.n3060 avdd.n3059 1.93672
R3945 avdd.n3045 avdd.n3044 1.93672
R3946 avdd.n3154 avdd.n2959 1.93672
R3947 avdd.n3329 avdd.n3328 1.93672
R3948 avdd.n3331 avdd.n3330 1.93672
R3949 avdd.n3339 avdd.n3266 1.93672
R3950 avdd.n3259 avdd.n3252 1.93672
R3951 avdd.n3350 avdd.n3260 1.93672
R3952 avdd.n3364 avdd.n3363 1.93672
R3953 avdd.n3235 avdd.n3176 1.93672
R3954 avdd.n3234 avdd.n3233 1.93672
R3955 avdd.n3222 avdd.n3221 1.93672
R3956 avdd.n3321 avdd.n3313 1.93672
R3957 avdd.n3544 avdd.n3543 1.93672
R3958 avdd.n3546 avdd.n3545 1.93672
R3959 avdd.n3554 avdd.n3481 1.93672
R3960 avdd.n3474 avdd.n3467 1.93672
R3961 avdd.n3565 avdd.n3475 1.93672
R3962 avdd.n3579 avdd.n3578 1.93672
R3963 avdd.n3450 avdd.n3391 1.93672
R3964 avdd.n3449 avdd.n3448 1.93672
R3965 avdd.n3437 avdd.n3436 1.93672
R3966 avdd.n3536 avdd.n3528 1.93672
R3967 avdd.n3759 avdd.n3758 1.93672
R3968 avdd.n3761 avdd.n3760 1.93672
R3969 avdd.n3769 avdd.n3696 1.93672
R3970 avdd.n3689 avdd.n3682 1.93672
R3971 avdd.n3780 avdd.n3690 1.93672
R3972 avdd.n3794 avdd.n3793 1.93672
R3973 avdd.n3665 avdd.n3606 1.93672
R3974 avdd.n3664 avdd.n3663 1.93672
R3975 avdd.n3652 avdd.n3651 1.93672
R3976 avdd.n3751 avdd.n3743 1.93672
R3977 avdd.n3974 avdd.n3973 1.93672
R3978 avdd.n3976 avdd.n3975 1.93672
R3979 avdd.n3984 avdd.n3911 1.93672
R3980 avdd.n3904 avdd.n3897 1.93672
R3981 avdd.n3995 avdd.n3905 1.93672
R3982 avdd.n4009 avdd.n4008 1.93672
R3983 avdd.n3880 avdd.n3821 1.93672
R3984 avdd.n3879 avdd.n3878 1.93672
R3985 avdd.n3867 avdd.n3866 1.93672
R3986 avdd.n3966 avdd.n3958 1.93672
R3987 avdd.n4189 avdd.n4188 1.93672
R3988 avdd.n4191 avdd.n4190 1.93672
R3989 avdd.n4199 avdd.n4126 1.93672
R3990 avdd.n4119 avdd.n4112 1.93672
R3991 avdd.n4210 avdd.n4120 1.93672
R3992 avdd.n4224 avdd.n4223 1.93672
R3993 avdd.n4095 avdd.n4036 1.93672
R3994 avdd.n4094 avdd.n4093 1.93672
R3995 avdd.n4082 avdd.n4081 1.93672
R3996 avdd.n4181 avdd.n4173 1.93672
R3997 avdd.n4404 avdd.n4403 1.93672
R3998 avdd.n4406 avdd.n4405 1.93672
R3999 avdd.n4414 avdd.n4341 1.93672
R4000 avdd.n4334 avdd.n4327 1.93672
R4001 avdd.n4425 avdd.n4335 1.93672
R4002 avdd.n4439 avdd.n4438 1.93672
R4003 avdd.n4310 avdd.n4251 1.93672
R4004 avdd.n4309 avdd.n4308 1.93672
R4005 avdd.n4297 avdd.n4296 1.93672
R4006 avdd.n4396 avdd.n4388 1.93672
R4007 avdd.n4908 avdd.n4907 1.93672
R4008 avdd.n4922 avdd.n4921 1.93672
R4009 avdd.n4924 avdd.n4923 1.93672
R4010 avdd.n4943 avdd.n4847 1.93672
R4011 avdd.n4955 avdd.n4839 1.93672
R4012 avdd.n4964 avdd.n4963 1.93672
R4013 avdd.n4983 avdd.n4982 1.93672
R4014 avdd.n4999 avdd.n4998 1.93672
R4015 avdd.n5002 avdd.n5000 1.93672
R4016 avdd.n5013 avdd.n5011 1.93672
R4017 avdd.n5124 avdd.n5123 1.93672
R4018 avdd.n5138 avdd.n5137 1.93672
R4019 avdd.n5140 avdd.n5139 1.93672
R4020 avdd.n5159 avdd.n5063 1.93672
R4021 avdd.n5171 avdd.n5055 1.93672
R4022 avdd.n5180 avdd.n5179 1.93672
R4023 avdd.n5199 avdd.n5198 1.93672
R4024 avdd.n5215 avdd.n5214 1.93672
R4025 avdd.n5218 avdd.n5216 1.93672
R4026 avdd.n5229 avdd.n5227 1.93672
R4027 avdd.n5340 avdd.n5339 1.93672
R4028 avdd.n5354 avdd.n5353 1.93672
R4029 avdd.n5356 avdd.n5355 1.93672
R4030 avdd.n5375 avdd.n5279 1.93672
R4031 avdd.n5387 avdd.n5271 1.93672
R4032 avdd.n5396 avdd.n5395 1.93672
R4033 avdd.n5415 avdd.n5414 1.93672
R4034 avdd.n5431 avdd.n5430 1.93672
R4035 avdd.n5434 avdd.n5432 1.93672
R4036 avdd.n5445 avdd.n5443 1.93672
R4037 avdd.n5556 avdd.n5555 1.93672
R4038 avdd.n5570 avdd.n5569 1.93672
R4039 avdd.n5572 avdd.n5571 1.93672
R4040 avdd.n5591 avdd.n5495 1.93672
R4041 avdd.n5603 avdd.n5487 1.93672
R4042 avdd.n5612 avdd.n5611 1.93672
R4043 avdd.n5631 avdd.n5630 1.93672
R4044 avdd.n5647 avdd.n5646 1.93672
R4045 avdd.n5650 avdd.n5648 1.93672
R4046 avdd.n5661 avdd.n5659 1.93672
R4047 avdd.n5772 avdd.n5771 1.93672
R4048 avdd.n5786 avdd.n5785 1.93672
R4049 avdd.n5788 avdd.n5787 1.93672
R4050 avdd.n5807 avdd.n5711 1.93672
R4051 avdd.n5819 avdd.n5703 1.93672
R4052 avdd.n5828 avdd.n5827 1.93672
R4053 avdd.n5847 avdd.n5846 1.93672
R4054 avdd.n5863 avdd.n5862 1.93672
R4055 avdd.n5866 avdd.n5864 1.93672
R4056 avdd.n5877 avdd.n5875 1.93672
R4057 avdd.n5988 avdd.n5987 1.93672
R4058 avdd.n6002 avdd.n6001 1.93672
R4059 avdd.n6004 avdd.n6003 1.93672
R4060 avdd.n6023 avdd.n5927 1.93672
R4061 avdd.n6035 avdd.n5919 1.93672
R4062 avdd.n6044 avdd.n6043 1.93672
R4063 avdd.n6063 avdd.n6062 1.93672
R4064 avdd.n6079 avdd.n6078 1.93672
R4065 avdd.n6082 avdd.n6080 1.93672
R4066 avdd.n6093 avdd.n6091 1.93672
R4067 avdd.n6204 avdd.n6203 1.93672
R4068 avdd.n6218 avdd.n6217 1.93672
R4069 avdd.n6220 avdd.n6219 1.93672
R4070 avdd.n6239 avdd.n6143 1.93672
R4071 avdd.n6251 avdd.n6135 1.93672
R4072 avdd.n6260 avdd.n6259 1.93672
R4073 avdd.n6279 avdd.n6278 1.93672
R4074 avdd.n6295 avdd.n6294 1.93672
R4075 avdd.n6298 avdd.n6296 1.93672
R4076 avdd.n6309 avdd.n6307 1.93672
R4077 avdd.n6420 avdd.n6419 1.93672
R4078 avdd.n6434 avdd.n6433 1.93672
R4079 avdd.n6436 avdd.n6435 1.93672
R4080 avdd.n6455 avdd.n6359 1.93672
R4081 avdd.n6467 avdd.n6351 1.93672
R4082 avdd.n6476 avdd.n6475 1.93672
R4083 avdd.n6495 avdd.n6494 1.93672
R4084 avdd.n6511 avdd.n6510 1.93672
R4085 avdd.n6514 avdd.n6512 1.93672
R4086 avdd.n6525 avdd.n6523 1.93672
R4087 avdd.n6636 avdd.n6635 1.93672
R4088 avdd.n6650 avdd.n6649 1.93672
R4089 avdd.n6652 avdd.n6651 1.93672
R4090 avdd.n6671 avdd.n6575 1.93672
R4091 avdd.n6683 avdd.n6567 1.93672
R4092 avdd.n6692 avdd.n6691 1.93672
R4093 avdd.n6711 avdd.n6710 1.93672
R4094 avdd.n6727 avdd.n6726 1.93672
R4095 avdd.n6730 avdd.n6728 1.93672
R4096 avdd.n6741 avdd.n6739 1.93672
R4097 avdd.n6852 avdd.n6851 1.93672
R4098 avdd.n6866 avdd.n6865 1.93672
R4099 avdd.n6868 avdd.n6867 1.93672
R4100 avdd.n6887 avdd.n6791 1.93672
R4101 avdd.n6899 avdd.n6783 1.93672
R4102 avdd.n6908 avdd.n6907 1.93672
R4103 avdd.n6927 avdd.n6926 1.93672
R4104 avdd.n6943 avdd.n6942 1.93672
R4105 avdd.n6946 avdd.n6944 1.93672
R4106 avdd.n6957 avdd.n6955 1.93672
R4107 avdd.n7068 avdd.n7067 1.93672
R4108 avdd.n7082 avdd.n7081 1.93672
R4109 avdd.n7084 avdd.n7083 1.93672
R4110 avdd.n7103 avdd.n7007 1.93672
R4111 avdd.n7115 avdd.n6999 1.93672
R4112 avdd.n7124 avdd.n7123 1.93672
R4113 avdd.n7143 avdd.n7142 1.93672
R4114 avdd.n7159 avdd.n7158 1.93672
R4115 avdd.n7162 avdd.n7160 1.93672
R4116 avdd.n7173 avdd.n7171 1.93672
R4117 avdd.n7284 avdd.n7283 1.93672
R4118 avdd.n7298 avdd.n7297 1.93672
R4119 avdd.n7300 avdd.n7299 1.93672
R4120 avdd.n7319 avdd.n7223 1.93672
R4121 avdd.n7331 avdd.n7215 1.93672
R4122 avdd.n7340 avdd.n7339 1.93672
R4123 avdd.n7359 avdd.n7358 1.93672
R4124 avdd.n7375 avdd.n7374 1.93672
R4125 avdd.n7378 avdd.n7376 1.93672
R4126 avdd.n7389 avdd.n7387 1.93672
R4127 avdd.n7713 avdd.n7712 1.93672
R4128 avdd.n7732 avdd.n7731 1.93672
R4129 avdd.n7691 avdd.n7690 1.93672
R4130 avdd.n7672 avdd.n7671 1.93672
R4131 avdd.n7657 avdd.n7656 1.93672
R4132 avdd.n7660 avdd.n7659 1.93672
R4133 avdd.n7802 avdd.n7801 1.93672
R4134 avdd.n7822 avdd.n7821 1.93672
R4135 avdd.n7838 avdd.n7837 1.93672
R4136 avdd.n7785 avdd.n7784 1.93672
R4137 avdd.n10192 avdd.n10191 1.93672
R4138 avdd.n10211 avdd.n10210 1.93672
R4139 avdd.n10170 avdd.n10169 1.93672
R4140 avdd.n10151 avdd.n10150 1.93672
R4141 avdd.n10135 avdd.n10134 1.93672
R4142 avdd.n10139 avdd.n10138 1.93672
R4143 avdd.n10060 avdd.n10059 1.93672
R4144 avdd.n10080 avdd.n10079 1.93672
R4145 avdd.n10096 avdd.n10095 1.93672
R4146 avdd.n10045 avdd.n10044 1.93672
R4147 avdd.n9996 avdd.n9995 1.93672
R4148 avdd.n10017 avdd.n10016 1.93672
R4149 avdd.n9954 avdd.n9953 1.93672
R4150 avdd.n9935 avdd.n9934 1.93672
R4151 avdd.n10275 avdd.n10274 1.93672
R4152 avdd.n10277 avdd.n10276 1.93672
R4153 avdd.n10292 avdd.n10291 1.93672
R4154 avdd.n10312 avdd.n10311 1.93672
R4155 avdd.n10328 avdd.n10327 1.93672
R4156 avdd.n10261 avdd.n10260 1.93672
R4157 avdd.n9882 avdd.n9881 1.93672
R4158 avdd.n9903 avdd.n9902 1.93672
R4159 avdd.n9840 avdd.n9839 1.93672
R4160 avdd.n9821 avdd.n9820 1.93672
R4161 avdd.n10377 avdd.n10376 1.93672
R4162 avdd.n10379 avdd.n10378 1.93672
R4163 avdd.n10394 avdd.n10393 1.93672
R4164 avdd.n10414 avdd.n10413 1.93672
R4165 avdd.n10430 avdd.n10429 1.93672
R4166 avdd.n10363 avdd.n10362 1.93672
R4167 avdd.n9768 avdd.n9767 1.93672
R4168 avdd.n9789 avdd.n9788 1.93672
R4169 avdd.n9726 avdd.n9725 1.93672
R4170 avdd.n9707 avdd.n9706 1.93672
R4171 avdd.n10479 avdd.n10478 1.93672
R4172 avdd.n10481 avdd.n10480 1.93672
R4173 avdd.n10496 avdd.n10495 1.93672
R4174 avdd.n10516 avdd.n10515 1.93672
R4175 avdd.n10532 avdd.n10531 1.93672
R4176 avdd.n10465 avdd.n10464 1.93672
R4177 avdd.n9655 avdd.n9654 1.93672
R4178 avdd.n9676 avdd.n9675 1.93672
R4179 avdd.n9613 avdd.n9612 1.93672
R4180 avdd.n9594 avdd.n9593 1.93672
R4181 avdd.n10581 avdd.n10580 1.93672
R4182 avdd.n10583 avdd.n10582 1.93672
R4183 avdd.n10598 avdd.n10597 1.93672
R4184 avdd.n10618 avdd.n10617 1.93672
R4185 avdd.n10634 avdd.n10633 1.93672
R4186 avdd.n10567 avdd.n10566 1.93672
R4187 avdd.n9540 avdd.n9539 1.93672
R4188 avdd.n9561 avdd.n9560 1.93672
R4189 avdd.n9498 avdd.n9497 1.93672
R4190 avdd.n9479 avdd.n9478 1.93672
R4191 avdd.n10683 avdd.n10682 1.93672
R4192 avdd.n10685 avdd.n10684 1.93672
R4193 avdd.n10700 avdd.n10699 1.93672
R4194 avdd.n10720 avdd.n10719 1.93672
R4195 avdd.n10736 avdd.n10735 1.93672
R4196 avdd.n10669 avdd.n10668 1.93672
R4197 avdd.n9426 avdd.n9425 1.93672
R4198 avdd.n9447 avdd.n9446 1.93672
R4199 avdd.n9384 avdd.n9383 1.93672
R4200 avdd.n9365 avdd.n9364 1.93672
R4201 avdd.n10785 avdd.n10784 1.93672
R4202 avdd.n10787 avdd.n10786 1.93672
R4203 avdd.n10802 avdd.n10801 1.93672
R4204 avdd.n10822 avdd.n10821 1.93672
R4205 avdd.n10838 avdd.n10837 1.93672
R4206 avdd.n10771 avdd.n10770 1.93672
R4207 avdd.n9312 avdd.n9311 1.93672
R4208 avdd.n9333 avdd.n9332 1.93672
R4209 avdd.n9270 avdd.n9269 1.93672
R4210 avdd.n9251 avdd.n9250 1.93672
R4211 avdd.n10887 avdd.n10886 1.93672
R4212 avdd.n10889 avdd.n10888 1.93672
R4213 avdd.n10904 avdd.n10903 1.93672
R4214 avdd.n10924 avdd.n10923 1.93672
R4215 avdd.n10940 avdd.n10939 1.93672
R4216 avdd.n10873 avdd.n10872 1.93672
R4217 avdd.n9198 avdd.n9197 1.93672
R4218 avdd.n9219 avdd.n9218 1.93672
R4219 avdd.n9156 avdd.n9155 1.93672
R4220 avdd.n9137 avdd.n9136 1.93672
R4221 avdd.n10989 avdd.n10988 1.93672
R4222 avdd.n10991 avdd.n10990 1.93672
R4223 avdd.n11006 avdd.n11005 1.93672
R4224 avdd.n11026 avdd.n11025 1.93672
R4225 avdd.n11042 avdd.n11041 1.93672
R4226 avdd.n10975 avdd.n10974 1.93672
R4227 avdd.n9084 avdd.n9083 1.93672
R4228 avdd.n9105 avdd.n9104 1.93672
R4229 avdd.n9042 avdd.n9041 1.93672
R4230 avdd.n9023 avdd.n9022 1.93672
R4231 avdd.n11091 avdd.n11090 1.93672
R4232 avdd.n11093 avdd.n11092 1.93672
R4233 avdd.n11108 avdd.n11107 1.93672
R4234 avdd.n11128 avdd.n11127 1.93672
R4235 avdd.n11144 avdd.n11143 1.93672
R4236 avdd.n11077 avdd.n11076 1.93672
R4237 avdd.n8970 avdd.n8969 1.93672
R4238 avdd.n8991 avdd.n8990 1.93672
R4239 avdd.n8928 avdd.n8927 1.93672
R4240 avdd.n8909 avdd.n8908 1.93672
R4241 avdd.n11193 avdd.n11192 1.93672
R4242 avdd.n11195 avdd.n11194 1.93672
R4243 avdd.n11210 avdd.n11209 1.93672
R4244 avdd.n11230 avdd.n11229 1.93672
R4245 avdd.n11246 avdd.n11245 1.93672
R4246 avdd.n11179 avdd.n11178 1.93672
R4247 avdd.n8859 avdd.n8858 1.93672
R4248 avdd.n8843 avdd.n8842 1.93672
R4249 avdd.n8823 avdd.n8822 1.93672
R4250 avdd.n139 avdd.n138 1.93672
R4251 avdd.n143 avdd.n142 1.93672
R4252 avdd.n155 avdd.n154 1.93672
R4253 avdd.n174 avdd.n173 1.93672
R4254 avdd.n127 avdd.n126 1.93672
R4255 avdd.n107 avdd.n106 1.93672
R4256 avdd.n8808 avdd.n8807 1.93672
R4257 avdd.n8773 avdd.n8772 1.93672
R4258 avdd.n8757 avdd.n8756 1.93672
R4259 avdd.n8737 avdd.n8736 1.93672
R4260 avdd.n269 avdd.n268 1.93672
R4261 avdd.n273 avdd.n272 1.93672
R4262 avdd.n285 avdd.n284 1.93672
R4263 avdd.n304 avdd.n303 1.93672
R4264 avdd.n257 avdd.n256 1.93672
R4265 avdd.n237 avdd.n236 1.93672
R4266 avdd.n8722 avdd.n8721 1.93672
R4267 avdd.n8687 avdd.n8686 1.93672
R4268 avdd.n8671 avdd.n8670 1.93672
R4269 avdd.n8651 avdd.n8650 1.93672
R4270 avdd.n399 avdd.n398 1.93672
R4271 avdd.n403 avdd.n402 1.93672
R4272 avdd.n415 avdd.n414 1.93672
R4273 avdd.n434 avdd.n433 1.93672
R4274 avdd.n387 avdd.n386 1.93672
R4275 avdd.n367 avdd.n366 1.93672
R4276 avdd.n8636 avdd.n8635 1.93672
R4277 avdd.n8601 avdd.n8600 1.93672
R4278 avdd.n8585 avdd.n8584 1.93672
R4279 avdd.n8565 avdd.n8564 1.93672
R4280 avdd.n529 avdd.n528 1.93672
R4281 avdd.n533 avdd.n532 1.93672
R4282 avdd.n545 avdd.n544 1.93672
R4283 avdd.n564 avdd.n563 1.93672
R4284 avdd.n517 avdd.n516 1.93672
R4285 avdd.n497 avdd.n496 1.93672
R4286 avdd.n8550 avdd.n8549 1.93672
R4287 avdd.n8515 avdd.n8514 1.93672
R4288 avdd.n8499 avdd.n8498 1.93672
R4289 avdd.n8479 avdd.n8478 1.93672
R4290 avdd.n659 avdd.n658 1.93672
R4291 avdd.n663 avdd.n662 1.93672
R4292 avdd.n675 avdd.n674 1.93672
R4293 avdd.n694 avdd.n693 1.93672
R4294 avdd.n647 avdd.n646 1.93672
R4295 avdd.n627 avdd.n626 1.93672
R4296 avdd.n8464 avdd.n8463 1.93672
R4297 avdd.n8429 avdd.n8428 1.93672
R4298 avdd.n8413 avdd.n8412 1.93672
R4299 avdd.n8393 avdd.n8392 1.93672
R4300 avdd.n789 avdd.n788 1.93672
R4301 avdd.n793 avdd.n792 1.93672
R4302 avdd.n805 avdd.n804 1.93672
R4303 avdd.n824 avdd.n823 1.93672
R4304 avdd.n777 avdd.n776 1.93672
R4305 avdd.n757 avdd.n756 1.93672
R4306 avdd.n8378 avdd.n8377 1.93672
R4307 avdd.n8343 avdd.n8342 1.93672
R4308 avdd.n8327 avdd.n8326 1.93672
R4309 avdd.n8307 avdd.n8306 1.93672
R4310 avdd.n919 avdd.n918 1.93672
R4311 avdd.n923 avdd.n922 1.93672
R4312 avdd.n935 avdd.n934 1.93672
R4313 avdd.n954 avdd.n953 1.93672
R4314 avdd.n907 avdd.n906 1.93672
R4315 avdd.n887 avdd.n886 1.93672
R4316 avdd.n8292 avdd.n8291 1.93672
R4317 avdd.n8257 avdd.n8256 1.93672
R4318 avdd.n8241 avdd.n8240 1.93672
R4319 avdd.n8221 avdd.n8220 1.93672
R4320 avdd.n1049 avdd.n1048 1.93672
R4321 avdd.n1053 avdd.n1052 1.93672
R4322 avdd.n1065 avdd.n1064 1.93672
R4323 avdd.n1084 avdd.n1083 1.93672
R4324 avdd.n1037 avdd.n1036 1.93672
R4325 avdd.n1017 avdd.n1016 1.93672
R4326 avdd.n8206 avdd.n8205 1.93672
R4327 avdd.n8171 avdd.n8170 1.93672
R4328 avdd.n8155 avdd.n8154 1.93672
R4329 avdd.n8135 avdd.n8134 1.93672
R4330 avdd.n1179 avdd.n1178 1.93672
R4331 avdd.n1183 avdd.n1182 1.93672
R4332 avdd.n1195 avdd.n1194 1.93672
R4333 avdd.n1214 avdd.n1213 1.93672
R4334 avdd.n1167 avdd.n1166 1.93672
R4335 avdd.n1147 avdd.n1146 1.93672
R4336 avdd.n8120 avdd.n8119 1.93672
R4337 avdd.n8085 avdd.n8084 1.93672
R4338 avdd.n8069 avdd.n8068 1.93672
R4339 avdd.n8049 avdd.n8048 1.93672
R4340 avdd.n1309 avdd.n1308 1.93672
R4341 avdd.n1313 avdd.n1312 1.93672
R4342 avdd.n1325 avdd.n1324 1.93672
R4343 avdd.n1344 avdd.n1343 1.93672
R4344 avdd.n1297 avdd.n1296 1.93672
R4345 avdd.n1277 avdd.n1276 1.93672
R4346 avdd.n8034 avdd.n8033 1.93672
R4347 avdd.n7999 avdd.n7998 1.93672
R4348 avdd.n7983 avdd.n7982 1.93672
R4349 avdd.n7963 avdd.n7962 1.93672
R4350 avdd.n1439 avdd.n1438 1.93672
R4351 avdd.n1443 avdd.n1442 1.93672
R4352 avdd.n1455 avdd.n1454 1.93672
R4353 avdd.n1474 avdd.n1473 1.93672
R4354 avdd.n1427 avdd.n1426 1.93672
R4355 avdd.n1407 avdd.n1406 1.93672
R4356 avdd.n7948 avdd.n7947 1.93672
R4357 avdd.n7913 avdd.n7912 1.93672
R4358 avdd.n7897 avdd.n7896 1.93672
R4359 avdd.n7877 avdd.n7876 1.93672
R4360 avdd.n1569 avdd.n1568 1.93672
R4361 avdd.n1573 avdd.n1572 1.93672
R4362 avdd.n1585 avdd.n1584 1.93672
R4363 avdd.n1604 avdd.n1603 1.93672
R4364 avdd.n1557 avdd.n1556 1.93672
R4365 avdd.n1537 avdd.n1536 1.93672
R4366 avdd.n7862 avdd.n7861 1.93672
R4367 avdd.n4596 avdd.n4515 1.88285
R4368 avdd.n4625 avdd.n4568 1.88285
R4369 avdd.n7630 avdd 1.88073
R4370 avdd.n1708 avdd.n1707 1.85582
R4371 avdd.n1743 avdd.n1741 1.85582
R4372 avdd.n1798 avdd.n1797 1.85582
R4373 avdd.n1833 avdd.n1831 1.85582
R4374 avdd.n7503 avdd.n7502 1.84013
R4375 avdd.n7571 avdd.n7570 1.84013
R4376 avdd.n7603 avdd.n7602 1.84013
R4377 avdd.n7472 avdd.n7471 1.84013
R4378 avdd.n2036 avdd.n2004 1.77885
R4379 avdd.n2296 avdd.n2093 1.77885
R4380 avdd.n2511 avdd.n2308 1.77885
R4381 avdd.n2726 avdd.n2523 1.77885
R4382 avdd.n2941 avdd.n2738 1.77885
R4383 avdd.n3156 avdd.n2953 1.77885
R4384 avdd.n3325 avdd.n3294 1.77885
R4385 avdd.n3540 avdd.n3509 1.77885
R4386 avdd.n3755 avdd.n3724 1.77885
R4387 avdd.n3970 avdd.n3939 1.77885
R4388 avdd.n4185 avdd.n4154 1.77885
R4389 avdd.n4400 avdd.n4369 1.77885
R4390 avdd.n5021 avdd.n5020 1.77885
R4391 avdd.n5237 avdd.n5236 1.77885
R4392 avdd.n5453 avdd.n5452 1.77885
R4393 avdd.n5669 avdd.n5668 1.77885
R4394 avdd.n5885 avdd.n5884 1.77885
R4395 avdd.n6101 avdd.n6100 1.77885
R4396 avdd.n6317 avdd.n6316 1.77885
R4397 avdd.n6533 avdd.n6532 1.77885
R4398 avdd.n6749 avdd.n6748 1.77885
R4399 avdd.n6965 avdd.n6964 1.77885
R4400 avdd.n7181 avdd.n7180 1.77885
R4401 avdd.n7397 avdd.n7396 1.77885
R4402 avdd.n4917 avdd.n4861 1.70675
R4403 avdd.n5133 avdd.n5077 1.70675
R4404 avdd.n5349 avdd.n5293 1.70675
R4405 avdd.n5565 avdd.n5509 1.70675
R4406 avdd.n5781 avdd.n5725 1.70675
R4407 avdd.n5997 avdd.n5941 1.70675
R4408 avdd.n6213 avdd.n6157 1.70675
R4409 avdd.n6429 avdd.n6373 1.70675
R4410 avdd.n6645 avdd.n6589 1.70675
R4411 avdd.n6861 avdd.n6805 1.70675
R4412 avdd.n7077 avdd.n7021 1.70675
R4413 avdd.n7293 avdd.n7237 1.70675
R4414 avdd.n4919 avdd.n4861 1.706
R4415 avdd.n5135 avdd.n5077 1.706
R4416 avdd.n5351 avdd.n5293 1.706
R4417 avdd.n5567 avdd.n5509 1.706
R4418 avdd.n5783 avdd.n5725 1.706
R4419 avdd.n5999 avdd.n5941 1.706
R4420 avdd.n6215 avdd.n6157 1.706
R4421 avdd.n6431 avdd.n6373 1.706
R4422 avdd.n6647 avdd.n6589 1.706
R4423 avdd.n6863 avdd.n6805 1.706
R4424 avdd.n7079 avdd.n7021 1.706
R4425 avdd.n7295 avdd.n7237 1.706
R4426 avdd.n1898 avdd.n1897 1.7055
R4427 avdd.n1925 avdd.n1924 1.7055
R4428 avdd.n1955 avdd.n1954 1.7055
R4429 avdd.n2069 avdd.n2068 1.7055
R4430 avdd.n2067 avdd.n1957 1.7055
R4431 avdd.n2057 avdd.n1971 1.7055
R4432 avdd.n2056 avdd.n2055 1.7055
R4433 avdd.n1990 avdd.n1981 1.7055
R4434 avdd.n2035 avdd.n2034 1.7055
R4435 avdd.n2152 avdd.n2151 1.7055
R4436 avdd.n2179 avdd.n2178 1.7055
R4437 avdd.n2213 avdd.n2209 1.7055
R4438 avdd.n2229 avdd.n2121 1.7055
R4439 avdd.n2231 avdd.n2230 1.7055
R4440 avdd.n2115 avdd.n2114 1.7055
R4441 avdd.n2250 avdd.n2249 1.7055
R4442 avdd.n2255 avdd.n2254 1.7055
R4443 avdd.n2274 avdd.n2273 1.7055
R4444 avdd.n2367 avdd.n2366 1.7055
R4445 avdd.n2394 avdd.n2393 1.7055
R4446 avdd.n2428 avdd.n2424 1.7055
R4447 avdd.n2444 avdd.n2336 1.7055
R4448 avdd.n2446 avdd.n2445 1.7055
R4449 avdd.n2330 avdd.n2329 1.7055
R4450 avdd.n2465 avdd.n2464 1.7055
R4451 avdd.n2470 avdd.n2469 1.7055
R4452 avdd.n2489 avdd.n2488 1.7055
R4453 avdd.n2582 avdd.n2581 1.7055
R4454 avdd.n2609 avdd.n2608 1.7055
R4455 avdd.n2643 avdd.n2639 1.7055
R4456 avdd.n2659 avdd.n2551 1.7055
R4457 avdd.n2661 avdd.n2660 1.7055
R4458 avdd.n2545 avdd.n2544 1.7055
R4459 avdd.n2680 avdd.n2679 1.7055
R4460 avdd.n2685 avdd.n2684 1.7055
R4461 avdd.n2704 avdd.n2703 1.7055
R4462 avdd.n2797 avdd.n2796 1.7055
R4463 avdd.n2824 avdd.n2823 1.7055
R4464 avdd.n2858 avdd.n2854 1.7055
R4465 avdd.n2874 avdd.n2766 1.7055
R4466 avdd.n2876 avdd.n2875 1.7055
R4467 avdd.n2760 avdd.n2759 1.7055
R4468 avdd.n2895 avdd.n2894 1.7055
R4469 avdd.n2900 avdd.n2899 1.7055
R4470 avdd.n2919 avdd.n2918 1.7055
R4471 avdd.n3012 avdd.n3011 1.7055
R4472 avdd.n3039 avdd.n3038 1.7055
R4473 avdd.n3073 avdd.n3069 1.7055
R4474 avdd.n3089 avdd.n2981 1.7055
R4475 avdd.n3091 avdd.n3090 1.7055
R4476 avdd.n2975 avdd.n2974 1.7055
R4477 avdd.n3110 avdd.n3109 1.7055
R4478 avdd.n3115 avdd.n3114 1.7055
R4479 avdd.n3134 avdd.n3133 1.7055
R4480 avdd.n3188 avdd.n3187 1.7055
R4481 avdd.n3215 avdd.n3214 1.7055
R4482 avdd.n3245 avdd.n3244 1.7055
R4483 avdd.n3358 avdd.n3357 1.7055
R4484 avdd.n3356 avdd.n3247 1.7055
R4485 avdd.n3346 avdd.n3261 1.7055
R4486 avdd.n3345 avdd.n3344 1.7055
R4487 avdd.n3280 avdd.n3271 1.7055
R4488 avdd.n3303 avdd.n3295 1.7055
R4489 avdd.n3403 avdd.n3402 1.7055
R4490 avdd.n3430 avdd.n3429 1.7055
R4491 avdd.n3460 avdd.n3459 1.7055
R4492 avdd.n3573 avdd.n3572 1.7055
R4493 avdd.n3571 avdd.n3462 1.7055
R4494 avdd.n3561 avdd.n3476 1.7055
R4495 avdd.n3560 avdd.n3559 1.7055
R4496 avdd.n3495 avdd.n3486 1.7055
R4497 avdd.n3518 avdd.n3510 1.7055
R4498 avdd.n3618 avdd.n3617 1.7055
R4499 avdd.n3645 avdd.n3644 1.7055
R4500 avdd.n3675 avdd.n3674 1.7055
R4501 avdd.n3788 avdd.n3787 1.7055
R4502 avdd.n3786 avdd.n3677 1.7055
R4503 avdd.n3776 avdd.n3691 1.7055
R4504 avdd.n3775 avdd.n3774 1.7055
R4505 avdd.n3710 avdd.n3701 1.7055
R4506 avdd.n3733 avdd.n3725 1.7055
R4507 avdd.n3833 avdd.n3832 1.7055
R4508 avdd.n3860 avdd.n3859 1.7055
R4509 avdd.n3890 avdd.n3889 1.7055
R4510 avdd.n4003 avdd.n4002 1.7055
R4511 avdd.n4001 avdd.n3892 1.7055
R4512 avdd.n3991 avdd.n3906 1.7055
R4513 avdd.n3990 avdd.n3989 1.7055
R4514 avdd.n3925 avdd.n3916 1.7055
R4515 avdd.n3948 avdd.n3940 1.7055
R4516 avdd.n4048 avdd.n4047 1.7055
R4517 avdd.n4075 avdd.n4074 1.7055
R4518 avdd.n4105 avdd.n4104 1.7055
R4519 avdd.n4218 avdd.n4217 1.7055
R4520 avdd.n4216 avdd.n4107 1.7055
R4521 avdd.n4206 avdd.n4121 1.7055
R4522 avdd.n4205 avdd.n4204 1.7055
R4523 avdd.n4140 avdd.n4131 1.7055
R4524 avdd.n4163 avdd.n4155 1.7055
R4525 avdd.n4263 avdd.n4262 1.7055
R4526 avdd.n4290 avdd.n4289 1.7055
R4527 avdd.n4320 avdd.n4319 1.7055
R4528 avdd.n4433 avdd.n4432 1.7055
R4529 avdd.n4431 avdd.n4322 1.7055
R4530 avdd.n4421 avdd.n4336 1.7055
R4531 avdd.n4420 avdd.n4419 1.7055
R4532 avdd.n4355 avdd.n4346 1.7055
R4533 avdd.n4378 avdd.n4370 1.7055
R4534 avdd.n4874 avdd.n4873 1.7055
R4535 avdd.n4901 avdd.n4900 1.7055
R4536 avdd.n4935 avdd.n4931 1.7055
R4537 avdd.n4951 avdd.n4843 1.7055
R4538 avdd.n4953 avdd.n4952 1.7055
R4539 avdd.n4837 avdd.n4836 1.7055
R4540 avdd.n4972 avdd.n4971 1.7055
R4541 avdd.n4977 avdd.n4976 1.7055
R4542 avdd.n4827 avdd.n4813 1.7055
R4543 avdd.n5090 avdd.n5089 1.7055
R4544 avdd.n5117 avdd.n5116 1.7055
R4545 avdd.n5151 avdd.n5147 1.7055
R4546 avdd.n5167 avdd.n5059 1.7055
R4547 avdd.n5169 avdd.n5168 1.7055
R4548 avdd.n5053 avdd.n5052 1.7055
R4549 avdd.n5188 avdd.n5187 1.7055
R4550 avdd.n5193 avdd.n5192 1.7055
R4551 avdd.n5043 avdd.n5029 1.7055
R4552 avdd.n5306 avdd.n5305 1.7055
R4553 avdd.n5333 avdd.n5332 1.7055
R4554 avdd.n5367 avdd.n5363 1.7055
R4555 avdd.n5383 avdd.n5275 1.7055
R4556 avdd.n5385 avdd.n5384 1.7055
R4557 avdd.n5269 avdd.n5268 1.7055
R4558 avdd.n5404 avdd.n5403 1.7055
R4559 avdd.n5409 avdd.n5408 1.7055
R4560 avdd.n5259 avdd.n5245 1.7055
R4561 avdd.n5522 avdd.n5521 1.7055
R4562 avdd.n5549 avdd.n5548 1.7055
R4563 avdd.n5583 avdd.n5579 1.7055
R4564 avdd.n5599 avdd.n5491 1.7055
R4565 avdd.n5601 avdd.n5600 1.7055
R4566 avdd.n5485 avdd.n5484 1.7055
R4567 avdd.n5620 avdd.n5619 1.7055
R4568 avdd.n5625 avdd.n5624 1.7055
R4569 avdd.n5475 avdd.n5461 1.7055
R4570 avdd.n5738 avdd.n5737 1.7055
R4571 avdd.n5765 avdd.n5764 1.7055
R4572 avdd.n5799 avdd.n5795 1.7055
R4573 avdd.n5815 avdd.n5707 1.7055
R4574 avdd.n5817 avdd.n5816 1.7055
R4575 avdd.n5701 avdd.n5700 1.7055
R4576 avdd.n5836 avdd.n5835 1.7055
R4577 avdd.n5841 avdd.n5840 1.7055
R4578 avdd.n5691 avdd.n5677 1.7055
R4579 avdd.n5954 avdd.n5953 1.7055
R4580 avdd.n5981 avdd.n5980 1.7055
R4581 avdd.n6015 avdd.n6011 1.7055
R4582 avdd.n6031 avdd.n5923 1.7055
R4583 avdd.n6033 avdd.n6032 1.7055
R4584 avdd.n5917 avdd.n5916 1.7055
R4585 avdd.n6052 avdd.n6051 1.7055
R4586 avdd.n6057 avdd.n6056 1.7055
R4587 avdd.n5907 avdd.n5893 1.7055
R4588 avdd.n6170 avdd.n6169 1.7055
R4589 avdd.n6197 avdd.n6196 1.7055
R4590 avdd.n6231 avdd.n6227 1.7055
R4591 avdd.n6247 avdd.n6139 1.7055
R4592 avdd.n6249 avdd.n6248 1.7055
R4593 avdd.n6133 avdd.n6132 1.7055
R4594 avdd.n6268 avdd.n6267 1.7055
R4595 avdd.n6273 avdd.n6272 1.7055
R4596 avdd.n6123 avdd.n6109 1.7055
R4597 avdd.n6386 avdd.n6385 1.7055
R4598 avdd.n6413 avdd.n6412 1.7055
R4599 avdd.n6447 avdd.n6443 1.7055
R4600 avdd.n6463 avdd.n6355 1.7055
R4601 avdd.n6465 avdd.n6464 1.7055
R4602 avdd.n6349 avdd.n6348 1.7055
R4603 avdd.n6484 avdd.n6483 1.7055
R4604 avdd.n6489 avdd.n6488 1.7055
R4605 avdd.n6339 avdd.n6325 1.7055
R4606 avdd.n6602 avdd.n6601 1.7055
R4607 avdd.n6629 avdd.n6628 1.7055
R4608 avdd.n6663 avdd.n6659 1.7055
R4609 avdd.n6679 avdd.n6571 1.7055
R4610 avdd.n6681 avdd.n6680 1.7055
R4611 avdd.n6565 avdd.n6564 1.7055
R4612 avdd.n6700 avdd.n6699 1.7055
R4613 avdd.n6705 avdd.n6704 1.7055
R4614 avdd.n6555 avdd.n6541 1.7055
R4615 avdd.n6818 avdd.n6817 1.7055
R4616 avdd.n6845 avdd.n6844 1.7055
R4617 avdd.n6879 avdd.n6875 1.7055
R4618 avdd.n6895 avdd.n6787 1.7055
R4619 avdd.n6897 avdd.n6896 1.7055
R4620 avdd.n6781 avdd.n6780 1.7055
R4621 avdd.n6916 avdd.n6915 1.7055
R4622 avdd.n6921 avdd.n6920 1.7055
R4623 avdd.n6771 avdd.n6757 1.7055
R4624 avdd.n7034 avdd.n7033 1.7055
R4625 avdd.n7061 avdd.n7060 1.7055
R4626 avdd.n7095 avdd.n7091 1.7055
R4627 avdd.n7111 avdd.n7003 1.7055
R4628 avdd.n7113 avdd.n7112 1.7055
R4629 avdd.n6997 avdd.n6996 1.7055
R4630 avdd.n7132 avdd.n7131 1.7055
R4631 avdd.n7137 avdd.n7136 1.7055
R4632 avdd.n6987 avdd.n6973 1.7055
R4633 avdd.n7250 avdd.n7249 1.7055
R4634 avdd.n7277 avdd.n7276 1.7055
R4635 avdd.n7311 avdd.n7307 1.7055
R4636 avdd.n7327 avdd.n7219 1.7055
R4637 avdd.n7329 avdd.n7328 1.7055
R4638 avdd.n7213 avdd.n7212 1.7055
R4639 avdd.n7348 avdd.n7347 1.7055
R4640 avdd.n7353 avdd.n7352 1.7055
R4641 avdd.n7203 avdd.n7189 1.7055
R4642 avdd.n2029 avdd.n2005 1.70483
R4643 avdd.n2304 avdd.n2303 1.70483
R4644 avdd.n2519 avdd.n2518 1.70483
R4645 avdd.n2734 avdd.n2733 1.70483
R4646 avdd.n2949 avdd.n2948 1.70483
R4647 avdd.n3164 avdd.n3163 1.70483
R4648 avdd.n3380 avdd.n3379 1.70483
R4649 avdd.n3595 avdd.n3594 1.70483
R4650 avdd.n3810 avdd.n3809 1.70483
R4651 avdd.n4025 avdd.n4024 1.70483
R4652 avdd.n4240 avdd.n4239 1.70483
R4653 avdd.n4455 avdd.n4454 1.70483
R4654 avdd.n5022 avdd.n4812 1.70483
R4655 avdd.n5238 avdd.n5028 1.70483
R4656 avdd.n5454 avdd.n5244 1.70483
R4657 avdd.n5670 avdd.n5460 1.70483
R4658 avdd.n5886 avdd.n5676 1.70483
R4659 avdd.n6102 avdd.n5892 1.70483
R4660 avdd.n6318 avdd.n6108 1.70483
R4661 avdd.n6534 avdd.n6324 1.70483
R4662 avdd.n6750 avdd.n6540 1.70483
R4663 avdd.n6966 avdd.n6756 1.70483
R4664 avdd.n7182 avdd.n6972 1.70483
R4665 avdd.n7398 avdd.n7188 1.70483
R4666 avdd.n3325 avdd.n3298 1.7044
R4667 avdd.n3540 avdd.n3513 1.7044
R4668 avdd.n3755 avdd.n3728 1.7044
R4669 avdd.n3970 avdd.n3943 1.7044
R4670 avdd.n4185 avdd.n4158 1.7044
R4671 avdd.n4400 avdd.n4373 1.7044
R4672 avdd.n5021 avdd.n4818 1.7044
R4673 avdd.n5237 avdd.n5034 1.7044
R4674 avdd.n5453 avdd.n5250 1.7044
R4675 avdd.n5669 avdd.n5466 1.7044
R4676 avdd.n5885 avdd.n5682 1.7044
R4677 avdd.n6101 avdd.n5898 1.7044
R4678 avdd.n6317 avdd.n6114 1.7044
R4679 avdd.n6533 avdd.n6330 1.7044
R4680 avdd.n6749 avdd.n6546 1.7044
R4681 avdd.n6965 avdd.n6762 1.7044
R4682 avdd.n7181 avdd.n6978 1.7044
R4683 avdd.n7397 avdd.n7194 1.7044
R4684 avdd.n2036 avdd.n2006 1.70333
R4685 avdd.n2272 avdd.n2093 1.70333
R4686 avdd.n2487 avdd.n2308 1.70333
R4687 avdd.n2702 avdd.n2523 1.70333
R4688 avdd.n2917 avdd.n2738 1.70333
R4689 avdd.n3132 avdd.n2953 1.70333
R4690 avdd.n3325 avdd.n3304 1.70333
R4691 avdd.n3540 avdd.n3519 1.70333
R4692 avdd.n3755 avdd.n3734 1.70333
R4693 avdd.n3970 avdd.n3949 1.70333
R4694 avdd.n4185 avdd.n4164 1.70333
R4695 avdd.n4400 avdd.n4379 1.70333
R4696 avdd.n1934 avdd.n1878 1.70156
R4697 avdd.n2195 avdd.n2194 1.70156
R4698 avdd.n2410 avdd.n2409 1.70156
R4699 avdd.n2625 avdd.n2624 1.70156
R4700 avdd.n2840 avdd.n2839 1.70156
R4701 avdd.n3055 avdd.n3054 1.70156
R4702 avdd.n3224 avdd.n3169 1.70156
R4703 avdd.n3439 avdd.n3384 1.70156
R4704 avdd.n3654 avdd.n3599 1.70156
R4705 avdd.n3869 avdd.n3814 1.70156
R4706 avdd.n4084 avdd.n4029 1.70156
R4707 avdd.n4299 avdd.n4244 1.70156
R4708 avdd.n2036 avdd.n2007 1.70121
R4709 avdd.n2290 avdd.n2093 1.70121
R4710 avdd.n2505 avdd.n2308 1.70121
R4711 avdd.n2720 avdd.n2523 1.70121
R4712 avdd.n2935 avdd.n2738 1.70121
R4713 avdd.n3150 avdd.n2953 1.70121
R4714 avdd.n5021 avdd.n4814 1.70121
R4715 avdd.n5237 avdd.n5030 1.70121
R4716 avdd.n5453 avdd.n5246 1.70121
R4717 avdd.n5669 avdd.n5462 1.70121
R4718 avdd.n5885 avdd.n5678 1.70121
R4719 avdd.n6101 avdd.n5894 1.70121
R4720 avdd.n6317 avdd.n6110 1.70121
R4721 avdd.n6533 avdd.n6326 1.70121
R4722 avdd.n6749 avdd.n6542 1.70121
R4723 avdd.n6965 avdd.n6758 1.70121
R4724 avdd.n7181 avdd.n6974 1.70121
R4725 avdd.n7397 avdd.n7190 1.70121
R4726 avdd.n7450 avdd.n7445 1.67304
R4727 avdd.n7489 avdd.n7484 1.67304
R4728 avdd.n7549 avdd.n7544 1.67304
R4729 avdd.n7589 avdd.n7584 1.67304
R4730 avdd.n1814 avdd.n1809 1.59114
R4731 avdd.n1640 avdd.n1635 1.59114
R4732 avdd.n1724 avdd.n1719 1.59114
R4733 avdd.n1676 avdd.n1671 1.59114
R4734 avdd.n4595 avdd.n4592 1.50638
R4735 avdd.n4527 avdd.n4526 1.41
R4736 avdd.n2086 avdd.n1882 1.13717
R4737 avdd.n1920 avdd.n1919 1.13717
R4738 avdd.n1940 avdd.n1890 1.13717
R4739 avdd.n2082 avdd.n1885 1.13717
R4740 avdd.n1964 avdd.n1963 1.13717
R4741 avdd.n1982 avdd.n1975 1.13717
R4742 avdd.n1999 avdd.n1995 1.13717
R4743 avdd.n2013 avdd.n2003 1.13717
R4744 avdd.n2025 avdd.n2024 1.13717
R4745 avdd.n1907 avdd.n1906 1.13717
R4746 avdd.n1929 avdd.n1928 1.13717
R4747 avdd.n1951 avdd.n1888 1.13717
R4748 avdd.n2072 avdd.n2071 1.13717
R4749 avdd.n1961 avdd.n1960 1.13717
R4750 avdd.n1987 avdd.n1986 1.13717
R4751 avdd.n1993 avdd.n1979 1.13717
R4752 avdd.n2032 avdd.n1994 1.13717
R4753 avdd.n2140 avdd.n2133 1.13717
R4754 avdd.n2174 avdd.n2173 1.13717
R4755 avdd.n2188 avdd.n2187 1.13717
R4756 avdd.n2205 avdd.n2135 1.13717
R4757 avdd.n2225 avdd.n2124 1.13717
R4758 avdd.n2245 avdd.n2244 1.13717
R4759 avdd.n2264 avdd.n2263 1.13717
R4760 avdd.n2286 avdd.n2102 1.13717
R4761 avdd.n2299 avdd.n2098 1.13717
R4762 avdd.n2161 avdd.n2160 1.13717
R4763 avdd.n2182 avdd.n2181 1.13717
R4764 avdd.n2216 avdd.n2132 1.13717
R4765 avdd.n2123 avdd.n2122 1.13717
R4766 avdd.n2237 avdd.n2119 1.13717
R4767 avdd.n2258 avdd.n2257 1.13717
R4768 avdd.n2108 avdd.n2107 1.13717
R4769 avdd.n2277 avdd.n2276 1.13717
R4770 avdd.n2355 avdd.n2348 1.13717
R4771 avdd.n2389 avdd.n2388 1.13717
R4772 avdd.n2403 avdd.n2402 1.13717
R4773 avdd.n2420 avdd.n2350 1.13717
R4774 avdd.n2440 avdd.n2339 1.13717
R4775 avdd.n2460 avdd.n2459 1.13717
R4776 avdd.n2479 avdd.n2478 1.13717
R4777 avdd.n2501 avdd.n2317 1.13717
R4778 avdd.n2514 avdd.n2313 1.13717
R4779 avdd.n2376 avdd.n2375 1.13717
R4780 avdd.n2397 avdd.n2396 1.13717
R4781 avdd.n2431 avdd.n2347 1.13717
R4782 avdd.n2338 avdd.n2337 1.13717
R4783 avdd.n2452 avdd.n2334 1.13717
R4784 avdd.n2473 avdd.n2472 1.13717
R4785 avdd.n2323 avdd.n2322 1.13717
R4786 avdd.n2492 avdd.n2491 1.13717
R4787 avdd.n2570 avdd.n2563 1.13717
R4788 avdd.n2604 avdd.n2603 1.13717
R4789 avdd.n2618 avdd.n2617 1.13717
R4790 avdd.n2635 avdd.n2565 1.13717
R4791 avdd.n2655 avdd.n2554 1.13717
R4792 avdd.n2675 avdd.n2674 1.13717
R4793 avdd.n2694 avdd.n2693 1.13717
R4794 avdd.n2716 avdd.n2532 1.13717
R4795 avdd.n2729 avdd.n2528 1.13717
R4796 avdd.n2591 avdd.n2590 1.13717
R4797 avdd.n2612 avdd.n2611 1.13717
R4798 avdd.n2646 avdd.n2562 1.13717
R4799 avdd.n2553 avdd.n2552 1.13717
R4800 avdd.n2667 avdd.n2549 1.13717
R4801 avdd.n2688 avdd.n2687 1.13717
R4802 avdd.n2538 avdd.n2537 1.13717
R4803 avdd.n2707 avdd.n2706 1.13717
R4804 avdd.n2785 avdd.n2778 1.13717
R4805 avdd.n2819 avdd.n2818 1.13717
R4806 avdd.n2833 avdd.n2832 1.13717
R4807 avdd.n2850 avdd.n2780 1.13717
R4808 avdd.n2870 avdd.n2769 1.13717
R4809 avdd.n2890 avdd.n2889 1.13717
R4810 avdd.n2909 avdd.n2908 1.13717
R4811 avdd.n2931 avdd.n2747 1.13717
R4812 avdd.n2944 avdd.n2743 1.13717
R4813 avdd.n2806 avdd.n2805 1.13717
R4814 avdd.n2827 avdd.n2826 1.13717
R4815 avdd.n2861 avdd.n2777 1.13717
R4816 avdd.n2768 avdd.n2767 1.13717
R4817 avdd.n2882 avdd.n2764 1.13717
R4818 avdd.n2903 avdd.n2902 1.13717
R4819 avdd.n2753 avdd.n2752 1.13717
R4820 avdd.n2922 avdd.n2921 1.13717
R4821 avdd.n3000 avdd.n2993 1.13717
R4822 avdd.n3034 avdd.n3033 1.13717
R4823 avdd.n3048 avdd.n3047 1.13717
R4824 avdd.n3065 avdd.n2995 1.13717
R4825 avdd.n3085 avdd.n2984 1.13717
R4826 avdd.n3105 avdd.n3104 1.13717
R4827 avdd.n3124 avdd.n3123 1.13717
R4828 avdd.n3146 avdd.n2962 1.13717
R4829 avdd.n3159 avdd.n2958 1.13717
R4830 avdd.n3021 avdd.n3020 1.13717
R4831 avdd.n3042 avdd.n3041 1.13717
R4832 avdd.n3076 avdd.n2992 1.13717
R4833 avdd.n2983 avdd.n2982 1.13717
R4834 avdd.n3097 avdd.n2979 1.13717
R4835 avdd.n3118 avdd.n3117 1.13717
R4836 avdd.n2968 avdd.n2967 1.13717
R4837 avdd.n3137 avdd.n3136 1.13717
R4838 avdd.n3210 avdd.n3209 1.13717
R4839 avdd.n3230 avdd.n3180 1.13717
R4840 avdd.n3371 avdd.n3175 1.13717
R4841 avdd.n3254 avdd.n3253 1.13717
R4842 avdd.n3272 avdd.n3265 1.13717
R4843 avdd.n3289 avdd.n3285 1.13717
R4844 avdd.n3306 avdd.n3293 1.13717
R4845 avdd.n3318 avdd.n3314 1.13717
R4846 avdd.n3197 avdd.n3196 1.13717
R4847 avdd.n3219 avdd.n3218 1.13717
R4848 avdd.n3375 avdd.n3172 1.13717
R4849 avdd.n3241 avdd.n3178 1.13717
R4850 avdd.n3361 avdd.n3360 1.13717
R4851 avdd.n3251 avdd.n3250 1.13717
R4852 avdd.n3277 avdd.n3276 1.13717
R4853 avdd.n3283 avdd.n3269 1.13717
R4854 avdd.n3300 avdd.n3284 1.13717
R4855 avdd.n3425 avdd.n3424 1.13717
R4856 avdd.n3445 avdd.n3395 1.13717
R4857 avdd.n3586 avdd.n3390 1.13717
R4858 avdd.n3469 avdd.n3468 1.13717
R4859 avdd.n3487 avdd.n3480 1.13717
R4860 avdd.n3504 avdd.n3500 1.13717
R4861 avdd.n3521 avdd.n3508 1.13717
R4862 avdd.n3533 avdd.n3529 1.13717
R4863 avdd.n3412 avdd.n3411 1.13717
R4864 avdd.n3434 avdd.n3433 1.13717
R4865 avdd.n3590 avdd.n3387 1.13717
R4866 avdd.n3456 avdd.n3393 1.13717
R4867 avdd.n3576 avdd.n3575 1.13717
R4868 avdd.n3466 avdd.n3465 1.13717
R4869 avdd.n3492 avdd.n3491 1.13717
R4870 avdd.n3498 avdd.n3484 1.13717
R4871 avdd.n3515 avdd.n3499 1.13717
R4872 avdd.n3640 avdd.n3639 1.13717
R4873 avdd.n3660 avdd.n3610 1.13717
R4874 avdd.n3801 avdd.n3605 1.13717
R4875 avdd.n3684 avdd.n3683 1.13717
R4876 avdd.n3702 avdd.n3695 1.13717
R4877 avdd.n3719 avdd.n3715 1.13717
R4878 avdd.n3736 avdd.n3723 1.13717
R4879 avdd.n3748 avdd.n3744 1.13717
R4880 avdd.n3627 avdd.n3626 1.13717
R4881 avdd.n3649 avdd.n3648 1.13717
R4882 avdd.n3805 avdd.n3602 1.13717
R4883 avdd.n3671 avdd.n3608 1.13717
R4884 avdd.n3791 avdd.n3790 1.13717
R4885 avdd.n3681 avdd.n3680 1.13717
R4886 avdd.n3707 avdd.n3706 1.13717
R4887 avdd.n3713 avdd.n3699 1.13717
R4888 avdd.n3730 avdd.n3714 1.13717
R4889 avdd.n3855 avdd.n3854 1.13717
R4890 avdd.n3875 avdd.n3825 1.13717
R4891 avdd.n4016 avdd.n3820 1.13717
R4892 avdd.n3899 avdd.n3898 1.13717
R4893 avdd.n3917 avdd.n3910 1.13717
R4894 avdd.n3934 avdd.n3930 1.13717
R4895 avdd.n3951 avdd.n3938 1.13717
R4896 avdd.n3963 avdd.n3959 1.13717
R4897 avdd.n3842 avdd.n3841 1.13717
R4898 avdd.n3864 avdd.n3863 1.13717
R4899 avdd.n4020 avdd.n3817 1.13717
R4900 avdd.n3886 avdd.n3823 1.13717
R4901 avdd.n4006 avdd.n4005 1.13717
R4902 avdd.n3896 avdd.n3895 1.13717
R4903 avdd.n3922 avdd.n3921 1.13717
R4904 avdd.n3928 avdd.n3914 1.13717
R4905 avdd.n3945 avdd.n3929 1.13717
R4906 avdd.n4070 avdd.n4069 1.13717
R4907 avdd.n4090 avdd.n4040 1.13717
R4908 avdd.n4231 avdd.n4035 1.13717
R4909 avdd.n4114 avdd.n4113 1.13717
R4910 avdd.n4132 avdd.n4125 1.13717
R4911 avdd.n4149 avdd.n4145 1.13717
R4912 avdd.n4166 avdd.n4153 1.13717
R4913 avdd.n4178 avdd.n4174 1.13717
R4914 avdd.n4057 avdd.n4056 1.13717
R4915 avdd.n4079 avdd.n4078 1.13717
R4916 avdd.n4235 avdd.n4032 1.13717
R4917 avdd.n4101 avdd.n4038 1.13717
R4918 avdd.n4221 avdd.n4220 1.13717
R4919 avdd.n4111 avdd.n4110 1.13717
R4920 avdd.n4137 avdd.n4136 1.13717
R4921 avdd.n4143 avdd.n4129 1.13717
R4922 avdd.n4160 avdd.n4144 1.13717
R4923 avdd.n4285 avdd.n4284 1.13717
R4924 avdd.n4305 avdd.n4255 1.13717
R4925 avdd.n4446 avdd.n4250 1.13717
R4926 avdd.n4329 avdd.n4328 1.13717
R4927 avdd.n4347 avdd.n4340 1.13717
R4928 avdd.n4364 avdd.n4360 1.13717
R4929 avdd.n4381 avdd.n4368 1.13717
R4930 avdd.n4393 avdd.n4389 1.13717
R4931 avdd.n4272 avdd.n4271 1.13717
R4932 avdd.n4294 avdd.n4293 1.13717
R4933 avdd.n4450 avdd.n4247 1.13717
R4934 avdd.n4316 avdd.n4253 1.13717
R4935 avdd.n4436 avdd.n4435 1.13717
R4936 avdd.n4326 avdd.n4325 1.13717
R4937 avdd.n4352 avdd.n4351 1.13717
R4938 avdd.n4358 avdd.n4344 1.13717
R4939 avdd.n4375 avdd.n4359 1.13717
R4940 avdd.n4883 avdd.n4882 1.13717
R4941 avdd.n4896 avdd.n4895 1.13717
R4942 avdd.n4905 avdd.n4904 1.13717
R4943 avdd.n4911 avdd.n4910 1.13717
R4944 avdd.n4927 avdd.n4857 1.13717
R4945 avdd.n4938 avdd.n4854 1.13717
R4946 avdd.n4863 avdd.n4855 1.13717
R4947 avdd.n4947 avdd.n4846 1.13717
R4948 avdd.n4845 avdd.n4844 1.13717
R4949 avdd.n4959 avdd.n4841 1.13717
R4950 avdd.n4967 avdd.n4966 1.13717
R4951 avdd.n4980 avdd.n4979 1.13717
R4952 avdd.n4986 avdd.n4985 1.13717
R4953 avdd.n4996 avdd.n4995 1.13717
R4954 avdd.n4830 avdd.n4829 1.13717
R4955 avdd.n5004 avdd.n4823 1.13717
R4956 avdd.n5017 avdd.n5016 1.13717
R4957 avdd.n5099 avdd.n5098 1.13717
R4958 avdd.n5112 avdd.n5111 1.13717
R4959 avdd.n5121 avdd.n5120 1.13717
R4960 avdd.n5127 avdd.n5126 1.13717
R4961 avdd.n5143 avdd.n5073 1.13717
R4962 avdd.n5154 avdd.n5070 1.13717
R4963 avdd.n5079 avdd.n5071 1.13717
R4964 avdd.n5163 avdd.n5062 1.13717
R4965 avdd.n5061 avdd.n5060 1.13717
R4966 avdd.n5175 avdd.n5057 1.13717
R4967 avdd.n5183 avdd.n5182 1.13717
R4968 avdd.n5196 avdd.n5195 1.13717
R4969 avdd.n5202 avdd.n5201 1.13717
R4970 avdd.n5212 avdd.n5211 1.13717
R4971 avdd.n5046 avdd.n5045 1.13717
R4972 avdd.n5220 avdd.n5039 1.13717
R4973 avdd.n5233 avdd.n5232 1.13717
R4974 avdd.n5315 avdd.n5314 1.13717
R4975 avdd.n5328 avdd.n5327 1.13717
R4976 avdd.n5337 avdd.n5336 1.13717
R4977 avdd.n5343 avdd.n5342 1.13717
R4978 avdd.n5359 avdd.n5289 1.13717
R4979 avdd.n5370 avdd.n5286 1.13717
R4980 avdd.n5295 avdd.n5287 1.13717
R4981 avdd.n5379 avdd.n5278 1.13717
R4982 avdd.n5277 avdd.n5276 1.13717
R4983 avdd.n5391 avdd.n5273 1.13717
R4984 avdd.n5399 avdd.n5398 1.13717
R4985 avdd.n5412 avdd.n5411 1.13717
R4986 avdd.n5418 avdd.n5417 1.13717
R4987 avdd.n5428 avdd.n5427 1.13717
R4988 avdd.n5262 avdd.n5261 1.13717
R4989 avdd.n5436 avdd.n5255 1.13717
R4990 avdd.n5449 avdd.n5448 1.13717
R4991 avdd.n5531 avdd.n5530 1.13717
R4992 avdd.n5544 avdd.n5543 1.13717
R4993 avdd.n5553 avdd.n5552 1.13717
R4994 avdd.n5559 avdd.n5558 1.13717
R4995 avdd.n5575 avdd.n5505 1.13717
R4996 avdd.n5586 avdd.n5502 1.13717
R4997 avdd.n5511 avdd.n5503 1.13717
R4998 avdd.n5595 avdd.n5494 1.13717
R4999 avdd.n5493 avdd.n5492 1.13717
R5000 avdd.n5607 avdd.n5489 1.13717
R5001 avdd.n5615 avdd.n5614 1.13717
R5002 avdd.n5628 avdd.n5627 1.13717
R5003 avdd.n5634 avdd.n5633 1.13717
R5004 avdd.n5644 avdd.n5643 1.13717
R5005 avdd.n5478 avdd.n5477 1.13717
R5006 avdd.n5652 avdd.n5471 1.13717
R5007 avdd.n5665 avdd.n5664 1.13717
R5008 avdd.n5747 avdd.n5746 1.13717
R5009 avdd.n5760 avdd.n5759 1.13717
R5010 avdd.n5769 avdd.n5768 1.13717
R5011 avdd.n5775 avdd.n5774 1.13717
R5012 avdd.n5791 avdd.n5721 1.13717
R5013 avdd.n5802 avdd.n5718 1.13717
R5014 avdd.n5727 avdd.n5719 1.13717
R5015 avdd.n5811 avdd.n5710 1.13717
R5016 avdd.n5709 avdd.n5708 1.13717
R5017 avdd.n5823 avdd.n5705 1.13717
R5018 avdd.n5831 avdd.n5830 1.13717
R5019 avdd.n5844 avdd.n5843 1.13717
R5020 avdd.n5850 avdd.n5849 1.13717
R5021 avdd.n5860 avdd.n5859 1.13717
R5022 avdd.n5694 avdd.n5693 1.13717
R5023 avdd.n5868 avdd.n5687 1.13717
R5024 avdd.n5881 avdd.n5880 1.13717
R5025 avdd.n5963 avdd.n5962 1.13717
R5026 avdd.n5976 avdd.n5975 1.13717
R5027 avdd.n5985 avdd.n5984 1.13717
R5028 avdd.n5991 avdd.n5990 1.13717
R5029 avdd.n6007 avdd.n5937 1.13717
R5030 avdd.n6018 avdd.n5934 1.13717
R5031 avdd.n5943 avdd.n5935 1.13717
R5032 avdd.n6027 avdd.n5926 1.13717
R5033 avdd.n5925 avdd.n5924 1.13717
R5034 avdd.n6039 avdd.n5921 1.13717
R5035 avdd.n6047 avdd.n6046 1.13717
R5036 avdd.n6060 avdd.n6059 1.13717
R5037 avdd.n6066 avdd.n6065 1.13717
R5038 avdd.n6076 avdd.n6075 1.13717
R5039 avdd.n5910 avdd.n5909 1.13717
R5040 avdd.n6084 avdd.n5903 1.13717
R5041 avdd.n6097 avdd.n6096 1.13717
R5042 avdd.n6179 avdd.n6178 1.13717
R5043 avdd.n6192 avdd.n6191 1.13717
R5044 avdd.n6201 avdd.n6200 1.13717
R5045 avdd.n6207 avdd.n6206 1.13717
R5046 avdd.n6223 avdd.n6153 1.13717
R5047 avdd.n6234 avdd.n6150 1.13717
R5048 avdd.n6159 avdd.n6151 1.13717
R5049 avdd.n6243 avdd.n6142 1.13717
R5050 avdd.n6141 avdd.n6140 1.13717
R5051 avdd.n6255 avdd.n6137 1.13717
R5052 avdd.n6263 avdd.n6262 1.13717
R5053 avdd.n6276 avdd.n6275 1.13717
R5054 avdd.n6282 avdd.n6281 1.13717
R5055 avdd.n6292 avdd.n6291 1.13717
R5056 avdd.n6126 avdd.n6125 1.13717
R5057 avdd.n6300 avdd.n6119 1.13717
R5058 avdd.n6313 avdd.n6312 1.13717
R5059 avdd.n6395 avdd.n6394 1.13717
R5060 avdd.n6408 avdd.n6407 1.13717
R5061 avdd.n6417 avdd.n6416 1.13717
R5062 avdd.n6423 avdd.n6422 1.13717
R5063 avdd.n6439 avdd.n6369 1.13717
R5064 avdd.n6450 avdd.n6366 1.13717
R5065 avdd.n6375 avdd.n6367 1.13717
R5066 avdd.n6459 avdd.n6358 1.13717
R5067 avdd.n6357 avdd.n6356 1.13717
R5068 avdd.n6471 avdd.n6353 1.13717
R5069 avdd.n6479 avdd.n6478 1.13717
R5070 avdd.n6492 avdd.n6491 1.13717
R5071 avdd.n6498 avdd.n6497 1.13717
R5072 avdd.n6508 avdd.n6507 1.13717
R5073 avdd.n6342 avdd.n6341 1.13717
R5074 avdd.n6516 avdd.n6335 1.13717
R5075 avdd.n6529 avdd.n6528 1.13717
R5076 avdd.n6611 avdd.n6610 1.13717
R5077 avdd.n6624 avdd.n6623 1.13717
R5078 avdd.n6633 avdd.n6632 1.13717
R5079 avdd.n6639 avdd.n6638 1.13717
R5080 avdd.n6655 avdd.n6585 1.13717
R5081 avdd.n6666 avdd.n6582 1.13717
R5082 avdd.n6591 avdd.n6583 1.13717
R5083 avdd.n6675 avdd.n6574 1.13717
R5084 avdd.n6573 avdd.n6572 1.13717
R5085 avdd.n6687 avdd.n6569 1.13717
R5086 avdd.n6695 avdd.n6694 1.13717
R5087 avdd.n6708 avdd.n6707 1.13717
R5088 avdd.n6714 avdd.n6713 1.13717
R5089 avdd.n6724 avdd.n6723 1.13717
R5090 avdd.n6558 avdd.n6557 1.13717
R5091 avdd.n6732 avdd.n6551 1.13717
R5092 avdd.n6745 avdd.n6744 1.13717
R5093 avdd.n6827 avdd.n6826 1.13717
R5094 avdd.n6840 avdd.n6839 1.13717
R5095 avdd.n6849 avdd.n6848 1.13717
R5096 avdd.n6855 avdd.n6854 1.13717
R5097 avdd.n6871 avdd.n6801 1.13717
R5098 avdd.n6882 avdd.n6798 1.13717
R5099 avdd.n6807 avdd.n6799 1.13717
R5100 avdd.n6891 avdd.n6790 1.13717
R5101 avdd.n6789 avdd.n6788 1.13717
R5102 avdd.n6903 avdd.n6785 1.13717
R5103 avdd.n6911 avdd.n6910 1.13717
R5104 avdd.n6924 avdd.n6923 1.13717
R5105 avdd.n6930 avdd.n6929 1.13717
R5106 avdd.n6940 avdd.n6939 1.13717
R5107 avdd.n6774 avdd.n6773 1.13717
R5108 avdd.n6948 avdd.n6767 1.13717
R5109 avdd.n6961 avdd.n6960 1.13717
R5110 avdd.n7043 avdd.n7042 1.13717
R5111 avdd.n7056 avdd.n7055 1.13717
R5112 avdd.n7065 avdd.n7064 1.13717
R5113 avdd.n7071 avdd.n7070 1.13717
R5114 avdd.n7087 avdd.n7017 1.13717
R5115 avdd.n7098 avdd.n7014 1.13717
R5116 avdd.n7023 avdd.n7015 1.13717
R5117 avdd.n7107 avdd.n7006 1.13717
R5118 avdd.n7005 avdd.n7004 1.13717
R5119 avdd.n7119 avdd.n7001 1.13717
R5120 avdd.n7127 avdd.n7126 1.13717
R5121 avdd.n7140 avdd.n7139 1.13717
R5122 avdd.n7146 avdd.n7145 1.13717
R5123 avdd.n7156 avdd.n7155 1.13717
R5124 avdd.n6990 avdd.n6989 1.13717
R5125 avdd.n7164 avdd.n6983 1.13717
R5126 avdd.n7177 avdd.n7176 1.13717
R5127 avdd.n7259 avdd.n7258 1.13717
R5128 avdd.n7272 avdd.n7271 1.13717
R5129 avdd.n7281 avdd.n7280 1.13717
R5130 avdd.n7287 avdd.n7286 1.13717
R5131 avdd.n7303 avdd.n7233 1.13717
R5132 avdd.n7314 avdd.n7230 1.13717
R5133 avdd.n7239 avdd.n7231 1.13717
R5134 avdd.n7323 avdd.n7222 1.13717
R5135 avdd.n7221 avdd.n7220 1.13717
R5136 avdd.n7335 avdd.n7217 1.13717
R5137 avdd.n7343 avdd.n7342 1.13717
R5138 avdd.n7356 avdd.n7355 1.13717
R5139 avdd.n7362 avdd.n7361 1.13717
R5140 avdd.n7372 avdd.n7371 1.13717
R5141 avdd.n7206 avdd.n7205 1.13717
R5142 avdd.n7380 avdd.n7199 1.13717
R5143 avdd.n7393 avdd.n7392 1.13717
R5144 avdd.n7716 avdd.n7715 1.13717
R5145 avdd.n7735 avdd.n7734 1.13717
R5146 avdd.n7697 avdd.n7696 1.13717
R5147 avdd.n7677 avdd.n7676 1.13717
R5148 avdd.n7805 avdd.n7804 1.13717
R5149 avdd.n7825 avdd.n7824 1.13717
R5150 avdd.n7844 avdd.n7843 1.13717
R5151 avdd.n7790 avdd.n7789 1.13717
R5152 avdd.n10195 avdd.n10194 1.13717
R5153 avdd.n10214 avdd.n10213 1.13717
R5154 avdd.n10176 avdd.n10175 1.13717
R5155 avdd.n10156 avdd.n10155 1.13717
R5156 avdd.n10063 avdd.n10062 1.13717
R5157 avdd.n10083 avdd.n10082 1.13717
R5158 avdd.n10102 avdd.n10101 1.13717
R5159 avdd.n10050 avdd.n10049 1.13717
R5160 avdd.n9999 avdd.n9998 1.13717
R5161 avdd.n10004 avdd.n10003 1.13717
R5162 avdd.n10020 avdd.n10019 1.13717
R5163 avdd.n9960 avdd.n9959 1.13717
R5164 avdd.n9964 avdd.n9963 1.13717
R5165 avdd.n9940 avdd.n9939 1.13717
R5166 avdd.n10295 avdd.n10294 1.13717
R5167 avdd.n10315 avdd.n10314 1.13717
R5168 avdd.n10334 avdd.n10333 1.13717
R5169 avdd.n10266 avdd.n10265 1.13717
R5170 avdd.n9885 avdd.n9884 1.13717
R5171 avdd.n9890 avdd.n9889 1.13717
R5172 avdd.n9906 avdd.n9905 1.13717
R5173 avdd.n9846 avdd.n9845 1.13717
R5174 avdd.n9850 avdd.n9849 1.13717
R5175 avdd.n9826 avdd.n9825 1.13717
R5176 avdd.n10397 avdd.n10396 1.13717
R5177 avdd.n10417 avdd.n10416 1.13717
R5178 avdd.n10436 avdd.n10435 1.13717
R5179 avdd.n10368 avdd.n10367 1.13717
R5180 avdd.n9771 avdd.n9770 1.13717
R5181 avdd.n9776 avdd.n9775 1.13717
R5182 avdd.n9792 avdd.n9791 1.13717
R5183 avdd.n9732 avdd.n9731 1.13717
R5184 avdd.n9736 avdd.n9735 1.13717
R5185 avdd.n9712 avdd.n9711 1.13717
R5186 avdd.n10499 avdd.n10498 1.13717
R5187 avdd.n10519 avdd.n10518 1.13717
R5188 avdd.n10538 avdd.n10537 1.13717
R5189 avdd.n10470 avdd.n10469 1.13717
R5190 avdd.n9658 avdd.n9657 1.13717
R5191 avdd.n9663 avdd.n9662 1.13717
R5192 avdd.n9679 avdd.n9678 1.13717
R5193 avdd.n9619 avdd.n9618 1.13717
R5194 avdd.n9623 avdd.n9622 1.13717
R5195 avdd.n9599 avdd.n9598 1.13717
R5196 avdd.n10601 avdd.n10600 1.13717
R5197 avdd.n10621 avdd.n10620 1.13717
R5198 avdd.n10640 avdd.n10639 1.13717
R5199 avdd.n10572 avdd.n10571 1.13717
R5200 avdd.n9543 avdd.n9542 1.13717
R5201 avdd.n9548 avdd.n9547 1.13717
R5202 avdd.n9564 avdd.n9563 1.13717
R5203 avdd.n9504 avdd.n9503 1.13717
R5204 avdd.n9508 avdd.n9507 1.13717
R5205 avdd.n9484 avdd.n9483 1.13717
R5206 avdd.n10703 avdd.n10702 1.13717
R5207 avdd.n10723 avdd.n10722 1.13717
R5208 avdd.n10742 avdd.n10741 1.13717
R5209 avdd.n10674 avdd.n10673 1.13717
R5210 avdd.n9429 avdd.n9428 1.13717
R5211 avdd.n9434 avdd.n9433 1.13717
R5212 avdd.n9450 avdd.n9449 1.13717
R5213 avdd.n9390 avdd.n9389 1.13717
R5214 avdd.n9394 avdd.n9393 1.13717
R5215 avdd.n9370 avdd.n9369 1.13717
R5216 avdd.n10805 avdd.n10804 1.13717
R5217 avdd.n10825 avdd.n10824 1.13717
R5218 avdd.n10844 avdd.n10843 1.13717
R5219 avdd.n10776 avdd.n10775 1.13717
R5220 avdd.n9315 avdd.n9314 1.13717
R5221 avdd.n9320 avdd.n9319 1.13717
R5222 avdd.n9336 avdd.n9335 1.13717
R5223 avdd.n9276 avdd.n9275 1.13717
R5224 avdd.n9280 avdd.n9279 1.13717
R5225 avdd.n9256 avdd.n9255 1.13717
R5226 avdd.n10907 avdd.n10906 1.13717
R5227 avdd.n10927 avdd.n10926 1.13717
R5228 avdd.n10946 avdd.n10945 1.13717
R5229 avdd.n10878 avdd.n10877 1.13717
R5230 avdd.n9201 avdd.n9200 1.13717
R5231 avdd.n9206 avdd.n9205 1.13717
R5232 avdd.n9222 avdd.n9221 1.13717
R5233 avdd.n9162 avdd.n9161 1.13717
R5234 avdd.n9166 avdd.n9165 1.13717
R5235 avdd.n9142 avdd.n9141 1.13717
R5236 avdd.n11009 avdd.n11008 1.13717
R5237 avdd.n11029 avdd.n11028 1.13717
R5238 avdd.n11048 avdd.n11047 1.13717
R5239 avdd.n10980 avdd.n10979 1.13717
R5240 avdd.n9087 avdd.n9086 1.13717
R5241 avdd.n9092 avdd.n9091 1.13717
R5242 avdd.n9108 avdd.n9107 1.13717
R5243 avdd.n9048 avdd.n9047 1.13717
R5244 avdd.n9052 avdd.n9051 1.13717
R5245 avdd.n9028 avdd.n9027 1.13717
R5246 avdd.n11111 avdd.n11110 1.13717
R5247 avdd.n11131 avdd.n11130 1.13717
R5248 avdd.n11150 avdd.n11149 1.13717
R5249 avdd.n11082 avdd.n11081 1.13717
R5250 avdd.n8973 avdd.n8972 1.13717
R5251 avdd.n8978 avdd.n8977 1.13717
R5252 avdd.n8994 avdd.n8993 1.13717
R5253 avdd.n8934 avdd.n8933 1.13717
R5254 avdd.n8938 avdd.n8937 1.13717
R5255 avdd.n8914 avdd.n8913 1.13717
R5256 avdd.n11213 avdd.n11212 1.13717
R5257 avdd.n11233 avdd.n11232 1.13717
R5258 avdd.n11252 avdd.n11251 1.13717
R5259 avdd.n11184 avdd.n11183 1.13717
R5260 avdd.n110 avdd.n109 1.13717
R5261 avdd.n130 avdd.n129 1.13717
R5262 avdd.n180 avdd.n179 1.13717
R5263 avdd.n160 avdd.n159 1.13717
R5264 avdd.n8826 avdd.n8825 1.13717
R5265 avdd.n8846 avdd.n8845 1.13717
R5266 avdd.n8865 avdd.n8864 1.13717
R5267 avdd.n8813 avdd.n8812 1.13717
R5268 avdd.n240 avdd.n239 1.13717
R5269 avdd.n260 avdd.n259 1.13717
R5270 avdd.n310 avdd.n309 1.13717
R5271 avdd.n290 avdd.n289 1.13717
R5272 avdd.n8740 avdd.n8739 1.13717
R5273 avdd.n8760 avdd.n8759 1.13717
R5274 avdd.n8779 avdd.n8778 1.13717
R5275 avdd.n8727 avdd.n8726 1.13717
R5276 avdd.n370 avdd.n369 1.13717
R5277 avdd.n390 avdd.n389 1.13717
R5278 avdd.n440 avdd.n439 1.13717
R5279 avdd.n420 avdd.n419 1.13717
R5280 avdd.n8654 avdd.n8653 1.13717
R5281 avdd.n8674 avdd.n8673 1.13717
R5282 avdd.n8693 avdd.n8692 1.13717
R5283 avdd.n8641 avdd.n8640 1.13717
R5284 avdd.n500 avdd.n499 1.13717
R5285 avdd.n520 avdd.n519 1.13717
R5286 avdd.n570 avdd.n569 1.13717
R5287 avdd.n550 avdd.n549 1.13717
R5288 avdd.n8568 avdd.n8567 1.13717
R5289 avdd.n8588 avdd.n8587 1.13717
R5290 avdd.n8607 avdd.n8606 1.13717
R5291 avdd.n8555 avdd.n8554 1.13717
R5292 avdd.n630 avdd.n629 1.13717
R5293 avdd.n650 avdd.n649 1.13717
R5294 avdd.n700 avdd.n699 1.13717
R5295 avdd.n680 avdd.n679 1.13717
R5296 avdd.n8482 avdd.n8481 1.13717
R5297 avdd.n8502 avdd.n8501 1.13717
R5298 avdd.n8521 avdd.n8520 1.13717
R5299 avdd.n8469 avdd.n8468 1.13717
R5300 avdd.n760 avdd.n759 1.13717
R5301 avdd.n780 avdd.n779 1.13717
R5302 avdd.n830 avdd.n829 1.13717
R5303 avdd.n810 avdd.n809 1.13717
R5304 avdd.n8396 avdd.n8395 1.13717
R5305 avdd.n8416 avdd.n8415 1.13717
R5306 avdd.n8435 avdd.n8434 1.13717
R5307 avdd.n8383 avdd.n8382 1.13717
R5308 avdd.n890 avdd.n889 1.13717
R5309 avdd.n910 avdd.n909 1.13717
R5310 avdd.n960 avdd.n959 1.13717
R5311 avdd.n940 avdd.n939 1.13717
R5312 avdd.n8310 avdd.n8309 1.13717
R5313 avdd.n8330 avdd.n8329 1.13717
R5314 avdd.n8349 avdd.n8348 1.13717
R5315 avdd.n8297 avdd.n8296 1.13717
R5316 avdd.n1020 avdd.n1019 1.13717
R5317 avdd.n1040 avdd.n1039 1.13717
R5318 avdd.n1090 avdd.n1089 1.13717
R5319 avdd.n1070 avdd.n1069 1.13717
R5320 avdd.n8224 avdd.n8223 1.13717
R5321 avdd.n8244 avdd.n8243 1.13717
R5322 avdd.n8263 avdd.n8262 1.13717
R5323 avdd.n8211 avdd.n8210 1.13717
R5324 avdd.n1150 avdd.n1149 1.13717
R5325 avdd.n1170 avdd.n1169 1.13717
R5326 avdd.n1220 avdd.n1219 1.13717
R5327 avdd.n1200 avdd.n1199 1.13717
R5328 avdd.n8138 avdd.n8137 1.13717
R5329 avdd.n8158 avdd.n8157 1.13717
R5330 avdd.n8177 avdd.n8176 1.13717
R5331 avdd.n8125 avdd.n8124 1.13717
R5332 avdd.n1280 avdd.n1279 1.13717
R5333 avdd.n1300 avdd.n1299 1.13717
R5334 avdd.n1350 avdd.n1349 1.13717
R5335 avdd.n1330 avdd.n1329 1.13717
R5336 avdd.n8052 avdd.n8051 1.13717
R5337 avdd.n8072 avdd.n8071 1.13717
R5338 avdd.n8091 avdd.n8090 1.13717
R5339 avdd.n8039 avdd.n8038 1.13717
R5340 avdd.n1410 avdd.n1409 1.13717
R5341 avdd.n1430 avdd.n1429 1.13717
R5342 avdd.n1480 avdd.n1479 1.13717
R5343 avdd.n1460 avdd.n1459 1.13717
R5344 avdd.n7966 avdd.n7965 1.13717
R5345 avdd.n7986 avdd.n7985 1.13717
R5346 avdd.n8005 avdd.n8004 1.13717
R5347 avdd.n7953 avdd.n7952 1.13717
R5348 avdd.n1540 avdd.n1539 1.13717
R5349 avdd.n1560 avdd.n1559 1.13717
R5350 avdd.n1610 avdd.n1609 1.13717
R5351 avdd.n1590 avdd.n1589 1.13717
R5352 avdd.n7880 avdd.n7879 1.13717
R5353 avdd.n7900 avdd.n7899 1.13717
R5354 avdd.n7919 avdd.n7918 1.13717
R5355 avdd.n7867 avdd.n7866 1.13717
R5356 avdd.n4603 avdd.n4589 1.12991
R5357 avdd.n4538 avdd.n4520 1.12991
R5358 avdd.n3378 avdd.n3169 1.12716
R5359 avdd.n3593 avdd.n3384 1.12716
R5360 avdd.n3808 avdd.n3599 1.12716
R5361 avdd.n4023 avdd.n3814 1.12716
R5362 avdd.n4238 avdd.n4029 1.12716
R5363 avdd.n4453 avdd.n4244 1.12716
R5364 avdd.n4866 avdd.n4862 1.12716
R5365 avdd.n5082 avdd.n5078 1.12716
R5366 avdd.n5298 avdd.n5294 1.12716
R5367 avdd.n5514 avdd.n5510 1.12716
R5368 avdd.n5730 avdd.n5726 1.12716
R5369 avdd.n5946 avdd.n5942 1.12716
R5370 avdd.n6162 avdd.n6158 1.12716
R5371 avdd.n6378 avdd.n6374 1.12716
R5372 avdd.n6594 avdd.n6590 1.12716
R5373 avdd.n6810 avdd.n6806 1.12716
R5374 avdd.n7026 avdd.n7022 1.12716
R5375 avdd.n7242 avdd.n7238 1.12716
R5376 avdd.n10027 avdd.n10025 1.12716
R5377 avdd.n9913 avdd.n9911 1.12716
R5378 avdd.n9799 avdd.n9797 1.12716
R5379 avdd.n9685 avdd.n9683 1.12716
R5380 avdd.n9571 avdd.n9569 1.12716
R5381 avdd.n9457 avdd.n9455 1.12716
R5382 avdd.n9343 avdd.n9341 1.12716
R5383 avdd.n9229 avdd.n9227 1.12716
R5384 avdd.n9115 avdd.n9113 1.12716
R5385 avdd.n9001 avdd.n8999 1.12716
R5386 avdd.n1895 avdd.n1878 1.12623
R5387 avdd.n2195 avdd.n2144 1.12623
R5388 avdd.n2410 avdd.n2359 1.12623
R5389 avdd.n2625 avdd.n2574 1.12623
R5390 avdd.n2840 avdd.n2789 1.12623
R5391 avdd.n3055 avdd.n3004 1.12623
R5392 avdd.n3185 avdd.n3169 1.12623
R5393 avdd.n3400 avdd.n3384 1.12623
R5394 avdd.n3615 avdd.n3599 1.12623
R5395 avdd.n3830 avdd.n3814 1.12623
R5396 avdd.n4045 avdd.n4029 1.12623
R5397 avdd.n4260 avdd.n4244 1.12623
R5398 avdd.n4867 avdd.n4866 1.12623
R5399 avdd.n5083 avdd.n5082 1.12623
R5400 avdd.n5299 avdd.n5298 1.12623
R5401 avdd.n5515 avdd.n5514 1.12623
R5402 avdd.n5731 avdd.n5730 1.12623
R5403 avdd.n5947 avdd.n5946 1.12623
R5404 avdd.n6163 avdd.n6162 1.12623
R5405 avdd.n6379 avdd.n6378 1.12623
R5406 avdd.n6595 avdd.n6594 1.12623
R5407 avdd.n6811 avdd.n6810 1.12623
R5408 avdd.n7027 avdd.n7026 1.12623
R5409 avdd.n7243 avdd.n7242 1.12623
R5410 avdd.n10027 avdd.n10010 1.12623
R5411 avdd.n9913 avdd.n9896 1.12623
R5412 avdd.n9799 avdd.n9782 1.12623
R5413 avdd.n9685 avdd.n9669 1.12623
R5414 avdd.n9571 avdd.n9554 1.12623
R5415 avdd.n9457 avdd.n9440 1.12623
R5416 avdd.n9343 avdd.n9326 1.12623
R5417 avdd.n9229 avdd.n9212 1.12623
R5418 avdd.n9115 avdd.n9098 1.12623
R5419 avdd.n9001 avdd.n8984 1.12623
R5420 avdd avdd.n4463 1.1018
R5421 avdd.n7504 avdd.n7503 1.09272
R5422 avdd.n7570 avdd.n7408 1.09272
R5423 avdd.n7604 avdd.n7603 1.09272
R5424 avdd.n7471 avdd.n7425 1.09216
R5425 avdd.n1707 avdd.n1659 1.09203
R5426 avdd.n1743 avdd.n1742 1.09203
R5427 avdd.n1797 avdd.n1623 1.09203
R5428 avdd.n1833 avdd.n1832 1.09203
R5429 avdd.n4808 avdd.n4457 1.08442
R5430 avdd.n7401 avdd.n1872 1.06427
R5431 avdd.n11265 avdd.n11264 1.05726
R5432 avdd.n4610 avdd.n4609 0.88175
R5433 avdd.n1909 avdd.n1906 0.874073
R5434 avdd.n2163 avdd.n2160 0.874073
R5435 avdd.n2378 avdd.n2375 0.874073
R5436 avdd.n2593 avdd.n2590 0.874073
R5437 avdd.n2808 avdd.n2805 0.874073
R5438 avdd.n3023 avdd.n3020 0.874073
R5439 avdd.n3199 avdd.n3196 0.874073
R5440 avdd.n3414 avdd.n3411 0.874073
R5441 avdd.n3629 avdd.n3626 0.874073
R5442 avdd.n3844 avdd.n3841 0.874073
R5443 avdd.n4059 avdd.n4056 0.874073
R5444 avdd.n4274 avdd.n4271 0.874073
R5445 avdd.n4885 avdd.n4882 0.874073
R5446 avdd.n5101 avdd.n5098 0.874073
R5447 avdd.n5317 avdd.n5314 0.874073
R5448 avdd.n5533 avdd.n5530 0.874073
R5449 avdd.n5749 avdd.n5746 0.874073
R5450 avdd.n5965 avdd.n5962 0.874073
R5451 avdd.n6181 avdd.n6178 0.874073
R5452 avdd.n6397 avdd.n6394 0.874073
R5453 avdd.n6613 avdd.n6610 0.874073
R5454 avdd.n6829 avdd.n6826 0.874073
R5455 avdd.n7045 avdd.n7042 0.874073
R5456 avdd.n7261 avdd.n7258 0.874073
R5457 avdd.n7755 avdd.n7754 0.874073
R5458 avdd.n10234 avdd.n10233 0.874073
R5459 avdd.n9988 avdd.n9987 0.874073
R5460 avdd.n9874 avdd.n9873 0.874073
R5461 avdd.n9760 avdd.n9759 0.874073
R5462 avdd.n9647 avdd.n9646 0.874073
R5463 avdd.n9532 avdd.n9531 0.874073
R5464 avdd.n9418 avdd.n9417 0.874073
R5465 avdd.n9304 avdd.n9303 0.874073
R5466 avdd.n9190 avdd.n9189 0.874073
R5467 avdd.n9076 avdd.n9075 0.874073
R5468 avdd.n8962 avdd.n8961 0.874073
R5469 avdd.n88 avdd.n87 0.874073
R5470 avdd.n218 avdd.n217 0.874073
R5471 avdd.n348 avdd.n347 0.874073
R5472 avdd.n478 avdd.n477 0.874073
R5473 avdd.n608 avdd.n607 0.874073
R5474 avdd.n738 avdd.n737 0.874073
R5475 avdd.n868 avdd.n867 0.874073
R5476 avdd.n998 avdd.n997 0.874073
R5477 avdd.n1128 avdd.n1127 0.874073
R5478 avdd.n1258 avdd.n1257 0.874073
R5479 avdd.n1388 avdd.n1387 0.874073
R5480 avdd.n1518 avdd.n1517 0.874073
R5481 avdd.n7579 avdd.n7578 0.863992
R5482 avdd.n7538 avdd.n7537 0.863992
R5483 avdd.n7479 avdd.n7478 0.863992
R5484 avdd.n7439 avdd.n7438 0.863992
R5485 avdd.n1686 avdd.n1685 0.863992
R5486 avdd.n1715 avdd.n1714 0.863992
R5487 avdd.n1776 avdd.n1775 0.863992
R5488 avdd.n1805 avdd.n1804 0.863992
R5489 avdd.n4614 avdd.n4613 0.853625
R5490 avdd.n2063 avdd.n2062 0.853
R5491 avdd.n1908 avdd.n1902 0.853
R5492 avdd.n2235 avdd.n2118 0.853
R5493 avdd.n2162 avdd.n2156 0.853
R5494 avdd.n2450 avdd.n2333 0.853
R5495 avdd.n2377 avdd.n2371 0.853
R5496 avdd.n2665 avdd.n2548 0.853
R5497 avdd.n2592 avdd.n2586 0.853
R5498 avdd.n2880 avdd.n2763 0.853
R5499 avdd.n2807 avdd.n2801 0.853
R5500 avdd.n3095 avdd.n2978 0.853
R5501 avdd.n3022 avdd.n3016 0.853
R5502 avdd.n3352 avdd.n3351 0.853
R5503 avdd.n3198 avdd.n3192 0.853
R5504 avdd.n3567 avdd.n3566 0.853
R5505 avdd.n3413 avdd.n3407 0.853
R5506 avdd.n3782 avdd.n3781 0.853
R5507 avdd.n3628 avdd.n3622 0.853
R5508 avdd.n3997 avdd.n3996 0.853
R5509 avdd.n3843 avdd.n3837 0.853
R5510 avdd.n4212 avdd.n4211 0.853
R5511 avdd.n4058 avdd.n4052 0.853
R5512 avdd.n4427 avdd.n4426 0.853
R5513 avdd.n4273 avdd.n4267 0.853
R5514 avdd.n4884 avdd.n4878 0.853
R5515 avdd.n4957 avdd.n4840 0.853
R5516 avdd.n5100 avdd.n5094 0.853
R5517 avdd.n5173 avdd.n5056 0.853
R5518 avdd.n5316 avdd.n5310 0.853
R5519 avdd.n5389 avdd.n5272 0.853
R5520 avdd.n5532 avdd.n5526 0.853
R5521 avdd.n5605 avdd.n5488 0.853
R5522 avdd.n5748 avdd.n5742 0.853
R5523 avdd.n5821 avdd.n5704 0.853
R5524 avdd.n5964 avdd.n5958 0.853
R5525 avdd.n6037 avdd.n5920 0.853
R5526 avdd.n6180 avdd.n6174 0.853
R5527 avdd.n6253 avdd.n6136 0.853
R5528 avdd.n6396 avdd.n6390 0.853
R5529 avdd.n6469 avdd.n6352 0.853
R5530 avdd.n6612 avdd.n6606 0.853
R5531 avdd.n6685 avdd.n6568 0.853
R5532 avdd.n6828 avdd.n6822 0.853
R5533 avdd.n6901 avdd.n6784 0.853
R5534 avdd.n7044 avdd.n7038 0.853
R5535 avdd.n7117 avdd.n7000 0.853
R5536 avdd.n7260 avdd.n7254 0.853
R5537 avdd.n7333 avdd.n7216 0.853
R5538 avdd.n7753 avdd.n7752 0.853
R5539 avdd.n7662 avdd.n7661 0.853
R5540 avdd.n10232 avdd.n10231 0.853
R5541 avdd.n10141 avdd.n10140 0.853
R5542 avdd.n9986 avdd.n9985 0.853
R5543 avdd.n10279 avdd.n10278 0.853
R5544 avdd.n9872 avdd.n9871 0.853
R5545 avdd.n10381 avdd.n10380 0.853
R5546 avdd.n9758 avdd.n9757 0.853
R5547 avdd.n10483 avdd.n10482 0.853
R5548 avdd.n9645 avdd.n9644 0.853
R5549 avdd.n10585 avdd.n10584 0.853
R5550 avdd.n9530 avdd.n9529 0.853
R5551 avdd.n10687 avdd.n10686 0.853
R5552 avdd.n9416 avdd.n9415 0.853
R5553 avdd.n10789 avdd.n10788 0.853
R5554 avdd.n9302 avdd.n9301 0.853
R5555 avdd.n10891 avdd.n10890 0.853
R5556 avdd.n9188 avdd.n9187 0.853
R5557 avdd.n10993 avdd.n10992 0.853
R5558 avdd.n9074 avdd.n9073 0.853
R5559 avdd.n11095 avdd.n11094 0.853
R5560 avdd.n8960 avdd.n8959 0.853
R5561 avdd.n11197 avdd.n11196 0.853
R5562 avdd.n145 avdd.n144 0.853
R5563 avdd.n86 avdd.n85 0.853
R5564 avdd.n275 avdd.n274 0.853
R5565 avdd.n216 avdd.n215 0.853
R5566 avdd.n405 avdd.n404 0.853
R5567 avdd.n346 avdd.n345 0.853
R5568 avdd.n535 avdd.n534 0.853
R5569 avdd.n476 avdd.n475 0.853
R5570 avdd.n665 avdd.n664 0.853
R5571 avdd.n606 avdd.n605 0.853
R5572 avdd.n795 avdd.n794 0.853
R5573 avdd.n736 avdd.n735 0.853
R5574 avdd.n925 avdd.n924 0.853
R5575 avdd.n866 avdd.n865 0.853
R5576 avdd.n1055 avdd.n1054 0.853
R5577 avdd.n996 avdd.n995 0.853
R5578 avdd.n1185 avdd.n1184 0.853
R5579 avdd.n1126 avdd.n1125 0.853
R5580 avdd.n1315 avdd.n1314 0.853
R5581 avdd.n1256 avdd.n1255 0.853
R5582 avdd.n1445 avdd.n1444 0.853
R5583 avdd.n1386 avdd.n1385 0.853
R5584 avdd.n1575 avdd.n1574 0.853
R5585 avdd.n1516 avdd.n1515 0.853
R5586 avdd.n2089 avdd.n1878 0.840229
R5587 avdd.n2196 avdd.n2195 0.840229
R5588 avdd.n2411 avdd.n2410 0.840229
R5589 avdd.n2626 avdd.n2625 0.840229
R5590 avdd.n2841 avdd.n2840 0.840229
R5591 avdd.n3056 avdd.n3055 0.840229
R5592 avdd.n186 avdd.n185 0.840229
R5593 avdd.n316 avdd.n315 0.840229
R5594 avdd.n446 avdd.n445 0.840229
R5595 avdd.n576 avdd.n575 0.840229
R5596 avdd.n706 avdd.n705 0.840229
R5597 avdd.n836 avdd.n835 0.840229
R5598 avdd.n966 avdd.n965 0.840229
R5599 avdd.n1096 avdd.n1095 0.840229
R5600 avdd.n1226 avdd.n1225 0.840229
R5601 avdd.n1356 avdd.n1355 0.840229
R5602 avdd.n1486 avdd.n1485 0.840229
R5603 avdd.n1616 avdd.n1615 0.840229
R5604 avdd.n7762 avdd.n7739 0.84004
R5605 avdd.n10241 avdd.n10218 0.84004
R5606 avdd.n2036 avdd.n2008 0.836345
R5607 avdd.n2096 avdd.n2093 0.836345
R5608 avdd.n2311 avdd.n2308 0.836345
R5609 avdd.n2526 avdd.n2523 0.836345
R5610 avdd.n2741 avdd.n2738 0.836345
R5611 avdd.n2956 avdd.n2953 0.836345
R5612 avdd.n5021 avdd.n4817 0.836345
R5613 avdd.n5237 avdd.n5033 0.836345
R5614 avdd.n5453 avdd.n5249 0.836345
R5615 avdd.n5669 avdd.n5465 0.836345
R5616 avdd.n5885 avdd.n5681 0.836345
R5617 avdd.n6101 avdd.n5897 0.836345
R5618 avdd.n6317 avdd.n6113 0.836345
R5619 avdd.n6533 avdd.n6329 0.836345
R5620 avdd.n6749 avdd.n6545 0.836345
R5621 avdd.n6965 avdd.n6761 0.836345
R5622 avdd.n7181 avdd.n6977 0.836345
R5623 avdd.n7397 avdd.n7193 0.836345
R5624 avdd.n7852 avdd.n7849 0.836345
R5625 avdd.n10110 avdd.n10107 0.836345
R5626 avdd.n10342 avdd.n10340 0.836345
R5627 avdd.n10444 avdd.n10442 0.836345
R5628 avdd.n10546 avdd.n10544 0.836345
R5629 avdd.n10648 avdd.n10646 0.836345
R5630 avdd.n10750 avdd.n10748 0.836345
R5631 avdd.n10852 avdd.n10850 0.836345
R5632 avdd.n10954 avdd.n10952 0.836345
R5633 avdd.n11056 avdd.n11054 0.836345
R5634 avdd.n11158 avdd.n11156 0.836345
R5635 avdd.n11260 avdd.n11258 0.836345
R5636 avdd.n8885 avdd.n8871 0.836345
R5637 avdd.n8799 avdd.n8785 0.836345
R5638 avdd.n8713 avdd.n8699 0.836345
R5639 avdd.n8627 avdd.n8613 0.836345
R5640 avdd.n8541 avdd.n8527 0.836345
R5641 avdd.n8455 avdd.n8441 0.836345
R5642 avdd.n8369 avdd.n8355 0.836345
R5643 avdd.n8283 avdd.n8269 0.836345
R5644 avdd.n8197 avdd.n8183 0.836345
R5645 avdd.n8111 avdd.n8097 0.836345
R5646 avdd.n8025 avdd.n8011 0.836345
R5647 avdd.n7939 avdd.n7925 0.836345
R5648 avdd.n7453 avdd.n7452 0.820933
R5649 avdd.n7492 avdd.n7491 0.820933
R5650 avdd.n7552 avdd.n7551 0.820933
R5651 avdd.n7592 avdd.n7591 0.820933
R5652 avdd.n1818 avdd.n1806 0.820933
R5653 avdd.n1644 avdd.n1632 0.820933
R5654 avdd.n1728 avdd.n1716 0.820933
R5655 avdd.n1680 avdd.n1668 0.820933
R5656 avdd.n1709 avdd.n1708 0.806383
R5657 avdd.n1741 avdd.n1740 0.806383
R5658 avdd.n1799 avdd.n1798 0.806383
R5659 avdd.n1831 avdd.n1830 0.806383
R5660 avdd.n7856 avdd.n7855 0.80544
R5661 avdd.n7502 avdd.n7501 0.79957
R5662 avdd.n7573 avdd.n7571 0.79957
R5663 avdd.n7602 avdd.n7601 0.79957
R5664 avdd.n7473 avdd.n7472 0.79957
R5665 avdd.n4605 avdd.n4504 0.753441
R5666 avdd.n4735 avdd.n4734 0.753441
R5667 avdd.n3325 avdd.n3324 0.66357
R5668 avdd.n3540 avdd.n3539 0.66357
R5669 avdd.n3755 avdd.n3754 0.66357
R5670 avdd.n3970 avdd.n3969 0.66357
R5671 avdd.n4185 avdd.n4184 0.66357
R5672 avdd.n4400 avdd.n4399 0.66357
R5673 avdd.n7532 avdd.n7531 0.467369
R5674 avdd.n7628 avdd.n7406 0.467369
R5675 avdd.n7633 avdd.n7632 0.467369
R5676 avdd.n7528 avdd.n7423 0.467369
R5677 avdd.n1766 avdd.n1657 0.467369
R5678 avdd.n1770 avdd.n1769 0.467369
R5679 avdd.n1856 avdd.n1621 0.467369
R5680 avdd.n1867 avdd.n1866 0.467369
R5681 avdd.n4644 avdd.n4643 0.425158
R5682 avdd.n4463 avdd.n4458 0.388379
R5683 avdd.n4524 avdd.n4519 0.376971
R5684 avdd.n1945 avdd.n1944 0.329317
R5685 avdd.n2041 avdd.n2040 0.329317
R5686 avdd.n2201 avdd.n2200 0.329317
R5687 avdd.n2281 avdd.n2280 0.329317
R5688 avdd.n2416 avdd.n2415 0.329317
R5689 avdd.n2496 avdd.n2495 0.329317
R5690 avdd.n2631 avdd.n2630 0.329317
R5691 avdd.n2711 avdd.n2710 0.329317
R5692 avdd.n2846 avdd.n2845 0.329317
R5693 avdd.n2926 avdd.n2925 0.329317
R5694 avdd.n3061 avdd.n3060 0.329317
R5695 avdd.n3141 avdd.n3140 0.329317
R5696 avdd.n3235 avdd.n3234 0.329317
R5697 avdd.n3330 avdd.n3329 0.329317
R5698 avdd.n3450 avdd.n3449 0.329317
R5699 avdd.n3545 avdd.n3544 0.329317
R5700 avdd.n3665 avdd.n3664 0.329317
R5701 avdd.n3760 avdd.n3759 0.329317
R5702 avdd.n3880 avdd.n3879 0.329317
R5703 avdd.n3975 avdd.n3974 0.329317
R5704 avdd.n4095 avdd.n4094 0.329317
R5705 avdd.n4190 avdd.n4189 0.329317
R5706 avdd.n4310 avdd.n4309 0.329317
R5707 avdd.n4405 avdd.n4404 0.329317
R5708 avdd.n4923 avdd.n4922 0.329317
R5709 avdd.n5000 avdd.n4999 0.329317
R5710 avdd.n5139 avdd.n5138 0.329317
R5711 avdd.n5216 avdd.n5215 0.329317
R5712 avdd.n5355 avdd.n5354 0.329317
R5713 avdd.n5432 avdd.n5431 0.329317
R5714 avdd.n5571 avdd.n5570 0.329317
R5715 avdd.n5648 avdd.n5647 0.329317
R5716 avdd.n5787 avdd.n5786 0.329317
R5717 avdd.n5864 avdd.n5863 0.329317
R5718 avdd.n6003 avdd.n6002 0.329317
R5719 avdd.n6080 avdd.n6079 0.329317
R5720 avdd.n6219 avdd.n6218 0.329317
R5721 avdd.n6296 avdd.n6295 0.329317
R5722 avdd.n6435 avdd.n6434 0.329317
R5723 avdd.n6512 avdd.n6511 0.329317
R5724 avdd.n6651 avdd.n6650 0.329317
R5725 avdd.n6728 avdd.n6727 0.329317
R5726 avdd.n6867 avdd.n6866 0.329317
R5727 avdd.n6944 avdd.n6943 0.329317
R5728 avdd.n7083 avdd.n7082 0.329317
R5729 avdd.n7160 avdd.n7159 0.329317
R5730 avdd.n7299 avdd.n7298 0.329317
R5731 avdd.n7376 avdd.n7375 0.329317
R5732 avdd.n1933 avdd.n1932 0.306507
R5733 avdd.n2076 avdd.n2075 0.306507
R5734 avdd.n1969 avdd.n1968 0.306507
R5735 avdd.n1974 avdd.n1970 0.306507
R5736 avdd.n2050 avdd.n2049 0.306507
R5737 avdd.n2020 avdd.n2019 0.306507
R5738 avdd.n2186 avdd.n2185 0.306507
R5739 avdd.n2221 avdd.n2220 0.306507
R5740 avdd.n2222 avdd.n2117 0.306507
R5741 avdd.n2243 avdd.n2242 0.306507
R5742 avdd.n2262 avdd.n2261 0.306507
R5743 avdd.n2294 avdd.n2293 0.306507
R5744 avdd.n2401 avdd.n2400 0.306507
R5745 avdd.n2436 avdd.n2435 0.306507
R5746 avdd.n2437 avdd.n2332 0.306507
R5747 avdd.n2458 avdd.n2457 0.306507
R5748 avdd.n2477 avdd.n2476 0.306507
R5749 avdd.n2509 avdd.n2508 0.306507
R5750 avdd.n2616 avdd.n2615 0.306507
R5751 avdd.n2651 avdd.n2650 0.306507
R5752 avdd.n2652 avdd.n2547 0.306507
R5753 avdd.n2673 avdd.n2672 0.306507
R5754 avdd.n2692 avdd.n2691 0.306507
R5755 avdd.n2724 avdd.n2723 0.306507
R5756 avdd.n2831 avdd.n2830 0.306507
R5757 avdd.n2866 avdd.n2865 0.306507
R5758 avdd.n2867 avdd.n2762 0.306507
R5759 avdd.n2888 avdd.n2887 0.306507
R5760 avdd.n2907 avdd.n2906 0.306507
R5761 avdd.n2939 avdd.n2938 0.306507
R5762 avdd.n3046 avdd.n3045 0.306507
R5763 avdd.n3081 avdd.n3080 0.306507
R5764 avdd.n3082 avdd.n2977 0.306507
R5765 avdd.n3103 avdd.n3102 0.306507
R5766 avdd.n3122 avdd.n3121 0.306507
R5767 avdd.n3154 avdd.n3153 0.306507
R5768 avdd.n3223 avdd.n3222 0.306507
R5769 avdd.n3365 avdd.n3364 0.306507
R5770 avdd.n3259 avdd.n3258 0.306507
R5771 avdd.n3264 avdd.n3260 0.306507
R5772 avdd.n3339 avdd.n3338 0.306507
R5773 avdd.n3313 avdd.n3312 0.306507
R5774 avdd.n3438 avdd.n3437 0.306507
R5775 avdd.n3580 avdd.n3579 0.306507
R5776 avdd.n3474 avdd.n3473 0.306507
R5777 avdd.n3479 avdd.n3475 0.306507
R5778 avdd.n3554 avdd.n3553 0.306507
R5779 avdd.n3528 avdd.n3527 0.306507
R5780 avdd.n3653 avdd.n3652 0.306507
R5781 avdd.n3795 avdd.n3794 0.306507
R5782 avdd.n3689 avdd.n3688 0.306507
R5783 avdd.n3694 avdd.n3690 0.306507
R5784 avdd.n3769 avdd.n3768 0.306507
R5785 avdd.n3743 avdd.n3742 0.306507
R5786 avdd.n3868 avdd.n3867 0.306507
R5787 avdd.n4010 avdd.n4009 0.306507
R5788 avdd.n3904 avdd.n3903 0.306507
R5789 avdd.n3909 avdd.n3905 0.306507
R5790 avdd.n3984 avdd.n3983 0.306507
R5791 avdd.n3958 avdd.n3957 0.306507
R5792 avdd.n4083 avdd.n4082 0.306507
R5793 avdd.n4225 avdd.n4224 0.306507
R5794 avdd.n4119 avdd.n4118 0.306507
R5795 avdd.n4124 avdd.n4120 0.306507
R5796 avdd.n4199 avdd.n4198 0.306507
R5797 avdd.n4173 avdd.n4172 0.306507
R5798 avdd.n4298 avdd.n4297 0.306507
R5799 avdd.n4440 avdd.n4439 0.306507
R5800 avdd.n4334 avdd.n4333 0.306507
R5801 avdd.n4339 avdd.n4335 0.306507
R5802 avdd.n4414 avdd.n4413 0.306507
R5803 avdd.n4388 avdd.n4387 0.306507
R5804 avdd.n4909 avdd.n4908 0.306507
R5805 avdd.n4943 avdd.n4942 0.306507
R5806 avdd.n4944 avdd.n4839 0.306507
R5807 avdd.n4965 avdd.n4964 0.306507
R5808 avdd.n4984 avdd.n4983 0.306507
R5809 avdd.n5011 avdd.n5010 0.306507
R5810 avdd.n5125 avdd.n5124 0.306507
R5811 avdd.n5159 avdd.n5158 0.306507
R5812 avdd.n5160 avdd.n5055 0.306507
R5813 avdd.n5181 avdd.n5180 0.306507
R5814 avdd.n5200 avdd.n5199 0.306507
R5815 avdd.n5227 avdd.n5226 0.306507
R5816 avdd.n5341 avdd.n5340 0.306507
R5817 avdd.n5375 avdd.n5374 0.306507
R5818 avdd.n5376 avdd.n5271 0.306507
R5819 avdd.n5397 avdd.n5396 0.306507
R5820 avdd.n5416 avdd.n5415 0.306507
R5821 avdd.n5443 avdd.n5442 0.306507
R5822 avdd.n5557 avdd.n5556 0.306507
R5823 avdd.n5591 avdd.n5590 0.306507
R5824 avdd.n5592 avdd.n5487 0.306507
R5825 avdd.n5613 avdd.n5612 0.306507
R5826 avdd.n5632 avdd.n5631 0.306507
R5827 avdd.n5659 avdd.n5658 0.306507
R5828 avdd.n5773 avdd.n5772 0.306507
R5829 avdd.n5807 avdd.n5806 0.306507
R5830 avdd.n5808 avdd.n5703 0.306507
R5831 avdd.n5829 avdd.n5828 0.306507
R5832 avdd.n5848 avdd.n5847 0.306507
R5833 avdd.n5875 avdd.n5874 0.306507
R5834 avdd.n5989 avdd.n5988 0.306507
R5835 avdd.n6023 avdd.n6022 0.306507
R5836 avdd.n6024 avdd.n5919 0.306507
R5837 avdd.n6045 avdd.n6044 0.306507
R5838 avdd.n6064 avdd.n6063 0.306507
R5839 avdd.n6091 avdd.n6090 0.306507
R5840 avdd.n6205 avdd.n6204 0.306507
R5841 avdd.n6239 avdd.n6238 0.306507
R5842 avdd.n6240 avdd.n6135 0.306507
R5843 avdd.n6261 avdd.n6260 0.306507
R5844 avdd.n6280 avdd.n6279 0.306507
R5845 avdd.n6307 avdd.n6306 0.306507
R5846 avdd.n6421 avdd.n6420 0.306507
R5847 avdd.n6455 avdd.n6454 0.306507
R5848 avdd.n6456 avdd.n6351 0.306507
R5849 avdd.n6477 avdd.n6476 0.306507
R5850 avdd.n6496 avdd.n6495 0.306507
R5851 avdd.n6523 avdd.n6522 0.306507
R5852 avdd.n6637 avdd.n6636 0.306507
R5853 avdd.n6671 avdd.n6670 0.306507
R5854 avdd.n6672 avdd.n6567 0.306507
R5855 avdd.n6693 avdd.n6692 0.306507
R5856 avdd.n6712 avdd.n6711 0.306507
R5857 avdd.n6739 avdd.n6738 0.306507
R5858 avdd.n6853 avdd.n6852 0.306507
R5859 avdd.n6887 avdd.n6886 0.306507
R5860 avdd.n6888 avdd.n6783 0.306507
R5861 avdd.n6909 avdd.n6908 0.306507
R5862 avdd.n6928 avdd.n6927 0.306507
R5863 avdd.n6955 avdd.n6954 0.306507
R5864 avdd.n7069 avdd.n7068 0.306507
R5865 avdd.n7103 avdd.n7102 0.306507
R5866 avdd.n7104 avdd.n6999 0.306507
R5867 avdd.n7125 avdd.n7124 0.306507
R5868 avdd.n7144 avdd.n7143 0.306507
R5869 avdd.n7171 avdd.n7170 0.306507
R5870 avdd.n7285 avdd.n7284 0.306507
R5871 avdd.n7319 avdd.n7318 0.306507
R5872 avdd.n7320 avdd.n7215 0.306507
R5873 avdd.n7341 avdd.n7340 0.306507
R5874 avdd.n7360 avdd.n7359 0.306507
R5875 avdd.n7387 avdd.n7386 0.306507
R5876 avdd.n7659 avdd.n7658 0.306507
R5877 avdd.n10138 avdd.n10137 0.306507
R5878 avdd.n10274 avdd.n10273 0.306507
R5879 avdd.n10376 avdd.n10375 0.306507
R5880 avdd.n10478 avdd.n10477 0.306507
R5881 avdd.n10580 avdd.n10579 0.306507
R5882 avdd.n10682 avdd.n10681 0.306507
R5883 avdd.n10784 avdd.n10783 0.306507
R5884 avdd.n10886 avdd.n10885 0.306507
R5885 avdd.n10988 avdd.n10987 0.306507
R5886 avdd.n11090 avdd.n11089 0.306507
R5887 avdd.n11192 avdd.n11191 0.306507
R5888 avdd.n142 avdd.n141 0.306507
R5889 avdd.n272 avdd.n271 0.306507
R5890 avdd.n402 avdd.n401 0.306507
R5891 avdd.n532 avdd.n531 0.306507
R5892 avdd.n662 avdd.n661 0.306507
R5893 avdd.n792 avdd.n791 0.306507
R5894 avdd.n922 avdd.n921 0.306507
R5895 avdd.n1052 avdd.n1051 0.306507
R5896 avdd.n1182 avdd.n1181 0.306507
R5897 avdd.n1312 avdd.n1311 0.306507
R5898 avdd.n1442 avdd.n1441 0.306507
R5899 avdd.n1572 avdd.n1571 0.306507
R5900 avdd.n7578 avdd.n7407 0.305262
R5901 avdd.n7621 avdd.n7620 0.305262
R5902 avdd.n7537 avdd.n7536 0.305262
R5903 avdd.n7555 avdd.n7417 0.305262
R5904 avdd.n7478 avdd.n7424 0.305262
R5905 avdd.n7521 avdd.n7520 0.305262
R5906 avdd.n7438 avdd.n7437 0.305262
R5907 avdd.n7456 avdd.n7435 0.305262
R5908 avdd.n1685 avdd.n1684 0.305262
R5909 avdd.n1689 avdd.n1688 0.305262
R5910 avdd.n1714 avdd.n1658 0.305262
R5911 avdd.n1759 avdd.n1758 0.305262
R5912 avdd.n1775 avdd.n1774 0.305262
R5913 avdd.n1779 avdd.n1778 0.305262
R5914 avdd.n1804 avdd.n1622 0.305262
R5915 avdd.n1849 avdd.n1848 0.305262
R5916 avdd.n4611 avdd.n4521 0.302583
R5917 avdd.n1832 avdd.n1619 0.295115
R5918 avdd.n1801 avdd.n1623 0.295115
R5919 avdd.n1742 avdd.n1648 0.295115
R5920 avdd.n1711 avdd.n1659 0.295115
R5921 avdd.n7504 avdd.n7420 0.294492
R5922 avdd.n7575 avdd.n7408 0.294492
R5923 avdd.n7604 avdd.n7404 0.294492
R5924 avdd.n7475 avdd.n7425 0.294041
R5925 avdd.n4807 avdd.n4806 0.292715
R5926 avdd.n4608 avdd.n4607 0.271333
R5927 avdd.n1914 avdd.n1900 0.261864
R5928 avdd.n1916 avdd.n1915 0.261864
R5929 avdd.n2168 avdd.n2154 0.261864
R5930 avdd.n2170 avdd.n2169 0.261864
R5931 avdd.n2383 avdd.n2369 0.261864
R5932 avdd.n2385 avdd.n2384 0.261864
R5933 avdd.n2598 avdd.n2584 0.261864
R5934 avdd.n2600 avdd.n2599 0.261864
R5935 avdd.n2813 avdd.n2799 0.261864
R5936 avdd.n2815 avdd.n2814 0.261864
R5937 avdd.n3028 avdd.n3014 0.261864
R5938 avdd.n3030 avdd.n3029 0.261864
R5939 avdd.n3204 avdd.n3190 0.261864
R5940 avdd.n3206 avdd.n3205 0.261864
R5941 avdd.n3419 avdd.n3405 0.261864
R5942 avdd.n3421 avdd.n3420 0.261864
R5943 avdd.n3634 avdd.n3620 0.261864
R5944 avdd.n3636 avdd.n3635 0.261864
R5945 avdd.n3849 avdd.n3835 0.261864
R5946 avdd.n3851 avdd.n3850 0.261864
R5947 avdd.n4064 avdd.n4050 0.261864
R5948 avdd.n4066 avdd.n4065 0.261864
R5949 avdd.n4279 avdd.n4265 0.261864
R5950 avdd.n4281 avdd.n4280 0.261864
R5951 avdd.n4890 avdd.n4876 0.261864
R5952 avdd.n4892 avdd.n4891 0.261864
R5953 avdd.n5106 avdd.n5092 0.261864
R5954 avdd.n5108 avdd.n5107 0.261864
R5955 avdd.n5322 avdd.n5308 0.261864
R5956 avdd.n5324 avdd.n5323 0.261864
R5957 avdd.n5538 avdd.n5524 0.261864
R5958 avdd.n5540 avdd.n5539 0.261864
R5959 avdd.n5754 avdd.n5740 0.261864
R5960 avdd.n5756 avdd.n5755 0.261864
R5961 avdd.n5970 avdd.n5956 0.261864
R5962 avdd.n5972 avdd.n5971 0.261864
R5963 avdd.n6186 avdd.n6172 0.261864
R5964 avdd.n6188 avdd.n6187 0.261864
R5965 avdd.n6402 avdd.n6388 0.261864
R5966 avdd.n6404 avdd.n6403 0.261864
R5967 avdd.n6618 avdd.n6604 0.261864
R5968 avdd.n6620 avdd.n6619 0.261864
R5969 avdd.n6834 avdd.n6820 0.261864
R5970 avdd.n6836 avdd.n6835 0.261864
R5971 avdd.n7050 avdd.n7036 0.261864
R5972 avdd.n7052 avdd.n7051 0.261864
R5973 avdd.n7266 avdd.n7252 0.261864
R5974 avdd.n7268 avdd.n7267 0.261864
R5975 avdd.n9982 avdd.n9981 0.261864
R5976 avdd.n9974 avdd.n9973 0.261864
R5977 avdd.n9868 avdd.n9867 0.261864
R5978 avdd.n9860 avdd.n9859 0.261864
R5979 avdd.n9754 avdd.n9753 0.261864
R5980 avdd.n9746 avdd.n9745 0.261864
R5981 avdd.n9641 avdd.n9640 0.261864
R5982 avdd.n9633 avdd.n9632 0.261864
R5983 avdd.n9526 avdd.n9525 0.261864
R5984 avdd.n9518 avdd.n9517 0.261864
R5985 avdd.n9412 avdd.n9411 0.261864
R5986 avdd.n9404 avdd.n9403 0.261864
R5987 avdd.n9298 avdd.n9297 0.261864
R5988 avdd.n9290 avdd.n9289 0.261864
R5989 avdd.n9184 avdd.n9183 0.261864
R5990 avdd.n9176 avdd.n9175 0.261864
R5991 avdd.n9070 avdd.n9069 0.261864
R5992 avdd.n9062 avdd.n9061 0.261864
R5993 avdd.n8956 avdd.n8955 0.261864
R5994 avdd.n8948 avdd.n8947 0.261864
R5995 avdd.n4628 avdd.n4627 0.240083
R5996 avdd.n4738 avdd.n4517 0.240083
R5997 avdd.n7445 avdd.n7443 0.237984
R5998 avdd.n7484 avdd.n7482 0.237984
R5999 avdd.n7544 avdd.n7542 0.237984
R6000 avdd.n7584 avdd.n7582 0.237984
R6001 avdd.n1814 avdd.n1813 0.237984
R6002 avdd.n1640 avdd.n1639 0.237984
R6003 avdd.n1724 avdd.n1723 0.237984
R6004 avdd.n1676 avdd.n1675 0.237984
R6005 avdd avdd.n7504 0.234
R6006 avdd avdd.n7408 0.234
R6007 avdd avdd.n7604 0.234
R6008 avdd avdd.n1659 0.232359
R6009 avdd.n1742 avdd 0.232359
R6010 avdd avdd.n1623 0.232359
R6011 avdd.n1832 avdd 0.232359
R6012 avdd avdd.n7425 0.231541
R6013 avdd.n7856 avdd.n7639 0.225822
R6014 avdd.n2030 avdd.n1872 0.210867
R6015 avdd.n2092 avdd.n2091 0.210867
R6016 avdd.n2306 avdd.n2305 0.210867
R6017 avdd.n2307 avdd.n1877 0.210867
R6018 avdd.n2521 avdd.n2520 0.210867
R6019 avdd.n2522 avdd.n1876 0.210867
R6020 avdd.n2736 avdd.n2735 0.210867
R6021 avdd.n2737 avdd.n1875 0.210867
R6022 avdd.n2951 avdd.n2950 0.210867
R6023 avdd.n2952 avdd.n1874 0.210867
R6024 avdd.n3166 avdd.n3165 0.210867
R6025 avdd.n3167 avdd.n1873 0.210867
R6026 avdd.n3382 avdd.n3381 0.210867
R6027 avdd.n3299 avdd.n3168 0.210867
R6028 avdd.n3597 avdd.n3596 0.210867
R6029 avdd.n3514 avdd.n3383 0.210867
R6030 avdd.n3812 avdd.n3811 0.210867
R6031 avdd.n3729 avdd.n3598 0.210867
R6032 avdd.n4027 avdd.n4026 0.210867
R6033 avdd.n3944 avdd.n3813 0.210867
R6034 avdd.n4242 avdd.n4241 0.210867
R6035 avdd.n4159 avdd.n4028 0.210867
R6036 avdd.n4457 avdd.n4456 0.210867
R6037 avdd.n4374 avdd.n4243 0.210867
R6038 avdd.n5024 avdd.n5023 0.210867
R6039 avdd.n4918 avdd.n4809 0.210867
R6040 avdd.n5240 avdd.n5239 0.210867
R6041 avdd.n5134 avdd.n5025 0.210867
R6042 avdd.n5456 avdd.n5455 0.210867
R6043 avdd.n5350 avdd.n5241 0.210867
R6044 avdd.n5672 avdd.n5671 0.210867
R6045 avdd.n5566 avdd.n5457 0.210867
R6046 avdd.n5888 avdd.n5887 0.210867
R6047 avdd.n5782 avdd.n5673 0.210867
R6048 avdd.n6104 avdd.n6103 0.210867
R6049 avdd.n5998 avdd.n5889 0.210867
R6050 avdd.n6320 avdd.n6319 0.210867
R6051 avdd.n6214 avdd.n6105 0.210867
R6052 avdd.n6536 avdd.n6535 0.210867
R6053 avdd.n6430 avdd.n6321 0.210867
R6054 avdd.n6752 avdd.n6751 0.210867
R6055 avdd.n6646 avdd.n6537 0.210867
R6056 avdd.n6968 avdd.n6967 0.210867
R6057 avdd.n6862 avdd.n6753 0.210867
R6058 avdd.n7184 avdd.n7183 0.210867
R6059 avdd.n7078 avdd.n6969 0.210867
R6060 avdd.n7400 avdd.n7399 0.210867
R6061 avdd.n7294 avdd.n7185 0.210867
R6062 avdd.n7765 avdd.n7764 0.210867
R6063 avdd.n7855 avdd.n7854 0.210867
R6064 avdd.n10244 avdd.n10243 0.210867
R6065 avdd.n10113 avdd.n10112 0.210867
R6066 avdd.n10345 avdd.n10344 0.210867
R6067 avdd.n10346 avdd.n10028 0.210867
R6068 avdd.n10447 avdd.n10446 0.210867
R6069 avdd.n10448 avdd.n9914 0.210867
R6070 avdd.n10549 avdd.n10548 0.210867
R6071 avdd.n10550 avdd.n9800 0.210867
R6072 avdd.n10651 avdd.n10650 0.210867
R6073 avdd.n10652 avdd.n9686 0.210867
R6074 avdd.n10753 avdd.n10752 0.210867
R6075 avdd.n10754 avdd.n9572 0.210867
R6076 avdd.n10855 avdd.n10854 0.210867
R6077 avdd.n10856 avdd.n9458 0.210867
R6078 avdd.n10957 avdd.n10956 0.210867
R6079 avdd.n10958 avdd.n9344 0.210867
R6080 avdd.n11059 avdd.n11058 0.210867
R6081 avdd.n11060 avdd.n9230 0.210867
R6082 avdd.n11161 avdd.n11160 0.210867
R6083 avdd.n11162 avdd.n9116 0.210867
R6084 avdd.n11263 avdd.n11262 0.210867
R6085 avdd.n11264 avdd.n9002 0.210867
R6086 avdd.n8887 avdd.n8886 0.210867
R6087 avdd.n8888 avdd.n187 0.210867
R6088 avdd.n8801 avdd.n8800 0.210867
R6089 avdd.n8802 avdd.n317 0.210867
R6090 avdd.n8715 avdd.n8714 0.210867
R6091 avdd.n8716 avdd.n447 0.210867
R6092 avdd.n8629 avdd.n8628 0.210867
R6093 avdd.n8630 avdd.n577 0.210867
R6094 avdd.n8543 avdd.n8542 0.210867
R6095 avdd.n8544 avdd.n707 0.210867
R6096 avdd.n8457 avdd.n8456 0.210867
R6097 avdd.n8458 avdd.n837 0.210867
R6098 avdd.n8371 avdd.n8370 0.210867
R6099 avdd.n8372 avdd.n967 0.210867
R6100 avdd.n8285 avdd.n8284 0.210867
R6101 avdd.n8286 avdd.n1097 0.210867
R6102 avdd.n8199 avdd.n8198 0.210867
R6103 avdd.n8200 avdd.n1227 0.210867
R6104 avdd.n8113 avdd.n8112 0.210867
R6105 avdd.n8114 avdd.n1357 0.210867
R6106 avdd.n8027 avdd.n8026 0.210867
R6107 avdd.n8028 avdd.n1487 0.210867
R6108 avdd.n7941 avdd.n7940 0.210867
R6109 avdd.n7942 avdd.n1617 0.210867
R6110 avdd.n4641 avdd.n4640 0.18175
R6111 avdd.n7525 avdd.n7476 0.180551
R6112 avdd.n7534 avdd.n7533 0.180551
R6113 avdd.n7625 avdd.n7576 0.180551
R6114 avdd.n7636 avdd.n7634 0.180551
R6115 avdd.n1763 avdd.n1712 0.180294
R6116 avdd.n1772 avdd.n1771 0.180294
R6117 avdd.n1853 avdd.n1802 0.180294
R6118 avdd.n1869 avdd.n1868 0.179926
R6119 avdd.n7402 avdd.n7401 0.151837
R6120 avdd avdd.n7638 0.137535
R6121 avdd avdd.n1871 0.137535
R6122 avdd.n7441 avdd.n7436 0.120292
R6123 avdd.n7455 avdd.n7441 0.120292
R6124 avdd.n7459 avdd.n7434 0.120292
R6125 avdd.n7460 avdd.n7459 0.120292
R6126 avdd.n7461 avdd.n7460 0.120292
R6127 avdd.n7461 avdd.n7431 0.120292
R6128 avdd.n7466 avdd.n7430 0.120292
R6129 avdd.n7467 avdd.n7466 0.120292
R6130 avdd.n7468 avdd.n7467 0.120292
R6131 avdd.n7468 avdd.n7427 0.120292
R6132 avdd.n7476 avdd.n7475 0.120292
R6133 avdd.n7524 avdd.n7523 0.120292
R6134 avdd.n7523 avdd.n7477 0.120292
R6135 avdd.n7518 avdd.n7517 0.120292
R6136 avdd.n7517 avdd.n7516 0.120292
R6137 avdd.n7516 avdd.n7494 0.120292
R6138 avdd.n7512 avdd.n7494 0.120292
R6139 avdd.n7511 avdd.n7510 0.120292
R6140 avdd.n7510 avdd.n7497 0.120292
R6141 avdd.n7506 avdd.n7497 0.120292
R6142 avdd.n7506 avdd.n7505 0.120292
R6143 avdd.n7533 avdd.n7420 0.120292
R6144 avdd.n7540 avdd.n7418 0.120292
R6145 avdd.n7554 avdd.n7540 0.120292
R6146 avdd.n7558 avdd.n7416 0.120292
R6147 avdd.n7559 avdd.n7558 0.120292
R6148 avdd.n7560 avdd.n7559 0.120292
R6149 avdd.n7560 avdd.n7413 0.120292
R6150 avdd.n7565 avdd.n7412 0.120292
R6151 avdd.n7566 avdd.n7565 0.120292
R6152 avdd.n7567 avdd.n7566 0.120292
R6153 avdd.n7567 avdd.n7409 0.120292
R6154 avdd.n7576 avdd.n7575 0.120292
R6155 avdd.n7624 avdd.n7623 0.120292
R6156 avdd.n7623 avdd.n7577 0.120292
R6157 avdd.n7618 avdd.n7617 0.120292
R6158 avdd.n7617 avdd.n7616 0.120292
R6159 avdd.n7616 avdd.n7594 0.120292
R6160 avdd.n7612 avdd.n7594 0.120292
R6161 avdd.n7611 avdd.n7610 0.120292
R6162 avdd.n7610 avdd.n7597 0.120292
R6163 avdd.n7606 avdd.n7597 0.120292
R6164 avdd.n7606 avdd.n7605 0.120292
R6165 avdd.n7634 avdd.n7404 0.120292
R6166 avdd.n1683 avdd.n1682 0.120292
R6167 avdd.n1690 avdd.n1682 0.120292
R6168 avdd.n1693 avdd.n1692 0.120292
R6169 avdd.n1693 avdd.n1665 0.120292
R6170 avdd.n1697 avdd.n1665 0.120292
R6171 avdd.n1698 avdd.n1697 0.120292
R6172 avdd.n1699 avdd.n1662 0.120292
R6173 avdd.n1703 avdd.n1662 0.120292
R6174 avdd.n1704 avdd.n1703 0.120292
R6175 avdd.n1705 avdd.n1704 0.120292
R6176 avdd.n1712 avdd.n1711 0.120292
R6177 avdd.n1762 avdd.n1761 0.120292
R6178 avdd.n1761 avdd.n1713 0.120292
R6179 avdd.n1755 avdd.n1731 0.120292
R6180 avdd.n1755 avdd.n1754 0.120292
R6181 avdd.n1754 avdd.n1753 0.120292
R6182 avdd.n1753 avdd.n1734 0.120292
R6183 avdd.n1748 avdd.n1735 0.120292
R6184 avdd.n1748 avdd.n1747 0.120292
R6185 avdd.n1747 avdd.n1746 0.120292
R6186 avdd.n1746 avdd.n1738 0.120292
R6187 avdd.n1771 avdd.n1648 0.120292
R6188 avdd.n1773 avdd.n1646 0.120292
R6189 avdd.n1780 avdd.n1646 0.120292
R6190 avdd.n1783 avdd.n1782 0.120292
R6191 avdd.n1783 avdd.n1629 0.120292
R6192 avdd.n1787 avdd.n1629 0.120292
R6193 avdd.n1788 avdd.n1787 0.120292
R6194 avdd.n1789 avdd.n1626 0.120292
R6195 avdd.n1793 avdd.n1626 0.120292
R6196 avdd.n1794 avdd.n1793 0.120292
R6197 avdd.n1795 avdd.n1794 0.120292
R6198 avdd.n1802 avdd.n1801 0.120292
R6199 avdd.n1852 avdd.n1851 0.120292
R6200 avdd.n1851 avdd.n1803 0.120292
R6201 avdd.n1845 avdd.n1821 0.120292
R6202 avdd.n1845 avdd.n1844 0.120292
R6203 avdd.n1844 avdd.n1843 0.120292
R6204 avdd.n1843 avdd.n1824 0.120292
R6205 avdd.n1838 avdd.n1825 0.120292
R6206 avdd.n1838 avdd.n1837 0.120292
R6207 avdd.n1837 avdd.n1836 0.120292
R6208 avdd.n1836 avdd.n1828 0.120292
R6209 avdd.n1868 avdd.n1619 0.120292
R6210 avdd.n4803 avdd.n4467 0.120292
R6211 avdd.n4798 avdd.n4797 0.120292
R6212 avdd.n4795 avdd.n4471 0.120292
R6213 avdd.n4790 avdd.n4789 0.120292
R6214 avdd.n4787 avdd.n4475 0.120292
R6215 avdd.n4782 avdd.n4781 0.120292
R6216 avdd.n4779 avdd.n4479 0.120292
R6217 avdd.n4774 avdd.n4773 0.120292
R6218 avdd.n4771 avdd.n4483 0.120292
R6219 avdd.n4767 avdd.n4766 0.120292
R6220 avdd.n13 avdd.n12 0.120292
R6221 avdd.n14 avdd.n13 0.120292
R6222 avdd.n18 avdd.n17 0.120292
R6223 avdd.n19 avdd.n18 0.120292
R6224 avdd.n23 avdd.n22 0.120292
R6225 avdd.n24 avdd.n23 0.120292
R6226 avdd.n28 avdd.n27 0.120292
R6227 avdd.n29 avdd.n28 0.120292
R6228 avdd.n33 avdd.n32 0.120292
R6229 avdd.n34 avdd.n33 0.120292
R6230 avdd.n38 avdd.n37 0.120292
R6231 avdd.n39 avdd.n38 0.120292
R6232 avdd.n43 avdd.n42 0.120292
R6233 avdd.n44 avdd.n43 0.120292
R6234 avdd.n48 avdd.n47 0.120292
R6235 avdd.n49 avdd.n48 0.120292
R6236 avdd.n53 avdd.n1 0.120292
R6237 avdd.n54 avdd.n53 0.120292
R6238 avdd.n4630 avdd.n4623 0.110917
R6239 avdd.n4624 avdd.n4574 0.110917
R6240 avdd.n4593 avdd.n4588 0.110917
R6241 avdd.n4737 avdd.n4736 0.110917
R6242 avdd avdd.n4805 0.102062
R6243 avdd.n4613 avdd.n4610 0.1005
R6244 avdd.n4642 avdd.n4614 0.1005
R6245 avdd.n1970 avdd.n1969 0.0994901
R6246 avdd.n2242 avdd.n2117 0.0994901
R6247 avdd.n2457 avdd.n2332 0.0994901
R6248 avdd.n2672 avdd.n2547 0.0994901
R6249 avdd.n2887 avdd.n2762 0.0994901
R6250 avdd.n3102 avdd.n2977 0.0994901
R6251 avdd.n3260 avdd.n3259 0.0994901
R6252 avdd.n3475 avdd.n3474 0.0994901
R6253 avdd.n3690 avdd.n3689 0.0994901
R6254 avdd.n3905 avdd.n3904 0.0994901
R6255 avdd.n4120 avdd.n4119 0.0994901
R6256 avdd.n4335 avdd.n4334 0.0994901
R6257 avdd.n4964 avdd.n4839 0.0994901
R6258 avdd.n5180 avdd.n5055 0.0994901
R6259 avdd.n5396 avdd.n5271 0.0994901
R6260 avdd.n5612 avdd.n5487 0.0994901
R6261 avdd.n5828 avdd.n5703 0.0994901
R6262 avdd.n6044 avdd.n5919 0.0994901
R6263 avdd.n6260 avdd.n6135 0.0994901
R6264 avdd.n6476 avdd.n6351 0.0994901
R6265 avdd.n6692 avdd.n6567 0.0994901
R6266 avdd.n6908 avdd.n6783 0.0994901
R6267 avdd.n7124 avdd.n6999 0.0994901
R6268 avdd.n7340 avdd.n7215 0.0994901
R6269 avdd avdd.n4803 0.0981562
R6270 avdd avdd.n4798 0.0981562
R6271 avdd avdd.n4795 0.0981562
R6272 avdd avdd.n4790 0.0981562
R6273 avdd avdd.n4787 0.0981562
R6274 avdd avdd.n4782 0.0981562
R6275 avdd avdd.n4779 0.0981562
R6276 avdd avdd.n4774 0.0981562
R6277 avdd avdd.n4771 0.0981562
R6278 avdd.n1819 avdd 0.0924118
R6279 avdd.n1645 avdd 0.0924118
R6280 avdd.n1729 avdd 0.0924118
R6281 avdd.n1681 avdd 0.0924118
R6282 avdd.n1815 avdd.n1807 0.083167
R6283 avdd.n1641 avdd.n1633 0.083167
R6284 avdd.n1725 avdd.n1717 0.083167
R6285 avdd.n1677 avdd.n1669 0.083167
R6286 avdd.n1853 avdd 0.0828946
R6287 avdd avdd.n1772 0.0828946
R6288 avdd.n1763 avdd 0.0828946
R6289 avdd.n7446 avdd.n7445 0.0827222
R6290 avdd.n7485 avdd.n7484 0.0827222
R6291 avdd.n7545 avdd.n7544 0.0827222
R6292 avdd.n7585 avdd.n7584 0.0827222
R6293 avdd.n7525 avdd 0.0826382
R6294 avdd.n7534 avdd 0.0826382
R6295 avdd.n7625 avdd 0.0826382
R6296 avdd.n7636 avdd 0.0826382
R6297 avdd.n57 avdd 0.0825312
R6298 avdd avdd.n1869 0.0822696
R6299 avdd.n1932 avdd.n1892 0.082192
R6300 avdd.n1944 avdd.n1889 0.082192
R6301 avdd.n1946 avdd.n1945 0.082192
R6302 avdd.n2075 avdd.n1947 0.082192
R6303 avdd.n2051 avdd.n2050 0.082192
R6304 avdd.n2041 avdd.n1977 0.082192
R6305 avdd.n2040 avdd.n2000 0.082192
R6306 avdd.n2185 avdd.n2147 0.082192
R6307 avdd.n2200 avdd.n2136 0.082192
R6308 avdd.n2201 avdd.n2129 0.082192
R6309 avdd.n2223 avdd.n2221 0.082192
R6310 avdd.n2261 avdd.n2110 0.082192
R6311 avdd.n2280 avdd.n2103 0.082192
R6312 avdd.n2281 avdd.n2100 0.082192
R6313 avdd.n2400 avdd.n2362 0.082192
R6314 avdd.n2415 avdd.n2351 0.082192
R6315 avdd.n2416 avdd.n2344 0.082192
R6316 avdd.n2438 avdd.n2436 0.082192
R6317 avdd.n2476 avdd.n2325 0.082192
R6318 avdd.n2495 avdd.n2318 0.082192
R6319 avdd.n2496 avdd.n2315 0.082192
R6320 avdd.n2615 avdd.n2577 0.082192
R6321 avdd.n2630 avdd.n2566 0.082192
R6322 avdd.n2631 avdd.n2559 0.082192
R6323 avdd.n2653 avdd.n2651 0.082192
R6324 avdd.n2691 avdd.n2540 0.082192
R6325 avdd.n2710 avdd.n2533 0.082192
R6326 avdd.n2711 avdd.n2530 0.082192
R6327 avdd.n2830 avdd.n2792 0.082192
R6328 avdd.n2845 avdd.n2781 0.082192
R6329 avdd.n2846 avdd.n2774 0.082192
R6330 avdd.n2868 avdd.n2866 0.082192
R6331 avdd.n2906 avdd.n2755 0.082192
R6332 avdd.n2925 avdd.n2748 0.082192
R6333 avdd.n2926 avdd.n2745 0.082192
R6334 avdd.n3045 avdd.n3007 0.082192
R6335 avdd.n3060 avdd.n2996 0.082192
R6336 avdd.n3061 avdd.n2989 0.082192
R6337 avdd.n3083 avdd.n3081 0.082192
R6338 avdd.n3121 avdd.n2970 0.082192
R6339 avdd.n3140 avdd.n2963 0.082192
R6340 avdd.n3141 avdd.n2960 0.082192
R6341 avdd.n3222 avdd.n3182 0.082192
R6342 avdd.n3234 avdd.n3179 0.082192
R6343 avdd.n3236 avdd.n3235 0.082192
R6344 avdd.n3364 avdd.n3237 0.082192
R6345 avdd.n3340 avdd.n3339 0.082192
R6346 avdd.n3330 avdd.n3267 0.082192
R6347 avdd.n3329 avdd.n3290 0.082192
R6348 avdd.n3437 avdd.n3397 0.082192
R6349 avdd.n3449 avdd.n3394 0.082192
R6350 avdd.n3451 avdd.n3450 0.082192
R6351 avdd.n3579 avdd.n3452 0.082192
R6352 avdd.n3555 avdd.n3554 0.082192
R6353 avdd.n3545 avdd.n3482 0.082192
R6354 avdd.n3544 avdd.n3505 0.082192
R6355 avdd.n3652 avdd.n3612 0.082192
R6356 avdd.n3664 avdd.n3609 0.082192
R6357 avdd.n3666 avdd.n3665 0.082192
R6358 avdd.n3794 avdd.n3667 0.082192
R6359 avdd.n3770 avdd.n3769 0.082192
R6360 avdd.n3760 avdd.n3697 0.082192
R6361 avdd.n3759 avdd.n3720 0.082192
R6362 avdd.n3867 avdd.n3827 0.082192
R6363 avdd.n3879 avdd.n3824 0.082192
R6364 avdd.n3881 avdd.n3880 0.082192
R6365 avdd.n4009 avdd.n3882 0.082192
R6366 avdd.n3985 avdd.n3984 0.082192
R6367 avdd.n3975 avdd.n3912 0.082192
R6368 avdd.n3974 avdd.n3935 0.082192
R6369 avdd.n4082 avdd.n4042 0.082192
R6370 avdd.n4094 avdd.n4039 0.082192
R6371 avdd.n4096 avdd.n4095 0.082192
R6372 avdd.n4224 avdd.n4097 0.082192
R6373 avdd.n4200 avdd.n4199 0.082192
R6374 avdd.n4190 avdd.n4127 0.082192
R6375 avdd.n4189 avdd.n4150 0.082192
R6376 avdd.n4297 avdd.n4257 0.082192
R6377 avdd.n4309 avdd.n4254 0.082192
R6378 avdd.n4311 avdd.n4310 0.082192
R6379 avdd.n4439 avdd.n4312 0.082192
R6380 avdd.n4415 avdd.n4414 0.082192
R6381 avdd.n4405 avdd.n4342 0.082192
R6382 avdd.n4404 avdd.n4365 0.082192
R6383 avdd.n4908 avdd.n4869 0.082192
R6384 avdd.n4922 avdd.n4858 0.082192
R6385 avdd.n4923 avdd.n4851 0.082192
R6386 avdd.n4945 avdd.n4943 0.082192
R6387 avdd.n4983 avdd.n4832 0.082192
R6388 avdd.n4999 avdd.n4824 0.082192
R6389 avdd.n5000 avdd.n4821 0.082192
R6390 avdd.n5124 avdd.n5085 0.082192
R6391 avdd.n5138 avdd.n5074 0.082192
R6392 avdd.n5139 avdd.n5067 0.082192
R6393 avdd.n5161 avdd.n5159 0.082192
R6394 avdd.n5199 avdd.n5048 0.082192
R6395 avdd.n5215 avdd.n5040 0.082192
R6396 avdd.n5216 avdd.n5037 0.082192
R6397 avdd.n5340 avdd.n5301 0.082192
R6398 avdd.n5354 avdd.n5290 0.082192
R6399 avdd.n5355 avdd.n5283 0.082192
R6400 avdd.n5377 avdd.n5375 0.082192
R6401 avdd.n5415 avdd.n5264 0.082192
R6402 avdd.n5431 avdd.n5256 0.082192
R6403 avdd.n5432 avdd.n5253 0.082192
R6404 avdd.n5556 avdd.n5517 0.082192
R6405 avdd.n5570 avdd.n5506 0.082192
R6406 avdd.n5571 avdd.n5499 0.082192
R6407 avdd.n5593 avdd.n5591 0.082192
R6408 avdd.n5631 avdd.n5480 0.082192
R6409 avdd.n5647 avdd.n5472 0.082192
R6410 avdd.n5648 avdd.n5469 0.082192
R6411 avdd.n5772 avdd.n5733 0.082192
R6412 avdd.n5786 avdd.n5722 0.082192
R6413 avdd.n5787 avdd.n5715 0.082192
R6414 avdd.n5809 avdd.n5807 0.082192
R6415 avdd.n5847 avdd.n5696 0.082192
R6416 avdd.n5863 avdd.n5688 0.082192
R6417 avdd.n5864 avdd.n5685 0.082192
R6418 avdd.n5988 avdd.n5949 0.082192
R6419 avdd.n6002 avdd.n5938 0.082192
R6420 avdd.n6003 avdd.n5931 0.082192
R6421 avdd.n6025 avdd.n6023 0.082192
R6422 avdd.n6063 avdd.n5912 0.082192
R6423 avdd.n6079 avdd.n5904 0.082192
R6424 avdd.n6080 avdd.n5901 0.082192
R6425 avdd.n6204 avdd.n6165 0.082192
R6426 avdd.n6218 avdd.n6154 0.082192
R6427 avdd.n6219 avdd.n6147 0.082192
R6428 avdd.n6241 avdd.n6239 0.082192
R6429 avdd.n6279 avdd.n6128 0.082192
R6430 avdd.n6295 avdd.n6120 0.082192
R6431 avdd.n6296 avdd.n6117 0.082192
R6432 avdd.n6420 avdd.n6381 0.082192
R6433 avdd.n6434 avdd.n6370 0.082192
R6434 avdd.n6435 avdd.n6363 0.082192
R6435 avdd.n6457 avdd.n6455 0.082192
R6436 avdd.n6495 avdd.n6344 0.082192
R6437 avdd.n6511 avdd.n6336 0.082192
R6438 avdd.n6512 avdd.n6333 0.082192
R6439 avdd.n6636 avdd.n6597 0.082192
R6440 avdd.n6650 avdd.n6586 0.082192
R6441 avdd.n6651 avdd.n6579 0.082192
R6442 avdd.n6673 avdd.n6671 0.082192
R6443 avdd.n6711 avdd.n6560 0.082192
R6444 avdd.n6727 avdd.n6552 0.082192
R6445 avdd.n6728 avdd.n6549 0.082192
R6446 avdd.n6852 avdd.n6813 0.082192
R6447 avdd.n6866 avdd.n6802 0.082192
R6448 avdd.n6867 avdd.n6795 0.082192
R6449 avdd.n6889 avdd.n6887 0.082192
R6450 avdd.n6927 avdd.n6776 0.082192
R6451 avdd.n6943 avdd.n6768 0.082192
R6452 avdd.n6944 avdd.n6765 0.082192
R6453 avdd.n7068 avdd.n7029 0.082192
R6454 avdd.n7082 avdd.n7018 0.082192
R6455 avdd.n7083 avdd.n7011 0.082192
R6456 avdd.n7105 avdd.n7103 0.082192
R6457 avdd.n7143 avdd.n6992 0.082192
R6458 avdd.n7159 avdd.n6984 0.082192
R6459 avdd.n7160 avdd.n6981 0.082192
R6460 avdd.n7284 avdd.n7245 0.082192
R6461 avdd.n7298 avdd.n7234 0.082192
R6462 avdd.n7299 avdd.n7227 0.082192
R6463 avdd.n7321 avdd.n7319 0.082192
R6464 avdd.n7359 avdd.n7208 0.082192
R6465 avdd.n7375 avdd.n7200 0.082192
R6466 avdd.n7376 avdd.n7197 0.082192
R6467 avdd.n7712 avdd.n7711 0.082192
R6468 avdd.n7731 avdd.n7730 0.082192
R6469 avdd.n7690 avdd.n7689 0.082192
R6470 avdd.n7671 avdd.n7670 0.082192
R6471 avdd.n7801 avdd.n7800 0.082192
R6472 avdd.n7821 avdd.n7820 0.082192
R6473 avdd.n7837 avdd.n7836 0.082192
R6474 avdd.n10191 avdd.n10190 0.082192
R6475 avdd.n10210 avdd.n10209 0.082192
R6476 avdd.n10169 avdd.n10168 0.082192
R6477 avdd.n10150 avdd.n10149 0.082192
R6478 avdd.n10079 avdd.n10078 0.082192
R6479 avdd.n10095 avdd.n10094 0.082192
R6480 avdd.n10016 avdd.n10015 0.082192
R6481 avdd.n9953 avdd.n9952 0.082192
R6482 avdd.n9934 avdd.n9933 0.082192
R6483 avdd.n10291 avdd.n10290 0.082192
R6484 avdd.n10311 avdd.n10310 0.082192
R6485 avdd.n10327 avdd.n10326 0.082192
R6486 avdd.n9902 avdd.n9901 0.082192
R6487 avdd.n9839 avdd.n9838 0.082192
R6488 avdd.n9820 avdd.n9819 0.082192
R6489 avdd.n10393 avdd.n10392 0.082192
R6490 avdd.n10413 avdd.n10412 0.082192
R6491 avdd.n10429 avdd.n10428 0.082192
R6492 avdd.n9788 avdd.n9787 0.082192
R6493 avdd.n9725 avdd.n9724 0.082192
R6494 avdd.n9706 avdd.n9705 0.082192
R6495 avdd.n10495 avdd.n10494 0.082192
R6496 avdd.n10515 avdd.n10514 0.082192
R6497 avdd.n10531 avdd.n10530 0.082192
R6498 avdd.n9675 avdd.n9674 0.082192
R6499 avdd.n9612 avdd.n9611 0.082192
R6500 avdd.n9593 avdd.n9592 0.082192
R6501 avdd.n10597 avdd.n10596 0.082192
R6502 avdd.n10617 avdd.n10616 0.082192
R6503 avdd.n10633 avdd.n10632 0.082192
R6504 avdd.n9560 avdd.n9559 0.082192
R6505 avdd.n9497 avdd.n9496 0.082192
R6506 avdd.n9478 avdd.n9477 0.082192
R6507 avdd.n10699 avdd.n10698 0.082192
R6508 avdd.n10719 avdd.n10718 0.082192
R6509 avdd.n10735 avdd.n10734 0.082192
R6510 avdd.n9446 avdd.n9445 0.082192
R6511 avdd.n9383 avdd.n9382 0.082192
R6512 avdd.n9364 avdd.n9363 0.082192
R6513 avdd.n10801 avdd.n10800 0.082192
R6514 avdd.n10821 avdd.n10820 0.082192
R6515 avdd.n10837 avdd.n10836 0.082192
R6516 avdd.n9332 avdd.n9331 0.082192
R6517 avdd.n9269 avdd.n9268 0.082192
R6518 avdd.n9250 avdd.n9249 0.082192
R6519 avdd.n10903 avdd.n10902 0.082192
R6520 avdd.n10923 avdd.n10922 0.082192
R6521 avdd.n10939 avdd.n10938 0.082192
R6522 avdd.n9218 avdd.n9217 0.082192
R6523 avdd.n9155 avdd.n9154 0.082192
R6524 avdd.n9136 avdd.n9135 0.082192
R6525 avdd.n11005 avdd.n11004 0.082192
R6526 avdd.n11025 avdd.n11024 0.082192
R6527 avdd.n11041 avdd.n11040 0.082192
R6528 avdd.n9104 avdd.n9103 0.082192
R6529 avdd.n9041 avdd.n9040 0.082192
R6530 avdd.n9022 avdd.n9021 0.082192
R6531 avdd.n11107 avdd.n11106 0.082192
R6532 avdd.n11127 avdd.n11126 0.082192
R6533 avdd.n11143 avdd.n11142 0.082192
R6534 avdd.n8990 avdd.n8989 0.082192
R6535 avdd.n8927 avdd.n8926 0.082192
R6536 avdd.n8908 avdd.n8907 0.082192
R6537 avdd.n11209 avdd.n11208 0.082192
R6538 avdd.n11229 avdd.n11228 0.082192
R6539 avdd.n11245 avdd.n11244 0.082192
R6540 avdd.n106 avdd.n105 0.082192
R6541 avdd.n126 avdd.n125 0.082192
R6542 avdd.n173 avdd.n172 0.082192
R6543 avdd.n154 avdd.n153 0.082192
R6544 avdd.n8842 avdd.n8841 0.082192
R6545 avdd.n8858 avdd.n8857 0.082192
R6546 avdd.n236 avdd.n235 0.082192
R6547 avdd.n256 avdd.n255 0.082192
R6548 avdd.n303 avdd.n302 0.082192
R6549 avdd.n284 avdd.n283 0.082192
R6550 avdd.n8756 avdd.n8755 0.082192
R6551 avdd.n8772 avdd.n8771 0.082192
R6552 avdd.n366 avdd.n365 0.082192
R6553 avdd.n386 avdd.n385 0.082192
R6554 avdd.n433 avdd.n432 0.082192
R6555 avdd.n414 avdd.n413 0.082192
R6556 avdd.n8670 avdd.n8669 0.082192
R6557 avdd.n8686 avdd.n8685 0.082192
R6558 avdd.n496 avdd.n495 0.082192
R6559 avdd.n516 avdd.n515 0.082192
R6560 avdd.n563 avdd.n562 0.082192
R6561 avdd.n544 avdd.n543 0.082192
R6562 avdd.n8584 avdd.n8583 0.082192
R6563 avdd.n8600 avdd.n8599 0.082192
R6564 avdd.n626 avdd.n625 0.082192
R6565 avdd.n646 avdd.n645 0.082192
R6566 avdd.n693 avdd.n692 0.082192
R6567 avdd.n674 avdd.n673 0.082192
R6568 avdd.n8498 avdd.n8497 0.082192
R6569 avdd.n8514 avdd.n8513 0.082192
R6570 avdd.n756 avdd.n755 0.082192
R6571 avdd.n776 avdd.n775 0.082192
R6572 avdd.n823 avdd.n822 0.082192
R6573 avdd.n804 avdd.n803 0.082192
R6574 avdd.n8412 avdd.n8411 0.082192
R6575 avdd.n8428 avdd.n8427 0.082192
R6576 avdd.n886 avdd.n885 0.082192
R6577 avdd.n906 avdd.n905 0.082192
R6578 avdd.n953 avdd.n952 0.082192
R6579 avdd.n934 avdd.n933 0.082192
R6580 avdd.n8326 avdd.n8325 0.082192
R6581 avdd.n8342 avdd.n8341 0.082192
R6582 avdd.n1016 avdd.n1015 0.082192
R6583 avdd.n1036 avdd.n1035 0.082192
R6584 avdd.n1083 avdd.n1082 0.082192
R6585 avdd.n1064 avdd.n1063 0.082192
R6586 avdd.n8240 avdd.n8239 0.082192
R6587 avdd.n8256 avdd.n8255 0.082192
R6588 avdd.n1146 avdd.n1145 0.082192
R6589 avdd.n1166 avdd.n1165 0.082192
R6590 avdd.n1213 avdd.n1212 0.082192
R6591 avdd.n1194 avdd.n1193 0.082192
R6592 avdd.n8154 avdd.n8153 0.082192
R6593 avdd.n8170 avdd.n8169 0.082192
R6594 avdd.n1276 avdd.n1275 0.082192
R6595 avdd.n1296 avdd.n1295 0.082192
R6596 avdd.n1343 avdd.n1342 0.082192
R6597 avdd.n1324 avdd.n1323 0.082192
R6598 avdd.n8068 avdd.n8067 0.082192
R6599 avdd.n8084 avdd.n8083 0.082192
R6600 avdd.n1406 avdd.n1405 0.082192
R6601 avdd.n1426 avdd.n1425 0.082192
R6602 avdd.n1473 avdd.n1472 0.082192
R6603 avdd.n1454 avdd.n1453 0.082192
R6604 avdd.n7982 avdd.n7981 0.082192
R6605 avdd.n7998 avdd.n7997 0.082192
R6606 avdd.n1536 avdd.n1535 0.082192
R6607 avdd.n1556 avdd.n1555 0.082192
R6608 avdd.n1603 avdd.n1602 0.082192
R6609 avdd.n1584 avdd.n1583 0.082192
R6610 avdd.n7896 avdd.n7895 0.082192
R6611 avdd.n7912 avdd.n7911 0.082192
R6612 avdd.n4609 avdd 0.0770625
R6613 avdd.n10 avdd 0.0742201
R6614 avdd.n4809 avdd.n4808 0.0740675
R6615 avdd.n2089 avdd.n2088 0.0736831
R6616 avdd.n2196 avdd.n2141 0.0736831
R6617 avdd.n2411 avdd.n2356 0.0736831
R6618 avdd.n2626 avdd.n2571 0.0736831
R6619 avdd.n2841 avdd.n2786 0.0736831
R6620 avdd.n3056 avdd.n3001 0.0736831
R6621 avdd.n185 avdd.n184 0.0736831
R6622 avdd.n315 avdd.n314 0.0736831
R6623 avdd.n445 avdd.n444 0.0736831
R6624 avdd.n575 avdd.n574 0.0736831
R6625 avdd.n705 avdd.n704 0.0736831
R6626 avdd.n835 avdd.n834 0.0736831
R6627 avdd.n965 avdd.n964 0.0736831
R6628 avdd.n1095 avdd.n1094 0.0736831
R6629 avdd.n1225 avdd.n1224 0.0736831
R6630 avdd.n1355 avdd.n1354 0.0736831
R6631 avdd.n1485 avdd.n1484 0.0736831
R6632 avdd.n1615 avdd.n1614 0.0736831
R6633 avdd.n7739 avdd.n7701 0.0733157
R6634 avdd.n10218 avdd.n10180 0.0733157
R6635 avdd.n7638 avdd 0.0720601
R6636 avdd.n1871 avdd 0.0720601
R6637 avdd.n3324 avdd.n3322 0.0704421
R6638 avdd.n3539 avdd.n3537 0.0704421
R6639 avdd.n3754 avdd.n3752 0.0704421
R6640 avdd.n3969 avdd.n3967 0.0704421
R6641 avdd.n4184 avdd.n4182 0.0704421
R6642 avdd.n4399 avdd.n4397 0.0704421
R6643 avdd.n10 avdd 0.0695542
R6644 avdd.n4641 avdd.n4615 0.0671667
R6645 avdd.n4608 avdd.n4587 0.0671667
R6646 avdd.n4612 avdd.n4611 0.0671667
R6647 avdd.n3378 avdd.n3377 0.0630449
R6648 avdd.n3593 avdd.n3592 0.0630449
R6649 avdd.n3808 avdd.n3807 0.0630449
R6650 avdd.n4023 avdd.n4022 0.0630449
R6651 avdd.n4238 avdd.n4237 0.0630449
R6652 avdd.n4453 avdd.n4452 0.0630449
R6653 avdd.n4864 avdd.n4862 0.0630449
R6654 avdd.n5080 avdd.n5078 0.0630449
R6655 avdd.n5296 avdd.n5294 0.0630449
R6656 avdd.n5512 avdd.n5510 0.0630449
R6657 avdd.n5728 avdd.n5726 0.0630449
R6658 avdd.n5944 avdd.n5942 0.0630449
R6659 avdd.n6160 avdd.n6158 0.0630449
R6660 avdd.n6376 avdd.n6374 0.0630449
R6661 avdd.n6592 avdd.n6590 0.0630449
R6662 avdd.n6808 avdd.n6806 0.0630449
R6663 avdd.n7024 avdd.n7022 0.0630449
R6664 avdd.n7240 avdd.n7238 0.0630449
R6665 avdd.n10025 avdd.n10024 0.0630449
R6666 avdd.n9911 avdd.n9910 0.0630449
R6667 avdd.n9797 avdd.n9796 0.0630449
R6668 avdd.n9569 avdd.n9568 0.0630449
R6669 avdd.n9455 avdd.n9454 0.0630449
R6670 avdd.n9341 avdd.n9340 0.0630449
R6671 avdd.n9227 avdd.n9226 0.0630449
R6672 avdd.n9113 avdd.n9112 0.0630449
R6673 avdd.n8999 avdd.n8998 0.0630449
R6674 avdd.n1819 avdd 0.063
R6675 avdd.n1645 avdd 0.063
R6676 avdd.n1729 avdd 0.063
R6677 avdd.n1681 avdd 0.063
R6678 avdd avdd.n11266 0.0616979
R6679 avdd.n11265 avdd.n8888 0.0609314
R6680 avdd avdd.n7436 0.0603958
R6681 avdd avdd.n7434 0.0603958
R6682 avdd avdd.n7524 0.0603958
R6683 avdd.n7518 avdd 0.0603958
R6684 avdd avdd.n7418 0.0603958
R6685 avdd avdd.n7416 0.0603958
R6686 avdd avdd.n7624 0.0603958
R6687 avdd.n7618 avdd 0.0603958
R6688 avdd.n1683 avdd 0.0603958
R6689 avdd.n1692 avdd 0.0603958
R6690 avdd avdd.n1762 0.0603958
R6691 avdd.n1731 avdd 0.0603958
R6692 avdd.n1773 avdd 0.0603958
R6693 avdd.n1782 avdd 0.0603958
R6694 avdd avdd.n1852 0.0603958
R6695 avdd.n1821 avdd 0.0603958
R6696 avdd avdd.n4467 0.0603958
R6697 avdd.n4797 avdd 0.0603958
R6698 avdd avdd.n4471 0.0603958
R6699 avdd.n4789 avdd 0.0603958
R6700 avdd avdd.n4788 0.0603958
R6701 avdd avdd.n4475 0.0603958
R6702 avdd.n4781 avdd 0.0603958
R6703 avdd avdd.n4479 0.0603958
R6704 avdd.n4773 avdd 0.0603958
R6705 avdd avdd.n4483 0.0603958
R6706 avdd.n37 avdd 0.0603958
R6707 avdd avdd.n57 0.0603958
R6708 avdd.n1896 avdd.n1895 0.0601691
R6709 avdd.n2150 avdd.n2144 0.0601691
R6710 avdd.n2365 avdd.n2359 0.0601691
R6711 avdd.n2580 avdd.n2574 0.0601691
R6712 avdd.n2795 avdd.n2789 0.0601691
R6713 avdd.n3010 avdd.n3004 0.0601691
R6714 avdd.n3186 avdd.n3185 0.0601691
R6715 avdd.n3401 avdd.n3400 0.0601691
R6716 avdd.n3616 avdd.n3615 0.0601691
R6717 avdd.n3831 avdd.n3830 0.0601691
R6718 avdd.n4046 avdd.n4045 0.0601691
R6719 avdd.n4261 avdd.n4260 0.0601691
R6720 avdd.n4872 avdd.n4867 0.0601691
R6721 avdd.n5088 avdd.n5083 0.0601691
R6722 avdd.n5304 avdd.n5299 0.0601691
R6723 avdd.n5520 avdd.n5515 0.0601691
R6724 avdd.n5736 avdd.n5731 0.0601691
R6725 avdd.n5952 avdd.n5947 0.0601691
R6726 avdd.n6168 avdd.n6163 0.0601691
R6727 avdd.n6384 avdd.n6379 0.0601691
R6728 avdd.n6600 avdd.n6595 0.0601691
R6729 avdd.n6816 avdd.n6811 0.0601691
R6730 avdd.n7032 avdd.n7027 0.0601691
R6731 avdd.n7248 avdd.n7243 0.0601691
R6732 avdd.n7721 avdd.n7720 0.0601691
R6733 avdd.n10200 avdd.n10199 0.0601691
R6734 avdd.n115 avdd.n114 0.0601691
R6735 avdd.n245 avdd.n244 0.0601691
R6736 avdd.n375 avdd.n374 0.0601691
R6737 avdd.n505 avdd.n504 0.0601691
R6738 avdd.n635 avdd.n634 0.0601691
R6739 avdd.n765 avdd.n764 0.0601691
R6740 avdd.n895 avdd.n894 0.0601691
R6741 avdd.n1025 avdd.n1024 0.0601691
R6742 avdd.n1155 avdd.n1154 0.0601691
R6743 avdd.n1285 avdd.n1284 0.0601691
R6744 avdd.n1415 avdd.n1414 0.0601691
R6745 avdd.n1545 avdd.n1544 0.0601691
R6746 avdd.n10244 avdd.n10113 0.0593999
R6747 avdd.n7855 avdd.n7765 0.0593999
R6748 avdd.n4799 avdd 0.0590938
R6749 avdd.n4791 avdd 0.0590938
R6750 avdd.n4783 avdd 0.0590938
R6751 avdd avdd.n4780 0.0590938
R6752 avdd avdd.n4772 0.0590938
R6753 avdd.n17 avdd 0.0590938
R6754 avdd.n27 avdd 0.0590938
R6755 avdd.n32 avdd 0.0590938
R6756 avdd.n42 avdd 0.0590938
R6757 avdd avdd.n1 0.0590938
R6758 avdd.n10652 avdd.n10651 0.0590694
R6759 avdd.n10550 avdd.n10549 0.0590694
R6760 avdd.n10448 avdd.n10447 0.0590694
R6761 avdd.n10346 avdd.n10345 0.0590694
R6762 avdd.n2028 avdd.n2008 0.05882
R6763 avdd.n2097 avdd.n2096 0.05882
R6764 avdd.n2312 avdd.n2311 0.05882
R6765 avdd.n2527 avdd.n2526 0.05882
R6766 avdd.n2742 avdd.n2741 0.05882
R6767 avdd.n2957 avdd.n2956 0.05882
R6768 avdd.n5012 avdd.n4817 0.05882
R6769 avdd.n5228 avdd.n5033 0.05882
R6770 avdd.n5444 avdd.n5249 0.05882
R6771 avdd.n5660 avdd.n5465 0.05882
R6772 avdd.n5876 avdd.n5681 0.05882
R6773 avdd.n6092 avdd.n5897 0.05882
R6774 avdd.n6308 avdd.n6113 0.05882
R6775 avdd.n6524 avdd.n6329 0.05882
R6776 avdd.n6740 avdd.n6545 0.05882
R6777 avdd.n6956 avdd.n6761 0.05882
R6778 avdd.n7172 avdd.n6977 0.05882
R6779 avdd.n7388 avdd.n7193 0.05882
R6780 avdd.n7849 avdd.n7793 0.05882
R6781 avdd.n10107 avdd.n10053 0.05882
R6782 avdd.n10340 avdd.n10270 0.05882
R6783 avdd.n10442 avdd.n10372 0.05882
R6784 avdd.n10544 avdd.n10474 0.05882
R6785 avdd.n10646 avdd.n10576 0.05882
R6786 avdd.n10748 avdd.n10678 0.05882
R6787 avdd.n10850 avdd.n10780 0.05882
R6788 avdd.n10952 avdd.n10882 0.05882
R6789 avdd.n11054 avdd.n10984 0.05882
R6790 avdd.n11156 avdd.n11086 0.05882
R6791 avdd.n11258 avdd.n11188 0.05882
R6792 avdd.n8871 avdd.n8816 0.05882
R6793 avdd.n8785 avdd.n8730 0.05882
R6794 avdd.n8699 avdd.n8644 0.05882
R6795 avdd.n8613 avdd.n8558 0.05882
R6796 avdd.n8527 avdd.n8472 0.05882
R6797 avdd.n8441 avdd.n8386 0.05882
R6798 avdd.n8355 avdd.n8300 0.05882
R6799 avdd.n8269 avdd.n8214 0.05882
R6800 avdd.n8183 avdd.n8128 0.05882
R6801 avdd.n8097 avdd.n8042 0.05882
R6802 avdd.n8011 avdd.n7956 0.05882
R6803 avdd.n7925 avdd.n7870 0.05882
R6804 avdd.n11060 avdd.n11059 0.0587427
R6805 avdd.n10958 avdd.n10957 0.0587427
R6806 avdd.n10856 avdd.n10855 0.0587427
R6807 avdd.n10754 avdd.n10753 0.0587427
R6808 avdd.n11264 avdd.n11263 0.0584196
R6809 avdd.n11162 avdd.n11161 0.0584196
R6810 avdd avdd.n4796 0.0577917
R6811 avdd.n4775 avdd 0.0577917
R6812 avdd.n22 avdd 0.0577917
R6813 avdd.n47 avdd 0.0577917
R6814 avdd.n2069 avdd.n1957 0.0574697
R6815 avdd.n2057 avdd.n2056 0.0574697
R6816 avdd.n1925 avdd.n1897 0.0574697
R6817 avdd.n1924 avdd.n1898 0.0574697
R6818 avdd.n2068 avdd.n2067 0.0574697
R6819 avdd.n2055 avdd.n1971 0.0574697
R6820 avdd.n2230 avdd.n2229 0.0574697
R6821 avdd.n2250 avdd.n2114 0.0574697
R6822 avdd.n2179 avdd.n2151 0.0574697
R6823 avdd.n2178 avdd.n2152 0.0574697
R6824 avdd.n2231 avdd.n2121 0.0574697
R6825 avdd.n2249 avdd.n2115 0.0574697
R6826 avdd.n2445 avdd.n2444 0.0574697
R6827 avdd.n2465 avdd.n2329 0.0574697
R6828 avdd.n2394 avdd.n2366 0.0574697
R6829 avdd.n2393 avdd.n2367 0.0574697
R6830 avdd.n2446 avdd.n2336 0.0574697
R6831 avdd.n2464 avdd.n2330 0.0574697
R6832 avdd.n2660 avdd.n2659 0.0574697
R6833 avdd.n2680 avdd.n2544 0.0574697
R6834 avdd.n2609 avdd.n2581 0.0574697
R6835 avdd.n2608 avdd.n2582 0.0574697
R6836 avdd.n2661 avdd.n2551 0.0574697
R6837 avdd.n2679 avdd.n2545 0.0574697
R6838 avdd.n2875 avdd.n2874 0.0574697
R6839 avdd.n2895 avdd.n2759 0.0574697
R6840 avdd.n2824 avdd.n2796 0.0574697
R6841 avdd.n2823 avdd.n2797 0.0574697
R6842 avdd.n2876 avdd.n2766 0.0574697
R6843 avdd.n2894 avdd.n2760 0.0574697
R6844 avdd.n3090 avdd.n3089 0.0574697
R6845 avdd.n3110 avdd.n2974 0.0574697
R6846 avdd.n3039 avdd.n3011 0.0574697
R6847 avdd.n3038 avdd.n3012 0.0574697
R6848 avdd.n3091 avdd.n2981 0.0574697
R6849 avdd.n3109 avdd.n2975 0.0574697
R6850 avdd.n3358 avdd.n3247 0.0574697
R6851 avdd.n3346 avdd.n3345 0.0574697
R6852 avdd.n3215 avdd.n3187 0.0574697
R6853 avdd.n3214 avdd.n3188 0.0574697
R6854 avdd.n3357 avdd.n3356 0.0574697
R6855 avdd.n3344 avdd.n3261 0.0574697
R6856 avdd.n3573 avdd.n3462 0.0574697
R6857 avdd.n3561 avdd.n3560 0.0574697
R6858 avdd.n3430 avdd.n3402 0.0574697
R6859 avdd.n3429 avdd.n3403 0.0574697
R6860 avdd.n3572 avdd.n3571 0.0574697
R6861 avdd.n3559 avdd.n3476 0.0574697
R6862 avdd.n3788 avdd.n3677 0.0574697
R6863 avdd.n3776 avdd.n3775 0.0574697
R6864 avdd.n3645 avdd.n3617 0.0574697
R6865 avdd.n3644 avdd.n3618 0.0574697
R6866 avdd.n3787 avdd.n3786 0.0574697
R6867 avdd.n3774 avdd.n3691 0.0574697
R6868 avdd.n4003 avdd.n3892 0.0574697
R6869 avdd.n3991 avdd.n3990 0.0574697
R6870 avdd.n3860 avdd.n3832 0.0574697
R6871 avdd.n3859 avdd.n3833 0.0574697
R6872 avdd.n4002 avdd.n4001 0.0574697
R6873 avdd.n3989 avdd.n3906 0.0574697
R6874 avdd.n4218 avdd.n4107 0.0574697
R6875 avdd.n4206 avdd.n4205 0.0574697
R6876 avdd.n4075 avdd.n4047 0.0574697
R6877 avdd.n4074 avdd.n4048 0.0574697
R6878 avdd.n4217 avdd.n4216 0.0574697
R6879 avdd.n4204 avdd.n4121 0.0574697
R6880 avdd.n4433 avdd.n4322 0.0574697
R6881 avdd.n4421 avdd.n4420 0.0574697
R6882 avdd.n4290 avdd.n4262 0.0574697
R6883 avdd.n4289 avdd.n4263 0.0574697
R6884 avdd.n4432 avdd.n4431 0.0574697
R6885 avdd.n4419 avdd.n4336 0.0574697
R6886 avdd.n4952 avdd.n4951 0.0574697
R6887 avdd.n4972 avdd.n4836 0.0574697
R6888 avdd.n4901 avdd.n4873 0.0574697
R6889 avdd.n4900 avdd.n4874 0.0574697
R6890 avdd.n4953 avdd.n4843 0.0574697
R6891 avdd.n4971 avdd.n4837 0.0574697
R6892 avdd.n5168 avdd.n5167 0.0574697
R6893 avdd.n5188 avdd.n5052 0.0574697
R6894 avdd.n5117 avdd.n5089 0.0574697
R6895 avdd.n5116 avdd.n5090 0.0574697
R6896 avdd.n5169 avdd.n5059 0.0574697
R6897 avdd.n5187 avdd.n5053 0.0574697
R6898 avdd.n5384 avdd.n5383 0.0574697
R6899 avdd.n5404 avdd.n5268 0.0574697
R6900 avdd.n5333 avdd.n5305 0.0574697
R6901 avdd.n5332 avdd.n5306 0.0574697
R6902 avdd.n5385 avdd.n5275 0.0574697
R6903 avdd.n5403 avdd.n5269 0.0574697
R6904 avdd.n5600 avdd.n5599 0.0574697
R6905 avdd.n5620 avdd.n5484 0.0574697
R6906 avdd.n5549 avdd.n5521 0.0574697
R6907 avdd.n5548 avdd.n5522 0.0574697
R6908 avdd.n5601 avdd.n5491 0.0574697
R6909 avdd.n5619 avdd.n5485 0.0574697
R6910 avdd.n5816 avdd.n5815 0.0574697
R6911 avdd.n5836 avdd.n5700 0.0574697
R6912 avdd.n5765 avdd.n5737 0.0574697
R6913 avdd.n5764 avdd.n5738 0.0574697
R6914 avdd.n5817 avdd.n5707 0.0574697
R6915 avdd.n5835 avdd.n5701 0.0574697
R6916 avdd.n6032 avdd.n6031 0.0574697
R6917 avdd.n6052 avdd.n5916 0.0574697
R6918 avdd.n5981 avdd.n5953 0.0574697
R6919 avdd.n5980 avdd.n5954 0.0574697
R6920 avdd.n6033 avdd.n5923 0.0574697
R6921 avdd.n6051 avdd.n5917 0.0574697
R6922 avdd.n6248 avdd.n6247 0.0574697
R6923 avdd.n6268 avdd.n6132 0.0574697
R6924 avdd.n6197 avdd.n6169 0.0574697
R6925 avdd.n6196 avdd.n6170 0.0574697
R6926 avdd.n6249 avdd.n6139 0.0574697
R6927 avdd.n6267 avdd.n6133 0.0574697
R6928 avdd.n6464 avdd.n6463 0.0574697
R6929 avdd.n6484 avdd.n6348 0.0574697
R6930 avdd.n6413 avdd.n6385 0.0574697
R6931 avdd.n6412 avdd.n6386 0.0574697
R6932 avdd.n6465 avdd.n6355 0.0574697
R6933 avdd.n6483 avdd.n6349 0.0574697
R6934 avdd.n6680 avdd.n6679 0.0574697
R6935 avdd.n6700 avdd.n6564 0.0574697
R6936 avdd.n6629 avdd.n6601 0.0574697
R6937 avdd.n6628 avdd.n6602 0.0574697
R6938 avdd.n6681 avdd.n6571 0.0574697
R6939 avdd.n6699 avdd.n6565 0.0574697
R6940 avdd.n6896 avdd.n6895 0.0574697
R6941 avdd.n6916 avdd.n6780 0.0574697
R6942 avdd.n6845 avdd.n6817 0.0574697
R6943 avdd.n6844 avdd.n6818 0.0574697
R6944 avdd.n6897 avdd.n6787 0.0574697
R6945 avdd.n6915 avdd.n6781 0.0574697
R6946 avdd.n7112 avdd.n7111 0.0574697
R6947 avdd.n7132 avdd.n6996 0.0574697
R6948 avdd.n7061 avdd.n7033 0.0574697
R6949 avdd.n7060 avdd.n7034 0.0574697
R6950 avdd.n7113 avdd.n7003 0.0574697
R6951 avdd.n7131 avdd.n6997 0.0574697
R6952 avdd.n7328 avdd.n7327 0.0574697
R6953 avdd.n7348 avdd.n7212 0.0574697
R6954 avdd.n7277 avdd.n7249 0.0574697
R6955 avdd.n7276 avdd.n7250 0.0574697
R6956 avdd.n7329 avdd.n7219 0.0574697
R6957 avdd.n7347 avdd.n7213 0.0574697
R6958 avdd.n7642 avdd.n7641 0.0574697
R6959 avdd.n7770 avdd.n7769 0.0574697
R6960 avdd.n7758 avdd.n7757 0.0574697
R6961 avdd.n7666 avdd.n7665 0.0574697
R6962 avdd.n7795 avdd.n7794 0.0574697
R6963 avdd.n10119 avdd.n10118 0.0574697
R6964 avdd.n10030 avdd.n10029 0.0574697
R6965 avdd.n10237 avdd.n10236 0.0574697
R6966 avdd.n10145 avdd.n10144 0.0574697
R6967 avdd.n9920 avdd.n9919 0.0574697
R6968 avdd.n10246 avdd.n10245 0.0574697
R6969 avdd.n9991 avdd.n9990 0.0574697
R6970 avdd.n9967 avdd.n9966 0.0574697
R6971 avdd.n9930 avdd.n9929 0.0574697
R6972 avdd.n10284 avdd.n10283 0.0574697
R6973 avdd.n9806 avdd.n9805 0.0574697
R6974 avdd.n10348 avdd.n10347 0.0574697
R6975 avdd.n9877 avdd.n9876 0.0574697
R6976 avdd.n9853 avdd.n9852 0.0574697
R6977 avdd.n9816 avdd.n9815 0.0574697
R6978 avdd.n10386 avdd.n10385 0.0574697
R6979 avdd.n9692 avdd.n9691 0.0574697
R6980 avdd.n10450 avdd.n10449 0.0574697
R6981 avdd.n9763 avdd.n9762 0.0574697
R6982 avdd.n9739 avdd.n9738 0.0574697
R6983 avdd.n9702 avdd.n9701 0.0574697
R6984 avdd.n10488 avdd.n10487 0.0574697
R6985 avdd.n9578 avdd.n9577 0.0574697
R6986 avdd.n10552 avdd.n10551 0.0574697
R6987 avdd.n9650 avdd.n9649 0.0574697
R6988 avdd.n9626 avdd.n9625 0.0574697
R6989 avdd.n9589 avdd.n9588 0.0574697
R6990 avdd.n10590 avdd.n10589 0.0574697
R6991 avdd.n9464 avdd.n9463 0.0574697
R6992 avdd.n10654 avdd.n10653 0.0574697
R6993 avdd.n9535 avdd.n9534 0.0574697
R6994 avdd.n9511 avdd.n9510 0.0574697
R6995 avdd.n9474 avdd.n9473 0.0574697
R6996 avdd.n10692 avdd.n10691 0.0574697
R6997 avdd.n9350 avdd.n9349 0.0574697
R6998 avdd.n10756 avdd.n10755 0.0574697
R6999 avdd.n9421 avdd.n9420 0.0574697
R7000 avdd.n9397 avdd.n9396 0.0574697
R7001 avdd.n9360 avdd.n9359 0.0574697
R7002 avdd.n10794 avdd.n10793 0.0574697
R7003 avdd.n9236 avdd.n9235 0.0574697
R7004 avdd.n10858 avdd.n10857 0.0574697
R7005 avdd.n9307 avdd.n9306 0.0574697
R7006 avdd.n9283 avdd.n9282 0.0574697
R7007 avdd.n9246 avdd.n9245 0.0574697
R7008 avdd.n10896 avdd.n10895 0.0574697
R7009 avdd.n9122 avdd.n9121 0.0574697
R7010 avdd.n10960 avdd.n10959 0.0574697
R7011 avdd.n9193 avdd.n9192 0.0574697
R7012 avdd.n9169 avdd.n9168 0.0574697
R7013 avdd.n9132 avdd.n9131 0.0574697
R7014 avdd.n10998 avdd.n10997 0.0574697
R7015 avdd.n9008 avdd.n9007 0.0574697
R7016 avdd.n11062 avdd.n11061 0.0574697
R7017 avdd.n9079 avdd.n9078 0.0574697
R7018 avdd.n9055 avdd.n9054 0.0574697
R7019 avdd.n9018 avdd.n9017 0.0574697
R7020 avdd.n11100 avdd.n11099 0.0574697
R7021 avdd.n8894 avdd.n8893 0.0574697
R7022 avdd.n11164 avdd.n11163 0.0574697
R7023 avdd.n8965 avdd.n8964 0.0574697
R7024 avdd.n8941 avdd.n8940 0.0574697
R7025 avdd.n8904 avdd.n8903 0.0574697
R7026 avdd.n11202 avdd.n11201 0.0574697
R7027 avdd.n63 avdd.n62 0.0574697
R7028 avdd.n8873 avdd.n8872 0.0574697
R7029 avdd.n91 avdd.n90 0.0574697
R7030 avdd.n149 avdd.n148 0.0574697
R7031 avdd.n193 avdd.n192 0.0574697
R7032 avdd.n8787 avdd.n8786 0.0574697
R7033 avdd.n221 avdd.n220 0.0574697
R7034 avdd.n279 avdd.n278 0.0574697
R7035 avdd.n323 avdd.n322 0.0574697
R7036 avdd.n8701 avdd.n8700 0.0574697
R7037 avdd.n351 avdd.n350 0.0574697
R7038 avdd.n409 avdd.n408 0.0574697
R7039 avdd.n453 avdd.n452 0.0574697
R7040 avdd.n8615 avdd.n8614 0.0574697
R7041 avdd.n481 avdd.n480 0.0574697
R7042 avdd.n539 avdd.n538 0.0574697
R7043 avdd.n583 avdd.n582 0.0574697
R7044 avdd.n8529 avdd.n8528 0.0574697
R7045 avdd.n611 avdd.n610 0.0574697
R7046 avdd.n669 avdd.n668 0.0574697
R7047 avdd.n713 avdd.n712 0.0574697
R7048 avdd.n8443 avdd.n8442 0.0574697
R7049 avdd.n741 avdd.n740 0.0574697
R7050 avdd.n799 avdd.n798 0.0574697
R7051 avdd.n843 avdd.n842 0.0574697
R7052 avdd.n8357 avdd.n8356 0.0574697
R7053 avdd.n871 avdd.n870 0.0574697
R7054 avdd.n929 avdd.n928 0.0574697
R7055 avdd.n973 avdd.n972 0.0574697
R7056 avdd.n8271 avdd.n8270 0.0574697
R7057 avdd.n1001 avdd.n1000 0.0574697
R7058 avdd.n1059 avdd.n1058 0.0574697
R7059 avdd.n1103 avdd.n1102 0.0574697
R7060 avdd.n8185 avdd.n8184 0.0574697
R7061 avdd.n1131 avdd.n1130 0.0574697
R7062 avdd.n1189 avdd.n1188 0.0574697
R7063 avdd.n1233 avdd.n1232 0.0574697
R7064 avdd.n8099 avdd.n8098 0.0574697
R7065 avdd.n1261 avdd.n1260 0.0574697
R7066 avdd.n1319 avdd.n1318 0.0574697
R7067 avdd.n1363 avdd.n1362 0.0574697
R7068 avdd.n8013 avdd.n8012 0.0574697
R7069 avdd.n1391 avdd.n1390 0.0574697
R7070 avdd.n1449 avdd.n1448 0.0574697
R7071 avdd.n1493 avdd.n1492 0.0574697
R7072 avdd.n7927 avdd.n7926 0.0574697
R7073 avdd.n1521 avdd.n1520 0.0574697
R7074 avdd.n1579 avdd.n1578 0.0574697
R7075 avdd.n7942 avdd.n7941 0.0568563
R7076 avdd.n8028 avdd.n8027 0.0568563
R7077 avdd.n8114 avdd.n8113 0.0565537
R7078 avdd.n8200 avdd.n8199 0.0565537
R7079 avdd.n8286 avdd.n8285 0.0565537
R7080 avdd.n8372 avdd.n8371 0.0565537
R7081 avdd avdd.n4804 0.0564896
R7082 avdd.n4767 avdd 0.0564896
R7083 avdd.n12 avdd 0.0564896
R7084 avdd.n55 avdd 0.0564896
R7085 avdd.n11266 avdd 0.0564896
R7086 avdd.n8458 avdd.n8457 0.0562543
R7087 avdd.n8544 avdd.n8543 0.0562543
R7088 avdd.n8630 avdd.n8629 0.0562543
R7089 avdd.n8716 avdd.n8715 0.0562543
R7090 avdd.n8802 avdd.n8801 0.0559582
R7091 avdd.n8888 avdd.n8887 0.0559582
R7092 avdd.n2011 avdd.n2008 0.0546809
R7093 avdd.n2096 avdd.n2094 0.0546809
R7094 avdd.n2311 avdd.n2309 0.0546809
R7095 avdd.n2526 avdd.n2524 0.0546809
R7096 avdd.n2741 avdd.n2739 0.0546809
R7097 avdd.n2956 avdd.n2954 0.0546809
R7098 avdd.n4817 avdd.n4810 0.0546809
R7099 avdd.n5033 avdd.n5026 0.0546809
R7100 avdd.n5249 avdd.n5242 0.0546809
R7101 avdd.n5465 avdd.n5458 0.0546809
R7102 avdd.n5681 avdd.n5674 0.0546809
R7103 avdd.n5897 avdd.n5890 0.0546809
R7104 avdd.n6113 avdd.n6106 0.0546809
R7105 avdd.n6329 avdd.n6322 0.0546809
R7106 avdd.n6545 avdd.n6538 0.0546809
R7107 avdd.n6761 avdd.n6754 0.0546809
R7108 avdd.n6977 avdd.n6970 0.0546809
R7109 avdd.n7193 avdd.n7186 0.0546809
R7110 avdd.n7849 avdd.n7848 0.0546809
R7111 avdd.n10107 avdd.n10106 0.0546809
R7112 avdd.n10340 avdd.n10339 0.0546809
R7113 avdd.n10442 avdd.n10441 0.0546809
R7114 avdd.n10544 avdd.n10543 0.0546809
R7115 avdd.n10646 avdd.n10645 0.0546809
R7116 avdd.n10748 avdd.n10747 0.0546809
R7117 avdd.n10850 avdd.n10849 0.0546809
R7118 avdd.n10952 avdd.n10951 0.0546809
R7119 avdd.n11054 avdd.n11053 0.0546809
R7120 avdd.n11156 avdd.n11155 0.0546809
R7121 avdd.n11258 avdd.n11257 0.0546809
R7122 avdd.n8871 avdd.n8870 0.0546809
R7123 avdd.n8785 avdd.n8784 0.0546809
R7124 avdd.n8699 avdd.n8698 0.0546809
R7125 avdd.n8613 avdd.n8612 0.0546809
R7126 avdd.n8527 avdd.n8526 0.0546809
R7127 avdd.n8441 avdd.n8440 0.0546809
R7128 avdd.n8355 avdd.n8354 0.0546809
R7129 avdd.n8269 avdd.n8268 0.0546809
R7130 avdd.n8183 avdd.n8182 0.0546809
R7131 avdd.n8097 avdd.n8096 0.0546809
R7132 avdd.n8011 avdd.n8010 0.0546809
R7133 avdd.n7925 avdd.n7924 0.0546809
R7134 avdd.n2307 avdd.n2306 0.0543839
R7135 avdd.n2092 avdd.n1872 0.0543839
R7136 avdd.n3167 avdd.n3166 0.0541072
R7137 avdd.n2952 avdd.n2951 0.0541072
R7138 avdd.n2737 avdd.n2736 0.0541072
R7139 avdd.n2522 avdd.n2521 0.0541072
R7140 avdd.n1955 avdd.n1952 0.0539091
R7141 avdd.n1954 avdd.n1953 0.0539091
R7142 avdd.n2215 avdd.n2209 0.0539091
R7143 avdd.n2214 avdd.n2213 0.0539091
R7144 avdd.n2430 avdd.n2424 0.0539091
R7145 avdd.n2429 avdd.n2428 0.0539091
R7146 avdd.n2645 avdd.n2639 0.0539091
R7147 avdd.n2644 avdd.n2643 0.0539091
R7148 avdd.n2860 avdd.n2854 0.0539091
R7149 avdd.n2859 avdd.n2858 0.0539091
R7150 avdd.n3075 avdd.n3069 0.0539091
R7151 avdd.n3074 avdd.n3073 0.0539091
R7152 avdd.n3245 avdd.n3242 0.0539091
R7153 avdd.n3244 avdd.n3243 0.0539091
R7154 avdd.n3460 avdd.n3457 0.0539091
R7155 avdd.n3459 avdd.n3458 0.0539091
R7156 avdd.n3675 avdd.n3672 0.0539091
R7157 avdd.n3674 avdd.n3673 0.0539091
R7158 avdd.n3890 avdd.n3887 0.0539091
R7159 avdd.n3889 avdd.n3888 0.0539091
R7160 avdd.n4105 avdd.n4102 0.0539091
R7161 avdd.n4104 avdd.n4103 0.0539091
R7162 avdd.n4320 avdd.n4317 0.0539091
R7163 avdd.n4319 avdd.n4318 0.0539091
R7164 avdd.n4937 avdd.n4931 0.0539091
R7165 avdd.n4936 avdd.n4935 0.0539091
R7166 avdd.n5153 avdd.n5147 0.0539091
R7167 avdd.n5152 avdd.n5151 0.0539091
R7168 avdd.n5369 avdd.n5363 0.0539091
R7169 avdd.n5368 avdd.n5367 0.0539091
R7170 avdd.n5585 avdd.n5579 0.0539091
R7171 avdd.n5584 avdd.n5583 0.0539091
R7172 avdd.n5801 avdd.n5795 0.0539091
R7173 avdd.n5800 avdd.n5799 0.0539091
R7174 avdd.n6017 avdd.n6011 0.0539091
R7175 avdd.n6016 avdd.n6015 0.0539091
R7176 avdd.n6233 avdd.n6227 0.0539091
R7177 avdd.n6232 avdd.n6231 0.0539091
R7178 avdd.n6449 avdd.n6443 0.0539091
R7179 avdd.n6448 avdd.n6447 0.0539091
R7180 avdd.n6665 avdd.n6659 0.0539091
R7181 avdd.n6664 avdd.n6663 0.0539091
R7182 avdd.n6881 avdd.n6875 0.0539091
R7183 avdd.n6880 avdd.n6879 0.0539091
R7184 avdd.n7097 avdd.n7091 0.0539091
R7185 avdd.n7096 avdd.n7095 0.0539091
R7186 avdd.n7313 avdd.n7307 0.0539091
R7187 avdd.n7312 avdd.n7311 0.0539091
R7188 avdd.n7647 avdd.n7646 0.0539091
R7189 avdd.n7683 avdd.n7682 0.0539091
R7190 avdd.n10124 avdd.n10123 0.0539091
R7191 avdd.n10162 avdd.n10161 0.0539091
R7192 avdd.n9925 avdd.n9924 0.0539091
R7193 avdd.n9946 avdd.n9945 0.0539091
R7194 avdd.n9811 avdd.n9810 0.0539091
R7195 avdd.n9832 avdd.n9831 0.0539091
R7196 avdd.n9697 avdd.n9696 0.0539091
R7197 avdd.n9718 avdd.n9717 0.0539091
R7198 avdd.n9583 avdd.n9582 0.0539091
R7199 avdd.n9605 avdd.n9604 0.0539091
R7200 avdd.n9469 avdd.n9468 0.0539091
R7201 avdd.n9490 avdd.n9489 0.0539091
R7202 avdd.n9355 avdd.n9354 0.0539091
R7203 avdd.n9376 avdd.n9375 0.0539091
R7204 avdd.n9241 avdd.n9240 0.0539091
R7205 avdd.n9262 avdd.n9261 0.0539091
R7206 avdd.n9127 avdd.n9126 0.0539091
R7207 avdd.n9148 avdd.n9147 0.0539091
R7208 avdd.n9013 avdd.n9012 0.0539091
R7209 avdd.n9034 avdd.n9033 0.0539091
R7210 avdd.n8899 avdd.n8898 0.0539091
R7211 avdd.n8920 avdd.n8919 0.0539091
R7212 avdd.n68 avdd.n67 0.0539091
R7213 avdd.n166 avdd.n165 0.0539091
R7214 avdd.n198 avdd.n197 0.0539091
R7215 avdd.n296 avdd.n295 0.0539091
R7216 avdd.n328 avdd.n327 0.0539091
R7217 avdd.n426 avdd.n425 0.0539091
R7218 avdd.n458 avdd.n457 0.0539091
R7219 avdd.n556 avdd.n555 0.0539091
R7220 avdd.n588 avdd.n587 0.0539091
R7221 avdd.n686 avdd.n685 0.0539091
R7222 avdd.n718 avdd.n717 0.0539091
R7223 avdd.n816 avdd.n815 0.0539091
R7224 avdd.n848 avdd.n847 0.0539091
R7225 avdd.n946 avdd.n945 0.0539091
R7226 avdd.n978 avdd.n977 0.0539091
R7227 avdd.n1076 avdd.n1075 0.0539091
R7228 avdd.n1108 avdd.n1107 0.0539091
R7229 avdd.n1206 avdd.n1205 0.0539091
R7230 avdd.n1238 avdd.n1237 0.0539091
R7231 avdd.n1336 avdd.n1335 0.0539091
R7232 avdd.n1368 avdd.n1367 0.0539091
R7233 avdd.n1466 avdd.n1465 0.0539091
R7234 avdd.n1498 avdd.n1497 0.0539091
R7235 avdd.n1596 avdd.n1595 0.0539091
R7236 avdd.n4027 avdd.n3813 0.0538333
R7237 avdd.n3812 avdd.n3598 0.0538333
R7238 avdd.n3597 avdd.n3383 0.0538333
R7239 avdd.n3382 avdd.n3168 0.0538333
R7240 avdd.n7444 avdd.n7442 0.0536084
R7241 avdd.n7483 avdd.n7481 0.0536084
R7242 avdd.n7543 avdd.n7541 0.0536084
R7243 avdd.n7583 avdd.n7581 0.0536084
R7244 avdd.n4457 avdd.n4243 0.0535623
R7245 avdd.n4242 avdd.n4028 0.0535623
R7246 avdd.n7400 avdd.n7185 0.0534278
R7247 avdd.n7184 avdd.n6969 0.0534278
R7248 avdd.n6968 avdd.n6753 0.0531608
R7249 avdd.n6752 avdd.n6537 0.0531608
R7250 avdd.n6536 avdd.n6321 0.0531608
R7251 avdd.n6320 avdd.n6105 0.0531608
R7252 avdd.n6104 avdd.n5889 0.0528965
R7253 avdd.n5888 avdd.n5673 0.0528965
R7254 avdd.n5672 avdd.n5457 0.0528965
R7255 avdd.n5456 avdd.n5241 0.0528965
R7256 avdd.n5240 avdd.n5025 0.0526348
R7257 avdd.n5024 avdd.n4809 0.0526348
R7258 avdd.n2034 avdd.n2006 0.0526204
R7259 avdd.n2273 avdd.n2272 0.0526204
R7260 avdd.n2488 avdd.n2487 0.0526204
R7261 avdd.n2703 avdd.n2702 0.0526204
R7262 avdd.n2918 avdd.n2917 0.0526204
R7263 avdd.n3133 avdd.n3132 0.0526204
R7264 avdd.n3304 avdd.n3303 0.0526204
R7265 avdd.n3519 avdd.n3518 0.0526204
R7266 avdd.n3734 avdd.n3733 0.0526204
R7267 avdd.n3949 avdd.n3948 0.0526204
R7268 avdd.n4164 avdd.n4163 0.0526204
R7269 avdd.n4379 avdd.n4378 0.0526204
R7270 avdd.n7831 avdd.n7830 0.0526204
R7271 avdd.n10089 avdd.n10088 0.0526204
R7272 avdd.n8852 avdd.n8851 0.0526204
R7273 avdd.n8766 avdd.n8765 0.0526204
R7274 avdd.n8680 avdd.n8679 0.0526204
R7275 avdd.n8594 avdd.n8593 0.0526204
R7276 avdd.n8508 avdd.n8507 0.0526204
R7277 avdd.n8422 avdd.n8421 0.0526204
R7278 avdd.n8336 avdd.n8335 0.0526204
R7279 avdd.n8250 avdd.n8249 0.0526204
R7280 avdd.n8164 avdd.n8163 0.0526204
R7281 avdd.n8078 avdd.n8077 0.0526204
R7282 avdd.n7992 avdd.n7991 0.0526204
R7283 avdd.n7906 avdd.n7905 0.0526204
R7284 avdd.n1992 avdd.n1981 0.0524848
R7285 avdd.n1991 avdd.n1990 0.0524848
R7286 avdd.n2255 avdd.n2252 0.0524848
R7287 avdd.n2254 avdd.n2253 0.0524848
R7288 avdd.n2470 avdd.n2467 0.0524848
R7289 avdd.n2469 avdd.n2468 0.0524848
R7290 avdd.n2685 avdd.n2682 0.0524848
R7291 avdd.n2684 avdd.n2683 0.0524848
R7292 avdd.n2900 avdd.n2897 0.0524848
R7293 avdd.n2899 avdd.n2898 0.0524848
R7294 avdd.n3115 avdd.n3112 0.0524848
R7295 avdd.n3114 avdd.n3113 0.0524848
R7296 avdd.n3282 avdd.n3271 0.0524848
R7297 avdd.n3281 avdd.n3280 0.0524848
R7298 avdd.n3497 avdd.n3486 0.0524848
R7299 avdd.n3496 avdd.n3495 0.0524848
R7300 avdd.n3712 avdd.n3701 0.0524848
R7301 avdd.n3711 avdd.n3710 0.0524848
R7302 avdd.n3927 avdd.n3916 0.0524848
R7303 avdd.n3926 avdd.n3925 0.0524848
R7304 avdd.n4142 avdd.n4131 0.0524848
R7305 avdd.n4141 avdd.n4140 0.0524848
R7306 avdd.n4357 avdd.n4346 0.0524848
R7307 avdd.n4356 avdd.n4355 0.0524848
R7308 avdd.n4977 avdd.n4974 0.0524848
R7309 avdd.n4976 avdd.n4975 0.0524848
R7310 avdd.n5193 avdd.n5190 0.0524848
R7311 avdd.n5192 avdd.n5191 0.0524848
R7312 avdd.n5409 avdd.n5406 0.0524848
R7313 avdd.n5408 avdd.n5407 0.0524848
R7314 avdd.n5625 avdd.n5622 0.0524848
R7315 avdd.n5624 avdd.n5623 0.0524848
R7316 avdd.n5841 avdd.n5838 0.0524848
R7317 avdd.n5840 avdd.n5839 0.0524848
R7318 avdd.n6057 avdd.n6054 0.0524848
R7319 avdd.n6056 avdd.n6055 0.0524848
R7320 avdd.n6273 avdd.n6270 0.0524848
R7321 avdd.n6272 avdd.n6271 0.0524848
R7322 avdd.n6489 avdd.n6486 0.0524848
R7323 avdd.n6488 avdd.n6487 0.0524848
R7324 avdd.n6705 avdd.n6702 0.0524848
R7325 avdd.n6704 avdd.n6703 0.0524848
R7326 avdd.n6921 avdd.n6918 0.0524848
R7327 avdd.n6920 avdd.n6919 0.0524848
R7328 avdd.n7137 avdd.n7134 0.0524848
R7329 avdd.n7136 avdd.n7135 0.0524848
R7330 avdd.n7353 avdd.n7350 0.0524848
R7331 avdd.n7352 avdd.n7351 0.0524848
R7332 avdd.n7775 avdd.n7774 0.0524848
R7333 avdd.n7811 avdd.n7810 0.0524848
R7334 avdd.n10035 avdd.n10034 0.0524848
R7335 avdd.n10069 avdd.n10068 0.0524848
R7336 avdd.n10251 avdd.n10250 0.0524848
R7337 avdd.n10301 avdd.n10300 0.0524848
R7338 avdd.n10353 avdd.n10352 0.0524848
R7339 avdd.n10403 avdd.n10402 0.0524848
R7340 avdd.n10455 avdd.n10454 0.0524848
R7341 avdd.n10505 avdd.n10504 0.0524848
R7342 avdd.n10557 avdd.n10556 0.0524848
R7343 avdd.n10607 avdd.n10606 0.0524848
R7344 avdd.n10659 avdd.n10658 0.0524848
R7345 avdd.n10709 avdd.n10708 0.0524848
R7346 avdd.n10761 avdd.n10760 0.0524848
R7347 avdd.n10811 avdd.n10810 0.0524848
R7348 avdd.n10863 avdd.n10862 0.0524848
R7349 avdd.n10913 avdd.n10912 0.0524848
R7350 avdd.n10965 avdd.n10964 0.0524848
R7351 avdd.n11015 avdd.n11014 0.0524848
R7352 avdd.n11067 avdd.n11066 0.0524848
R7353 avdd.n11117 avdd.n11116 0.0524848
R7354 avdd.n11169 avdd.n11168 0.0524848
R7355 avdd.n11219 avdd.n11218 0.0524848
R7356 avdd.n8878 avdd.n8877 0.0524848
R7357 avdd.n8832 avdd.n8831 0.0524848
R7358 avdd.n8792 avdd.n8791 0.0524848
R7359 avdd.n8746 avdd.n8745 0.0524848
R7360 avdd.n8706 avdd.n8705 0.0524848
R7361 avdd.n8660 avdd.n8659 0.0524848
R7362 avdd.n8620 avdd.n8619 0.0524848
R7363 avdd.n8574 avdd.n8573 0.0524848
R7364 avdd.n8534 avdd.n8533 0.0524848
R7365 avdd.n8488 avdd.n8487 0.0524848
R7366 avdd.n8448 avdd.n8447 0.0524848
R7367 avdd.n8402 avdd.n8401 0.0524848
R7368 avdd.n8362 avdd.n8361 0.0524848
R7369 avdd.n8316 avdd.n8315 0.0524848
R7370 avdd.n8276 avdd.n8275 0.0524848
R7371 avdd.n8230 avdd.n8229 0.0524848
R7372 avdd.n8190 avdd.n8189 0.0524848
R7373 avdd.n8144 avdd.n8143 0.0524848
R7374 avdd.n8104 avdd.n8103 0.0524848
R7375 avdd.n8058 avdd.n8057 0.0524848
R7376 avdd.n8018 avdd.n8017 0.0524848
R7377 avdd.n7972 avdd.n7971 0.0524848
R7378 avdd.n7932 avdd.n7931 0.0524848
R7379 avdd.n7886 avdd.n7885 0.0524848
R7380 avdd avdd.n7430 0.0512812
R7381 avdd avdd.n7511 0.0512812
R7382 avdd avdd.n7412 0.0512812
R7383 avdd avdd.n7611 0.0512812
R7384 avdd.n1699 avdd 0.0512812
R7385 avdd.n1735 avdd 0.0512812
R7386 avdd.n1789 avdd 0.0512812
R7387 avdd.n1825 avdd 0.0512812
R7388 avdd.n2070 avdd.n2069 0.0510606
R7389 avdd.n2229 avdd.n2228 0.0510606
R7390 avdd.n2444 avdd.n2443 0.0510606
R7391 avdd.n2659 avdd.n2658 0.0510606
R7392 avdd.n2874 avdd.n2873 0.0510606
R7393 avdd.n3089 avdd.n3088 0.0510606
R7394 avdd.n3359 avdd.n3358 0.0510606
R7395 avdd.n3574 avdd.n3573 0.0510606
R7396 avdd.n3789 avdd.n3788 0.0510606
R7397 avdd.n4004 avdd.n4003 0.0510606
R7398 avdd.n4219 avdd.n4218 0.0510606
R7399 avdd.n4434 avdd.n4433 0.0510606
R7400 avdd.n4951 avdd.n4950 0.0510606
R7401 avdd.n5167 avdd.n5166 0.0510606
R7402 avdd.n5383 avdd.n5382 0.0510606
R7403 avdd.n5599 avdd.n5598 0.0510606
R7404 avdd.n5815 avdd.n5814 0.0510606
R7405 avdd.n6031 avdd.n6030 0.0510606
R7406 avdd.n6247 avdd.n6246 0.0510606
R7407 avdd.n6463 avdd.n6462 0.0510606
R7408 avdd.n6679 avdd.n6678 0.0510606
R7409 avdd.n6895 avdd.n6894 0.0510606
R7410 avdd.n7111 avdd.n7110 0.0510606
R7411 avdd.n7327 avdd.n7326 0.0510606
R7412 avdd.n7643 avdd.n7642 0.0510606
R7413 avdd.n10120 avdd.n10119 0.0510606
R7414 avdd.n9921 avdd.n9920 0.0510606
R7415 avdd.n9807 avdd.n9806 0.0510606
R7416 avdd.n9693 avdd.n9692 0.0510606
R7417 avdd.n9579 avdd.n9578 0.0510606
R7418 avdd.n9465 avdd.n9464 0.0510606
R7419 avdd.n9351 avdd.n9350 0.0510606
R7420 avdd.n9237 avdd.n9236 0.0510606
R7421 avdd.n9123 avdd.n9122 0.0510606
R7422 avdd.n9009 avdd.n9008 0.0510606
R7423 avdd.n8895 avdd.n8894 0.0510606
R7424 avdd.n64 avdd.n63 0.0510606
R7425 avdd.n194 avdd.n193 0.0510606
R7426 avdd.n324 avdd.n323 0.0510606
R7427 avdd.n454 avdd.n453 0.0510606
R7428 avdd.n584 avdd.n583 0.0510606
R7429 avdd.n714 avdd.n713 0.0510606
R7430 avdd.n844 avdd.n843 0.0510606
R7431 avdd.n974 avdd.n973 0.0510606
R7432 avdd.n1104 avdd.n1103 0.0510606
R7433 avdd.n1234 avdd.n1233 0.0510606
R7434 avdd.n1364 avdd.n1363 0.0510606
R7435 avdd.n1494 avdd.n1493 0.0510606
R7436 avdd.n2056 avdd.n1972 0.0496364
R7437 avdd.n1926 avdd.n1925 0.0496364
R7438 avdd.n2251 avdd.n2250 0.0496364
R7439 avdd.n2180 avdd.n2179 0.0496364
R7440 avdd.n2466 avdd.n2465 0.0496364
R7441 avdd.n2395 avdd.n2394 0.0496364
R7442 avdd.n2681 avdd.n2680 0.0496364
R7443 avdd.n2610 avdd.n2609 0.0496364
R7444 avdd.n2896 avdd.n2895 0.0496364
R7445 avdd.n2825 avdd.n2824 0.0496364
R7446 avdd.n3111 avdd.n3110 0.0496364
R7447 avdd.n3040 avdd.n3039 0.0496364
R7448 avdd.n3345 avdd.n3262 0.0496364
R7449 avdd.n3216 avdd.n3215 0.0496364
R7450 avdd.n3560 avdd.n3477 0.0496364
R7451 avdd.n3431 avdd.n3430 0.0496364
R7452 avdd.n3775 avdd.n3692 0.0496364
R7453 avdd.n3646 avdd.n3645 0.0496364
R7454 avdd.n3990 avdd.n3907 0.0496364
R7455 avdd.n3861 avdd.n3860 0.0496364
R7456 avdd.n4205 avdd.n4122 0.0496364
R7457 avdd.n4076 avdd.n4075 0.0496364
R7458 avdd.n4420 avdd.n4337 0.0496364
R7459 avdd.n4291 avdd.n4290 0.0496364
R7460 avdd.n4973 avdd.n4972 0.0496364
R7461 avdd.n4902 avdd.n4901 0.0496364
R7462 avdd.n5189 avdd.n5188 0.0496364
R7463 avdd.n5118 avdd.n5117 0.0496364
R7464 avdd.n5405 avdd.n5404 0.0496364
R7465 avdd.n5334 avdd.n5333 0.0496364
R7466 avdd.n5621 avdd.n5620 0.0496364
R7467 avdd.n5550 avdd.n5549 0.0496364
R7468 avdd.n5837 avdd.n5836 0.0496364
R7469 avdd.n5766 avdd.n5765 0.0496364
R7470 avdd.n6053 avdd.n6052 0.0496364
R7471 avdd.n5982 avdd.n5981 0.0496364
R7472 avdd.n6269 avdd.n6268 0.0496364
R7473 avdd.n6198 avdd.n6197 0.0496364
R7474 avdd.n6485 avdd.n6484 0.0496364
R7475 avdd.n6414 avdd.n6413 0.0496364
R7476 avdd.n6701 avdd.n6700 0.0496364
R7477 avdd.n6630 avdd.n6629 0.0496364
R7478 avdd.n6917 avdd.n6916 0.0496364
R7479 avdd.n6846 avdd.n6845 0.0496364
R7480 avdd.n7133 avdd.n7132 0.0496364
R7481 avdd.n7062 avdd.n7061 0.0496364
R7482 avdd.n7349 avdd.n7348 0.0496364
R7483 avdd.n7278 avdd.n7277 0.0496364
R7484 avdd.n7771 avdd.n7770 0.0496364
R7485 avdd.n7759 avdd.n7758 0.0496364
R7486 avdd.n10031 avdd.n10030 0.0496364
R7487 avdd.n10238 avdd.n10237 0.0496364
R7488 avdd.n10247 avdd.n10246 0.0496364
R7489 avdd.n9992 avdd.n9991 0.0496364
R7490 avdd.n10349 avdd.n10348 0.0496364
R7491 avdd.n9878 avdd.n9877 0.0496364
R7492 avdd.n10451 avdd.n10450 0.0496364
R7493 avdd.n9764 avdd.n9763 0.0496364
R7494 avdd.n10553 avdd.n10552 0.0496364
R7495 avdd.n9651 avdd.n9650 0.0496364
R7496 avdd.n10655 avdd.n10654 0.0496364
R7497 avdd.n9536 avdd.n9535 0.0496364
R7498 avdd.n10757 avdd.n10756 0.0496364
R7499 avdd.n9422 avdd.n9421 0.0496364
R7500 avdd.n10859 avdd.n10858 0.0496364
R7501 avdd.n9308 avdd.n9307 0.0496364
R7502 avdd.n10961 avdd.n10960 0.0496364
R7503 avdd.n9194 avdd.n9193 0.0496364
R7504 avdd.n11063 avdd.n11062 0.0496364
R7505 avdd.n9080 avdd.n9079 0.0496364
R7506 avdd.n11165 avdd.n11164 0.0496364
R7507 avdd.n8966 avdd.n8965 0.0496364
R7508 avdd.n8874 avdd.n8873 0.0496364
R7509 avdd.n92 avdd.n91 0.0496364
R7510 avdd.n8788 avdd.n8787 0.0496364
R7511 avdd.n222 avdd.n221 0.0496364
R7512 avdd.n8702 avdd.n8701 0.0496364
R7513 avdd.n352 avdd.n351 0.0496364
R7514 avdd.n8616 avdd.n8615 0.0496364
R7515 avdd.n482 avdd.n481 0.0496364
R7516 avdd.n8530 avdd.n8529 0.0496364
R7517 avdd.n612 avdd.n611 0.0496364
R7518 avdd.n8444 avdd.n8443 0.0496364
R7519 avdd.n742 avdd.n741 0.0496364
R7520 avdd.n8358 avdd.n8357 0.0496364
R7521 avdd.n872 avdd.n871 0.0496364
R7522 avdd.n8272 avdd.n8271 0.0496364
R7523 avdd.n1002 avdd.n1001 0.0496364
R7524 avdd.n8186 avdd.n8185 0.0496364
R7525 avdd.n1132 avdd.n1131 0.0496364
R7526 avdd.n8100 avdd.n8099 0.0496364
R7527 avdd.n1262 avdd.n1261 0.0496364
R7528 avdd.n8014 avdd.n8013 0.0496364
R7529 avdd.n1392 avdd.n1391 0.0496364
R7530 avdd.n7928 avdd.n7927 0.0496364
R7531 avdd.n1522 avdd.n1521 0.0496364
R7532 avdd.n10345 avdd.n10244 0.0495971
R7533 avdd.n7941 avdd.n7856 0.049469
R7534 avdd.n10651 avdd.n10550 0.0494659
R7535 avdd.n10447 avdd.n10346 0.0494659
R7536 avdd.n10753 avdd.n10652 0.0494046
R7537 avdd.n11059 avdd.n10958 0.0492748
R7538 avdd.n10957 avdd.n10856 0.0492748
R7539 avdd.n10855 avdd.n10754 0.0492748
R7540 avdd.n11161 avdd.n11060 0.0492142
R7541 avdd.n10549 avdd.n10448 0.0491154
R7542 avdd.n11263 avdd.n11162 0.0490859
R7543 avdd.n2035 avdd.n2031 0.0482121
R7544 avdd.n2034 avdd.n2033 0.0482121
R7545 avdd.n2275 avdd.n2274 0.0482121
R7546 avdd.n2273 avdd.n2106 0.0482121
R7547 avdd.n2490 avdd.n2489 0.0482121
R7548 avdd.n2488 avdd.n2321 0.0482121
R7549 avdd.n2705 avdd.n2704 0.0482121
R7550 avdd.n2703 avdd.n2536 0.0482121
R7551 avdd.n2920 avdd.n2919 0.0482121
R7552 avdd.n2918 avdd.n2751 0.0482121
R7553 avdd.n3135 avdd.n3134 0.0482121
R7554 avdd.n3133 avdd.n2966 0.0482121
R7555 avdd.n3301 avdd.n3295 0.0482121
R7556 avdd.n3303 avdd.n3302 0.0482121
R7557 avdd.n3516 avdd.n3510 0.0482121
R7558 avdd.n3518 avdd.n3517 0.0482121
R7559 avdd.n3731 avdd.n3725 0.0482121
R7560 avdd.n3733 avdd.n3732 0.0482121
R7561 avdd.n3946 avdd.n3940 0.0482121
R7562 avdd.n3948 avdd.n3947 0.0482121
R7563 avdd.n4161 avdd.n4155 0.0482121
R7564 avdd.n4163 avdd.n4162 0.0482121
R7565 avdd.n4376 avdd.n4370 0.0482121
R7566 avdd.n4378 avdd.n4377 0.0482121
R7567 avdd.n4994 avdd.n4813 0.0482121
R7568 avdd.n4828 avdd.n4827 0.0482121
R7569 avdd.n5210 avdd.n5029 0.0482121
R7570 avdd.n5044 avdd.n5043 0.0482121
R7571 avdd.n5426 avdd.n5245 0.0482121
R7572 avdd.n5260 avdd.n5259 0.0482121
R7573 avdd.n5642 avdd.n5461 0.0482121
R7574 avdd.n5476 avdd.n5475 0.0482121
R7575 avdd.n5858 avdd.n5677 0.0482121
R7576 avdd.n5692 avdd.n5691 0.0482121
R7577 avdd.n6074 avdd.n5893 0.0482121
R7578 avdd.n5908 avdd.n5907 0.0482121
R7579 avdd.n6290 avdd.n6109 0.0482121
R7580 avdd.n6124 avdd.n6123 0.0482121
R7581 avdd.n6506 avdd.n6325 0.0482121
R7582 avdd.n6340 avdd.n6339 0.0482121
R7583 avdd.n6722 avdd.n6541 0.0482121
R7584 avdd.n6556 avdd.n6555 0.0482121
R7585 avdd.n6938 avdd.n6757 0.0482121
R7586 avdd.n6772 avdd.n6771 0.0482121
R7587 avdd.n7154 avdd.n6973 0.0482121
R7588 avdd.n6988 avdd.n6987 0.0482121
R7589 avdd.n7370 avdd.n7189 0.0482121
R7590 avdd.n7204 avdd.n7203 0.0482121
R7591 avdd.n7781 avdd.n7780 0.0482121
R7592 avdd.n7830 avdd.n7829 0.0482121
R7593 avdd.n10041 avdd.n10040 0.0482121
R7594 avdd.n10088 avdd.n10087 0.0482121
R7595 avdd.n10257 avdd.n10256 0.0482121
R7596 avdd.n10320 avdd.n10319 0.0482121
R7597 avdd.n10359 avdd.n10358 0.0482121
R7598 avdd.n10422 avdd.n10421 0.0482121
R7599 avdd.n10461 avdd.n10460 0.0482121
R7600 avdd.n10524 avdd.n10523 0.0482121
R7601 avdd.n10563 avdd.n10562 0.0482121
R7602 avdd.n10626 avdd.n10625 0.0482121
R7603 avdd.n10665 avdd.n10664 0.0482121
R7604 avdd.n10728 avdd.n10727 0.0482121
R7605 avdd.n10767 avdd.n10766 0.0482121
R7606 avdd.n10830 avdd.n10829 0.0482121
R7607 avdd.n10869 avdd.n10868 0.0482121
R7608 avdd.n10932 avdd.n10931 0.0482121
R7609 avdd.n10971 avdd.n10970 0.0482121
R7610 avdd.n11034 avdd.n11033 0.0482121
R7611 avdd.n11073 avdd.n11072 0.0482121
R7612 avdd.n11136 avdd.n11135 0.0482121
R7613 avdd.n11175 avdd.n11174 0.0482121
R7614 avdd.n11238 avdd.n11237 0.0482121
R7615 avdd.n8884 avdd.n8883 0.0482121
R7616 avdd.n8851 avdd.n8850 0.0482121
R7617 avdd.n8798 avdd.n8797 0.0482121
R7618 avdd.n8765 avdd.n8764 0.0482121
R7619 avdd.n8712 avdd.n8711 0.0482121
R7620 avdd.n8679 avdd.n8678 0.0482121
R7621 avdd.n8626 avdd.n8625 0.0482121
R7622 avdd.n8593 avdd.n8592 0.0482121
R7623 avdd.n8540 avdd.n8539 0.0482121
R7624 avdd.n8507 avdd.n8506 0.0482121
R7625 avdd.n8454 avdd.n8453 0.0482121
R7626 avdd.n8421 avdd.n8420 0.0482121
R7627 avdd.n8368 avdd.n8367 0.0482121
R7628 avdd.n8335 avdd.n8334 0.0482121
R7629 avdd.n8282 avdd.n8281 0.0482121
R7630 avdd.n8249 avdd.n8248 0.0482121
R7631 avdd.n8196 avdd.n8195 0.0482121
R7632 avdd.n8163 avdd.n8162 0.0482121
R7633 avdd.n8110 avdd.n8109 0.0482121
R7634 avdd.n8077 avdd.n8076 0.0482121
R7635 avdd.n8024 avdd.n8023 0.0482121
R7636 avdd.n7991 avdd.n7990 0.0482121
R7637 avdd.n7938 avdd.n7937 0.0482121
R7638 avdd.n7905 avdd.n7904 0.0482121
R7639 avdd.n8027 avdd.n7942 0.0481718
R7640 avdd.n8113 avdd.n8028 0.0481151
R7641 avdd.n8199 avdd.n8114 0.0479949
R7642 avdd.n8371 avdd.n8286 0.0479949
R7643 avdd.n8457 avdd.n8372 0.0479387
R7644 avdd.n8543 avdd.n8458 0.0478198
R7645 avdd.n8629 avdd.n8544 0.0478198
R7646 avdd.n8715 avdd.n8630 0.0478198
R7647 avdd.n8801 avdd.n8716 0.0477643
R7648 avdd.n8887 avdd.n8802 0.0476467
R7649 avdd.n8285 avdd.n8200 0.0476444
R7650 avdd.n4827 avdd.n4816 0.0467879
R7651 avdd.n5043 avdd.n5032 0.0467879
R7652 avdd.n5259 avdd.n5248 0.0467879
R7653 avdd.n5475 avdd.n5464 0.0467879
R7654 avdd.n5691 avdd.n5680 0.0467879
R7655 avdd.n5907 avdd.n5896 0.0467879
R7656 avdd.n6123 avdd.n6112 0.0467879
R7657 avdd.n6339 avdd.n6328 0.0467879
R7658 avdd.n6555 avdd.n6544 0.0467879
R7659 avdd.n6771 avdd.n6760 0.0467879
R7660 avdd.n6987 avdd.n6976 0.0467879
R7661 avdd.n7203 avdd.n7192 0.0467879
R7662 avdd.n10321 avdd.n10320 0.0467879
R7663 avdd.n10423 avdd.n10422 0.0467879
R7664 avdd.n10525 avdd.n10524 0.0467879
R7665 avdd.n10627 avdd.n10626 0.0467879
R7666 avdd.n10729 avdd.n10728 0.0467879
R7667 avdd.n10831 avdd.n10830 0.0467879
R7668 avdd.n10933 avdd.n10932 0.0467879
R7669 avdd.n11035 avdd.n11034 0.0467879
R7670 avdd.n11137 avdd.n11136 0.0467879
R7671 avdd.n11239 avdd.n11238 0.0467879
R7672 avdd.n2306 avdd.n2092 0.0467261
R7673 avdd.n2521 avdd.n2307 0.0466743
R7674 avdd.n3166 avdd.n2952 0.0465643
R7675 avdd.n2736 avdd.n2522 0.0465643
R7676 avdd.n3168 avdd.n3167 0.046513
R7677 avdd.n3813 avdd.n3812 0.0464042
R7678 avdd.n3598 avdd.n3597 0.0464042
R7679 avdd.n3383 avdd.n3382 0.0464042
R7680 avdd.n4028 avdd.n4027 0.0463534
R7681 avdd.n4243 avdd.n4242 0.0462457
R7682 avdd.n2951 avdd.n2737 0.0462139
R7683 avdd.n7185 avdd.n7184 0.0461671
R7684 avdd.n6969 avdd.n6968 0.046117
R7685 avdd.n6753 avdd.n6752 0.046011
R7686 avdd.n6321 avdd.n6320 0.046011
R7687 avdd.n6105 avdd.n6104 0.0459614
R7688 avdd.n5889 avdd.n5888 0.0458564
R7689 avdd.n5673 avdd.n5672 0.0458564
R7690 avdd.n5457 avdd.n5456 0.0458564
R7691 avdd.n5241 avdd.n5240 0.0458074
R7692 avdd.n5025 avdd.n5024 0.0457034
R7693 avdd.n6537 avdd.n6536 0.0456605
R7694 avdd.n7401 avdd.n7400 0.045234
R7695 avdd.n3324 avdd.n3323 0.0443504
R7696 avdd.n3539 avdd.n3538 0.0443504
R7697 avdd.n3754 avdd.n3753 0.0443504
R7698 avdd.n3969 avdd.n3968 0.0443504
R7699 avdd.n4184 avdd.n4183 0.0443504
R7700 avdd.n4399 avdd.n4398 0.0443504
R7701 avdd.n1988 avdd.n1981 0.0425152
R7702 avdd.n1990 avdd.n1989 0.0425152
R7703 avdd.n2256 avdd.n2255 0.0425152
R7704 avdd.n2254 avdd.n2113 0.0425152
R7705 avdd.n2471 avdd.n2470 0.0425152
R7706 avdd.n2469 avdd.n2328 0.0425152
R7707 avdd.n2686 avdd.n2685 0.0425152
R7708 avdd.n2684 avdd.n2543 0.0425152
R7709 avdd.n2901 avdd.n2900 0.0425152
R7710 avdd.n2899 avdd.n2758 0.0425152
R7711 avdd.n3116 avdd.n3115 0.0425152
R7712 avdd.n3114 avdd.n2973 0.0425152
R7713 avdd.n3278 avdd.n3271 0.0425152
R7714 avdd.n3280 avdd.n3279 0.0425152
R7715 avdd.n3493 avdd.n3486 0.0425152
R7716 avdd.n3495 avdd.n3494 0.0425152
R7717 avdd.n3708 avdd.n3701 0.0425152
R7718 avdd.n3710 avdd.n3709 0.0425152
R7719 avdd.n3923 avdd.n3916 0.0425152
R7720 avdd.n3925 avdd.n3924 0.0425152
R7721 avdd.n4138 avdd.n4131 0.0425152
R7722 avdd.n4140 avdd.n4139 0.0425152
R7723 avdd.n4353 avdd.n4346 0.0425152
R7724 avdd.n4355 avdd.n4354 0.0425152
R7725 avdd.n4978 avdd.n4977 0.0425152
R7726 avdd.n4976 avdd.n4835 0.0425152
R7727 avdd.n5194 avdd.n5193 0.0425152
R7728 avdd.n5192 avdd.n5051 0.0425152
R7729 avdd.n5410 avdd.n5409 0.0425152
R7730 avdd.n5408 avdd.n5267 0.0425152
R7731 avdd.n5626 avdd.n5625 0.0425152
R7732 avdd.n5624 avdd.n5483 0.0425152
R7733 avdd.n5842 avdd.n5841 0.0425152
R7734 avdd.n5840 avdd.n5699 0.0425152
R7735 avdd.n6058 avdd.n6057 0.0425152
R7736 avdd.n6056 avdd.n5915 0.0425152
R7737 avdd.n6274 avdd.n6273 0.0425152
R7738 avdd.n6272 avdd.n6131 0.0425152
R7739 avdd.n6490 avdd.n6489 0.0425152
R7740 avdd.n6488 avdd.n6347 0.0425152
R7741 avdd.n6706 avdd.n6705 0.0425152
R7742 avdd.n6704 avdd.n6563 0.0425152
R7743 avdd.n6922 avdd.n6921 0.0425152
R7744 avdd.n6920 avdd.n6779 0.0425152
R7745 avdd.n7138 avdd.n7137 0.0425152
R7746 avdd.n7136 avdd.n6995 0.0425152
R7747 avdd.n7354 avdd.n7353 0.0425152
R7748 avdd.n7352 avdd.n7211 0.0425152
R7749 avdd.n7774 avdd.n7773 0.0425152
R7750 avdd.n7810 avdd.n7809 0.0425152
R7751 avdd.n10034 avdd.n10033 0.0425152
R7752 avdd.n10068 avdd.n10067 0.0425152
R7753 avdd.n10250 avdd.n10249 0.0425152
R7754 avdd.n10300 avdd.n10299 0.0425152
R7755 avdd.n10352 avdd.n10351 0.0425152
R7756 avdd.n10402 avdd.n10401 0.0425152
R7757 avdd.n10454 avdd.n10453 0.0425152
R7758 avdd.n10504 avdd.n10503 0.0425152
R7759 avdd.n10556 avdd.n10555 0.0425152
R7760 avdd.n10606 avdd.n10605 0.0425152
R7761 avdd.n10658 avdd.n10657 0.0425152
R7762 avdd.n10708 avdd.n10707 0.0425152
R7763 avdd.n10760 avdd.n10759 0.0425152
R7764 avdd.n10810 avdd.n10809 0.0425152
R7765 avdd.n10862 avdd.n10861 0.0425152
R7766 avdd.n10912 avdd.n10911 0.0425152
R7767 avdd.n10964 avdd.n10963 0.0425152
R7768 avdd.n11014 avdd.n11013 0.0425152
R7769 avdd.n11066 avdd.n11065 0.0425152
R7770 avdd.n11116 avdd.n11115 0.0425152
R7771 avdd.n11168 avdd.n11167 0.0425152
R7772 avdd.n11218 avdd.n11217 0.0425152
R7773 avdd.n8877 avdd.n8876 0.0425152
R7774 avdd.n8831 avdd.n8830 0.0425152
R7775 avdd.n8791 avdd.n8790 0.0425152
R7776 avdd.n8745 avdd.n8744 0.0425152
R7777 avdd.n8705 avdd.n8704 0.0425152
R7778 avdd.n8659 avdd.n8658 0.0425152
R7779 avdd.n8619 avdd.n8618 0.0425152
R7780 avdd.n8573 avdd.n8572 0.0425152
R7781 avdd.n8533 avdd.n8532 0.0425152
R7782 avdd.n8487 avdd.n8486 0.0425152
R7783 avdd.n8447 avdd.n8446 0.0425152
R7784 avdd.n8401 avdd.n8400 0.0425152
R7785 avdd.n8361 avdd.n8360 0.0425152
R7786 avdd.n8315 avdd.n8314 0.0425152
R7787 avdd.n8275 avdd.n8274 0.0425152
R7788 avdd.n8229 avdd.n8228 0.0425152
R7789 avdd.n8189 avdd.n8188 0.0425152
R7790 avdd.n8143 avdd.n8142 0.0425152
R7791 avdd.n8103 avdd.n8102 0.0425152
R7792 avdd.n8057 avdd.n8056 0.0425152
R7793 avdd.n8017 avdd.n8016 0.0425152
R7794 avdd.n7971 avdd.n7970 0.0425152
R7795 avdd.n7931 avdd.n7930 0.0425152
R7796 avdd.n7885 avdd.n7884 0.0425152
R7797 avdd.n1816 avdd.n1815 0.0420926
R7798 avdd.n1642 avdd.n1641 0.0420926
R7799 avdd.n1726 avdd.n1725 0.0420926
R7800 avdd.n1678 avdd.n1677 0.0420926
R7801 avdd.n3380 avdd.n3378 0.0417717
R7802 avdd.n3595 avdd.n3593 0.0417717
R7803 avdd.n3810 avdd.n3808 0.0417717
R7804 avdd.n4025 avdd.n4023 0.0417717
R7805 avdd.n4240 avdd.n4238 0.0417717
R7806 avdd.n4455 avdd.n4453 0.0417717
R7807 avdd.n4919 avdd.n4862 0.0417717
R7808 avdd.n5135 avdd.n5078 0.0417717
R7809 avdd.n5351 avdd.n5294 0.0417717
R7810 avdd.n5567 avdd.n5510 0.0417717
R7811 avdd.n5783 avdd.n5726 0.0417717
R7812 avdd.n5999 avdd.n5942 0.0417717
R7813 avdd.n6215 avdd.n6158 0.0417717
R7814 avdd.n6431 avdd.n6374 0.0417717
R7815 avdd.n6647 avdd.n6590 0.0417717
R7816 avdd.n6863 avdd.n6806 0.0417717
R7817 avdd.n7079 avdd.n7022 0.0417717
R7818 avdd.n7295 avdd.n7238 0.0417717
R7819 avdd.n10025 avdd.n10023 0.0417717
R7820 avdd.n9911 avdd.n9909 0.0417717
R7821 avdd.n9797 avdd.n9795 0.0417717
R7822 avdd.n9683 avdd.n9682 0.0417717
R7823 avdd.n9569 avdd.n9567 0.0417717
R7824 avdd.n9455 avdd.n9453 0.0417717
R7825 avdd.n9341 avdd.n9339 0.0417717
R7826 avdd.n9227 avdd.n9225 0.0417717
R7827 avdd.n9113 avdd.n9111 0.0417717
R7828 avdd.n8999 avdd.n8997 0.0417717
R7829 avdd.n1817 avdd.n1816 0.0416202
R7830 avdd.n1643 avdd.n1642 0.0416202
R7831 avdd.n1727 avdd.n1726 0.0416202
R7832 avdd.n1679 avdd.n1678 0.0416202
R7833 avdd.n1956 avdd.n1955 0.0410909
R7834 avdd.n1954 avdd.n1949 0.0410909
R7835 avdd.n2211 avdd.n2209 0.0410909
R7836 avdd.n2213 avdd.n2212 0.0410909
R7837 avdd.n2426 avdd.n2424 0.0410909
R7838 avdd.n2428 avdd.n2427 0.0410909
R7839 avdd.n2641 avdd.n2639 0.0410909
R7840 avdd.n2643 avdd.n2642 0.0410909
R7841 avdd.n2856 avdd.n2854 0.0410909
R7842 avdd.n2858 avdd.n2857 0.0410909
R7843 avdd.n3071 avdd.n3069 0.0410909
R7844 avdd.n3073 avdd.n3072 0.0410909
R7845 avdd.n3246 avdd.n3245 0.0410909
R7846 avdd.n3244 avdd.n3239 0.0410909
R7847 avdd.n3461 avdd.n3460 0.0410909
R7848 avdd.n3459 avdd.n3454 0.0410909
R7849 avdd.n3676 avdd.n3675 0.0410909
R7850 avdd.n3674 avdd.n3669 0.0410909
R7851 avdd.n3891 avdd.n3890 0.0410909
R7852 avdd.n3889 avdd.n3884 0.0410909
R7853 avdd.n4106 avdd.n4105 0.0410909
R7854 avdd.n4104 avdd.n4099 0.0410909
R7855 avdd.n4321 avdd.n4320 0.0410909
R7856 avdd.n4319 avdd.n4314 0.0410909
R7857 avdd.n4933 avdd.n4931 0.0410909
R7858 avdd.n4935 avdd.n4934 0.0410909
R7859 avdd.n5149 avdd.n5147 0.0410909
R7860 avdd.n5151 avdd.n5150 0.0410909
R7861 avdd.n5365 avdd.n5363 0.0410909
R7862 avdd.n5367 avdd.n5366 0.0410909
R7863 avdd.n5581 avdd.n5579 0.0410909
R7864 avdd.n5583 avdd.n5582 0.0410909
R7865 avdd.n5797 avdd.n5795 0.0410909
R7866 avdd.n5799 avdd.n5798 0.0410909
R7867 avdd.n6013 avdd.n6011 0.0410909
R7868 avdd.n6015 avdd.n6014 0.0410909
R7869 avdd.n6229 avdd.n6227 0.0410909
R7870 avdd.n6231 avdd.n6230 0.0410909
R7871 avdd.n6445 avdd.n6443 0.0410909
R7872 avdd.n6447 avdd.n6446 0.0410909
R7873 avdd.n6661 avdd.n6659 0.0410909
R7874 avdd.n6663 avdd.n6662 0.0410909
R7875 avdd.n6877 avdd.n6875 0.0410909
R7876 avdd.n6879 avdd.n6878 0.0410909
R7877 avdd.n7093 avdd.n7091 0.0410909
R7878 avdd.n7095 avdd.n7094 0.0410909
R7879 avdd.n7309 avdd.n7307 0.0410909
R7880 avdd.n7311 avdd.n7310 0.0410909
R7881 avdd.n7646 avdd.n7645 0.0410909
R7882 avdd.n7682 avdd.n7681 0.0410909
R7883 avdd.n10123 avdd.n10122 0.0410909
R7884 avdd.n10161 avdd.n10160 0.0410909
R7885 avdd.n9924 avdd.n9923 0.0410909
R7886 avdd.n9945 avdd.n9944 0.0410909
R7887 avdd.n9810 avdd.n9809 0.0410909
R7888 avdd.n9831 avdd.n9830 0.0410909
R7889 avdd.n9696 avdd.n9695 0.0410909
R7890 avdd.n9717 avdd.n9716 0.0410909
R7891 avdd.n9582 avdd.n9581 0.0410909
R7892 avdd.n9604 avdd.n9603 0.0410909
R7893 avdd.n9468 avdd.n9467 0.0410909
R7894 avdd.n9489 avdd.n9488 0.0410909
R7895 avdd.n9354 avdd.n9353 0.0410909
R7896 avdd.n9375 avdd.n9374 0.0410909
R7897 avdd.n9240 avdd.n9239 0.0410909
R7898 avdd.n9261 avdd.n9260 0.0410909
R7899 avdd.n9126 avdd.n9125 0.0410909
R7900 avdd.n9147 avdd.n9146 0.0410909
R7901 avdd.n9012 avdd.n9011 0.0410909
R7902 avdd.n9033 avdd.n9032 0.0410909
R7903 avdd.n8898 avdd.n8897 0.0410909
R7904 avdd.n8919 avdd.n8918 0.0410909
R7905 avdd.n67 avdd.n66 0.0410909
R7906 avdd.n165 avdd.n164 0.0410909
R7907 avdd.n197 avdd.n196 0.0410909
R7908 avdd.n295 avdd.n294 0.0410909
R7909 avdd.n327 avdd.n326 0.0410909
R7910 avdd.n425 avdd.n424 0.0410909
R7911 avdd.n457 avdd.n456 0.0410909
R7912 avdd.n555 avdd.n554 0.0410909
R7913 avdd.n587 avdd.n586 0.0410909
R7914 avdd.n685 avdd.n684 0.0410909
R7915 avdd.n717 avdd.n716 0.0410909
R7916 avdd.n815 avdd.n814 0.0410909
R7917 avdd.n847 avdd.n846 0.0410909
R7918 avdd.n945 avdd.n944 0.0410909
R7919 avdd.n977 avdd.n976 0.0410909
R7920 avdd.n1075 avdd.n1074 0.0410909
R7921 avdd.n1107 avdd.n1106 0.0410909
R7922 avdd.n1205 avdd.n1204 0.0410909
R7923 avdd.n1237 avdd.n1236 0.0410909
R7924 avdd.n1335 avdd.n1334 0.0410909
R7925 avdd.n1367 avdd.n1366 0.0410909
R7926 avdd.n1465 avdd.n1464 0.0410909
R7927 avdd.n1497 avdd.n1496 0.0410909
R7928 avdd.n1595 avdd.n1594 0.0410909
R7929 avdd.n1895 avdd.n1879 0.0402927
R7930 avdd.n2145 avdd.n2144 0.0402927
R7931 avdd.n2360 avdd.n2359 0.0402927
R7932 avdd.n2575 avdd.n2574 0.0402927
R7933 avdd.n2790 avdd.n2789 0.0402927
R7934 avdd.n3005 avdd.n3004 0.0402927
R7935 avdd.n3185 avdd.n3170 0.0402927
R7936 avdd.n3400 avdd.n3385 0.0402927
R7937 avdd.n3615 avdd.n3600 0.0402927
R7938 avdd.n3830 avdd.n3815 0.0402927
R7939 avdd.n4045 avdd.n4030 0.0402927
R7940 avdd.n4260 avdd.n4245 0.0402927
R7941 avdd.n4917 avdd.n4867 0.0402927
R7942 avdd.n5133 avdd.n5083 0.0402927
R7943 avdd.n5349 avdd.n5299 0.0402927
R7944 avdd.n5565 avdd.n5515 0.0402927
R7945 avdd.n5781 avdd.n5731 0.0402927
R7946 avdd.n5997 avdd.n5947 0.0402927
R7947 avdd.n6213 avdd.n6163 0.0402927
R7948 avdd.n6429 avdd.n6379 0.0402927
R7949 avdd.n6645 avdd.n6595 0.0402927
R7950 avdd.n6861 avdd.n6811 0.0402927
R7951 avdd.n7077 avdd.n7027 0.0402927
R7952 avdd.n7293 avdd.n7243 0.0402927
R7953 avdd.n7722 avdd.n7721 0.0402927
R7954 avdd.n10201 avdd.n10200 0.0402927
R7955 avdd.n10010 avdd.n10009 0.0402927
R7956 avdd.n9896 avdd.n9895 0.0402927
R7957 avdd.n9782 avdd.n9781 0.0402927
R7958 avdd.n9669 avdd.n9668 0.0402927
R7959 avdd.n9554 avdd.n9553 0.0402927
R7960 avdd.n9440 avdd.n9439 0.0402927
R7961 avdd.n9326 avdd.n9325 0.0402927
R7962 avdd.n9212 avdd.n9211 0.0402927
R7963 avdd.n9098 avdd.n9097 0.0402927
R7964 avdd.n8984 avdd.n8983 0.0402927
R7965 avdd.n116 avdd.n115 0.0402927
R7966 avdd.n246 avdd.n245 0.0402927
R7967 avdd.n376 avdd.n375 0.0402927
R7968 avdd.n506 avdd.n505 0.0402927
R7969 avdd.n636 avdd.n635 0.0402927
R7970 avdd.n766 avdd.n765 0.0402927
R7971 avdd.n896 avdd.n895 0.0402927
R7972 avdd.n1026 avdd.n1025 0.0402927
R7973 avdd.n1156 avdd.n1155 0.0402927
R7974 avdd.n1286 avdd.n1285 0.0402927
R7975 avdd.n1416 avdd.n1415 0.0402927
R7976 avdd.n1546 avdd.n1545 0.0402927
R7977 avdd.n1933 avdd.n1889 0.0398017
R7978 avdd.n2076 avdd.n1946 0.0398017
R7979 avdd.n1968 avdd.n1947 0.0398017
R7980 avdd.n2051 avdd.n1974 0.0398017
R7981 avdd.n2049 avdd.n1977 0.0398017
R7982 avdd.n2019 avdd.n2000 0.0398017
R7983 avdd.n2186 avdd.n2136 0.0398017
R7984 avdd.n2220 avdd.n2129 0.0398017
R7985 avdd.n2223 avdd.n2222 0.0398017
R7986 avdd.n2243 avdd.n2110 0.0398017
R7987 avdd.n2262 avdd.n2103 0.0398017
R7988 avdd.n2293 avdd.n2100 0.0398017
R7989 avdd.n2401 avdd.n2351 0.0398017
R7990 avdd.n2435 avdd.n2344 0.0398017
R7991 avdd.n2438 avdd.n2437 0.0398017
R7992 avdd.n2458 avdd.n2325 0.0398017
R7993 avdd.n2477 avdd.n2318 0.0398017
R7994 avdd.n2508 avdd.n2315 0.0398017
R7995 avdd.n2616 avdd.n2566 0.0398017
R7996 avdd.n2650 avdd.n2559 0.0398017
R7997 avdd.n2653 avdd.n2652 0.0398017
R7998 avdd.n2673 avdd.n2540 0.0398017
R7999 avdd.n2692 avdd.n2533 0.0398017
R8000 avdd.n2723 avdd.n2530 0.0398017
R8001 avdd.n2831 avdd.n2781 0.0398017
R8002 avdd.n2865 avdd.n2774 0.0398017
R8003 avdd.n2868 avdd.n2867 0.0398017
R8004 avdd.n2888 avdd.n2755 0.0398017
R8005 avdd.n2907 avdd.n2748 0.0398017
R8006 avdd.n2938 avdd.n2745 0.0398017
R8007 avdd.n3046 avdd.n2996 0.0398017
R8008 avdd.n3080 avdd.n2989 0.0398017
R8009 avdd.n3083 avdd.n3082 0.0398017
R8010 avdd.n3103 avdd.n2970 0.0398017
R8011 avdd.n3122 avdd.n2963 0.0398017
R8012 avdd.n3153 avdd.n2960 0.0398017
R8013 avdd.n3223 avdd.n3179 0.0398017
R8014 avdd.n3365 avdd.n3236 0.0398017
R8015 avdd.n3258 avdd.n3237 0.0398017
R8016 avdd.n3340 avdd.n3264 0.0398017
R8017 avdd.n3338 avdd.n3267 0.0398017
R8018 avdd.n3312 avdd.n3290 0.0398017
R8019 avdd.n3438 avdd.n3394 0.0398017
R8020 avdd.n3580 avdd.n3451 0.0398017
R8021 avdd.n3473 avdd.n3452 0.0398017
R8022 avdd.n3555 avdd.n3479 0.0398017
R8023 avdd.n3553 avdd.n3482 0.0398017
R8024 avdd.n3527 avdd.n3505 0.0398017
R8025 avdd.n3653 avdd.n3609 0.0398017
R8026 avdd.n3795 avdd.n3666 0.0398017
R8027 avdd.n3688 avdd.n3667 0.0398017
R8028 avdd.n3770 avdd.n3694 0.0398017
R8029 avdd.n3768 avdd.n3697 0.0398017
R8030 avdd.n3742 avdd.n3720 0.0398017
R8031 avdd.n3868 avdd.n3824 0.0398017
R8032 avdd.n4010 avdd.n3881 0.0398017
R8033 avdd.n3903 avdd.n3882 0.0398017
R8034 avdd.n3985 avdd.n3909 0.0398017
R8035 avdd.n3983 avdd.n3912 0.0398017
R8036 avdd.n3957 avdd.n3935 0.0398017
R8037 avdd.n4083 avdd.n4039 0.0398017
R8038 avdd.n4225 avdd.n4096 0.0398017
R8039 avdd.n4118 avdd.n4097 0.0398017
R8040 avdd.n4200 avdd.n4124 0.0398017
R8041 avdd.n4198 avdd.n4127 0.0398017
R8042 avdd.n4172 avdd.n4150 0.0398017
R8043 avdd.n4298 avdd.n4254 0.0398017
R8044 avdd.n4440 avdd.n4311 0.0398017
R8045 avdd.n4333 avdd.n4312 0.0398017
R8046 avdd.n4415 avdd.n4339 0.0398017
R8047 avdd.n4413 avdd.n4342 0.0398017
R8048 avdd.n4387 avdd.n4365 0.0398017
R8049 avdd.n4909 avdd.n4858 0.0398017
R8050 avdd.n4942 avdd.n4851 0.0398017
R8051 avdd.n4945 avdd.n4944 0.0398017
R8052 avdd.n4965 avdd.n4832 0.0398017
R8053 avdd.n4984 avdd.n4824 0.0398017
R8054 avdd.n5010 avdd.n4821 0.0398017
R8055 avdd.n5125 avdd.n5074 0.0398017
R8056 avdd.n5158 avdd.n5067 0.0398017
R8057 avdd.n5161 avdd.n5160 0.0398017
R8058 avdd.n5181 avdd.n5048 0.0398017
R8059 avdd.n5200 avdd.n5040 0.0398017
R8060 avdd.n5226 avdd.n5037 0.0398017
R8061 avdd.n5341 avdd.n5290 0.0398017
R8062 avdd.n5374 avdd.n5283 0.0398017
R8063 avdd.n5377 avdd.n5376 0.0398017
R8064 avdd.n5397 avdd.n5264 0.0398017
R8065 avdd.n5416 avdd.n5256 0.0398017
R8066 avdd.n5442 avdd.n5253 0.0398017
R8067 avdd.n5557 avdd.n5506 0.0398017
R8068 avdd.n5590 avdd.n5499 0.0398017
R8069 avdd.n5593 avdd.n5592 0.0398017
R8070 avdd.n5613 avdd.n5480 0.0398017
R8071 avdd.n5632 avdd.n5472 0.0398017
R8072 avdd.n5658 avdd.n5469 0.0398017
R8073 avdd.n5773 avdd.n5722 0.0398017
R8074 avdd.n5806 avdd.n5715 0.0398017
R8075 avdd.n5809 avdd.n5808 0.0398017
R8076 avdd.n5829 avdd.n5696 0.0398017
R8077 avdd.n5848 avdd.n5688 0.0398017
R8078 avdd.n5874 avdd.n5685 0.0398017
R8079 avdd.n5989 avdd.n5938 0.0398017
R8080 avdd.n6022 avdd.n5931 0.0398017
R8081 avdd.n6025 avdd.n6024 0.0398017
R8082 avdd.n6045 avdd.n5912 0.0398017
R8083 avdd.n6064 avdd.n5904 0.0398017
R8084 avdd.n6090 avdd.n5901 0.0398017
R8085 avdd.n6205 avdd.n6154 0.0398017
R8086 avdd.n6238 avdd.n6147 0.0398017
R8087 avdd.n6241 avdd.n6240 0.0398017
R8088 avdd.n6261 avdd.n6128 0.0398017
R8089 avdd.n6280 avdd.n6120 0.0398017
R8090 avdd.n6306 avdd.n6117 0.0398017
R8091 avdd.n6421 avdd.n6370 0.0398017
R8092 avdd.n6454 avdd.n6363 0.0398017
R8093 avdd.n6457 avdd.n6456 0.0398017
R8094 avdd.n6477 avdd.n6344 0.0398017
R8095 avdd.n6496 avdd.n6336 0.0398017
R8096 avdd.n6522 avdd.n6333 0.0398017
R8097 avdd.n6637 avdd.n6586 0.0398017
R8098 avdd.n6670 avdd.n6579 0.0398017
R8099 avdd.n6673 avdd.n6672 0.0398017
R8100 avdd.n6693 avdd.n6560 0.0398017
R8101 avdd.n6712 avdd.n6552 0.0398017
R8102 avdd.n6738 avdd.n6549 0.0398017
R8103 avdd.n6853 avdd.n6802 0.0398017
R8104 avdd.n6886 avdd.n6795 0.0398017
R8105 avdd.n6889 avdd.n6888 0.0398017
R8106 avdd.n6909 avdd.n6776 0.0398017
R8107 avdd.n6928 avdd.n6768 0.0398017
R8108 avdd.n6954 avdd.n6765 0.0398017
R8109 avdd.n7069 avdd.n7018 0.0398017
R8110 avdd.n7102 avdd.n7011 0.0398017
R8111 avdd.n7105 avdd.n7104 0.0398017
R8112 avdd.n7125 avdd.n6992 0.0398017
R8113 avdd.n7144 avdd.n6984 0.0398017
R8114 avdd.n7170 avdd.n6981 0.0398017
R8115 avdd.n7285 avdd.n7234 0.0398017
R8116 avdd.n7318 avdd.n7227 0.0398017
R8117 avdd.n7321 avdd.n7320 0.0398017
R8118 avdd.n7341 avdd.n7208 0.0398017
R8119 avdd.n7360 avdd.n7200 0.0398017
R8120 avdd.n7386 avdd.n7197 0.0398017
R8121 avdd.n7730 avdd.n7729 0.0398017
R8122 avdd.n7689 avdd.n7688 0.0398017
R8123 avdd.n7670 avdd.n7669 0.0398017
R8124 avdd.n7820 avdd.n7819 0.0398017
R8125 avdd.n7836 avdd.n7835 0.0398017
R8126 avdd.n10209 avdd.n10208 0.0398017
R8127 avdd.n10168 avdd.n10167 0.0398017
R8128 avdd.n10149 avdd.n10148 0.0398017
R8129 avdd.n10137 avdd.n10136 0.0398017
R8130 avdd.n10078 avdd.n10077 0.0398017
R8131 avdd.n10094 avdd.n10093 0.0398017
R8132 avdd.n10015 avdd.n10014 0.0398017
R8133 avdd.n9952 avdd.n9951 0.0398017
R8134 avdd.n10290 avdd.n10289 0.0398017
R8135 avdd.n10310 avdd.n10309 0.0398017
R8136 avdd.n10326 avdd.n10325 0.0398017
R8137 avdd.n9901 avdd.n9900 0.0398017
R8138 avdd.n9838 avdd.n9837 0.0398017
R8139 avdd.n10392 avdd.n10391 0.0398017
R8140 avdd.n10412 avdd.n10411 0.0398017
R8141 avdd.n10428 avdd.n10427 0.0398017
R8142 avdd.n9787 avdd.n9786 0.0398017
R8143 avdd.n9724 avdd.n9723 0.0398017
R8144 avdd.n10494 avdd.n10493 0.0398017
R8145 avdd.n10514 avdd.n10513 0.0398017
R8146 avdd.n10530 avdd.n10529 0.0398017
R8147 avdd.n9674 avdd.n9673 0.0398017
R8148 avdd.n9611 avdd.n9610 0.0398017
R8149 avdd.n10596 avdd.n10595 0.0398017
R8150 avdd.n10616 avdd.n10615 0.0398017
R8151 avdd.n10632 avdd.n10631 0.0398017
R8152 avdd.n9559 avdd.n9558 0.0398017
R8153 avdd.n9496 avdd.n9495 0.0398017
R8154 avdd.n10698 avdd.n10697 0.0398017
R8155 avdd.n10718 avdd.n10717 0.0398017
R8156 avdd.n10734 avdd.n10733 0.0398017
R8157 avdd.n9445 avdd.n9444 0.0398017
R8158 avdd.n9382 avdd.n9381 0.0398017
R8159 avdd.n10800 avdd.n10799 0.0398017
R8160 avdd.n10820 avdd.n10819 0.0398017
R8161 avdd.n10836 avdd.n10835 0.0398017
R8162 avdd.n9331 avdd.n9330 0.0398017
R8163 avdd.n9268 avdd.n9267 0.0398017
R8164 avdd.n10902 avdd.n10901 0.0398017
R8165 avdd.n10922 avdd.n10921 0.0398017
R8166 avdd.n10938 avdd.n10937 0.0398017
R8167 avdd.n9217 avdd.n9216 0.0398017
R8168 avdd.n9154 avdd.n9153 0.0398017
R8169 avdd.n11004 avdd.n11003 0.0398017
R8170 avdd.n11024 avdd.n11023 0.0398017
R8171 avdd.n11040 avdd.n11039 0.0398017
R8172 avdd.n9103 avdd.n9102 0.0398017
R8173 avdd.n9040 avdd.n9039 0.0398017
R8174 avdd.n11106 avdd.n11105 0.0398017
R8175 avdd.n11126 avdd.n11125 0.0398017
R8176 avdd.n11142 avdd.n11141 0.0398017
R8177 avdd.n8989 avdd.n8988 0.0398017
R8178 avdd.n8926 avdd.n8925 0.0398017
R8179 avdd.n11208 avdd.n11207 0.0398017
R8180 avdd.n11228 avdd.n11227 0.0398017
R8181 avdd.n11244 avdd.n11243 0.0398017
R8182 avdd.n125 avdd.n124 0.0398017
R8183 avdd.n172 avdd.n171 0.0398017
R8184 avdd.n153 avdd.n152 0.0398017
R8185 avdd.n141 avdd.n140 0.0398017
R8186 avdd.n8841 avdd.n8840 0.0398017
R8187 avdd.n8857 avdd.n8856 0.0398017
R8188 avdd.n255 avdd.n254 0.0398017
R8189 avdd.n302 avdd.n301 0.0398017
R8190 avdd.n283 avdd.n282 0.0398017
R8191 avdd.n271 avdd.n270 0.0398017
R8192 avdd.n8755 avdd.n8754 0.0398017
R8193 avdd.n8771 avdd.n8770 0.0398017
R8194 avdd.n385 avdd.n384 0.0398017
R8195 avdd.n432 avdd.n431 0.0398017
R8196 avdd.n413 avdd.n412 0.0398017
R8197 avdd.n401 avdd.n400 0.0398017
R8198 avdd.n8669 avdd.n8668 0.0398017
R8199 avdd.n8685 avdd.n8684 0.0398017
R8200 avdd.n515 avdd.n514 0.0398017
R8201 avdd.n562 avdd.n561 0.0398017
R8202 avdd.n543 avdd.n542 0.0398017
R8203 avdd.n531 avdd.n530 0.0398017
R8204 avdd.n8583 avdd.n8582 0.0398017
R8205 avdd.n8599 avdd.n8598 0.0398017
R8206 avdd.n645 avdd.n644 0.0398017
R8207 avdd.n692 avdd.n691 0.0398017
R8208 avdd.n673 avdd.n672 0.0398017
R8209 avdd.n661 avdd.n660 0.0398017
R8210 avdd.n8497 avdd.n8496 0.0398017
R8211 avdd.n8513 avdd.n8512 0.0398017
R8212 avdd.n775 avdd.n774 0.0398017
R8213 avdd.n822 avdd.n821 0.0398017
R8214 avdd.n803 avdd.n802 0.0398017
R8215 avdd.n791 avdd.n790 0.0398017
R8216 avdd.n8411 avdd.n8410 0.0398017
R8217 avdd.n8427 avdd.n8426 0.0398017
R8218 avdd.n905 avdd.n904 0.0398017
R8219 avdd.n952 avdd.n951 0.0398017
R8220 avdd.n933 avdd.n932 0.0398017
R8221 avdd.n921 avdd.n920 0.0398017
R8222 avdd.n8325 avdd.n8324 0.0398017
R8223 avdd.n8341 avdd.n8340 0.0398017
R8224 avdd.n1035 avdd.n1034 0.0398017
R8225 avdd.n1082 avdd.n1081 0.0398017
R8226 avdd.n1063 avdd.n1062 0.0398017
R8227 avdd.n1051 avdd.n1050 0.0398017
R8228 avdd.n8239 avdd.n8238 0.0398017
R8229 avdd.n8255 avdd.n8254 0.0398017
R8230 avdd.n1165 avdd.n1164 0.0398017
R8231 avdd.n1212 avdd.n1211 0.0398017
R8232 avdd.n1193 avdd.n1192 0.0398017
R8233 avdd.n1181 avdd.n1180 0.0398017
R8234 avdd.n8153 avdd.n8152 0.0398017
R8235 avdd.n8169 avdd.n8168 0.0398017
R8236 avdd.n1295 avdd.n1294 0.0398017
R8237 avdd.n1342 avdd.n1341 0.0398017
R8238 avdd.n1323 avdd.n1322 0.0398017
R8239 avdd.n1311 avdd.n1310 0.0398017
R8240 avdd.n8067 avdd.n8066 0.0398017
R8241 avdd.n8083 avdd.n8082 0.0398017
R8242 avdd.n1425 avdd.n1424 0.0398017
R8243 avdd.n1472 avdd.n1471 0.0398017
R8244 avdd.n1453 avdd.n1452 0.0398017
R8245 avdd.n1441 avdd.n1440 0.0398017
R8246 avdd.n7981 avdd.n7980 0.0398017
R8247 avdd.n7997 avdd.n7996 0.0398017
R8248 avdd.n1555 avdd.n1554 0.0398017
R8249 avdd.n1602 avdd.n1601 0.0398017
R8250 avdd.n1583 avdd.n1582 0.0398017
R8251 avdd.n1571 avdd.n1570 0.0398017
R8252 avdd.n7895 avdd.n7894 0.0398017
R8253 avdd.n7911 avdd.n7910 0.0398017
R8254 avdd.n55 avdd 0.0382604
R8255 avdd.n1905 avdd.n1897 0.0368182
R8256 avdd.n2159 avdd.n2151 0.0368182
R8257 avdd.n2374 avdd.n2366 0.0368182
R8258 avdd.n2589 avdd.n2581 0.0368182
R8259 avdd.n2804 avdd.n2796 0.0368182
R8260 avdd.n3019 avdd.n3011 0.0368182
R8261 avdd.n3195 avdd.n3187 0.0368182
R8262 avdd.n3410 avdd.n3402 0.0368182
R8263 avdd.n3625 avdd.n3617 0.0368182
R8264 avdd.n3840 avdd.n3832 0.0368182
R8265 avdd.n4055 avdd.n4047 0.0368182
R8266 avdd.n4270 avdd.n4262 0.0368182
R8267 avdd.n4881 avdd.n4873 0.0368182
R8268 avdd.n5097 avdd.n5089 0.0368182
R8269 avdd.n5313 avdd.n5305 0.0368182
R8270 avdd.n5529 avdd.n5521 0.0368182
R8271 avdd.n5745 avdd.n5737 0.0368182
R8272 avdd.n5961 avdd.n5953 0.0368182
R8273 avdd.n6177 avdd.n6169 0.0368182
R8274 avdd.n6393 avdd.n6385 0.0368182
R8275 avdd.n6609 avdd.n6601 0.0368182
R8276 avdd.n6825 avdd.n6817 0.0368182
R8277 avdd.n7041 avdd.n7033 0.0368182
R8278 avdd.n7257 avdd.n7249 0.0368182
R8279 avdd.n7757 avdd.n7756 0.0368182
R8280 avdd.n10236 avdd.n10235 0.0368182
R8281 avdd.n9990 avdd.n9989 0.0368182
R8282 avdd.n9876 avdd.n9875 0.0368182
R8283 avdd.n9762 avdd.n9761 0.0368182
R8284 avdd.n9649 avdd.n9648 0.0368182
R8285 avdd.n9534 avdd.n9533 0.0368182
R8286 avdd.n9420 avdd.n9419 0.0368182
R8287 avdd.n9306 avdd.n9305 0.0368182
R8288 avdd.n9192 avdd.n9191 0.0368182
R8289 avdd.n9078 avdd.n9077 0.0368182
R8290 avdd.n8964 avdd.n8963 0.0368182
R8291 avdd.n90 avdd.n89 0.0368182
R8292 avdd.n220 avdd.n219 0.0368182
R8293 avdd.n350 avdd.n349 0.0368182
R8294 avdd.n480 avdd.n479 0.0368182
R8295 avdd.n610 avdd.n609 0.0368182
R8296 avdd.n740 avdd.n739 0.0368182
R8297 avdd.n870 avdd.n869 0.0368182
R8298 avdd.n1000 avdd.n999 0.0368182
R8299 avdd.n1130 avdd.n1129 0.0368182
R8300 avdd.n1260 avdd.n1259 0.0368182
R8301 avdd.n1390 avdd.n1389 0.0368182
R8302 avdd.n1520 avdd.n1519 0.0368182
R8303 avdd.n2058 avdd.n2057 0.0368182
R8304 avdd.n1904 avdd.n1898 0.0368182
R8305 avdd.n2059 avdd.n1971 0.0368182
R8306 avdd.n2238 avdd.n2114 0.0368182
R8307 avdd.n2158 avdd.n2152 0.0368182
R8308 avdd.n2239 avdd.n2115 0.0368182
R8309 avdd.n2453 avdd.n2329 0.0368182
R8310 avdd.n2373 avdd.n2367 0.0368182
R8311 avdd.n2454 avdd.n2330 0.0368182
R8312 avdd.n2668 avdd.n2544 0.0368182
R8313 avdd.n2588 avdd.n2582 0.0368182
R8314 avdd.n2669 avdd.n2545 0.0368182
R8315 avdd.n2883 avdd.n2759 0.0368182
R8316 avdd.n2803 avdd.n2797 0.0368182
R8317 avdd.n2884 avdd.n2760 0.0368182
R8318 avdd.n3098 avdd.n2974 0.0368182
R8319 avdd.n3018 avdd.n3012 0.0368182
R8320 avdd.n3099 avdd.n2975 0.0368182
R8321 avdd.n3347 avdd.n3346 0.0368182
R8322 avdd.n3194 avdd.n3188 0.0368182
R8323 avdd.n3348 avdd.n3261 0.0368182
R8324 avdd.n3562 avdd.n3561 0.0368182
R8325 avdd.n3409 avdd.n3403 0.0368182
R8326 avdd.n3563 avdd.n3476 0.0368182
R8327 avdd.n3777 avdd.n3776 0.0368182
R8328 avdd.n3624 avdd.n3618 0.0368182
R8329 avdd.n3778 avdd.n3691 0.0368182
R8330 avdd.n3992 avdd.n3991 0.0368182
R8331 avdd.n3839 avdd.n3833 0.0368182
R8332 avdd.n3993 avdd.n3906 0.0368182
R8333 avdd.n4207 avdd.n4206 0.0368182
R8334 avdd.n4054 avdd.n4048 0.0368182
R8335 avdd.n4208 avdd.n4121 0.0368182
R8336 avdd.n4422 avdd.n4421 0.0368182
R8337 avdd.n4269 avdd.n4263 0.0368182
R8338 avdd.n4423 avdd.n4336 0.0368182
R8339 avdd.n4960 avdd.n4836 0.0368182
R8340 avdd.n4880 avdd.n4874 0.0368182
R8341 avdd.n4961 avdd.n4837 0.0368182
R8342 avdd.n5176 avdd.n5052 0.0368182
R8343 avdd.n5096 avdd.n5090 0.0368182
R8344 avdd.n5177 avdd.n5053 0.0368182
R8345 avdd.n5392 avdd.n5268 0.0368182
R8346 avdd.n5312 avdd.n5306 0.0368182
R8347 avdd.n5393 avdd.n5269 0.0368182
R8348 avdd.n5608 avdd.n5484 0.0368182
R8349 avdd.n5528 avdd.n5522 0.0368182
R8350 avdd.n5609 avdd.n5485 0.0368182
R8351 avdd.n5824 avdd.n5700 0.0368182
R8352 avdd.n5744 avdd.n5738 0.0368182
R8353 avdd.n5825 avdd.n5701 0.0368182
R8354 avdd.n6040 avdd.n5916 0.0368182
R8355 avdd.n5960 avdd.n5954 0.0368182
R8356 avdd.n6041 avdd.n5917 0.0368182
R8357 avdd.n6256 avdd.n6132 0.0368182
R8358 avdd.n6176 avdd.n6170 0.0368182
R8359 avdd.n6257 avdd.n6133 0.0368182
R8360 avdd.n6472 avdd.n6348 0.0368182
R8361 avdd.n6392 avdd.n6386 0.0368182
R8362 avdd.n6473 avdd.n6349 0.0368182
R8363 avdd.n6688 avdd.n6564 0.0368182
R8364 avdd.n6608 avdd.n6602 0.0368182
R8365 avdd.n6689 avdd.n6565 0.0368182
R8366 avdd.n6904 avdd.n6780 0.0368182
R8367 avdd.n6824 avdd.n6818 0.0368182
R8368 avdd.n6905 avdd.n6781 0.0368182
R8369 avdd.n7120 avdd.n6996 0.0368182
R8370 avdd.n7040 avdd.n7034 0.0368182
R8371 avdd.n7121 avdd.n6997 0.0368182
R8372 avdd.n7336 avdd.n7212 0.0368182
R8373 avdd.n7256 avdd.n7250 0.0368182
R8374 avdd.n7337 avdd.n7213 0.0368182
R8375 avdd.n7769 avdd.n7768 0.0368182
R8376 avdd.n7742 avdd.n7741 0.0368182
R8377 avdd.n10221 avdd.n10220 0.0368182
R8378 avdd.n10131 avdd.n10130 0.0368182
R8379 avdd.n9968 avdd.n9967 0.0368182
R8380 avdd.n10283 avdd.n10282 0.0368182
R8381 avdd.n9854 avdd.n9853 0.0368182
R8382 avdd.n10385 avdd.n10384 0.0368182
R8383 avdd.n9740 avdd.n9739 0.0368182
R8384 avdd.n10487 avdd.n10486 0.0368182
R8385 avdd.n9627 avdd.n9626 0.0368182
R8386 avdd.n10589 avdd.n10588 0.0368182
R8387 avdd.n9512 avdd.n9511 0.0368182
R8388 avdd.n10691 avdd.n10690 0.0368182
R8389 avdd.n9398 avdd.n9397 0.0368182
R8390 avdd.n10793 avdd.n10792 0.0368182
R8391 avdd.n9284 avdd.n9283 0.0368182
R8392 avdd.n10895 avdd.n10894 0.0368182
R8393 avdd.n9170 avdd.n9169 0.0368182
R8394 avdd.n10997 avdd.n10996 0.0368182
R8395 avdd.n9056 avdd.n9055 0.0368182
R8396 avdd.n11099 avdd.n11098 0.0368182
R8397 avdd.n8942 avdd.n8941 0.0368182
R8398 avdd.n11201 avdd.n11200 0.0368182
R8399 avdd.n75 avdd.n74 0.0368182
R8400 avdd.n135 avdd.n134 0.0368182
R8401 avdd.n205 avdd.n204 0.0368182
R8402 avdd.n265 avdd.n264 0.0368182
R8403 avdd.n335 avdd.n334 0.0368182
R8404 avdd.n395 avdd.n394 0.0368182
R8405 avdd.n465 avdd.n464 0.0368182
R8406 avdd.n525 avdd.n524 0.0368182
R8407 avdd.n595 avdd.n594 0.0368182
R8408 avdd.n655 avdd.n654 0.0368182
R8409 avdd.n725 avdd.n724 0.0368182
R8410 avdd.n785 avdd.n784 0.0368182
R8411 avdd.n855 avdd.n854 0.0368182
R8412 avdd.n915 avdd.n914 0.0368182
R8413 avdd.n985 avdd.n984 0.0368182
R8414 avdd.n1045 avdd.n1044 0.0368182
R8415 avdd.n1115 avdd.n1114 0.0368182
R8416 avdd.n1175 avdd.n1174 0.0368182
R8417 avdd.n1245 avdd.n1244 0.0368182
R8418 avdd.n1305 avdd.n1304 0.0368182
R8419 avdd.n1375 avdd.n1374 0.0368182
R8420 avdd.n1435 avdd.n1434 0.0368182
R8421 avdd.n1505 avdd.n1504 0.0368182
R8422 avdd.n1565 avdd.n1564 0.0368182
R8423 avdd.n4738 avdd.n4737 0.0359167
R8424 avdd.n2065 avdd.n1957 0.0353939
R8425 avdd.n2067 avdd.n2066 0.0353939
R8426 avdd.n2230 avdd.n2120 0.0353939
R8427 avdd.n2232 avdd.n2231 0.0353939
R8428 avdd.n2445 avdd.n2335 0.0353939
R8429 avdd.n2447 avdd.n2446 0.0353939
R8430 avdd.n2660 avdd.n2550 0.0353939
R8431 avdd.n2662 avdd.n2661 0.0353939
R8432 avdd.n2875 avdd.n2765 0.0353939
R8433 avdd.n2877 avdd.n2876 0.0353939
R8434 avdd.n3090 avdd.n2980 0.0353939
R8435 avdd.n3092 avdd.n3091 0.0353939
R8436 avdd.n3354 avdd.n3247 0.0353939
R8437 avdd.n3356 avdd.n3355 0.0353939
R8438 avdd.n3569 avdd.n3462 0.0353939
R8439 avdd.n3571 avdd.n3570 0.0353939
R8440 avdd.n3784 avdd.n3677 0.0353939
R8441 avdd.n3786 avdd.n3785 0.0353939
R8442 avdd.n3999 avdd.n3892 0.0353939
R8443 avdd.n4001 avdd.n4000 0.0353939
R8444 avdd.n4214 avdd.n4107 0.0353939
R8445 avdd.n4216 avdd.n4215 0.0353939
R8446 avdd.n4429 avdd.n4322 0.0353939
R8447 avdd.n4431 avdd.n4430 0.0353939
R8448 avdd.n4952 avdd.n4842 0.0353939
R8449 avdd.n4954 avdd.n4953 0.0353939
R8450 avdd.n5168 avdd.n5058 0.0353939
R8451 avdd.n5170 avdd.n5169 0.0353939
R8452 avdd.n5384 avdd.n5274 0.0353939
R8453 avdd.n5386 avdd.n5385 0.0353939
R8454 avdd.n5600 avdd.n5490 0.0353939
R8455 avdd.n5602 avdd.n5601 0.0353939
R8456 avdd.n5816 avdd.n5706 0.0353939
R8457 avdd.n5818 avdd.n5817 0.0353939
R8458 avdd.n6032 avdd.n5922 0.0353939
R8459 avdd.n6034 avdd.n6033 0.0353939
R8460 avdd.n6248 avdd.n6138 0.0353939
R8461 avdd.n6250 avdd.n6249 0.0353939
R8462 avdd.n6464 avdd.n6354 0.0353939
R8463 avdd.n6466 avdd.n6465 0.0353939
R8464 avdd.n6680 avdd.n6570 0.0353939
R8465 avdd.n6682 avdd.n6681 0.0353939
R8466 avdd.n6896 avdd.n6786 0.0353939
R8467 avdd.n6898 avdd.n6897 0.0353939
R8468 avdd.n7112 avdd.n7002 0.0353939
R8469 avdd.n7114 avdd.n7113 0.0353939
R8470 avdd.n7328 avdd.n7218 0.0353939
R8471 avdd.n7330 avdd.n7329 0.0353939
R8472 avdd.n7641 avdd.n7640 0.0353939
R8473 avdd.n7665 avdd.n7664 0.0353939
R8474 avdd.n10118 avdd.n10117 0.0353939
R8475 avdd.n10144 avdd.n10143 0.0353939
R8476 avdd.n9919 avdd.n9918 0.0353939
R8477 avdd.n9805 avdd.n9804 0.0353939
R8478 avdd.n9691 avdd.n9690 0.0353939
R8479 avdd.n9577 avdd.n9576 0.0353939
R8480 avdd.n9463 avdd.n9462 0.0353939
R8481 avdd.n9349 avdd.n9348 0.0353939
R8482 avdd.n9235 avdd.n9234 0.0353939
R8483 avdd.n9121 avdd.n9120 0.0353939
R8484 avdd.n9007 avdd.n9006 0.0353939
R8485 avdd.n8893 avdd.n8892 0.0353939
R8486 avdd.n62 avdd.n61 0.0353939
R8487 avdd.n148 avdd.n147 0.0353939
R8488 avdd.n192 avdd.n191 0.0353939
R8489 avdd.n278 avdd.n277 0.0353939
R8490 avdd.n322 avdd.n321 0.0353939
R8491 avdd.n408 avdd.n407 0.0353939
R8492 avdd.n452 avdd.n451 0.0353939
R8493 avdd.n538 avdd.n537 0.0353939
R8494 avdd.n582 avdd.n581 0.0353939
R8495 avdd.n668 avdd.n667 0.0353939
R8496 avdd.n712 avdd.n711 0.0353939
R8497 avdd.n798 avdd.n797 0.0353939
R8498 avdd.n842 avdd.n841 0.0353939
R8499 avdd.n928 avdd.n927 0.0353939
R8500 avdd.n972 avdd.n971 0.0353939
R8501 avdd.n1058 avdd.n1057 0.0353939
R8502 avdd.n1102 avdd.n1101 0.0353939
R8503 avdd.n1188 avdd.n1187 0.0353939
R8504 avdd.n1232 avdd.n1231 0.0353939
R8505 avdd.n1318 avdd.n1317 0.0353939
R8506 avdd.n1362 avdd.n1361 0.0353939
R8507 avdd.n1448 avdd.n1447 0.0353939
R8508 avdd.n1492 avdd.n1491 0.0353939
R8509 avdd.n1578 avdd.n1577 0.0353939
R8510 avdd.n4805 avdd 0.0330521
R8511 avdd.n4766 avdd 0.0330521
R8512 avdd.n2090 avdd.n2089 0.0327477
R8513 avdd.n2197 avdd.n2196 0.0327477
R8514 avdd.n2412 avdd.n2411 0.0327477
R8515 avdd.n2627 avdd.n2626 0.0327477
R8516 avdd.n2842 avdd.n2841 0.0327477
R8517 avdd.n3057 avdd.n3056 0.0327477
R8518 avdd.n185 avdd.n133 0.0327477
R8519 avdd.n315 avdd.n263 0.0327477
R8520 avdd.n445 avdd.n393 0.0327477
R8521 avdd.n575 avdd.n523 0.0327477
R8522 avdd.n705 avdd.n653 0.0327477
R8523 avdd.n835 avdd.n783 0.0327477
R8524 avdd.n965 avdd.n913 0.0327477
R8525 avdd.n1095 avdd.n1043 0.0327477
R8526 avdd.n1225 avdd.n1173 0.0327477
R8527 avdd.n1355 avdd.n1303 0.0327477
R8528 avdd.n1485 avdd.n1433 0.0327477
R8529 avdd.n1615 avdd.n1563 0.0327477
R8530 avdd.n2052 avdd.n1975 0.032697
R8531 avdd.n2062 avdd.n1962 0.032697
R8532 avdd.n2062 avdd.n2061 0.032697
R8533 avdd.n1966 avdd.n1963 0.032697
R8534 avdd.n1910 avdd.n1902 0.032697
R8535 avdd.n1912 avdd.n1902 0.032697
R8536 avdd.n1921 avdd.n1920 0.032697
R8537 avdd.n2025 avdd.n2022 0.032697
R8538 avdd.n2246 avdd.n2245 0.032697
R8539 avdd.n2233 avdd.n2118 0.032697
R8540 avdd.n2241 avdd.n2118 0.032697
R8541 avdd.n2225 avdd.n2224 0.032697
R8542 avdd.n2164 avdd.n2156 0.032697
R8543 avdd.n2166 avdd.n2156 0.032697
R8544 avdd.n2175 avdd.n2174 0.032697
R8545 avdd.n2299 avdd.n2298 0.032697
R8546 avdd.n2461 avdd.n2460 0.032697
R8547 avdd.n2448 avdd.n2333 0.032697
R8548 avdd.n2456 avdd.n2333 0.032697
R8549 avdd.n2440 avdd.n2439 0.032697
R8550 avdd.n2379 avdd.n2371 0.032697
R8551 avdd.n2381 avdd.n2371 0.032697
R8552 avdd.n2390 avdd.n2389 0.032697
R8553 avdd.n2514 avdd.n2513 0.032697
R8554 avdd.n2676 avdd.n2675 0.032697
R8555 avdd.n2663 avdd.n2548 0.032697
R8556 avdd.n2671 avdd.n2548 0.032697
R8557 avdd.n2655 avdd.n2654 0.032697
R8558 avdd.n2594 avdd.n2586 0.032697
R8559 avdd.n2596 avdd.n2586 0.032697
R8560 avdd.n2605 avdd.n2604 0.032697
R8561 avdd.n2729 avdd.n2728 0.032697
R8562 avdd.n2891 avdd.n2890 0.032697
R8563 avdd.n2878 avdd.n2763 0.032697
R8564 avdd.n2886 avdd.n2763 0.032697
R8565 avdd.n2870 avdd.n2869 0.032697
R8566 avdd.n2809 avdd.n2801 0.032697
R8567 avdd.n2811 avdd.n2801 0.032697
R8568 avdd.n2820 avdd.n2819 0.032697
R8569 avdd.n2944 avdd.n2943 0.032697
R8570 avdd.n3106 avdd.n3105 0.032697
R8571 avdd.n3093 avdd.n2978 0.032697
R8572 avdd.n3101 avdd.n2978 0.032697
R8573 avdd.n3085 avdd.n3084 0.032697
R8574 avdd.n3024 avdd.n3016 0.032697
R8575 avdd.n3026 avdd.n3016 0.032697
R8576 avdd.n3035 avdd.n3034 0.032697
R8577 avdd.n3159 avdd.n3158 0.032697
R8578 avdd.n3341 avdd.n3265 0.032697
R8579 avdd.n3351 avdd.n3252 0.032697
R8580 avdd.n3351 avdd.n3350 0.032697
R8581 avdd.n3256 avdd.n3253 0.032697
R8582 avdd.n3200 avdd.n3192 0.032697
R8583 avdd.n3202 avdd.n3192 0.032697
R8584 avdd.n3211 avdd.n3210 0.032697
R8585 avdd.n3316 avdd.n3314 0.032697
R8586 avdd.n3556 avdd.n3480 0.032697
R8587 avdd.n3566 avdd.n3467 0.032697
R8588 avdd.n3566 avdd.n3565 0.032697
R8589 avdd.n3471 avdd.n3468 0.032697
R8590 avdd.n3415 avdd.n3407 0.032697
R8591 avdd.n3417 avdd.n3407 0.032697
R8592 avdd.n3426 avdd.n3425 0.032697
R8593 avdd.n3531 avdd.n3529 0.032697
R8594 avdd.n3771 avdd.n3695 0.032697
R8595 avdd.n3781 avdd.n3682 0.032697
R8596 avdd.n3781 avdd.n3780 0.032697
R8597 avdd.n3686 avdd.n3683 0.032697
R8598 avdd.n3630 avdd.n3622 0.032697
R8599 avdd.n3632 avdd.n3622 0.032697
R8600 avdd.n3641 avdd.n3640 0.032697
R8601 avdd.n3746 avdd.n3744 0.032697
R8602 avdd.n3986 avdd.n3910 0.032697
R8603 avdd.n3996 avdd.n3897 0.032697
R8604 avdd.n3996 avdd.n3995 0.032697
R8605 avdd.n3901 avdd.n3898 0.032697
R8606 avdd.n3845 avdd.n3837 0.032697
R8607 avdd.n3847 avdd.n3837 0.032697
R8608 avdd.n3856 avdd.n3855 0.032697
R8609 avdd.n3961 avdd.n3959 0.032697
R8610 avdd.n4201 avdd.n4125 0.032697
R8611 avdd.n4211 avdd.n4112 0.032697
R8612 avdd.n4211 avdd.n4210 0.032697
R8613 avdd.n4116 avdd.n4113 0.032697
R8614 avdd.n4060 avdd.n4052 0.032697
R8615 avdd.n4062 avdd.n4052 0.032697
R8616 avdd.n4071 avdd.n4070 0.032697
R8617 avdd.n4176 avdd.n4174 0.032697
R8618 avdd.n4416 avdd.n4340 0.032697
R8619 avdd.n4426 avdd.n4327 0.032697
R8620 avdd.n4426 avdd.n4425 0.032697
R8621 avdd.n4331 avdd.n4328 0.032697
R8622 avdd.n4275 avdd.n4267 0.032697
R8623 avdd.n4277 avdd.n4267 0.032697
R8624 avdd.n4286 avdd.n4285 0.032697
R8625 avdd.n4391 avdd.n4389 0.032697
R8626 avdd.n4886 avdd.n4878 0.032697
R8627 avdd.n4888 avdd.n4878 0.032697
R8628 avdd.n4897 avdd.n4896 0.032697
R8629 avdd.n4947 avdd.n4946 0.032697
R8630 avdd.n4955 avdd.n4840 0.032697
R8631 avdd.n4963 avdd.n4840 0.032697
R8632 avdd.n4968 avdd.n4967 0.032697
R8633 avdd.n5018 avdd.n5017 0.032697
R8634 avdd.n5102 avdd.n5094 0.032697
R8635 avdd.n5104 avdd.n5094 0.032697
R8636 avdd.n5113 avdd.n5112 0.032697
R8637 avdd.n5163 avdd.n5162 0.032697
R8638 avdd.n5171 avdd.n5056 0.032697
R8639 avdd.n5179 avdd.n5056 0.032697
R8640 avdd.n5184 avdd.n5183 0.032697
R8641 avdd.n5234 avdd.n5233 0.032697
R8642 avdd.n5318 avdd.n5310 0.032697
R8643 avdd.n5320 avdd.n5310 0.032697
R8644 avdd.n5329 avdd.n5328 0.032697
R8645 avdd.n5379 avdd.n5378 0.032697
R8646 avdd.n5387 avdd.n5272 0.032697
R8647 avdd.n5395 avdd.n5272 0.032697
R8648 avdd.n5400 avdd.n5399 0.032697
R8649 avdd.n5450 avdd.n5449 0.032697
R8650 avdd.n5534 avdd.n5526 0.032697
R8651 avdd.n5536 avdd.n5526 0.032697
R8652 avdd.n5545 avdd.n5544 0.032697
R8653 avdd.n5595 avdd.n5594 0.032697
R8654 avdd.n5603 avdd.n5488 0.032697
R8655 avdd.n5611 avdd.n5488 0.032697
R8656 avdd.n5616 avdd.n5615 0.032697
R8657 avdd.n5666 avdd.n5665 0.032697
R8658 avdd.n5750 avdd.n5742 0.032697
R8659 avdd.n5752 avdd.n5742 0.032697
R8660 avdd.n5761 avdd.n5760 0.032697
R8661 avdd.n5811 avdd.n5810 0.032697
R8662 avdd.n5819 avdd.n5704 0.032697
R8663 avdd.n5827 avdd.n5704 0.032697
R8664 avdd.n5832 avdd.n5831 0.032697
R8665 avdd.n5882 avdd.n5881 0.032697
R8666 avdd.n5966 avdd.n5958 0.032697
R8667 avdd.n5968 avdd.n5958 0.032697
R8668 avdd.n5977 avdd.n5976 0.032697
R8669 avdd.n6027 avdd.n6026 0.032697
R8670 avdd.n6035 avdd.n5920 0.032697
R8671 avdd.n6043 avdd.n5920 0.032697
R8672 avdd.n6048 avdd.n6047 0.032697
R8673 avdd.n6098 avdd.n6097 0.032697
R8674 avdd.n6182 avdd.n6174 0.032697
R8675 avdd.n6184 avdd.n6174 0.032697
R8676 avdd.n6193 avdd.n6192 0.032697
R8677 avdd.n6243 avdd.n6242 0.032697
R8678 avdd.n6251 avdd.n6136 0.032697
R8679 avdd.n6259 avdd.n6136 0.032697
R8680 avdd.n6264 avdd.n6263 0.032697
R8681 avdd.n6314 avdd.n6313 0.032697
R8682 avdd.n6398 avdd.n6390 0.032697
R8683 avdd.n6400 avdd.n6390 0.032697
R8684 avdd.n6409 avdd.n6408 0.032697
R8685 avdd.n6459 avdd.n6458 0.032697
R8686 avdd.n6467 avdd.n6352 0.032697
R8687 avdd.n6475 avdd.n6352 0.032697
R8688 avdd.n6480 avdd.n6479 0.032697
R8689 avdd.n6530 avdd.n6529 0.032697
R8690 avdd.n6614 avdd.n6606 0.032697
R8691 avdd.n6616 avdd.n6606 0.032697
R8692 avdd.n6625 avdd.n6624 0.032697
R8693 avdd.n6675 avdd.n6674 0.032697
R8694 avdd.n6683 avdd.n6568 0.032697
R8695 avdd.n6691 avdd.n6568 0.032697
R8696 avdd.n6696 avdd.n6695 0.032697
R8697 avdd.n6746 avdd.n6745 0.032697
R8698 avdd.n6830 avdd.n6822 0.032697
R8699 avdd.n6832 avdd.n6822 0.032697
R8700 avdd.n6841 avdd.n6840 0.032697
R8701 avdd.n6891 avdd.n6890 0.032697
R8702 avdd.n6899 avdd.n6784 0.032697
R8703 avdd.n6907 avdd.n6784 0.032697
R8704 avdd.n6912 avdd.n6911 0.032697
R8705 avdd.n6962 avdd.n6961 0.032697
R8706 avdd.n7046 avdd.n7038 0.032697
R8707 avdd.n7048 avdd.n7038 0.032697
R8708 avdd.n7057 avdd.n7056 0.032697
R8709 avdd.n7107 avdd.n7106 0.032697
R8710 avdd.n7115 avdd.n7000 0.032697
R8711 avdd.n7123 avdd.n7000 0.032697
R8712 avdd.n7128 avdd.n7127 0.032697
R8713 avdd.n7178 avdd.n7177 0.032697
R8714 avdd.n7262 avdd.n7254 0.032697
R8715 avdd.n7264 avdd.n7254 0.032697
R8716 avdd.n7273 avdd.n7272 0.032697
R8717 avdd.n7323 avdd.n7322 0.032697
R8718 avdd.n7331 avdd.n7216 0.032697
R8719 avdd.n7339 avdd.n7216 0.032697
R8720 avdd.n7344 avdd.n7343 0.032697
R8721 avdd.n7394 avdd.n7393 0.032697
R8722 avdd.n7752 avdd.n7748 0.032697
R8723 avdd.n7752 avdd.n7751 0.032697
R8724 avdd.n7715 avdd.n7708 0.032697
R8725 avdd.n7676 avdd.n7675 0.032697
R8726 avdd.n7661 avdd.n7657 0.032697
R8727 avdd.n7661 avdd.n7660 0.032697
R8728 avdd.n7804 avdd.n7799 0.032697
R8729 avdd.n7789 avdd.n7788 0.032697
R8730 avdd.n10231 avdd.n10227 0.032697
R8731 avdd.n10231 avdd.n10230 0.032697
R8732 avdd.n10194 avdd.n10187 0.032697
R8733 avdd.n10155 avdd.n10154 0.032697
R8734 avdd.n10140 avdd.n10135 0.032697
R8735 avdd.n10140 avdd.n10139 0.032697
R8736 avdd.n10062 avdd.n10058 0.032697
R8737 avdd.n10049 avdd.n10048 0.032697
R8738 avdd.n9985 avdd.n9977 0.032697
R8739 avdd.n9985 avdd.n9984 0.032697
R8740 avdd.n9939 avdd.n9938 0.032697
R8741 avdd.n10278 avdd.n10275 0.032697
R8742 avdd.n10278 avdd.n10277 0.032697
R8743 avdd.n10294 avdd.n10288 0.032697
R8744 avdd.n10265 avdd.n10264 0.032697
R8745 avdd.n9871 avdd.n9863 0.032697
R8746 avdd.n9871 avdd.n9870 0.032697
R8747 avdd.n9825 avdd.n9824 0.032697
R8748 avdd.n10380 avdd.n10377 0.032697
R8749 avdd.n10380 avdd.n10379 0.032697
R8750 avdd.n10396 avdd.n10390 0.032697
R8751 avdd.n10367 avdd.n10366 0.032697
R8752 avdd.n9757 avdd.n9749 0.032697
R8753 avdd.n9757 avdd.n9756 0.032697
R8754 avdd.n9711 avdd.n9710 0.032697
R8755 avdd.n10482 avdd.n10479 0.032697
R8756 avdd.n10482 avdd.n10481 0.032697
R8757 avdd.n10498 avdd.n10492 0.032697
R8758 avdd.n10469 avdd.n10468 0.032697
R8759 avdd.n9644 avdd.n9636 0.032697
R8760 avdd.n9644 avdd.n9643 0.032697
R8761 avdd.n9598 avdd.n9597 0.032697
R8762 avdd.n10584 avdd.n10581 0.032697
R8763 avdd.n10584 avdd.n10583 0.032697
R8764 avdd.n10600 avdd.n10594 0.032697
R8765 avdd.n10571 avdd.n10570 0.032697
R8766 avdd.n9529 avdd.n9521 0.032697
R8767 avdd.n9529 avdd.n9528 0.032697
R8768 avdd.n9483 avdd.n9482 0.032697
R8769 avdd.n10686 avdd.n10683 0.032697
R8770 avdd.n10686 avdd.n10685 0.032697
R8771 avdd.n10702 avdd.n10696 0.032697
R8772 avdd.n10673 avdd.n10672 0.032697
R8773 avdd.n9415 avdd.n9407 0.032697
R8774 avdd.n9415 avdd.n9414 0.032697
R8775 avdd.n9369 avdd.n9368 0.032697
R8776 avdd.n10788 avdd.n10785 0.032697
R8777 avdd.n10788 avdd.n10787 0.032697
R8778 avdd.n10804 avdd.n10798 0.032697
R8779 avdd.n10775 avdd.n10774 0.032697
R8780 avdd.n9301 avdd.n9293 0.032697
R8781 avdd.n9301 avdd.n9300 0.032697
R8782 avdd.n9255 avdd.n9254 0.032697
R8783 avdd.n10890 avdd.n10887 0.032697
R8784 avdd.n10890 avdd.n10889 0.032697
R8785 avdd.n10906 avdd.n10900 0.032697
R8786 avdd.n10877 avdd.n10876 0.032697
R8787 avdd.n9187 avdd.n9179 0.032697
R8788 avdd.n9187 avdd.n9186 0.032697
R8789 avdd.n9141 avdd.n9140 0.032697
R8790 avdd.n10992 avdd.n10989 0.032697
R8791 avdd.n10992 avdd.n10991 0.032697
R8792 avdd.n11008 avdd.n11002 0.032697
R8793 avdd.n10979 avdd.n10978 0.032697
R8794 avdd.n9073 avdd.n9065 0.032697
R8795 avdd.n9073 avdd.n9072 0.032697
R8796 avdd.n9027 avdd.n9026 0.032697
R8797 avdd.n11094 avdd.n11091 0.032697
R8798 avdd.n11094 avdd.n11093 0.032697
R8799 avdd.n11110 avdd.n11104 0.032697
R8800 avdd.n11081 avdd.n11080 0.032697
R8801 avdd.n8959 avdd.n8951 0.032697
R8802 avdd.n8959 avdd.n8958 0.032697
R8803 avdd.n8913 avdd.n8912 0.032697
R8804 avdd.n11196 avdd.n11193 0.032697
R8805 avdd.n11196 avdd.n11195 0.032697
R8806 avdd.n11212 avdd.n11206 0.032697
R8807 avdd.n11183 avdd.n11182 0.032697
R8808 avdd.n8825 avdd.n8821 0.032697
R8809 avdd.n144 avdd.n139 0.032697
R8810 avdd.n144 avdd.n143 0.032697
R8811 avdd.n159 avdd.n158 0.032697
R8812 avdd.n85 avdd.n81 0.032697
R8813 avdd.n85 avdd.n84 0.032697
R8814 avdd.n109 avdd.n102 0.032697
R8815 avdd.n8812 avdd.n8811 0.032697
R8816 avdd.n8739 avdd.n8735 0.032697
R8817 avdd.n274 avdd.n269 0.032697
R8818 avdd.n274 avdd.n273 0.032697
R8819 avdd.n289 avdd.n288 0.032697
R8820 avdd.n215 avdd.n211 0.032697
R8821 avdd.n215 avdd.n214 0.032697
R8822 avdd.n239 avdd.n232 0.032697
R8823 avdd.n8726 avdd.n8725 0.032697
R8824 avdd.n8653 avdd.n8649 0.032697
R8825 avdd.n404 avdd.n399 0.032697
R8826 avdd.n404 avdd.n403 0.032697
R8827 avdd.n419 avdd.n418 0.032697
R8828 avdd.n345 avdd.n341 0.032697
R8829 avdd.n345 avdd.n344 0.032697
R8830 avdd.n369 avdd.n362 0.032697
R8831 avdd.n8640 avdd.n8639 0.032697
R8832 avdd.n8567 avdd.n8563 0.032697
R8833 avdd.n534 avdd.n529 0.032697
R8834 avdd.n534 avdd.n533 0.032697
R8835 avdd.n549 avdd.n548 0.032697
R8836 avdd.n475 avdd.n471 0.032697
R8837 avdd.n475 avdd.n474 0.032697
R8838 avdd.n499 avdd.n492 0.032697
R8839 avdd.n8554 avdd.n8553 0.032697
R8840 avdd.n8481 avdd.n8477 0.032697
R8841 avdd.n664 avdd.n659 0.032697
R8842 avdd.n664 avdd.n663 0.032697
R8843 avdd.n679 avdd.n678 0.032697
R8844 avdd.n605 avdd.n601 0.032697
R8845 avdd.n605 avdd.n604 0.032697
R8846 avdd.n629 avdd.n622 0.032697
R8847 avdd.n8468 avdd.n8467 0.032697
R8848 avdd.n8395 avdd.n8391 0.032697
R8849 avdd.n794 avdd.n789 0.032697
R8850 avdd.n794 avdd.n793 0.032697
R8851 avdd.n809 avdd.n808 0.032697
R8852 avdd.n735 avdd.n731 0.032697
R8853 avdd.n735 avdd.n734 0.032697
R8854 avdd.n759 avdd.n752 0.032697
R8855 avdd.n8382 avdd.n8381 0.032697
R8856 avdd.n8309 avdd.n8305 0.032697
R8857 avdd.n924 avdd.n919 0.032697
R8858 avdd.n924 avdd.n923 0.032697
R8859 avdd.n939 avdd.n938 0.032697
R8860 avdd.n865 avdd.n861 0.032697
R8861 avdd.n865 avdd.n864 0.032697
R8862 avdd.n889 avdd.n882 0.032697
R8863 avdd.n8296 avdd.n8295 0.032697
R8864 avdd.n8223 avdd.n8219 0.032697
R8865 avdd.n1054 avdd.n1049 0.032697
R8866 avdd.n1054 avdd.n1053 0.032697
R8867 avdd.n1069 avdd.n1068 0.032697
R8868 avdd.n995 avdd.n991 0.032697
R8869 avdd.n995 avdd.n994 0.032697
R8870 avdd.n1019 avdd.n1012 0.032697
R8871 avdd.n8210 avdd.n8209 0.032697
R8872 avdd.n8137 avdd.n8133 0.032697
R8873 avdd.n1184 avdd.n1179 0.032697
R8874 avdd.n1184 avdd.n1183 0.032697
R8875 avdd.n1199 avdd.n1198 0.032697
R8876 avdd.n1125 avdd.n1121 0.032697
R8877 avdd.n1125 avdd.n1124 0.032697
R8878 avdd.n1149 avdd.n1142 0.032697
R8879 avdd.n8124 avdd.n8123 0.032697
R8880 avdd.n8051 avdd.n8047 0.032697
R8881 avdd.n1314 avdd.n1309 0.032697
R8882 avdd.n1314 avdd.n1313 0.032697
R8883 avdd.n1329 avdd.n1328 0.032697
R8884 avdd.n1255 avdd.n1251 0.032697
R8885 avdd.n1255 avdd.n1254 0.032697
R8886 avdd.n1279 avdd.n1272 0.032697
R8887 avdd.n8038 avdd.n8037 0.032697
R8888 avdd.n7965 avdd.n7961 0.032697
R8889 avdd.n1444 avdd.n1439 0.032697
R8890 avdd.n1444 avdd.n1443 0.032697
R8891 avdd.n1459 avdd.n1458 0.032697
R8892 avdd.n1385 avdd.n1381 0.032697
R8893 avdd.n1385 avdd.n1384 0.032697
R8894 avdd.n1409 avdd.n1402 0.032697
R8895 avdd.n7952 avdd.n7951 0.032697
R8896 avdd.n7879 avdd.n7875 0.032697
R8897 avdd.n1574 avdd.n1569 0.032697
R8898 avdd.n1574 avdd.n1573 0.032697
R8899 avdd.n1589 avdd.n1588 0.032697
R8900 avdd.n1515 avdd.n1511 0.032697
R8901 avdd.n1515 avdd.n1514 0.032697
R8902 avdd.n1539 avdd.n1532 0.032697
R8903 avdd.n7866 avdd.n7865 0.032697
R8904 avdd.n2087 avdd.n1878 0.0325455
R8905 avdd.n2195 avdd.n2142 0.0325455
R8906 avdd.n2410 avdd.n2357 0.0325455
R8907 avdd.n2625 avdd.n2572 0.0325455
R8908 avdd.n2840 avdd.n2787 0.0325455
R8909 avdd.n3055 avdd.n3002 0.0325455
R8910 avdd.n3376 avdd.n3169 0.0325455
R8911 avdd.n3591 avdd.n3384 0.0325455
R8912 avdd.n3806 avdd.n3599 0.0325455
R8913 avdd.n4021 avdd.n3814 0.0325455
R8914 avdd.n4236 avdd.n4029 0.0325455
R8915 avdd.n4451 avdd.n4244 0.0325455
R8916 avdd.n4866 avdd.n4865 0.0325455
R8917 avdd.n5082 avdd.n5081 0.0325455
R8918 avdd.n5298 avdd.n5297 0.0325455
R8919 avdd.n5514 avdd.n5513 0.0325455
R8920 avdd.n5730 avdd.n5729 0.0325455
R8921 avdd.n5946 avdd.n5945 0.0325455
R8922 avdd.n6162 avdd.n6161 0.0325455
R8923 avdd.n6378 avdd.n6377 0.0325455
R8924 avdd.n6594 avdd.n6593 0.0325455
R8925 avdd.n6810 avdd.n6809 0.0325455
R8926 avdd.n7026 avdd.n7025 0.0325455
R8927 avdd.n7242 avdd.n7241 0.0325455
R8928 avdd.n7762 avdd.n7652 0.0325455
R8929 avdd.n10241 avdd.n10129 0.0325455
R8930 avdd.n10027 avdd.n9965 0.0325455
R8931 avdd.n9913 avdd.n9851 0.0325455
R8932 avdd.n9799 avdd.n9737 0.0325455
R8933 avdd.n9685 avdd.n9624 0.0325455
R8934 avdd.n9571 avdd.n9509 0.0325455
R8935 avdd.n9457 avdd.n9395 0.0325455
R8936 avdd.n9343 avdd.n9281 0.0325455
R8937 avdd.n9229 avdd.n9167 0.0325455
R8938 avdd.n9115 avdd.n9053 0.0325455
R8939 avdd.n9001 avdd.n8939 0.0325455
R8940 avdd.n186 avdd.n73 0.0325455
R8941 avdd.n316 avdd.n203 0.0325455
R8942 avdd.n446 avdd.n333 0.0325455
R8943 avdd.n576 avdd.n463 0.0325455
R8944 avdd.n706 avdd.n593 0.0325455
R8945 avdd.n836 avdd.n723 0.0325455
R8946 avdd.n966 avdd.n853 0.0325455
R8947 avdd.n1096 avdd.n983 0.0325455
R8948 avdd.n1226 avdd.n1113 0.0325455
R8949 avdd.n1356 avdd.n1243 0.0325455
R8950 avdd.n1486 avdd.n1373 0.0325455
R8951 avdd.n1616 avdd.n1503 0.0325455
R8952 avdd.n7739 avdd.n7738 0.0321227
R8953 avdd.n10218 avdd.n10217 0.0321227
R8954 avdd.n4606 avdd.n4588 0.03175
R8955 avdd.n4521 avdd.n4518 0.03175
R8956 avdd.n2068 avdd.n1958 0.0311212
R8957 avdd.n2127 avdd.n2121 0.0311212
R8958 avdd.n2342 avdd.n2336 0.0311212
R8959 avdd.n2557 avdd.n2551 0.0311212
R8960 avdd.n2772 avdd.n2766 0.0311212
R8961 avdd.n2987 avdd.n2981 0.0311212
R8962 avdd.n3357 avdd.n3248 0.0311212
R8963 avdd.n3572 avdd.n3463 0.0311212
R8964 avdd.n3787 avdd.n3678 0.0311212
R8965 avdd.n4002 avdd.n3893 0.0311212
R8966 avdd.n4217 avdd.n4108 0.0311212
R8967 avdd.n4432 avdd.n4323 0.0311212
R8968 avdd.n4849 avdd.n4843 0.0311212
R8969 avdd.n5065 avdd.n5059 0.0311212
R8970 avdd.n5281 avdd.n5275 0.0311212
R8971 avdd.n5497 avdd.n5491 0.0311212
R8972 avdd.n5713 avdd.n5707 0.0311212
R8973 avdd.n5929 avdd.n5923 0.0311212
R8974 avdd.n6145 avdd.n6139 0.0311212
R8975 avdd.n6361 avdd.n6355 0.0311212
R8976 avdd.n6577 avdd.n6571 0.0311212
R8977 avdd.n6793 avdd.n6787 0.0311212
R8978 avdd.n7009 avdd.n7003 0.0311212
R8979 avdd.n7225 avdd.n7219 0.0311212
R8980 avdd.n7667 avdd.n7666 0.0311212
R8981 avdd.n10146 avdd.n10145 0.0311212
R8982 avdd.n9931 avdd.n9930 0.0311212
R8983 avdd.n9817 avdd.n9816 0.0311212
R8984 avdd.n9703 avdd.n9702 0.0311212
R8985 avdd.n9590 avdd.n9589 0.0311212
R8986 avdd.n9475 avdd.n9474 0.0311212
R8987 avdd.n9361 avdd.n9360 0.0311212
R8988 avdd.n9247 avdd.n9246 0.0311212
R8989 avdd.n9133 avdd.n9132 0.0311212
R8990 avdd.n9019 avdd.n9018 0.0311212
R8991 avdd.n8905 avdd.n8904 0.0311212
R8992 avdd.n150 avdd.n149 0.0311212
R8993 avdd.n280 avdd.n279 0.0311212
R8994 avdd.n410 avdd.n409 0.0311212
R8995 avdd.n540 avdd.n539 0.0311212
R8996 avdd.n670 avdd.n669 0.0311212
R8997 avdd.n800 avdd.n799 0.0311212
R8998 avdd.n930 avdd.n929 0.0311212
R8999 avdd.n1060 avdd.n1059 0.0311212
R9000 avdd.n1190 avdd.n1189 0.0311212
R9001 avdd.n1320 avdd.n1319 0.0311212
R9002 avdd.n1450 avdd.n1449 0.0311212
R9003 avdd.n1580 avdd.n1579 0.0311212
R9004 avdd.n1924 avdd.n1923 0.029697
R9005 avdd.n2055 avdd.n2054 0.029697
R9006 avdd.n2178 avdd.n2177 0.029697
R9007 avdd.n2249 avdd.n2248 0.029697
R9008 avdd.n2393 avdd.n2392 0.029697
R9009 avdd.n2464 avdd.n2463 0.029697
R9010 avdd.n2608 avdd.n2607 0.029697
R9011 avdd.n2679 avdd.n2678 0.029697
R9012 avdd.n2823 avdd.n2822 0.029697
R9013 avdd.n2894 avdd.n2893 0.029697
R9014 avdd.n3038 avdd.n3037 0.029697
R9015 avdd.n3109 avdd.n3108 0.029697
R9016 avdd.n3214 avdd.n3213 0.029697
R9017 avdd.n3344 avdd.n3343 0.029697
R9018 avdd.n3429 avdd.n3428 0.029697
R9019 avdd.n3559 avdd.n3558 0.029697
R9020 avdd.n3644 avdd.n3643 0.029697
R9021 avdd.n3774 avdd.n3773 0.029697
R9022 avdd.n3859 avdd.n3858 0.029697
R9023 avdd.n3989 avdd.n3988 0.029697
R9024 avdd.n4074 avdd.n4073 0.029697
R9025 avdd.n4204 avdd.n4203 0.029697
R9026 avdd.n4289 avdd.n4288 0.029697
R9027 avdd.n4419 avdd.n4418 0.029697
R9028 avdd.n4900 avdd.n4899 0.029697
R9029 avdd.n4971 avdd.n4970 0.029697
R9030 avdd.n5116 avdd.n5115 0.029697
R9031 avdd.n5187 avdd.n5186 0.029697
R9032 avdd.n5332 avdd.n5331 0.029697
R9033 avdd.n5403 avdd.n5402 0.029697
R9034 avdd.n5548 avdd.n5547 0.029697
R9035 avdd.n5619 avdd.n5618 0.029697
R9036 avdd.n5764 avdd.n5763 0.029697
R9037 avdd.n5835 avdd.n5834 0.029697
R9038 avdd.n5980 avdd.n5979 0.029697
R9039 avdd.n6051 avdd.n6050 0.029697
R9040 avdd.n6196 avdd.n6195 0.029697
R9041 avdd.n6267 avdd.n6266 0.029697
R9042 avdd.n6412 avdd.n6411 0.029697
R9043 avdd.n6483 avdd.n6482 0.029697
R9044 avdd.n6628 avdd.n6627 0.029697
R9045 avdd.n6699 avdd.n6698 0.029697
R9046 avdd.n6844 avdd.n6843 0.029697
R9047 avdd.n6915 avdd.n6914 0.029697
R9048 avdd.n7060 avdd.n7059 0.029697
R9049 avdd.n7131 avdd.n7130 0.029697
R9050 avdd.n7276 avdd.n7275 0.029697
R9051 avdd.n7347 avdd.n7346 0.029697
R9052 avdd.n7703 avdd.n7702 0.029697
R9053 avdd.n7796 avdd.n7795 0.029697
R9054 avdd.n10182 avdd.n10181 0.029697
R9055 avdd.n10055 avdd.n10054 0.029697
R9056 avdd.n10285 avdd.n10284 0.029697
R9057 avdd.n10387 avdd.n10386 0.029697
R9058 avdd.n10489 avdd.n10488 0.029697
R9059 avdd.n10591 avdd.n10590 0.029697
R9060 avdd.n10693 avdd.n10692 0.029697
R9061 avdd.n10795 avdd.n10794 0.029697
R9062 avdd.n10897 avdd.n10896 0.029697
R9063 avdd.n10999 avdd.n10998 0.029697
R9064 avdd.n11101 avdd.n11100 0.029697
R9065 avdd.n11203 avdd.n11202 0.029697
R9066 avdd.n97 avdd.n96 0.029697
R9067 avdd.n8818 avdd.n8817 0.029697
R9068 avdd.n227 avdd.n226 0.029697
R9069 avdd.n8732 avdd.n8731 0.029697
R9070 avdd.n357 avdd.n356 0.029697
R9071 avdd.n8646 avdd.n8645 0.029697
R9072 avdd.n487 avdd.n486 0.029697
R9073 avdd.n8560 avdd.n8559 0.029697
R9074 avdd.n617 avdd.n616 0.029697
R9075 avdd.n8474 avdd.n8473 0.029697
R9076 avdd.n747 avdd.n746 0.029697
R9077 avdd.n8388 avdd.n8387 0.029697
R9078 avdd.n877 avdd.n876 0.029697
R9079 avdd.n8302 avdd.n8301 0.029697
R9080 avdd.n1007 avdd.n1006 0.029697
R9081 avdd.n8216 avdd.n8215 0.029697
R9082 avdd.n1137 avdd.n1136 0.029697
R9083 avdd.n8130 avdd.n8129 0.029697
R9084 avdd.n1267 avdd.n1266 0.029697
R9085 avdd.n8044 avdd.n8043 0.029697
R9086 avdd.n1397 avdd.n1396 0.029697
R9087 avdd.n7958 avdd.n7957 0.029697
R9088 avdd.n1527 avdd.n1526 0.029697
R9089 avdd.n7872 avdd.n7871 0.029697
R9090 avdd.n2036 avdd.n2035 0.0289848
R9091 avdd.n2274 avdd.n2093 0.0289848
R9092 avdd.n2489 avdd.n2308 0.0289848
R9093 avdd.n2704 avdd.n2523 0.0289848
R9094 avdd.n2919 avdd.n2738 0.0289848
R9095 avdd.n3134 avdd.n2953 0.0289848
R9096 avdd.n3325 avdd.n3295 0.0289848
R9097 avdd.n3540 avdd.n3510 0.0289848
R9098 avdd.n3755 avdd.n3725 0.0289848
R9099 avdd.n3970 avdd.n3940 0.0289848
R9100 avdd.n4185 avdd.n4155 0.0289848
R9101 avdd.n4400 avdd.n4370 0.0289848
R9102 avdd.n5021 avdd.n4813 0.0289848
R9103 avdd.n5237 avdd.n5029 0.0289848
R9104 avdd.n5453 avdd.n5245 0.0289848
R9105 avdd.n5669 avdd.n5461 0.0289848
R9106 avdd.n5885 avdd.n5677 0.0289848
R9107 avdd.n6101 avdd.n5893 0.0289848
R9108 avdd.n6317 avdd.n6109 0.0289848
R9109 avdd.n6533 avdd.n6325 0.0289848
R9110 avdd.n6749 avdd.n6541 0.0289848
R9111 avdd.n6965 avdd.n6757 0.0289848
R9112 avdd.n7181 avdd.n6973 0.0289848
R9113 avdd.n7397 avdd.n7189 0.0289848
R9114 avdd.n7852 avdd.n7781 0.0289848
R9115 avdd.n10110 avdd.n10041 0.0289848
R9116 avdd.n10342 avdd.n10257 0.0289848
R9117 avdd.n10444 avdd.n10359 0.0289848
R9118 avdd.n10546 avdd.n10461 0.0289848
R9119 avdd.n10648 avdd.n10563 0.0289848
R9120 avdd.n10750 avdd.n10665 0.0289848
R9121 avdd.n10852 avdd.n10767 0.0289848
R9122 avdd.n10954 avdd.n10869 0.0289848
R9123 avdd.n11056 avdd.n10971 0.0289848
R9124 avdd.n11158 avdd.n11073 0.0289848
R9125 avdd.n11260 avdd.n11175 0.0289848
R9126 avdd.n8885 avdd.n8884 0.0289848
R9127 avdd.n8799 avdd.n8798 0.0289848
R9128 avdd.n8713 avdd.n8712 0.0289848
R9129 avdd.n8627 avdd.n8626 0.0289848
R9130 avdd.n8541 avdd.n8540 0.0289848
R9131 avdd.n8455 avdd.n8454 0.0289848
R9132 avdd.n8369 avdd.n8368 0.0289848
R9133 avdd.n8283 avdd.n8282 0.0289848
R9134 avdd.n8197 avdd.n8196 0.0289848
R9135 avdd.n8111 avdd.n8110 0.0289848
R9136 avdd.n8025 avdd.n8024 0.0289848
R9137 avdd.n7939 avdd.n7938 0.0289848
R9138 avdd.n2043 avdd.n1999 0.0289091
R9139 avdd.n1942 avdd.n1890 0.0289091
R9140 avdd.n1913 avdd.n1912 0.0289091
R9141 avdd.n1911 avdd.n1901 0.0289091
R9142 avdd.n1917 avdd.n1892 0.0289091
R9143 avdd.n2263 avdd.n2104 0.0289091
R9144 avdd.n2187 avdd.n2137 0.0289091
R9145 avdd.n2167 avdd.n2166 0.0289091
R9146 avdd.n2165 avdd.n2155 0.0289091
R9147 avdd.n2171 avdd.n2147 0.0289091
R9148 avdd.n2478 avdd.n2319 0.0289091
R9149 avdd.n2402 avdd.n2352 0.0289091
R9150 avdd.n2382 avdd.n2381 0.0289091
R9151 avdd.n2380 avdd.n2370 0.0289091
R9152 avdd.n2386 avdd.n2362 0.0289091
R9153 avdd.n2693 avdd.n2534 0.0289091
R9154 avdd.n2617 avdd.n2567 0.0289091
R9155 avdd.n2597 avdd.n2596 0.0289091
R9156 avdd.n2595 avdd.n2585 0.0289091
R9157 avdd.n2601 avdd.n2577 0.0289091
R9158 avdd.n2908 avdd.n2749 0.0289091
R9159 avdd.n2832 avdd.n2782 0.0289091
R9160 avdd.n2812 avdd.n2811 0.0289091
R9161 avdd.n2810 avdd.n2800 0.0289091
R9162 avdd.n2816 avdd.n2792 0.0289091
R9163 avdd.n3123 avdd.n2964 0.0289091
R9164 avdd.n3047 avdd.n2997 0.0289091
R9165 avdd.n3027 avdd.n3026 0.0289091
R9166 avdd.n3025 avdd.n3015 0.0289091
R9167 avdd.n3031 avdd.n3007 0.0289091
R9168 avdd.n3332 avdd.n3289 0.0289091
R9169 avdd.n3232 avdd.n3180 0.0289091
R9170 avdd.n3203 avdd.n3202 0.0289091
R9171 avdd.n3201 avdd.n3191 0.0289091
R9172 avdd.n3207 avdd.n3182 0.0289091
R9173 avdd.n3547 avdd.n3504 0.0289091
R9174 avdd.n3447 avdd.n3395 0.0289091
R9175 avdd.n3418 avdd.n3417 0.0289091
R9176 avdd.n3416 avdd.n3406 0.0289091
R9177 avdd.n3422 avdd.n3397 0.0289091
R9178 avdd.n3762 avdd.n3719 0.0289091
R9179 avdd.n3662 avdd.n3610 0.0289091
R9180 avdd.n3633 avdd.n3632 0.0289091
R9181 avdd.n3631 avdd.n3621 0.0289091
R9182 avdd.n3637 avdd.n3612 0.0289091
R9183 avdd.n3977 avdd.n3934 0.0289091
R9184 avdd.n3877 avdd.n3825 0.0289091
R9185 avdd.n3848 avdd.n3847 0.0289091
R9186 avdd.n3846 avdd.n3836 0.0289091
R9187 avdd.n3852 avdd.n3827 0.0289091
R9188 avdd.n4192 avdd.n4149 0.0289091
R9189 avdd.n4092 avdd.n4040 0.0289091
R9190 avdd.n4063 avdd.n4062 0.0289091
R9191 avdd.n4061 avdd.n4051 0.0289091
R9192 avdd.n4067 avdd.n4042 0.0289091
R9193 avdd.n4407 avdd.n4364 0.0289091
R9194 avdd.n4307 avdd.n4255 0.0289091
R9195 avdd.n4278 avdd.n4277 0.0289091
R9196 avdd.n4276 avdd.n4266 0.0289091
R9197 avdd.n4282 avdd.n4257 0.0289091
R9198 avdd.n4889 avdd.n4888 0.0289091
R9199 avdd.n4910 avdd.n4859 0.0289091
R9200 avdd.n4985 avdd.n4825 0.0289091
R9201 avdd.n4887 avdd.n4877 0.0289091
R9202 avdd.n4893 avdd.n4869 0.0289091
R9203 avdd.n5105 avdd.n5104 0.0289091
R9204 avdd.n5126 avdd.n5075 0.0289091
R9205 avdd.n5201 avdd.n5041 0.0289091
R9206 avdd.n5103 avdd.n5093 0.0289091
R9207 avdd.n5109 avdd.n5085 0.0289091
R9208 avdd.n5321 avdd.n5320 0.0289091
R9209 avdd.n5342 avdd.n5291 0.0289091
R9210 avdd.n5417 avdd.n5257 0.0289091
R9211 avdd.n5319 avdd.n5309 0.0289091
R9212 avdd.n5325 avdd.n5301 0.0289091
R9213 avdd.n5537 avdd.n5536 0.0289091
R9214 avdd.n5558 avdd.n5507 0.0289091
R9215 avdd.n5633 avdd.n5473 0.0289091
R9216 avdd.n5535 avdd.n5525 0.0289091
R9217 avdd.n5541 avdd.n5517 0.0289091
R9218 avdd.n5753 avdd.n5752 0.0289091
R9219 avdd.n5774 avdd.n5723 0.0289091
R9220 avdd.n5849 avdd.n5689 0.0289091
R9221 avdd.n5751 avdd.n5741 0.0289091
R9222 avdd.n5757 avdd.n5733 0.0289091
R9223 avdd.n5969 avdd.n5968 0.0289091
R9224 avdd.n5990 avdd.n5939 0.0289091
R9225 avdd.n6065 avdd.n5905 0.0289091
R9226 avdd.n5967 avdd.n5957 0.0289091
R9227 avdd.n5973 avdd.n5949 0.0289091
R9228 avdd.n6185 avdd.n6184 0.0289091
R9229 avdd.n6206 avdd.n6155 0.0289091
R9230 avdd.n6281 avdd.n6121 0.0289091
R9231 avdd.n6183 avdd.n6173 0.0289091
R9232 avdd.n6189 avdd.n6165 0.0289091
R9233 avdd.n6401 avdd.n6400 0.0289091
R9234 avdd.n6422 avdd.n6371 0.0289091
R9235 avdd.n6497 avdd.n6337 0.0289091
R9236 avdd.n6399 avdd.n6389 0.0289091
R9237 avdd.n6405 avdd.n6381 0.0289091
R9238 avdd.n6617 avdd.n6616 0.0289091
R9239 avdd.n6638 avdd.n6587 0.0289091
R9240 avdd.n6713 avdd.n6553 0.0289091
R9241 avdd.n6615 avdd.n6605 0.0289091
R9242 avdd.n6621 avdd.n6597 0.0289091
R9243 avdd.n6833 avdd.n6832 0.0289091
R9244 avdd.n6854 avdd.n6803 0.0289091
R9245 avdd.n6929 avdd.n6769 0.0289091
R9246 avdd.n6831 avdd.n6821 0.0289091
R9247 avdd.n6837 avdd.n6813 0.0289091
R9248 avdd.n7049 avdd.n7048 0.0289091
R9249 avdd.n7070 avdd.n7019 0.0289091
R9250 avdd.n7145 avdd.n6985 0.0289091
R9251 avdd.n7047 avdd.n7037 0.0289091
R9252 avdd.n7053 avdd.n7029 0.0289091
R9253 avdd.n7265 avdd.n7264 0.0289091
R9254 avdd.n7286 avdd.n7235 0.0289091
R9255 avdd.n7361 avdd.n7201 0.0289091
R9256 avdd.n7263 avdd.n7253 0.0289091
R9257 avdd.n7269 avdd.n7245 0.0289091
R9258 avdd.n7751 avdd.n7750 0.0289091
R9259 avdd.n7734 avdd.n7733 0.0289091
R9260 avdd.n7824 avdd.n7823 0.0289091
R9261 avdd.n7747 avdd.n7746 0.0289091
R9262 avdd.n7711 avdd.n7710 0.0289091
R9263 avdd.n10230 avdd.n10229 0.0289091
R9264 avdd.n10213 avdd.n10212 0.0289091
R9265 avdd.n10082 avdd.n10081 0.0289091
R9266 avdd.n10226 avdd.n10225 0.0289091
R9267 avdd.n10190 avdd.n10189 0.0289091
R9268 avdd.n9984 avdd.n9983 0.0289091
R9269 avdd.n10019 avdd.n10018 0.0289091
R9270 avdd.n10314 avdd.n10313 0.0289091
R9271 avdd.n9976 avdd.n9975 0.0289091
R9272 avdd.n9972 avdd.n9971 0.0289091
R9273 avdd.n9870 avdd.n9869 0.0289091
R9274 avdd.n9905 avdd.n9904 0.0289091
R9275 avdd.n10416 avdd.n10415 0.0289091
R9276 avdd.n9862 avdd.n9861 0.0289091
R9277 avdd.n9858 avdd.n9857 0.0289091
R9278 avdd.n9756 avdd.n9755 0.0289091
R9279 avdd.n9791 avdd.n9790 0.0289091
R9280 avdd.n10518 avdd.n10517 0.0289091
R9281 avdd.n9748 avdd.n9747 0.0289091
R9282 avdd.n9744 avdd.n9743 0.0289091
R9283 avdd.n9643 avdd.n9642 0.0289091
R9284 avdd.n9678 avdd.n9677 0.0289091
R9285 avdd.n10620 avdd.n10619 0.0289091
R9286 avdd.n9635 avdd.n9634 0.0289091
R9287 avdd.n9631 avdd.n9630 0.0289091
R9288 avdd.n9528 avdd.n9527 0.0289091
R9289 avdd.n9563 avdd.n9562 0.0289091
R9290 avdd.n10722 avdd.n10721 0.0289091
R9291 avdd.n9520 avdd.n9519 0.0289091
R9292 avdd.n9516 avdd.n9515 0.0289091
R9293 avdd.n9414 avdd.n9413 0.0289091
R9294 avdd.n9449 avdd.n9448 0.0289091
R9295 avdd.n10824 avdd.n10823 0.0289091
R9296 avdd.n9406 avdd.n9405 0.0289091
R9297 avdd.n9402 avdd.n9401 0.0289091
R9298 avdd.n9300 avdd.n9299 0.0289091
R9299 avdd.n9335 avdd.n9334 0.0289091
R9300 avdd.n10926 avdd.n10925 0.0289091
R9301 avdd.n9292 avdd.n9291 0.0289091
R9302 avdd.n9288 avdd.n9287 0.0289091
R9303 avdd.n9186 avdd.n9185 0.0289091
R9304 avdd.n9221 avdd.n9220 0.0289091
R9305 avdd.n11028 avdd.n11027 0.0289091
R9306 avdd.n9178 avdd.n9177 0.0289091
R9307 avdd.n9174 avdd.n9173 0.0289091
R9308 avdd.n9072 avdd.n9071 0.0289091
R9309 avdd.n9107 avdd.n9106 0.0289091
R9310 avdd.n11130 avdd.n11129 0.0289091
R9311 avdd.n9064 avdd.n9063 0.0289091
R9312 avdd.n9060 avdd.n9059 0.0289091
R9313 avdd.n8958 avdd.n8957 0.0289091
R9314 avdd.n8993 avdd.n8992 0.0289091
R9315 avdd.n11232 avdd.n11231 0.0289091
R9316 avdd.n8950 avdd.n8949 0.0289091
R9317 avdd.n8946 avdd.n8945 0.0289091
R9318 avdd.n8845 avdd.n8844 0.0289091
R9319 avdd.n129 avdd.n128 0.0289091
R9320 avdd.n84 avdd.n83 0.0289091
R9321 avdd.n80 avdd.n79 0.0289091
R9322 avdd.n105 avdd.n104 0.0289091
R9323 avdd.n8759 avdd.n8758 0.0289091
R9324 avdd.n259 avdd.n258 0.0289091
R9325 avdd.n214 avdd.n213 0.0289091
R9326 avdd.n210 avdd.n209 0.0289091
R9327 avdd.n235 avdd.n234 0.0289091
R9328 avdd.n8673 avdd.n8672 0.0289091
R9329 avdd.n389 avdd.n388 0.0289091
R9330 avdd.n344 avdd.n343 0.0289091
R9331 avdd.n340 avdd.n339 0.0289091
R9332 avdd.n365 avdd.n364 0.0289091
R9333 avdd.n8587 avdd.n8586 0.0289091
R9334 avdd.n519 avdd.n518 0.0289091
R9335 avdd.n474 avdd.n473 0.0289091
R9336 avdd.n470 avdd.n469 0.0289091
R9337 avdd.n495 avdd.n494 0.0289091
R9338 avdd.n8501 avdd.n8500 0.0289091
R9339 avdd.n649 avdd.n648 0.0289091
R9340 avdd.n604 avdd.n603 0.0289091
R9341 avdd.n600 avdd.n599 0.0289091
R9342 avdd.n625 avdd.n624 0.0289091
R9343 avdd.n8415 avdd.n8414 0.0289091
R9344 avdd.n779 avdd.n778 0.0289091
R9345 avdd.n734 avdd.n733 0.0289091
R9346 avdd.n730 avdd.n729 0.0289091
R9347 avdd.n755 avdd.n754 0.0289091
R9348 avdd.n8329 avdd.n8328 0.0289091
R9349 avdd.n909 avdd.n908 0.0289091
R9350 avdd.n864 avdd.n863 0.0289091
R9351 avdd.n860 avdd.n859 0.0289091
R9352 avdd.n885 avdd.n884 0.0289091
R9353 avdd.n8243 avdd.n8242 0.0289091
R9354 avdd.n1039 avdd.n1038 0.0289091
R9355 avdd.n994 avdd.n993 0.0289091
R9356 avdd.n990 avdd.n989 0.0289091
R9357 avdd.n1015 avdd.n1014 0.0289091
R9358 avdd.n8157 avdd.n8156 0.0289091
R9359 avdd.n1169 avdd.n1168 0.0289091
R9360 avdd.n1124 avdd.n1123 0.0289091
R9361 avdd.n1120 avdd.n1119 0.0289091
R9362 avdd.n1145 avdd.n1144 0.0289091
R9363 avdd.n8071 avdd.n8070 0.0289091
R9364 avdd.n1299 avdd.n1298 0.0289091
R9365 avdd.n1254 avdd.n1253 0.0289091
R9366 avdd.n1250 avdd.n1249 0.0289091
R9367 avdd.n1275 avdd.n1274 0.0289091
R9368 avdd.n7985 avdd.n7984 0.0289091
R9369 avdd.n1429 avdd.n1428 0.0289091
R9370 avdd.n1384 avdd.n1383 0.0289091
R9371 avdd.n1380 avdd.n1379 0.0289091
R9372 avdd.n1405 avdd.n1404 0.0289091
R9373 avdd.n7899 avdd.n7898 0.0289091
R9374 avdd.n1559 avdd.n1558 0.0289091
R9375 avdd.n1514 avdd.n1513 0.0289091
R9376 avdd.n1510 avdd.n1509 0.0289091
R9377 avdd.n1535 avdd.n1534 0.0289091
R9378 avdd.n4594 avdd.n4517 0.0275833
R9379 avdd.n7445 avdd.n7444 0.0272435
R9380 avdd.n7484 avdd.n7483 0.0272435
R9381 avdd.n7544 avdd.n7543 0.0272435
R9382 avdd.n7584 avdd.n7583 0.0272435
R9383 avdd.n2085 avdd.n1883 0.0261364
R9384 avdd.n2046 avdd.n2045 0.0261364
R9385 avdd.n2217 avdd.n2208 0.0261364
R9386 avdd.n2271 avdd.n2270 0.0261364
R9387 avdd.n2432 avdd.n2423 0.0261364
R9388 avdd.n2486 avdd.n2485 0.0261364
R9389 avdd.n2647 avdd.n2638 0.0261364
R9390 avdd.n2701 avdd.n2700 0.0261364
R9391 avdd.n2862 avdd.n2853 0.0261364
R9392 avdd.n2916 avdd.n2915 0.0261364
R9393 avdd.n3077 avdd.n3068 0.0261364
R9394 avdd.n3131 avdd.n3130 0.0261364
R9395 avdd.n3374 avdd.n3173 0.0261364
R9396 avdd.n3335 avdd.n3334 0.0261364
R9397 avdd.n3589 avdd.n3388 0.0261364
R9398 avdd.n3550 avdd.n3549 0.0261364
R9399 avdd.n3804 avdd.n3603 0.0261364
R9400 avdd.n3765 avdd.n3764 0.0261364
R9401 avdd.n4019 avdd.n3818 0.0261364
R9402 avdd.n3980 avdd.n3979 0.0261364
R9403 avdd.n4234 avdd.n4033 0.0261364
R9404 avdd.n4195 avdd.n4194 0.0261364
R9405 avdd.n4449 avdd.n4248 0.0261364
R9406 avdd.n4410 avdd.n4409 0.0261364
R9407 avdd.n4939 avdd.n4930 0.0261364
R9408 avdd.n4993 avdd.n4992 0.0261364
R9409 avdd.n5155 avdd.n5146 0.0261364
R9410 avdd.n5209 avdd.n5208 0.0261364
R9411 avdd.n5371 avdd.n5362 0.0261364
R9412 avdd.n5425 avdd.n5424 0.0261364
R9413 avdd.n5587 avdd.n5578 0.0261364
R9414 avdd.n5641 avdd.n5640 0.0261364
R9415 avdd.n5803 avdd.n5794 0.0261364
R9416 avdd.n5857 avdd.n5856 0.0261364
R9417 avdd.n6019 avdd.n6010 0.0261364
R9418 avdd.n6073 avdd.n6072 0.0261364
R9419 avdd.n6235 avdd.n6226 0.0261364
R9420 avdd.n6289 avdd.n6288 0.0261364
R9421 avdd.n6451 avdd.n6442 0.0261364
R9422 avdd.n6505 avdd.n6504 0.0261364
R9423 avdd.n6667 avdd.n6658 0.0261364
R9424 avdd.n6721 avdd.n6720 0.0261364
R9425 avdd.n6883 avdd.n6874 0.0261364
R9426 avdd.n6937 avdd.n6936 0.0261364
R9427 avdd.n7099 avdd.n7090 0.0261364
R9428 avdd.n7153 avdd.n7152 0.0261364
R9429 avdd.n7315 avdd.n7306 0.0261364
R9430 avdd.n7369 avdd.n7368 0.0261364
R9431 avdd.n7650 avdd.n7649 0.0261364
R9432 avdd.n7778 avdd.n7777 0.0261364
R9433 avdd.n10127 avdd.n10126 0.0261364
R9434 avdd.n10038 avdd.n10037 0.0261364
R9435 avdd.n9928 avdd.n9927 0.0261364
R9436 avdd.n10254 avdd.n10253 0.0261364
R9437 avdd.n9814 avdd.n9813 0.0261364
R9438 avdd.n10356 avdd.n10355 0.0261364
R9439 avdd.n9700 avdd.n9699 0.0261364
R9440 avdd.n10458 avdd.n10457 0.0261364
R9441 avdd.n9586 avdd.n9585 0.0261364
R9442 avdd.n10560 avdd.n10559 0.0261364
R9443 avdd.n9472 avdd.n9471 0.0261364
R9444 avdd.n10662 avdd.n10661 0.0261364
R9445 avdd.n9358 avdd.n9357 0.0261364
R9446 avdd.n10764 avdd.n10763 0.0261364
R9447 avdd.n9244 avdd.n9243 0.0261364
R9448 avdd.n10866 avdd.n10865 0.0261364
R9449 avdd.n9130 avdd.n9129 0.0261364
R9450 avdd.n10968 avdd.n10967 0.0261364
R9451 avdd.n9016 avdd.n9015 0.0261364
R9452 avdd.n11070 avdd.n11069 0.0261364
R9453 avdd.n8902 avdd.n8901 0.0261364
R9454 avdd.n11172 avdd.n11171 0.0261364
R9455 avdd.n71 avdd.n70 0.0261364
R9456 avdd.n8881 avdd.n8880 0.0261364
R9457 avdd.n201 avdd.n200 0.0261364
R9458 avdd.n8795 avdd.n8794 0.0261364
R9459 avdd.n331 avdd.n330 0.0261364
R9460 avdd.n8709 avdd.n8708 0.0261364
R9461 avdd.n461 avdd.n460 0.0261364
R9462 avdd.n8623 avdd.n8622 0.0261364
R9463 avdd.n591 avdd.n590 0.0261364
R9464 avdd.n8537 avdd.n8536 0.0261364
R9465 avdd.n721 avdd.n720 0.0261364
R9466 avdd.n8451 avdd.n8450 0.0261364
R9467 avdd.n851 avdd.n850 0.0261364
R9468 avdd.n8365 avdd.n8364 0.0261364
R9469 avdd.n981 avdd.n980 0.0261364
R9470 avdd.n8279 avdd.n8278 0.0261364
R9471 avdd.n1111 avdd.n1110 0.0261364
R9472 avdd.n8193 avdd.n8192 0.0261364
R9473 avdd.n1241 avdd.n1240 0.0261364
R9474 avdd.n8107 avdd.n8106 0.0261364
R9475 avdd.n1371 avdd.n1370 0.0261364
R9476 avdd.n8021 avdd.n8020 0.0261364
R9477 avdd.n1501 avdd.n1500 0.0261364
R9478 avdd.n7935 avdd.n7934 0.0261364
R9479 avdd.n4626 avdd.n4624 0.0255
R9480 avdd.n2013 avdd.n2001 0.0251212
R9481 avdd.n2083 avdd.n2082 0.0251212
R9482 avdd.n2286 avdd.n2285 0.0251212
R9483 avdd.n2206 avdd.n2205 0.0251212
R9484 avdd.n2501 avdd.n2500 0.0251212
R9485 avdd.n2421 avdd.n2420 0.0251212
R9486 avdd.n2716 avdd.n2715 0.0251212
R9487 avdd.n2636 avdd.n2635 0.0251212
R9488 avdd.n2931 avdd.n2930 0.0251212
R9489 avdd.n2851 avdd.n2850 0.0251212
R9490 avdd.n3146 avdd.n3145 0.0251212
R9491 avdd.n3066 avdd.n3065 0.0251212
R9492 avdd.n3306 avdd.n3291 0.0251212
R9493 avdd.n3372 avdd.n3371 0.0251212
R9494 avdd.n3521 avdd.n3506 0.0251212
R9495 avdd.n3587 avdd.n3586 0.0251212
R9496 avdd.n3736 avdd.n3721 0.0251212
R9497 avdd.n3802 avdd.n3801 0.0251212
R9498 avdd.n3951 avdd.n3936 0.0251212
R9499 avdd.n4017 avdd.n4016 0.0251212
R9500 avdd.n4166 avdd.n4151 0.0251212
R9501 avdd.n4232 avdd.n4231 0.0251212
R9502 avdd.n4381 avdd.n4366 0.0251212
R9503 avdd.n4447 avdd.n4446 0.0251212
R9504 avdd.n4928 avdd.n4927 0.0251212
R9505 avdd.n5004 avdd.n5003 0.0251212
R9506 avdd.n5144 avdd.n5143 0.0251212
R9507 avdd.n5220 avdd.n5219 0.0251212
R9508 avdd.n5360 avdd.n5359 0.0251212
R9509 avdd.n5436 avdd.n5435 0.0251212
R9510 avdd.n5576 avdd.n5575 0.0251212
R9511 avdd.n5652 avdd.n5651 0.0251212
R9512 avdd.n5792 avdd.n5791 0.0251212
R9513 avdd.n5868 avdd.n5867 0.0251212
R9514 avdd.n6008 avdd.n6007 0.0251212
R9515 avdd.n6084 avdd.n6083 0.0251212
R9516 avdd.n6224 avdd.n6223 0.0251212
R9517 avdd.n6300 avdd.n6299 0.0251212
R9518 avdd.n6440 avdd.n6439 0.0251212
R9519 avdd.n6516 avdd.n6515 0.0251212
R9520 avdd.n6656 avdd.n6655 0.0251212
R9521 avdd.n6732 avdd.n6731 0.0251212
R9522 avdd.n6872 avdd.n6871 0.0251212
R9523 avdd.n6948 avdd.n6947 0.0251212
R9524 avdd.n7088 avdd.n7087 0.0251212
R9525 avdd.n7164 avdd.n7163 0.0251212
R9526 avdd.n7304 avdd.n7303 0.0251212
R9527 avdd.n7380 avdd.n7379 0.0251212
R9528 avdd.n7696 avdd.n7692 0.0251212
R9529 avdd.n7843 avdd.n7839 0.0251212
R9530 avdd.n10175 avdd.n10171 0.0251212
R9531 avdd.n10101 avdd.n10097 0.0251212
R9532 avdd.n9959 avdd.n9955 0.0251212
R9533 avdd.n10333 avdd.n10329 0.0251212
R9534 avdd.n9845 avdd.n9841 0.0251212
R9535 avdd.n10435 avdd.n10431 0.0251212
R9536 avdd.n9731 avdd.n9727 0.0251212
R9537 avdd.n10537 avdd.n10533 0.0251212
R9538 avdd.n9618 avdd.n9614 0.0251212
R9539 avdd.n10639 avdd.n10635 0.0251212
R9540 avdd.n9503 avdd.n9499 0.0251212
R9541 avdd.n10741 avdd.n10737 0.0251212
R9542 avdd.n9389 avdd.n9385 0.0251212
R9543 avdd.n10843 avdd.n10839 0.0251212
R9544 avdd.n9275 avdd.n9271 0.0251212
R9545 avdd.n10945 avdd.n10941 0.0251212
R9546 avdd.n9161 avdd.n9157 0.0251212
R9547 avdd.n11047 avdd.n11043 0.0251212
R9548 avdd.n9047 avdd.n9043 0.0251212
R9549 avdd.n11149 avdd.n11145 0.0251212
R9550 avdd.n8933 avdd.n8929 0.0251212
R9551 avdd.n11251 avdd.n11247 0.0251212
R9552 avdd.n8864 avdd.n8860 0.0251212
R9553 avdd.n179 avdd.n175 0.0251212
R9554 avdd.n8778 avdd.n8774 0.0251212
R9555 avdd.n309 avdd.n305 0.0251212
R9556 avdd.n8692 avdd.n8688 0.0251212
R9557 avdd.n439 avdd.n435 0.0251212
R9558 avdd.n8606 avdd.n8602 0.0251212
R9559 avdd.n569 avdd.n565 0.0251212
R9560 avdd.n8520 avdd.n8516 0.0251212
R9561 avdd.n699 avdd.n695 0.0251212
R9562 avdd.n8434 avdd.n8430 0.0251212
R9563 avdd.n829 avdd.n825 0.0251212
R9564 avdd.n8348 avdd.n8344 0.0251212
R9565 avdd.n959 avdd.n955 0.0251212
R9566 avdd.n8262 avdd.n8258 0.0251212
R9567 avdd.n1089 avdd.n1085 0.0251212
R9568 avdd.n8176 avdd.n8172 0.0251212
R9569 avdd.n1219 avdd.n1215 0.0251212
R9570 avdd.n8090 avdd.n8086 0.0251212
R9571 avdd.n1349 avdd.n1345 0.0251212
R9572 avdd.n8004 avdd.n8000 0.0251212
R9573 avdd.n1479 avdd.n1475 0.0251212
R9574 avdd.n7918 avdd.n7914 0.0251212
R9575 avdd.n1609 avdd.n1605 0.0251212
R9576 avdd.n2074 avdd.n1948 0.0232273
R9577 avdd.n2027 avdd.n2026 0.0232273
R9578 avdd.n2226 avdd.n2125 0.0232273
R9579 avdd.n2300 avdd.n2099 0.0232273
R9580 avdd.n2441 avdd.n2340 0.0232273
R9581 avdd.n2515 avdd.n2314 0.0232273
R9582 avdd.n2656 avdd.n2555 0.0232273
R9583 avdd.n2730 avdd.n2529 0.0232273
R9584 avdd.n2871 avdd.n2770 0.0232273
R9585 avdd.n2945 avdd.n2744 0.0232273
R9586 avdd.n3086 avdd.n2985 0.0232273
R9587 avdd.n3160 avdd.n2959 0.0232273
R9588 avdd.n3363 avdd.n3238 0.0232273
R9589 avdd.n3321 avdd.n3320 0.0232273
R9590 avdd.n3578 avdd.n3453 0.0232273
R9591 avdd.n3536 avdd.n3535 0.0232273
R9592 avdd.n3793 avdd.n3668 0.0232273
R9593 avdd.n3751 avdd.n3750 0.0232273
R9594 avdd.n4008 avdd.n3883 0.0232273
R9595 avdd.n3966 avdd.n3965 0.0232273
R9596 avdd.n4223 avdd.n4098 0.0232273
R9597 avdd.n4181 avdd.n4180 0.0232273
R9598 avdd.n4438 avdd.n4313 0.0232273
R9599 avdd.n4396 avdd.n4395 0.0232273
R9600 avdd.n4948 avdd.n4847 0.0232273
R9601 avdd.n5014 avdd.n5013 0.0232273
R9602 avdd.n5164 avdd.n5063 0.0232273
R9603 avdd.n5230 avdd.n5229 0.0232273
R9604 avdd.n5380 avdd.n5279 0.0232273
R9605 avdd.n5446 avdd.n5445 0.0232273
R9606 avdd.n5596 avdd.n5495 0.0232273
R9607 avdd.n5662 avdd.n5661 0.0232273
R9608 avdd.n5812 avdd.n5711 0.0232273
R9609 avdd.n5878 avdd.n5877 0.0232273
R9610 avdd.n6028 avdd.n5927 0.0232273
R9611 avdd.n6094 avdd.n6093 0.0232273
R9612 avdd.n6244 avdd.n6143 0.0232273
R9613 avdd.n6310 avdd.n6309 0.0232273
R9614 avdd.n6460 avdd.n6359 0.0232273
R9615 avdd.n6526 avdd.n6525 0.0232273
R9616 avdd.n6676 avdd.n6575 0.0232273
R9617 avdd.n6742 avdd.n6741 0.0232273
R9618 avdd.n6892 avdd.n6791 0.0232273
R9619 avdd.n6958 avdd.n6957 0.0232273
R9620 avdd.n7108 avdd.n7007 0.0232273
R9621 avdd.n7174 avdd.n7173 0.0232273
R9622 avdd.n7324 avdd.n7223 0.0232273
R9623 avdd.n7390 avdd.n7389 0.0232273
R9624 avdd.n7673 avdd.n7672 0.0232273
R9625 avdd.n7786 avdd.n7785 0.0232273
R9626 avdd.n10152 avdd.n10151 0.0232273
R9627 avdd.n10046 avdd.n10045 0.0232273
R9628 avdd.n9936 avdd.n9935 0.0232273
R9629 avdd.n10262 avdd.n10261 0.0232273
R9630 avdd.n9822 avdd.n9821 0.0232273
R9631 avdd.n10364 avdd.n10363 0.0232273
R9632 avdd.n9708 avdd.n9707 0.0232273
R9633 avdd.n10466 avdd.n10465 0.0232273
R9634 avdd.n9595 avdd.n9594 0.0232273
R9635 avdd.n10568 avdd.n10567 0.0232273
R9636 avdd.n9480 avdd.n9479 0.0232273
R9637 avdd.n10670 avdd.n10669 0.0232273
R9638 avdd.n9366 avdd.n9365 0.0232273
R9639 avdd.n10772 avdd.n10771 0.0232273
R9640 avdd.n9252 avdd.n9251 0.0232273
R9641 avdd.n10874 avdd.n10873 0.0232273
R9642 avdd.n9138 avdd.n9137 0.0232273
R9643 avdd.n10976 avdd.n10975 0.0232273
R9644 avdd.n9024 avdd.n9023 0.0232273
R9645 avdd.n11078 avdd.n11077 0.0232273
R9646 avdd.n8910 avdd.n8909 0.0232273
R9647 avdd.n11180 avdd.n11179 0.0232273
R9648 avdd.n156 avdd.n155 0.0232273
R9649 avdd.n8809 avdd.n8808 0.0232273
R9650 avdd.n286 avdd.n285 0.0232273
R9651 avdd.n8723 avdd.n8722 0.0232273
R9652 avdd.n416 avdd.n415 0.0232273
R9653 avdd.n8637 avdd.n8636 0.0232273
R9654 avdd.n546 avdd.n545 0.0232273
R9655 avdd.n8551 avdd.n8550 0.0232273
R9656 avdd.n676 avdd.n675 0.0232273
R9657 avdd.n8465 avdd.n8464 0.0232273
R9658 avdd.n806 avdd.n805 0.0232273
R9659 avdd.n8379 avdd.n8378 0.0232273
R9660 avdd.n936 avdd.n935 0.0232273
R9661 avdd.n8293 avdd.n8292 0.0232273
R9662 avdd.n1066 avdd.n1065 0.0232273
R9663 avdd.n8207 avdd.n8206 0.0232273
R9664 avdd.n1196 avdd.n1195 0.0232273
R9665 avdd.n8121 avdd.n8120 0.0232273
R9666 avdd.n1326 avdd.n1325 0.0232273
R9667 avdd.n8035 avdd.n8034 0.0232273
R9668 avdd.n1456 avdd.n1455 0.0232273
R9669 avdd.n7949 avdd.n7948 0.0232273
R9670 avdd.n1586 avdd.n1585 0.0232273
R9671 avdd.n7863 avdd.n7862 0.0232273
R9672 avdd.n7431 avdd 0.0226354
R9673 avdd.n7427 avdd 0.0226354
R9674 avdd.n7512 avdd 0.0226354
R9675 avdd.n7505 avdd 0.0226354
R9676 avdd.n7413 avdd 0.0226354
R9677 avdd.n7409 avdd 0.0226354
R9678 avdd.n7612 avdd 0.0226354
R9679 avdd.n7605 avdd 0.0226354
R9680 avdd avdd.n1698 0.0226354
R9681 avdd.n1705 avdd 0.0226354
R9682 avdd avdd.n1734 0.0226354
R9683 avdd avdd.n1738 0.0226354
R9684 avdd avdd.n1788 0.0226354
R9685 avdd.n1795 avdd 0.0226354
R9686 avdd avdd.n1824 0.0226354
R9687 avdd avdd.n1828 0.0226354
R9688 avdd.n4804 avdd 0.0226354
R9689 avdd.n4799 avdd 0.0226354
R9690 avdd.n4796 avdd 0.0226354
R9691 avdd.n4791 avdd 0.0226354
R9692 avdd.n4788 avdd 0.0226354
R9693 avdd.n4783 avdd 0.0226354
R9694 avdd.n4780 avdd 0.0226354
R9695 avdd.n4775 avdd 0.0226354
R9696 avdd.n4772 avdd 0.0226354
R9697 avdd.n14 avdd 0.0226354
R9698 avdd.n19 avdd 0.0226354
R9699 avdd.n24 avdd 0.0226354
R9700 avdd.n29 avdd 0.0226354
R9701 avdd.n34 avdd 0.0226354
R9702 avdd.n39 avdd 0.0226354
R9703 avdd.n44 avdd 0.0226354
R9704 avdd.n49 avdd 0.0226354
R9705 avdd avdd.n54 0.0226354
R9706 avdd.n4464 avdd 0.0225588
R9707 avdd.n1998 avdd.n1978 0.0213333
R9708 avdd.n1938 avdd.n1937 0.0213333
R9709 avdd.n1914 avdd.n1913 0.0213333
R9710 avdd.n1918 avdd.n1900 0.0213333
R9711 avdd.n1922 avdd.n1918 0.0213333
R9712 avdd.n1915 avdd.n1901 0.0213333
R9713 avdd.n1917 avdd.n1916 0.0213333
R9714 avdd.n2267 avdd.n2266 0.0213333
R9715 avdd.n2191 avdd.n2190 0.0213333
R9716 avdd.n2168 avdd.n2167 0.0213333
R9717 avdd.n2172 avdd.n2154 0.0213333
R9718 avdd.n2176 avdd.n2172 0.0213333
R9719 avdd.n2169 avdd.n2155 0.0213333
R9720 avdd.n2171 avdd.n2170 0.0213333
R9721 avdd.n2482 avdd.n2481 0.0213333
R9722 avdd.n2406 avdd.n2405 0.0213333
R9723 avdd.n2383 avdd.n2382 0.0213333
R9724 avdd.n2387 avdd.n2369 0.0213333
R9725 avdd.n2391 avdd.n2387 0.0213333
R9726 avdd.n2384 avdd.n2370 0.0213333
R9727 avdd.n2386 avdd.n2385 0.0213333
R9728 avdd.n2697 avdd.n2696 0.0213333
R9729 avdd.n2621 avdd.n2620 0.0213333
R9730 avdd.n2598 avdd.n2597 0.0213333
R9731 avdd.n2602 avdd.n2584 0.0213333
R9732 avdd.n2606 avdd.n2602 0.0213333
R9733 avdd.n2599 avdd.n2585 0.0213333
R9734 avdd.n2601 avdd.n2600 0.0213333
R9735 avdd.n2912 avdd.n2911 0.0213333
R9736 avdd.n2836 avdd.n2835 0.0213333
R9737 avdd.n2813 avdd.n2812 0.0213333
R9738 avdd.n2817 avdd.n2799 0.0213333
R9739 avdd.n2821 avdd.n2817 0.0213333
R9740 avdd.n2814 avdd.n2800 0.0213333
R9741 avdd.n2816 avdd.n2815 0.0213333
R9742 avdd.n3127 avdd.n3126 0.0213333
R9743 avdd.n3051 avdd.n3050 0.0213333
R9744 avdd.n3028 avdd.n3027 0.0213333
R9745 avdd.n3032 avdd.n3014 0.0213333
R9746 avdd.n3036 avdd.n3032 0.0213333
R9747 avdd.n3029 avdd.n3015 0.0213333
R9748 avdd.n3031 avdd.n3030 0.0213333
R9749 avdd.n3288 avdd.n3268 0.0213333
R9750 avdd.n3228 avdd.n3227 0.0213333
R9751 avdd.n3204 avdd.n3203 0.0213333
R9752 avdd.n3208 avdd.n3190 0.0213333
R9753 avdd.n3212 avdd.n3208 0.0213333
R9754 avdd.n3205 avdd.n3191 0.0213333
R9755 avdd.n3207 avdd.n3206 0.0213333
R9756 avdd.n3503 avdd.n3483 0.0213333
R9757 avdd.n3443 avdd.n3442 0.0213333
R9758 avdd.n3419 avdd.n3418 0.0213333
R9759 avdd.n3423 avdd.n3405 0.0213333
R9760 avdd.n3427 avdd.n3423 0.0213333
R9761 avdd.n3420 avdd.n3406 0.0213333
R9762 avdd.n3422 avdd.n3421 0.0213333
R9763 avdd.n3718 avdd.n3698 0.0213333
R9764 avdd.n3658 avdd.n3657 0.0213333
R9765 avdd.n3634 avdd.n3633 0.0213333
R9766 avdd.n3638 avdd.n3620 0.0213333
R9767 avdd.n3642 avdd.n3638 0.0213333
R9768 avdd.n3635 avdd.n3621 0.0213333
R9769 avdd.n3637 avdd.n3636 0.0213333
R9770 avdd.n3933 avdd.n3913 0.0213333
R9771 avdd.n3873 avdd.n3872 0.0213333
R9772 avdd.n3849 avdd.n3848 0.0213333
R9773 avdd.n3853 avdd.n3835 0.0213333
R9774 avdd.n3857 avdd.n3853 0.0213333
R9775 avdd.n3850 avdd.n3836 0.0213333
R9776 avdd.n3852 avdd.n3851 0.0213333
R9777 avdd.n4148 avdd.n4128 0.0213333
R9778 avdd.n4088 avdd.n4087 0.0213333
R9779 avdd.n4064 avdd.n4063 0.0213333
R9780 avdd.n4068 avdd.n4050 0.0213333
R9781 avdd.n4072 avdd.n4068 0.0213333
R9782 avdd.n4065 avdd.n4051 0.0213333
R9783 avdd.n4067 avdd.n4066 0.0213333
R9784 avdd.n4363 avdd.n4343 0.0213333
R9785 avdd.n4303 avdd.n4302 0.0213333
R9786 avdd.n4279 avdd.n4278 0.0213333
R9787 avdd.n4283 avdd.n4265 0.0213333
R9788 avdd.n4287 avdd.n4283 0.0213333
R9789 avdd.n4280 avdd.n4266 0.0213333
R9790 avdd.n4282 avdd.n4281 0.0213333
R9791 avdd.n4890 avdd.n4889 0.0213333
R9792 avdd.n4894 avdd.n4876 0.0213333
R9793 avdd.n4898 avdd.n4894 0.0213333
R9794 avdd.n4914 avdd.n4913 0.0213333
R9795 avdd.n4989 avdd.n4988 0.0213333
R9796 avdd.n4891 avdd.n4877 0.0213333
R9797 avdd.n4893 avdd.n4892 0.0213333
R9798 avdd.n5106 avdd.n5105 0.0213333
R9799 avdd.n5110 avdd.n5092 0.0213333
R9800 avdd.n5114 avdd.n5110 0.0213333
R9801 avdd.n5130 avdd.n5129 0.0213333
R9802 avdd.n5205 avdd.n5204 0.0213333
R9803 avdd.n5107 avdd.n5093 0.0213333
R9804 avdd.n5109 avdd.n5108 0.0213333
R9805 avdd.n5322 avdd.n5321 0.0213333
R9806 avdd.n5326 avdd.n5308 0.0213333
R9807 avdd.n5330 avdd.n5326 0.0213333
R9808 avdd.n5346 avdd.n5345 0.0213333
R9809 avdd.n5421 avdd.n5420 0.0213333
R9810 avdd.n5323 avdd.n5309 0.0213333
R9811 avdd.n5325 avdd.n5324 0.0213333
R9812 avdd.n5538 avdd.n5537 0.0213333
R9813 avdd.n5542 avdd.n5524 0.0213333
R9814 avdd.n5546 avdd.n5542 0.0213333
R9815 avdd.n5562 avdd.n5561 0.0213333
R9816 avdd.n5637 avdd.n5636 0.0213333
R9817 avdd.n5539 avdd.n5525 0.0213333
R9818 avdd.n5541 avdd.n5540 0.0213333
R9819 avdd.n5754 avdd.n5753 0.0213333
R9820 avdd.n5758 avdd.n5740 0.0213333
R9821 avdd.n5762 avdd.n5758 0.0213333
R9822 avdd.n5778 avdd.n5777 0.0213333
R9823 avdd.n5853 avdd.n5852 0.0213333
R9824 avdd.n5755 avdd.n5741 0.0213333
R9825 avdd.n5757 avdd.n5756 0.0213333
R9826 avdd.n5970 avdd.n5969 0.0213333
R9827 avdd.n5974 avdd.n5956 0.0213333
R9828 avdd.n5978 avdd.n5974 0.0213333
R9829 avdd.n5994 avdd.n5993 0.0213333
R9830 avdd.n6069 avdd.n6068 0.0213333
R9831 avdd.n5971 avdd.n5957 0.0213333
R9832 avdd.n5973 avdd.n5972 0.0213333
R9833 avdd.n6186 avdd.n6185 0.0213333
R9834 avdd.n6190 avdd.n6172 0.0213333
R9835 avdd.n6194 avdd.n6190 0.0213333
R9836 avdd.n6210 avdd.n6209 0.0213333
R9837 avdd.n6285 avdd.n6284 0.0213333
R9838 avdd.n6187 avdd.n6173 0.0213333
R9839 avdd.n6189 avdd.n6188 0.0213333
R9840 avdd.n6402 avdd.n6401 0.0213333
R9841 avdd.n6406 avdd.n6388 0.0213333
R9842 avdd.n6410 avdd.n6406 0.0213333
R9843 avdd.n6426 avdd.n6425 0.0213333
R9844 avdd.n6501 avdd.n6500 0.0213333
R9845 avdd.n6403 avdd.n6389 0.0213333
R9846 avdd.n6405 avdd.n6404 0.0213333
R9847 avdd.n6618 avdd.n6617 0.0213333
R9848 avdd.n6622 avdd.n6604 0.0213333
R9849 avdd.n6626 avdd.n6622 0.0213333
R9850 avdd.n6642 avdd.n6641 0.0213333
R9851 avdd.n6717 avdd.n6716 0.0213333
R9852 avdd.n6619 avdd.n6605 0.0213333
R9853 avdd.n6621 avdd.n6620 0.0213333
R9854 avdd.n6834 avdd.n6833 0.0213333
R9855 avdd.n6838 avdd.n6820 0.0213333
R9856 avdd.n6842 avdd.n6838 0.0213333
R9857 avdd.n6858 avdd.n6857 0.0213333
R9858 avdd.n6933 avdd.n6932 0.0213333
R9859 avdd.n6835 avdd.n6821 0.0213333
R9860 avdd.n6837 avdd.n6836 0.0213333
R9861 avdd.n7050 avdd.n7049 0.0213333
R9862 avdd.n7054 avdd.n7036 0.0213333
R9863 avdd.n7058 avdd.n7054 0.0213333
R9864 avdd.n7074 avdd.n7073 0.0213333
R9865 avdd.n7149 avdd.n7148 0.0213333
R9866 avdd.n7051 avdd.n7037 0.0213333
R9867 avdd.n7053 avdd.n7052 0.0213333
R9868 avdd.n7266 avdd.n7265 0.0213333
R9869 avdd.n7270 avdd.n7252 0.0213333
R9870 avdd.n7274 avdd.n7270 0.0213333
R9871 avdd.n7290 avdd.n7289 0.0213333
R9872 avdd.n7365 avdd.n7364 0.0213333
R9873 avdd.n7267 avdd.n7253 0.0213333
R9874 avdd.n7269 avdd.n7268 0.0213333
R9875 avdd.n4623 avdd.n4616 0.0213333
R9876 avdd.n4644 avdd.n4586 0.0213333
R9877 avdd.n7750 avdd.n7749 0.0213333
R9878 avdd.n7706 avdd.n7705 0.0213333
R9879 avdd.n7707 avdd.n7706 0.0213333
R9880 avdd.n7728 avdd.n7727 0.0213333
R9881 avdd.n7818 avdd.n7817 0.0213333
R9882 avdd.n7746 avdd.n7745 0.0213333
R9883 avdd.n7710 avdd.n7709 0.0213333
R9884 avdd.n10229 avdd.n10228 0.0213333
R9885 avdd.n10185 avdd.n10184 0.0213333
R9886 avdd.n10186 avdd.n10185 0.0213333
R9887 avdd.n10207 avdd.n10206 0.0213333
R9888 avdd.n10076 avdd.n10075 0.0213333
R9889 avdd.n10225 avdd.n10224 0.0213333
R9890 avdd.n10189 avdd.n10188 0.0213333
R9891 avdd.n9983 avdd.n9982 0.0213333
R9892 avdd.n9981 avdd.n9980 0.0213333
R9893 avdd.n9980 avdd.n9979 0.0213333
R9894 avdd.n10013 avdd.n10012 0.0213333
R9895 avdd.n10308 avdd.n10307 0.0213333
R9896 avdd.n9975 avdd.n9974 0.0213333
R9897 avdd.n9973 avdd.n9972 0.0213333
R9898 avdd.n9869 avdd.n9868 0.0213333
R9899 avdd.n9867 avdd.n9866 0.0213333
R9900 avdd.n9866 avdd.n9865 0.0213333
R9901 avdd.n9899 avdd.n9898 0.0213333
R9902 avdd.n10410 avdd.n10409 0.0213333
R9903 avdd.n9861 avdd.n9860 0.0213333
R9904 avdd.n9859 avdd.n9858 0.0213333
R9905 avdd.n9755 avdd.n9754 0.0213333
R9906 avdd.n9753 avdd.n9752 0.0213333
R9907 avdd.n9752 avdd.n9751 0.0213333
R9908 avdd.n9785 avdd.n9784 0.0213333
R9909 avdd.n10512 avdd.n10511 0.0213333
R9910 avdd.n9747 avdd.n9746 0.0213333
R9911 avdd.n9745 avdd.n9744 0.0213333
R9912 avdd.n9642 avdd.n9641 0.0213333
R9913 avdd.n9640 avdd.n9639 0.0213333
R9914 avdd.n9639 avdd.n9638 0.0213333
R9915 avdd.n9672 avdd.n9671 0.0213333
R9916 avdd.n10614 avdd.n10613 0.0213333
R9917 avdd.n9634 avdd.n9633 0.0213333
R9918 avdd.n9632 avdd.n9631 0.0213333
R9919 avdd.n9527 avdd.n9526 0.0213333
R9920 avdd.n9525 avdd.n9524 0.0213333
R9921 avdd.n9524 avdd.n9523 0.0213333
R9922 avdd.n9557 avdd.n9556 0.0213333
R9923 avdd.n10716 avdd.n10715 0.0213333
R9924 avdd.n9519 avdd.n9518 0.0213333
R9925 avdd.n9517 avdd.n9516 0.0213333
R9926 avdd.n9413 avdd.n9412 0.0213333
R9927 avdd.n9411 avdd.n9410 0.0213333
R9928 avdd.n9410 avdd.n9409 0.0213333
R9929 avdd.n9443 avdd.n9442 0.0213333
R9930 avdd.n10818 avdd.n10817 0.0213333
R9931 avdd.n9405 avdd.n9404 0.0213333
R9932 avdd.n9403 avdd.n9402 0.0213333
R9933 avdd.n9299 avdd.n9298 0.0213333
R9934 avdd.n9297 avdd.n9296 0.0213333
R9935 avdd.n9296 avdd.n9295 0.0213333
R9936 avdd.n9329 avdd.n9328 0.0213333
R9937 avdd.n10920 avdd.n10919 0.0213333
R9938 avdd.n9291 avdd.n9290 0.0213333
R9939 avdd.n9289 avdd.n9288 0.0213333
R9940 avdd.n9185 avdd.n9184 0.0213333
R9941 avdd.n9183 avdd.n9182 0.0213333
R9942 avdd.n9182 avdd.n9181 0.0213333
R9943 avdd.n9215 avdd.n9214 0.0213333
R9944 avdd.n11022 avdd.n11021 0.0213333
R9945 avdd.n9177 avdd.n9176 0.0213333
R9946 avdd.n9175 avdd.n9174 0.0213333
R9947 avdd.n9071 avdd.n9070 0.0213333
R9948 avdd.n9069 avdd.n9068 0.0213333
R9949 avdd.n9068 avdd.n9067 0.0213333
R9950 avdd.n9101 avdd.n9100 0.0213333
R9951 avdd.n11124 avdd.n11123 0.0213333
R9952 avdd.n9063 avdd.n9062 0.0213333
R9953 avdd.n9061 avdd.n9060 0.0213333
R9954 avdd.n8957 avdd.n8956 0.0213333
R9955 avdd.n8955 avdd.n8954 0.0213333
R9956 avdd.n8954 avdd.n8953 0.0213333
R9957 avdd.n8987 avdd.n8986 0.0213333
R9958 avdd.n11226 avdd.n11225 0.0213333
R9959 avdd.n8949 avdd.n8948 0.0213333
R9960 avdd.n8947 avdd.n8946 0.0213333
R9961 avdd.n8839 avdd.n8838 0.0213333
R9962 avdd.n123 avdd.n122 0.0213333
R9963 avdd.n83 avdd.n82 0.0213333
R9964 avdd.n100 avdd.n99 0.0213333
R9965 avdd.n101 avdd.n100 0.0213333
R9966 avdd.n79 avdd.n78 0.0213333
R9967 avdd.n104 avdd.n103 0.0213333
R9968 avdd.n8753 avdd.n8752 0.0213333
R9969 avdd.n253 avdd.n252 0.0213333
R9970 avdd.n213 avdd.n212 0.0213333
R9971 avdd.n230 avdd.n229 0.0213333
R9972 avdd.n231 avdd.n230 0.0213333
R9973 avdd.n209 avdd.n208 0.0213333
R9974 avdd.n234 avdd.n233 0.0213333
R9975 avdd.n8667 avdd.n8666 0.0213333
R9976 avdd.n383 avdd.n382 0.0213333
R9977 avdd.n343 avdd.n342 0.0213333
R9978 avdd.n360 avdd.n359 0.0213333
R9979 avdd.n361 avdd.n360 0.0213333
R9980 avdd.n339 avdd.n338 0.0213333
R9981 avdd.n364 avdd.n363 0.0213333
R9982 avdd.n8581 avdd.n8580 0.0213333
R9983 avdd.n513 avdd.n512 0.0213333
R9984 avdd.n473 avdd.n472 0.0213333
R9985 avdd.n490 avdd.n489 0.0213333
R9986 avdd.n491 avdd.n490 0.0213333
R9987 avdd.n469 avdd.n468 0.0213333
R9988 avdd.n494 avdd.n493 0.0213333
R9989 avdd.n8495 avdd.n8494 0.0213333
R9990 avdd.n643 avdd.n642 0.0213333
R9991 avdd.n603 avdd.n602 0.0213333
R9992 avdd.n620 avdd.n619 0.0213333
R9993 avdd.n621 avdd.n620 0.0213333
R9994 avdd.n599 avdd.n598 0.0213333
R9995 avdd.n624 avdd.n623 0.0213333
R9996 avdd.n8409 avdd.n8408 0.0213333
R9997 avdd.n773 avdd.n772 0.0213333
R9998 avdd.n733 avdd.n732 0.0213333
R9999 avdd.n750 avdd.n749 0.0213333
R10000 avdd.n751 avdd.n750 0.0213333
R10001 avdd.n729 avdd.n728 0.0213333
R10002 avdd.n754 avdd.n753 0.0213333
R10003 avdd.n8323 avdd.n8322 0.0213333
R10004 avdd.n903 avdd.n902 0.0213333
R10005 avdd.n863 avdd.n862 0.0213333
R10006 avdd.n880 avdd.n879 0.0213333
R10007 avdd.n881 avdd.n880 0.0213333
R10008 avdd.n859 avdd.n858 0.0213333
R10009 avdd.n884 avdd.n883 0.0213333
R10010 avdd.n8237 avdd.n8236 0.0213333
R10011 avdd.n1033 avdd.n1032 0.0213333
R10012 avdd.n993 avdd.n992 0.0213333
R10013 avdd.n1010 avdd.n1009 0.0213333
R10014 avdd.n1011 avdd.n1010 0.0213333
R10015 avdd.n989 avdd.n988 0.0213333
R10016 avdd.n1014 avdd.n1013 0.0213333
R10017 avdd.n8151 avdd.n8150 0.0213333
R10018 avdd.n1163 avdd.n1162 0.0213333
R10019 avdd.n1123 avdd.n1122 0.0213333
R10020 avdd.n1140 avdd.n1139 0.0213333
R10021 avdd.n1141 avdd.n1140 0.0213333
R10022 avdd.n1119 avdd.n1118 0.0213333
R10023 avdd.n1144 avdd.n1143 0.0213333
R10024 avdd.n8065 avdd.n8064 0.0213333
R10025 avdd.n1293 avdd.n1292 0.0213333
R10026 avdd.n1253 avdd.n1252 0.0213333
R10027 avdd.n1270 avdd.n1269 0.0213333
R10028 avdd.n1271 avdd.n1270 0.0213333
R10029 avdd.n1249 avdd.n1248 0.0213333
R10030 avdd.n1274 avdd.n1273 0.0213333
R10031 avdd.n7979 avdd.n7978 0.0213333
R10032 avdd.n1423 avdd.n1422 0.0213333
R10033 avdd.n1383 avdd.n1382 0.0213333
R10034 avdd.n1400 avdd.n1399 0.0213333
R10035 avdd.n1401 avdd.n1400 0.0213333
R10036 avdd.n1379 avdd.n1378 0.0213333
R10037 avdd.n1404 avdd.n1403 0.0213333
R10038 avdd.n7893 avdd.n7892 0.0213333
R10039 avdd.n1553 avdd.n1552 0.0213333
R10040 avdd.n1513 avdd.n1512 0.0213333
R10041 avdd.n1530 avdd.n1529 0.0213333
R10042 avdd.n1531 avdd.n1530 0.0213333
R10043 avdd.n1509 avdd.n1508 0.0213333
R10044 avdd.n1534 avdd.n1533 0.0213333
R10045 avdd.n2065 avdd.n2064 0.0211515
R10046 avdd.n2058 avdd.n1960 0.0211515
R10047 avdd.n1906 avdd.n1905 0.0211515
R10048 avdd.n2236 avdd.n2120 0.0211515
R10049 avdd.n2238 avdd.n2237 0.0211515
R10050 avdd.n2160 avdd.n2159 0.0211515
R10051 avdd.n2451 avdd.n2335 0.0211515
R10052 avdd.n2453 avdd.n2452 0.0211515
R10053 avdd.n2375 avdd.n2374 0.0211515
R10054 avdd.n2666 avdd.n2550 0.0211515
R10055 avdd.n2668 avdd.n2667 0.0211515
R10056 avdd.n2590 avdd.n2589 0.0211515
R10057 avdd.n2881 avdd.n2765 0.0211515
R10058 avdd.n2883 avdd.n2882 0.0211515
R10059 avdd.n2805 avdd.n2804 0.0211515
R10060 avdd.n3096 avdd.n2980 0.0211515
R10061 avdd.n3098 avdd.n3097 0.0211515
R10062 avdd.n3020 avdd.n3019 0.0211515
R10063 avdd.n3354 avdd.n3353 0.0211515
R10064 avdd.n3347 avdd.n3250 0.0211515
R10065 avdd.n3196 avdd.n3195 0.0211515
R10066 avdd.n3569 avdd.n3568 0.0211515
R10067 avdd.n3562 avdd.n3465 0.0211515
R10068 avdd.n3411 avdd.n3410 0.0211515
R10069 avdd.n3784 avdd.n3783 0.0211515
R10070 avdd.n3777 avdd.n3680 0.0211515
R10071 avdd.n3626 avdd.n3625 0.0211515
R10072 avdd.n3999 avdd.n3998 0.0211515
R10073 avdd.n3992 avdd.n3895 0.0211515
R10074 avdd.n3841 avdd.n3840 0.0211515
R10075 avdd.n4214 avdd.n4213 0.0211515
R10076 avdd.n4207 avdd.n4110 0.0211515
R10077 avdd.n4056 avdd.n4055 0.0211515
R10078 avdd.n4429 avdd.n4428 0.0211515
R10079 avdd.n4422 avdd.n4325 0.0211515
R10080 avdd.n4271 avdd.n4270 0.0211515
R10081 avdd.n4958 avdd.n4842 0.0211515
R10082 avdd.n4960 avdd.n4959 0.0211515
R10083 avdd.n4882 avdd.n4881 0.0211515
R10084 avdd.n5174 avdd.n5058 0.0211515
R10085 avdd.n5176 avdd.n5175 0.0211515
R10086 avdd.n5098 avdd.n5097 0.0211515
R10087 avdd.n5390 avdd.n5274 0.0211515
R10088 avdd.n5392 avdd.n5391 0.0211515
R10089 avdd.n5314 avdd.n5313 0.0211515
R10090 avdd.n5606 avdd.n5490 0.0211515
R10091 avdd.n5608 avdd.n5607 0.0211515
R10092 avdd.n5530 avdd.n5529 0.0211515
R10093 avdd.n5822 avdd.n5706 0.0211515
R10094 avdd.n5824 avdd.n5823 0.0211515
R10095 avdd.n5746 avdd.n5745 0.0211515
R10096 avdd.n6038 avdd.n5922 0.0211515
R10097 avdd.n6040 avdd.n6039 0.0211515
R10098 avdd.n5962 avdd.n5961 0.0211515
R10099 avdd.n6254 avdd.n6138 0.0211515
R10100 avdd.n6256 avdd.n6255 0.0211515
R10101 avdd.n6178 avdd.n6177 0.0211515
R10102 avdd.n6470 avdd.n6354 0.0211515
R10103 avdd.n6472 avdd.n6471 0.0211515
R10104 avdd.n6394 avdd.n6393 0.0211515
R10105 avdd.n6686 avdd.n6570 0.0211515
R10106 avdd.n6688 avdd.n6687 0.0211515
R10107 avdd.n6610 avdd.n6609 0.0211515
R10108 avdd.n6902 avdd.n6786 0.0211515
R10109 avdd.n6904 avdd.n6903 0.0211515
R10110 avdd.n6826 avdd.n6825 0.0211515
R10111 avdd.n7118 avdd.n7002 0.0211515
R10112 avdd.n7120 avdd.n7119 0.0211515
R10113 avdd.n7042 avdd.n7041 0.0211515
R10114 avdd.n7334 avdd.n7218 0.0211515
R10115 avdd.n7336 avdd.n7335 0.0211515
R10116 avdd.n7258 avdd.n7257 0.0211515
R10117 avdd.n7768 avdd.n7767 0.0211515
R10118 avdd.n7756 avdd.n7755 0.0211515
R10119 avdd.n10117 avdd.n10116 0.0211515
R10120 avdd.n10115 avdd.n10114 0.0211515
R10121 avdd.n10235 avdd.n10234 0.0211515
R10122 avdd.n9918 avdd.n9917 0.0211515
R10123 avdd.n9916 avdd.n9915 0.0211515
R10124 avdd.n9989 avdd.n9988 0.0211515
R10125 avdd.n9804 avdd.n9803 0.0211515
R10126 avdd.n9802 avdd.n9801 0.0211515
R10127 avdd.n9875 avdd.n9874 0.0211515
R10128 avdd.n9690 avdd.n9689 0.0211515
R10129 avdd.n9688 avdd.n9687 0.0211515
R10130 avdd.n9761 avdd.n9760 0.0211515
R10131 avdd.n9576 avdd.n9575 0.0211515
R10132 avdd.n9574 avdd.n9573 0.0211515
R10133 avdd.n9648 avdd.n9647 0.0211515
R10134 avdd.n9462 avdd.n9461 0.0211515
R10135 avdd.n9460 avdd.n9459 0.0211515
R10136 avdd.n9533 avdd.n9532 0.0211515
R10137 avdd.n9348 avdd.n9347 0.0211515
R10138 avdd.n9346 avdd.n9345 0.0211515
R10139 avdd.n9419 avdd.n9418 0.0211515
R10140 avdd.n9234 avdd.n9233 0.0211515
R10141 avdd.n9232 avdd.n9231 0.0211515
R10142 avdd.n9305 avdd.n9304 0.0211515
R10143 avdd.n9120 avdd.n9119 0.0211515
R10144 avdd.n9118 avdd.n9117 0.0211515
R10145 avdd.n9191 avdd.n9190 0.0211515
R10146 avdd.n9006 avdd.n9005 0.0211515
R10147 avdd.n9004 avdd.n9003 0.0211515
R10148 avdd.n9077 avdd.n9076 0.0211515
R10149 avdd.n8892 avdd.n8891 0.0211515
R10150 avdd.n8890 avdd.n8889 0.0211515
R10151 avdd.n8963 avdd.n8962 0.0211515
R10152 avdd.n61 avdd.n60 0.0211515
R10153 avdd.n59 avdd.n58 0.0211515
R10154 avdd.n89 avdd.n88 0.0211515
R10155 avdd.n191 avdd.n190 0.0211515
R10156 avdd.n189 avdd.n188 0.0211515
R10157 avdd.n219 avdd.n218 0.0211515
R10158 avdd.n321 avdd.n320 0.0211515
R10159 avdd.n319 avdd.n318 0.0211515
R10160 avdd.n349 avdd.n348 0.0211515
R10161 avdd.n451 avdd.n450 0.0211515
R10162 avdd.n449 avdd.n448 0.0211515
R10163 avdd.n479 avdd.n478 0.0211515
R10164 avdd.n581 avdd.n580 0.0211515
R10165 avdd.n579 avdd.n578 0.0211515
R10166 avdd.n609 avdd.n608 0.0211515
R10167 avdd.n711 avdd.n710 0.0211515
R10168 avdd.n709 avdd.n708 0.0211515
R10169 avdd.n739 avdd.n738 0.0211515
R10170 avdd.n841 avdd.n840 0.0211515
R10171 avdd.n839 avdd.n838 0.0211515
R10172 avdd.n869 avdd.n868 0.0211515
R10173 avdd.n971 avdd.n970 0.0211515
R10174 avdd.n969 avdd.n968 0.0211515
R10175 avdd.n999 avdd.n998 0.0211515
R10176 avdd.n1101 avdd.n1100 0.0211515
R10177 avdd.n1099 avdd.n1098 0.0211515
R10178 avdd.n1129 avdd.n1128 0.0211515
R10179 avdd.n1231 avdd.n1230 0.0211515
R10180 avdd.n1229 avdd.n1228 0.0211515
R10181 avdd.n1259 avdd.n1258 0.0211515
R10182 avdd.n1361 avdd.n1360 0.0211515
R10183 avdd.n1359 avdd.n1358 0.0211515
R10184 avdd.n1389 avdd.n1388 0.0211515
R10185 avdd.n1491 avdd.n1490 0.0211515
R10186 avdd.n1489 avdd.n1488 0.0211515
R10187 avdd.n1519 avdd.n1518 0.0211515
R10188 avdd.n7454 avdd 0.0200312
R10189 avdd avdd.n7493 0.0200312
R10190 avdd.n7553 avdd 0.0200312
R10191 avdd avdd.n7593 0.0200312
R10192 avdd avdd.n7635 0.0200312
R10193 avdd avdd.n1691 0.0200312
R10194 avdd avdd.n1730 0.0200312
R10195 avdd avdd.n1781 0.0200312
R10196 avdd avdd.n1820 0.0200312
R10197 avdd.n1870 avdd 0.0200312
R10198 avdd.n1951 avdd.n1883 0.0197273
R10199 avdd.n2078 avdd.n1888 0.0197273
R10200 avdd.n2217 avdd.n2216 0.0197273
R10201 avdd.n2218 avdd.n2132 0.0197273
R10202 avdd.n2432 avdd.n2431 0.0197273
R10203 avdd.n2433 avdd.n2347 0.0197273
R10204 avdd.n2647 avdd.n2646 0.0197273
R10205 avdd.n2648 avdd.n2562 0.0197273
R10206 avdd.n2862 avdd.n2861 0.0197273
R10207 avdd.n2863 avdd.n2777 0.0197273
R10208 avdd.n3077 avdd.n3076 0.0197273
R10209 avdd.n3078 avdd.n2992 0.0197273
R10210 avdd.n3241 avdd.n3173 0.0197273
R10211 avdd.n3367 avdd.n3178 0.0197273
R10212 avdd.n3323 avdd.n3297 0.0197273
R10213 avdd.n3456 avdd.n3388 0.0197273
R10214 avdd.n3582 avdd.n3393 0.0197273
R10215 avdd.n3538 avdd.n3512 0.0197273
R10216 avdd.n3671 avdd.n3603 0.0197273
R10217 avdd.n3797 avdd.n3608 0.0197273
R10218 avdd.n3753 avdd.n3727 0.0197273
R10219 avdd.n3886 avdd.n3818 0.0197273
R10220 avdd.n4012 avdd.n3823 0.0197273
R10221 avdd.n3968 avdd.n3942 0.0197273
R10222 avdd.n4101 avdd.n4033 0.0197273
R10223 avdd.n4227 avdd.n4038 0.0197273
R10224 avdd.n4183 avdd.n4157 0.0197273
R10225 avdd.n4316 avdd.n4248 0.0197273
R10226 avdd.n4442 avdd.n4253 0.0197273
R10227 avdd.n4398 avdd.n4372 0.0197273
R10228 avdd.n4939 avdd.n4938 0.0197273
R10229 avdd.n4940 avdd.n4854 0.0197273
R10230 avdd.n5155 avdd.n5154 0.0197273
R10231 avdd.n5156 avdd.n5070 0.0197273
R10232 avdd.n5371 avdd.n5370 0.0197273
R10233 avdd.n5372 avdd.n5286 0.0197273
R10234 avdd.n5587 avdd.n5586 0.0197273
R10235 avdd.n5588 avdd.n5502 0.0197273
R10236 avdd.n5803 avdd.n5802 0.0197273
R10237 avdd.n5804 avdd.n5718 0.0197273
R10238 avdd.n6019 avdd.n6018 0.0197273
R10239 avdd.n6020 avdd.n5934 0.0197273
R10240 avdd.n6235 avdd.n6234 0.0197273
R10241 avdd.n6236 avdd.n6150 0.0197273
R10242 avdd.n6451 avdd.n6450 0.0197273
R10243 avdd.n6452 avdd.n6366 0.0197273
R10244 avdd.n6667 avdd.n6666 0.0197273
R10245 avdd.n6668 avdd.n6582 0.0197273
R10246 avdd.n6883 avdd.n6882 0.0197273
R10247 avdd.n6884 avdd.n6798 0.0197273
R10248 avdd.n7099 avdd.n7098 0.0197273
R10249 avdd.n7100 avdd.n7014 0.0197273
R10250 avdd.n7315 avdd.n7314 0.0197273
R10251 avdd.n7316 avdd.n7230 0.0197273
R10252 avdd.n7649 avdd.n7648 0.0197273
R10253 avdd.n7685 avdd.n7684 0.0197273
R10254 avdd.n7848 avdd.n7847 0.0197273
R10255 avdd.n10126 avdd.n10125 0.0197273
R10256 avdd.n10164 avdd.n10163 0.0197273
R10257 avdd.n10106 avdd.n10105 0.0197273
R10258 avdd.n9927 avdd.n9926 0.0197273
R10259 avdd.n9948 avdd.n9947 0.0197273
R10260 avdd.n9813 avdd.n9812 0.0197273
R10261 avdd.n9834 avdd.n9833 0.0197273
R10262 avdd.n9699 avdd.n9698 0.0197273
R10263 avdd.n9720 avdd.n9719 0.0197273
R10264 avdd.n9585 avdd.n9584 0.0197273
R10265 avdd.n9607 avdd.n9606 0.0197273
R10266 avdd.n9471 avdd.n9470 0.0197273
R10267 avdd.n9492 avdd.n9491 0.0197273
R10268 avdd.n9357 avdd.n9356 0.0197273
R10269 avdd.n9378 avdd.n9377 0.0197273
R10270 avdd.n9243 avdd.n9242 0.0197273
R10271 avdd.n9264 avdd.n9263 0.0197273
R10272 avdd.n9129 avdd.n9128 0.0197273
R10273 avdd.n9150 avdd.n9149 0.0197273
R10274 avdd.n9015 avdd.n9014 0.0197273
R10275 avdd.n9036 avdd.n9035 0.0197273
R10276 avdd.n8901 avdd.n8900 0.0197273
R10277 avdd.n8922 avdd.n8921 0.0197273
R10278 avdd.n70 avdd.n69 0.0197273
R10279 avdd.n168 avdd.n167 0.0197273
R10280 avdd.n200 avdd.n199 0.0197273
R10281 avdd.n298 avdd.n297 0.0197273
R10282 avdd.n330 avdd.n329 0.0197273
R10283 avdd.n428 avdd.n427 0.0197273
R10284 avdd.n460 avdd.n459 0.0197273
R10285 avdd.n558 avdd.n557 0.0197273
R10286 avdd.n590 avdd.n589 0.0197273
R10287 avdd.n688 avdd.n687 0.0197273
R10288 avdd.n720 avdd.n719 0.0197273
R10289 avdd.n818 avdd.n817 0.0197273
R10290 avdd.n850 avdd.n849 0.0197273
R10291 avdd.n948 avdd.n947 0.0197273
R10292 avdd.n980 avdd.n979 0.0197273
R10293 avdd.n1078 avdd.n1077 0.0197273
R10294 avdd.n1110 avdd.n1109 0.0197273
R10295 avdd.n1208 avdd.n1207 0.0197273
R10296 avdd.n1240 avdd.n1239 0.0197273
R10297 avdd.n1338 avdd.n1337 0.0197273
R10298 avdd.n1370 avdd.n1369 0.0197273
R10299 avdd.n1468 avdd.n1467 0.0197273
R10300 avdd.n1500 avdd.n1499 0.0197273
R10301 avdd.n1598 avdd.n1597 0.0197273
R10302 avdd.n2014 avdd.n2013 0.0194394
R10303 avdd.n1983 avdd.n1976 0.0194394
R10304 avdd.n2082 avdd.n2081 0.0194394
R10305 avdd.n1931 avdd.n1893 0.0194394
R10306 avdd.n2287 avdd.n2286 0.0194394
R10307 avdd.n2260 avdd.n2111 0.0194394
R10308 avdd.n2205 avdd.n2204 0.0194394
R10309 avdd.n2184 avdd.n2148 0.0194394
R10310 avdd.n2502 avdd.n2501 0.0194394
R10311 avdd.n2475 avdd.n2326 0.0194394
R10312 avdd.n2420 avdd.n2419 0.0194394
R10313 avdd.n2399 avdd.n2363 0.0194394
R10314 avdd.n2717 avdd.n2716 0.0194394
R10315 avdd.n2690 avdd.n2541 0.0194394
R10316 avdd.n2635 avdd.n2634 0.0194394
R10317 avdd.n2614 avdd.n2578 0.0194394
R10318 avdd.n2932 avdd.n2931 0.0194394
R10319 avdd.n2905 avdd.n2756 0.0194394
R10320 avdd.n2850 avdd.n2849 0.0194394
R10321 avdd.n2829 avdd.n2793 0.0194394
R10322 avdd.n3147 avdd.n3146 0.0194394
R10323 avdd.n3120 avdd.n2971 0.0194394
R10324 avdd.n3065 avdd.n3064 0.0194394
R10325 avdd.n3044 avdd.n3008 0.0194394
R10326 avdd.n3307 avdd.n3306 0.0194394
R10327 avdd.n3273 avdd.n3266 0.0194394
R10328 avdd.n3371 avdd.n3370 0.0194394
R10329 avdd.n3221 avdd.n3183 0.0194394
R10330 avdd.n3522 avdd.n3521 0.0194394
R10331 avdd.n3488 avdd.n3481 0.0194394
R10332 avdd.n3586 avdd.n3585 0.0194394
R10333 avdd.n3436 avdd.n3398 0.0194394
R10334 avdd.n3737 avdd.n3736 0.0194394
R10335 avdd.n3703 avdd.n3696 0.0194394
R10336 avdd.n3801 avdd.n3800 0.0194394
R10337 avdd.n3651 avdd.n3613 0.0194394
R10338 avdd.n3952 avdd.n3951 0.0194394
R10339 avdd.n3918 avdd.n3911 0.0194394
R10340 avdd.n4016 avdd.n4015 0.0194394
R10341 avdd.n3866 avdd.n3828 0.0194394
R10342 avdd.n4167 avdd.n4166 0.0194394
R10343 avdd.n4133 avdd.n4126 0.0194394
R10344 avdd.n4231 avdd.n4230 0.0194394
R10345 avdd.n4081 avdd.n4043 0.0194394
R10346 avdd.n4382 avdd.n4381 0.0194394
R10347 avdd.n4348 avdd.n4341 0.0194394
R10348 avdd.n4446 avdd.n4445 0.0194394
R10349 avdd.n4296 avdd.n4258 0.0194394
R10350 avdd.n4907 avdd.n4870 0.0194394
R10351 avdd.n4927 avdd.n4926 0.0194394
R10352 avdd.n4982 avdd.n4833 0.0194394
R10353 avdd.n5005 avdd.n5004 0.0194394
R10354 avdd.n5123 avdd.n5086 0.0194394
R10355 avdd.n5143 avdd.n5142 0.0194394
R10356 avdd.n5198 avdd.n5049 0.0194394
R10357 avdd.n5221 avdd.n5220 0.0194394
R10358 avdd.n5339 avdd.n5302 0.0194394
R10359 avdd.n5359 avdd.n5358 0.0194394
R10360 avdd.n5414 avdd.n5265 0.0194394
R10361 avdd.n5437 avdd.n5436 0.0194394
R10362 avdd.n5555 avdd.n5518 0.0194394
R10363 avdd.n5575 avdd.n5574 0.0194394
R10364 avdd.n5630 avdd.n5481 0.0194394
R10365 avdd.n5653 avdd.n5652 0.0194394
R10366 avdd.n5771 avdd.n5734 0.0194394
R10367 avdd.n5791 avdd.n5790 0.0194394
R10368 avdd.n5846 avdd.n5697 0.0194394
R10369 avdd.n5869 avdd.n5868 0.0194394
R10370 avdd.n5987 avdd.n5950 0.0194394
R10371 avdd.n6007 avdd.n6006 0.0194394
R10372 avdd.n6062 avdd.n5913 0.0194394
R10373 avdd.n6085 avdd.n6084 0.0194394
R10374 avdd.n6203 avdd.n6166 0.0194394
R10375 avdd.n6223 avdd.n6222 0.0194394
R10376 avdd.n6278 avdd.n6129 0.0194394
R10377 avdd.n6301 avdd.n6300 0.0194394
R10378 avdd.n6419 avdd.n6382 0.0194394
R10379 avdd.n6439 avdd.n6438 0.0194394
R10380 avdd.n6494 avdd.n6345 0.0194394
R10381 avdd.n6517 avdd.n6516 0.0194394
R10382 avdd.n6635 avdd.n6598 0.0194394
R10383 avdd.n6655 avdd.n6654 0.0194394
R10384 avdd.n6710 avdd.n6561 0.0194394
R10385 avdd.n6733 avdd.n6732 0.0194394
R10386 avdd.n6851 avdd.n6814 0.0194394
R10387 avdd.n6871 avdd.n6870 0.0194394
R10388 avdd.n6926 avdd.n6777 0.0194394
R10389 avdd.n6949 avdd.n6948 0.0194394
R10390 avdd.n7067 avdd.n7030 0.0194394
R10391 avdd.n7087 avdd.n7086 0.0194394
R10392 avdd.n7142 avdd.n6993 0.0194394
R10393 avdd.n7165 avdd.n7164 0.0194394
R10394 avdd.n7283 avdd.n7246 0.0194394
R10395 avdd.n7303 avdd.n7302 0.0194394
R10396 avdd.n7358 avdd.n7209 0.0194394
R10397 avdd.n7381 avdd.n7380 0.0194394
R10398 avdd.n7714 avdd.n7713 0.0194394
R10399 avdd.n7696 avdd.n7695 0.0194394
R10400 avdd.n7803 avdd.n7802 0.0194394
R10401 avdd.n7843 avdd.n7842 0.0194394
R10402 avdd.n10193 avdd.n10192 0.0194394
R10403 avdd.n10175 avdd.n10174 0.0194394
R10404 avdd.n10061 avdd.n10060 0.0194394
R10405 avdd.n10101 avdd.n10100 0.0194394
R10406 avdd.n9997 avdd.n9996 0.0194394
R10407 avdd.n9959 avdd.n9958 0.0194394
R10408 avdd.n10293 avdd.n10292 0.0194394
R10409 avdd.n10333 avdd.n10332 0.0194394
R10410 avdd.n9883 avdd.n9882 0.0194394
R10411 avdd.n9845 avdd.n9844 0.0194394
R10412 avdd.n10395 avdd.n10394 0.0194394
R10413 avdd.n10435 avdd.n10434 0.0194394
R10414 avdd.n9769 avdd.n9768 0.0194394
R10415 avdd.n9731 avdd.n9730 0.0194394
R10416 avdd.n10497 avdd.n10496 0.0194394
R10417 avdd.n10537 avdd.n10536 0.0194394
R10418 avdd.n9656 avdd.n9655 0.0194394
R10419 avdd.n9618 avdd.n9617 0.0194394
R10420 avdd.n10599 avdd.n10598 0.0194394
R10421 avdd.n10639 avdd.n10638 0.0194394
R10422 avdd.n9541 avdd.n9540 0.0194394
R10423 avdd.n9503 avdd.n9502 0.0194394
R10424 avdd.n10701 avdd.n10700 0.0194394
R10425 avdd.n10741 avdd.n10740 0.0194394
R10426 avdd.n9427 avdd.n9426 0.0194394
R10427 avdd.n9389 avdd.n9388 0.0194394
R10428 avdd.n10803 avdd.n10802 0.0194394
R10429 avdd.n10843 avdd.n10842 0.0194394
R10430 avdd.n9313 avdd.n9312 0.0194394
R10431 avdd.n9275 avdd.n9274 0.0194394
R10432 avdd.n10905 avdd.n10904 0.0194394
R10433 avdd.n10945 avdd.n10944 0.0194394
R10434 avdd.n9199 avdd.n9198 0.0194394
R10435 avdd.n9161 avdd.n9160 0.0194394
R10436 avdd.n11007 avdd.n11006 0.0194394
R10437 avdd.n11047 avdd.n11046 0.0194394
R10438 avdd.n9085 avdd.n9084 0.0194394
R10439 avdd.n9047 avdd.n9046 0.0194394
R10440 avdd.n11109 avdd.n11108 0.0194394
R10441 avdd.n11149 avdd.n11148 0.0194394
R10442 avdd.n8971 avdd.n8970 0.0194394
R10443 avdd.n8933 avdd.n8932 0.0194394
R10444 avdd.n11211 avdd.n11210 0.0194394
R10445 avdd.n11251 avdd.n11250 0.0194394
R10446 avdd.n8864 avdd.n8863 0.0194394
R10447 avdd.n8824 avdd.n8823 0.0194394
R10448 avdd.n179 avdd.n178 0.0194394
R10449 avdd.n108 avdd.n107 0.0194394
R10450 avdd.n8778 avdd.n8777 0.0194394
R10451 avdd.n8738 avdd.n8737 0.0194394
R10452 avdd.n309 avdd.n308 0.0194394
R10453 avdd.n238 avdd.n237 0.0194394
R10454 avdd.n8692 avdd.n8691 0.0194394
R10455 avdd.n8652 avdd.n8651 0.0194394
R10456 avdd.n439 avdd.n438 0.0194394
R10457 avdd.n368 avdd.n367 0.0194394
R10458 avdd.n8606 avdd.n8605 0.0194394
R10459 avdd.n8566 avdd.n8565 0.0194394
R10460 avdd.n569 avdd.n568 0.0194394
R10461 avdd.n498 avdd.n497 0.0194394
R10462 avdd.n8520 avdd.n8519 0.0194394
R10463 avdd.n8480 avdd.n8479 0.0194394
R10464 avdd.n699 avdd.n698 0.0194394
R10465 avdd.n628 avdd.n627 0.0194394
R10466 avdd.n8434 avdd.n8433 0.0194394
R10467 avdd.n8394 avdd.n8393 0.0194394
R10468 avdd.n829 avdd.n828 0.0194394
R10469 avdd.n758 avdd.n757 0.0194394
R10470 avdd.n8348 avdd.n8347 0.0194394
R10471 avdd.n8308 avdd.n8307 0.0194394
R10472 avdd.n959 avdd.n958 0.0194394
R10473 avdd.n888 avdd.n887 0.0194394
R10474 avdd.n8262 avdd.n8261 0.0194394
R10475 avdd.n8222 avdd.n8221 0.0194394
R10476 avdd.n1089 avdd.n1088 0.0194394
R10477 avdd.n1018 avdd.n1017 0.0194394
R10478 avdd.n8176 avdd.n8175 0.0194394
R10479 avdd.n8136 avdd.n8135 0.0194394
R10480 avdd.n1219 avdd.n1218 0.0194394
R10481 avdd.n1148 avdd.n1147 0.0194394
R10482 avdd.n8090 avdd.n8089 0.0194394
R10483 avdd.n8050 avdd.n8049 0.0194394
R10484 avdd.n1349 avdd.n1348 0.0194394
R10485 avdd.n1278 avdd.n1277 0.0194394
R10486 avdd.n8004 avdd.n8003 0.0194394
R10487 avdd.n7964 avdd.n7963 0.0194394
R10488 avdd.n1479 avdd.n1478 0.0194394
R10489 avdd.n1408 avdd.n1407 0.0194394
R10490 avdd.n7918 avdd.n7917 0.0194394
R10491 avdd.n7878 avdd.n7877 0.0194394
R10492 avdd.n1609 avdd.n1608 0.0194394
R10493 avdd.n1538 avdd.n1537 0.0194394
R10494 avdd.n4630 avdd.n4629 0.01925
R10495 avdd.n7635 avdd 0.0187292
R10496 avdd.n1870 avdd 0.0187292
R10497 avdd.n4806 avdd 0.0187292
R10498 avdd.n7635 avdd 0.0183571
R10499 avdd avdd.n1870 0.0183571
R10500 avdd.n2046 avdd.n1993 0.018303
R10501 avdd.n2047 avdd.n1979 0.018303
R10502 avdd.n2270 avdd.n2107 0.018303
R10503 avdd.n2269 avdd.n2108 0.018303
R10504 avdd.n2485 avdd.n2322 0.018303
R10505 avdd.n2484 avdd.n2323 0.018303
R10506 avdd.n2700 avdd.n2537 0.018303
R10507 avdd.n2699 avdd.n2538 0.018303
R10508 avdd.n2915 avdd.n2752 0.018303
R10509 avdd.n2914 avdd.n2753 0.018303
R10510 avdd.n3130 avdd.n2967 0.018303
R10511 avdd.n3129 avdd.n2968 0.018303
R10512 avdd.n3335 avdd.n3283 0.018303
R10513 avdd.n3336 avdd.n3269 0.018303
R10514 avdd.n3550 avdd.n3498 0.018303
R10515 avdd.n3551 avdd.n3484 0.018303
R10516 avdd.n3765 avdd.n3713 0.018303
R10517 avdd.n3766 avdd.n3699 0.018303
R10518 avdd.n3980 avdd.n3928 0.018303
R10519 avdd.n3981 avdd.n3914 0.018303
R10520 avdd.n4195 avdd.n4143 0.018303
R10521 avdd.n4196 avdd.n4129 0.018303
R10522 avdd.n4410 avdd.n4358 0.018303
R10523 avdd.n4411 avdd.n4344 0.018303
R10524 avdd.n4992 avdd.n4829 0.018303
R10525 avdd.n4917 avdd.n4916 0.018303
R10526 avdd.n4991 avdd.n4830 0.018303
R10527 avdd.n5208 avdd.n5045 0.018303
R10528 avdd.n5133 avdd.n5132 0.018303
R10529 avdd.n5207 avdd.n5046 0.018303
R10530 avdd.n5424 avdd.n5261 0.018303
R10531 avdd.n5349 avdd.n5348 0.018303
R10532 avdd.n5423 avdd.n5262 0.018303
R10533 avdd.n5640 avdd.n5477 0.018303
R10534 avdd.n5565 avdd.n5564 0.018303
R10535 avdd.n5639 avdd.n5478 0.018303
R10536 avdd.n5856 avdd.n5693 0.018303
R10537 avdd.n5781 avdd.n5780 0.018303
R10538 avdd.n5855 avdd.n5694 0.018303
R10539 avdd.n6072 avdd.n5909 0.018303
R10540 avdd.n5997 avdd.n5996 0.018303
R10541 avdd.n6071 avdd.n5910 0.018303
R10542 avdd.n6288 avdd.n6125 0.018303
R10543 avdd.n6213 avdd.n6212 0.018303
R10544 avdd.n6287 avdd.n6126 0.018303
R10545 avdd.n6504 avdd.n6341 0.018303
R10546 avdd.n6429 avdd.n6428 0.018303
R10547 avdd.n6503 avdd.n6342 0.018303
R10548 avdd.n6720 avdd.n6557 0.018303
R10549 avdd.n6645 avdd.n6644 0.018303
R10550 avdd.n6719 avdd.n6558 0.018303
R10551 avdd.n6936 avdd.n6773 0.018303
R10552 avdd.n6861 avdd.n6860 0.018303
R10553 avdd.n6935 avdd.n6774 0.018303
R10554 avdd.n7152 avdd.n6989 0.018303
R10555 avdd.n7077 avdd.n7076 0.018303
R10556 avdd.n7151 avdd.n6990 0.018303
R10557 avdd.n7368 avdd.n7205 0.018303
R10558 avdd.n7293 avdd.n7292 0.018303
R10559 avdd.n7367 avdd.n7206 0.018303
R10560 avdd.n7777 avdd.n7776 0.018303
R10561 avdd.n7723 avdd.n7722 0.018303
R10562 avdd.n7813 avdd.n7812 0.018303
R10563 avdd.n10037 avdd.n10036 0.018303
R10564 avdd.n10202 avdd.n10201 0.018303
R10565 avdd.n10071 avdd.n10070 0.018303
R10566 avdd.n10253 avdd.n10252 0.018303
R10567 avdd.n10009 avdd.n10008 0.018303
R10568 avdd.n10303 avdd.n10302 0.018303
R10569 avdd.n10355 avdd.n10354 0.018303
R10570 avdd.n9895 avdd.n9894 0.018303
R10571 avdd.n10405 avdd.n10404 0.018303
R10572 avdd.n10457 avdd.n10456 0.018303
R10573 avdd.n9781 avdd.n9780 0.018303
R10574 avdd.n10507 avdd.n10506 0.018303
R10575 avdd.n10559 avdd.n10558 0.018303
R10576 avdd.n9668 avdd.n9667 0.018303
R10577 avdd.n10609 avdd.n10608 0.018303
R10578 avdd.n10661 avdd.n10660 0.018303
R10579 avdd.n9553 avdd.n9552 0.018303
R10580 avdd.n10711 avdd.n10710 0.018303
R10581 avdd.n10763 avdd.n10762 0.018303
R10582 avdd.n9439 avdd.n9438 0.018303
R10583 avdd.n10813 avdd.n10812 0.018303
R10584 avdd.n10865 avdd.n10864 0.018303
R10585 avdd.n9325 avdd.n9324 0.018303
R10586 avdd.n10915 avdd.n10914 0.018303
R10587 avdd.n10967 avdd.n10966 0.018303
R10588 avdd.n9211 avdd.n9210 0.018303
R10589 avdd.n11017 avdd.n11016 0.018303
R10590 avdd.n11069 avdd.n11068 0.018303
R10591 avdd.n9097 avdd.n9096 0.018303
R10592 avdd.n11119 avdd.n11118 0.018303
R10593 avdd.n11171 avdd.n11170 0.018303
R10594 avdd.n8983 avdd.n8982 0.018303
R10595 avdd.n11221 avdd.n11220 0.018303
R10596 avdd.n8880 avdd.n8879 0.018303
R10597 avdd.n8834 avdd.n8833 0.018303
R10598 avdd.n8794 avdd.n8793 0.018303
R10599 avdd.n8748 avdd.n8747 0.018303
R10600 avdd.n8708 avdd.n8707 0.018303
R10601 avdd.n8662 avdd.n8661 0.018303
R10602 avdd.n8622 avdd.n8621 0.018303
R10603 avdd.n8576 avdd.n8575 0.018303
R10604 avdd.n8536 avdd.n8535 0.018303
R10605 avdd.n8490 avdd.n8489 0.018303
R10606 avdd.n8450 avdd.n8449 0.018303
R10607 avdd.n8404 avdd.n8403 0.018303
R10608 avdd.n8364 avdd.n8363 0.018303
R10609 avdd.n8318 avdd.n8317 0.018303
R10610 avdd.n8278 avdd.n8277 0.018303
R10611 avdd.n8232 avdd.n8231 0.018303
R10612 avdd.n8192 avdd.n8191 0.018303
R10613 avdd.n8146 avdd.n8145 0.018303
R10614 avdd.n8106 avdd.n8105 0.018303
R10615 avdd.n8060 avdd.n8059 0.018303
R10616 avdd.n8020 avdd.n8019 0.018303
R10617 avdd.n7974 avdd.n7973 0.018303
R10618 avdd.n7934 avdd.n7933 0.018303
R10619 avdd.n7888 avdd.n7887 0.018303
R10620 avdd.n4629 avdd.n4628 0.0171667
R10621 avdd.n2071 avdd.n1956 0.0168788
R10622 avdd.n2211 avdd.n2122 0.0168788
R10623 avdd.n2426 avdd.n2337 0.0168788
R10624 avdd.n2641 avdd.n2552 0.0168788
R10625 avdd.n2856 avdd.n2767 0.0168788
R10626 avdd.n3071 avdd.n2982 0.0168788
R10627 avdd.n3360 avdd.n3246 0.0168788
R10628 avdd.n3575 avdd.n3461 0.0168788
R10629 avdd.n3790 avdd.n3676 0.0168788
R10630 avdd.n4005 avdd.n3891 0.0168788
R10631 avdd.n4220 avdd.n4106 0.0168788
R10632 avdd.n4435 avdd.n4321 0.0168788
R10633 avdd.n4933 avdd.n4844 0.0168788
R10634 avdd.n5149 avdd.n5060 0.0168788
R10635 avdd.n5365 avdd.n5276 0.0168788
R10636 avdd.n5581 avdd.n5492 0.0168788
R10637 avdd.n5797 avdd.n5708 0.0168788
R10638 avdd.n6013 avdd.n5924 0.0168788
R10639 avdd.n6229 avdd.n6140 0.0168788
R10640 avdd.n6445 avdd.n6356 0.0168788
R10641 avdd.n6661 avdd.n6572 0.0168788
R10642 avdd.n6877 avdd.n6788 0.0168788
R10643 avdd.n7093 avdd.n7004 0.0168788
R10644 avdd.n7309 avdd.n7220 0.0168788
R10645 avdd.n7645 avdd.n7644 0.0168788
R10646 avdd.n10122 avdd.n10121 0.0168788
R10647 avdd.n9923 avdd.n9922 0.0168788
R10648 avdd.n9809 avdd.n9808 0.0168788
R10649 avdd.n9695 avdd.n9694 0.0168788
R10650 avdd.n9581 avdd.n9580 0.0168788
R10651 avdd.n9467 avdd.n9466 0.0168788
R10652 avdd.n9353 avdd.n9352 0.0168788
R10653 avdd.n9239 avdd.n9238 0.0168788
R10654 avdd.n9125 avdd.n9124 0.0168788
R10655 avdd.n9011 avdd.n9010 0.0168788
R10656 avdd.n8897 avdd.n8896 0.0168788
R10657 avdd.n66 avdd.n65 0.0168788
R10658 avdd.n196 avdd.n195 0.0168788
R10659 avdd.n326 avdd.n325 0.0168788
R10660 avdd.n456 avdd.n455 0.0168788
R10661 avdd.n586 avdd.n585 0.0168788
R10662 avdd.n716 avdd.n715 0.0168788
R10663 avdd.n846 avdd.n845 0.0168788
R10664 avdd.n976 avdd.n975 0.0168788
R10665 avdd.n1106 avdd.n1105 0.0168788
R10666 avdd.n1236 avdd.n1235 0.0168788
R10667 avdd.n1366 avdd.n1365 0.0168788
R10668 avdd.n1496 avdd.n1495 0.0168788
R10669 avdd.n1988 avdd.n1987 0.0154545
R10670 avdd.n1928 avdd.n1927 0.0154545
R10671 avdd.n1929 avdd.n1896 0.0154545
R10672 avdd.n1989 avdd.n1986 0.0154545
R10673 avdd.n2257 avdd.n2256 0.0154545
R10674 avdd.n2181 avdd.n2143 0.0154545
R10675 avdd.n2182 avdd.n2150 0.0154545
R10676 avdd.n2258 avdd.n2113 0.0154545
R10677 avdd.n2472 avdd.n2471 0.0154545
R10678 avdd.n2396 avdd.n2358 0.0154545
R10679 avdd.n2397 avdd.n2365 0.0154545
R10680 avdd.n2473 avdd.n2328 0.0154545
R10681 avdd.n2687 avdd.n2686 0.0154545
R10682 avdd.n2611 avdd.n2573 0.0154545
R10683 avdd.n2612 avdd.n2580 0.0154545
R10684 avdd.n2688 avdd.n2543 0.0154545
R10685 avdd.n2902 avdd.n2901 0.0154545
R10686 avdd.n2826 avdd.n2788 0.0154545
R10687 avdd.n2827 avdd.n2795 0.0154545
R10688 avdd.n2903 avdd.n2758 0.0154545
R10689 avdd.n3117 avdd.n3116 0.0154545
R10690 avdd.n3041 avdd.n3003 0.0154545
R10691 avdd.n3042 avdd.n3010 0.0154545
R10692 avdd.n3118 avdd.n2973 0.0154545
R10693 avdd.n3278 avdd.n3277 0.0154545
R10694 avdd.n3218 avdd.n3217 0.0154545
R10695 avdd.n3219 avdd.n3186 0.0154545
R10696 avdd.n3279 avdd.n3276 0.0154545
R10697 avdd.n3493 avdd.n3492 0.0154545
R10698 avdd.n3433 avdd.n3432 0.0154545
R10699 avdd.n3434 avdd.n3401 0.0154545
R10700 avdd.n3494 avdd.n3491 0.0154545
R10701 avdd.n3708 avdd.n3707 0.0154545
R10702 avdd.n3648 avdd.n3647 0.0154545
R10703 avdd.n3649 avdd.n3616 0.0154545
R10704 avdd.n3709 avdd.n3706 0.0154545
R10705 avdd.n3923 avdd.n3922 0.0154545
R10706 avdd.n3863 avdd.n3862 0.0154545
R10707 avdd.n3864 avdd.n3831 0.0154545
R10708 avdd.n3924 avdd.n3921 0.0154545
R10709 avdd.n4138 avdd.n4137 0.0154545
R10710 avdd.n4078 avdd.n4077 0.0154545
R10711 avdd.n4079 avdd.n4046 0.0154545
R10712 avdd.n4139 avdd.n4136 0.0154545
R10713 avdd.n4353 avdd.n4352 0.0154545
R10714 avdd.n4293 avdd.n4292 0.0154545
R10715 avdd.n4294 avdd.n4261 0.0154545
R10716 avdd.n4354 avdd.n4351 0.0154545
R10717 avdd.n4979 avdd.n4978 0.0154545
R10718 avdd.n4904 avdd.n4903 0.0154545
R10719 avdd.n4905 avdd.n4872 0.0154545
R10720 avdd.n4980 avdd.n4835 0.0154545
R10721 avdd.n5195 avdd.n5194 0.0154545
R10722 avdd.n5120 avdd.n5119 0.0154545
R10723 avdd.n5121 avdd.n5088 0.0154545
R10724 avdd.n5196 avdd.n5051 0.0154545
R10725 avdd.n5411 avdd.n5410 0.0154545
R10726 avdd.n5336 avdd.n5335 0.0154545
R10727 avdd.n5337 avdd.n5304 0.0154545
R10728 avdd.n5412 avdd.n5267 0.0154545
R10729 avdd.n5627 avdd.n5626 0.0154545
R10730 avdd.n5552 avdd.n5551 0.0154545
R10731 avdd.n5553 avdd.n5520 0.0154545
R10732 avdd.n5628 avdd.n5483 0.0154545
R10733 avdd.n5843 avdd.n5842 0.0154545
R10734 avdd.n5768 avdd.n5767 0.0154545
R10735 avdd.n5769 avdd.n5736 0.0154545
R10736 avdd.n5844 avdd.n5699 0.0154545
R10737 avdd.n6059 avdd.n6058 0.0154545
R10738 avdd.n5984 avdd.n5983 0.0154545
R10739 avdd.n5985 avdd.n5952 0.0154545
R10740 avdd.n6060 avdd.n5915 0.0154545
R10741 avdd.n6275 avdd.n6274 0.0154545
R10742 avdd.n6200 avdd.n6199 0.0154545
R10743 avdd.n6201 avdd.n6168 0.0154545
R10744 avdd.n6276 avdd.n6131 0.0154545
R10745 avdd.n6491 avdd.n6490 0.0154545
R10746 avdd.n6416 avdd.n6415 0.0154545
R10747 avdd.n6417 avdd.n6384 0.0154545
R10748 avdd.n6492 avdd.n6347 0.0154545
R10749 avdd.n6707 avdd.n6706 0.0154545
R10750 avdd.n6632 avdd.n6631 0.0154545
R10751 avdd.n6633 avdd.n6600 0.0154545
R10752 avdd.n6708 avdd.n6563 0.0154545
R10753 avdd.n6923 avdd.n6922 0.0154545
R10754 avdd.n6848 avdd.n6847 0.0154545
R10755 avdd.n6849 avdd.n6816 0.0154545
R10756 avdd.n6924 avdd.n6779 0.0154545
R10757 avdd.n7139 avdd.n7138 0.0154545
R10758 avdd.n7064 avdd.n7063 0.0154545
R10759 avdd.n7065 avdd.n7032 0.0154545
R10760 avdd.n7140 avdd.n6995 0.0154545
R10761 avdd.n7355 avdd.n7354 0.0154545
R10762 avdd.n7280 avdd.n7279 0.0154545
R10763 avdd.n7281 avdd.n7248 0.0154545
R10764 avdd.n7356 avdd.n7211 0.0154545
R10765 avdd.n7773 avdd.n7772 0.0154545
R10766 avdd.n7761 avdd.n7760 0.0154545
R10767 avdd.n7720 avdd.n7719 0.0154545
R10768 avdd.n7809 avdd.n7808 0.0154545
R10769 avdd.n10033 avdd.n10032 0.0154545
R10770 avdd.n10240 avdd.n10239 0.0154545
R10771 avdd.n10199 avdd.n10198 0.0154545
R10772 avdd.n10067 avdd.n10066 0.0154545
R10773 avdd.n10249 avdd.n10248 0.0154545
R10774 avdd.n10005 avdd.n10004 0.0154545
R10775 avdd.n10003 avdd.n10002 0.0154545
R10776 avdd.n10299 avdd.n10298 0.0154545
R10777 avdd.n10351 avdd.n10350 0.0154545
R10778 avdd.n9891 avdd.n9890 0.0154545
R10779 avdd.n9889 avdd.n9888 0.0154545
R10780 avdd.n10401 avdd.n10400 0.0154545
R10781 avdd.n10453 avdd.n10452 0.0154545
R10782 avdd.n9777 avdd.n9776 0.0154545
R10783 avdd.n9775 avdd.n9774 0.0154545
R10784 avdd.n10503 avdd.n10502 0.0154545
R10785 avdd.n10555 avdd.n10554 0.0154545
R10786 avdd.n9664 avdd.n9663 0.0154545
R10787 avdd.n9662 avdd.n9661 0.0154545
R10788 avdd.n10605 avdd.n10604 0.0154545
R10789 avdd.n10657 avdd.n10656 0.0154545
R10790 avdd.n9549 avdd.n9548 0.0154545
R10791 avdd.n9547 avdd.n9546 0.0154545
R10792 avdd.n10707 avdd.n10706 0.0154545
R10793 avdd.n10759 avdd.n10758 0.0154545
R10794 avdd.n9435 avdd.n9434 0.0154545
R10795 avdd.n9433 avdd.n9432 0.0154545
R10796 avdd.n10809 avdd.n10808 0.0154545
R10797 avdd.n10861 avdd.n10860 0.0154545
R10798 avdd.n9321 avdd.n9320 0.0154545
R10799 avdd.n9319 avdd.n9318 0.0154545
R10800 avdd.n10911 avdd.n10910 0.0154545
R10801 avdd.n10963 avdd.n10962 0.0154545
R10802 avdd.n9207 avdd.n9206 0.0154545
R10803 avdd.n9205 avdd.n9204 0.0154545
R10804 avdd.n11013 avdd.n11012 0.0154545
R10805 avdd.n11065 avdd.n11064 0.0154545
R10806 avdd.n9093 avdd.n9092 0.0154545
R10807 avdd.n9091 avdd.n9090 0.0154545
R10808 avdd.n11115 avdd.n11114 0.0154545
R10809 avdd.n11167 avdd.n11166 0.0154545
R10810 avdd.n8979 avdd.n8978 0.0154545
R10811 avdd.n8977 avdd.n8976 0.0154545
R10812 avdd.n11217 avdd.n11216 0.0154545
R10813 avdd.n8876 avdd.n8875 0.0154545
R10814 avdd.n94 avdd.n93 0.0154545
R10815 avdd.n114 avdd.n113 0.0154545
R10816 avdd.n8830 avdd.n8829 0.0154545
R10817 avdd.n8790 avdd.n8789 0.0154545
R10818 avdd.n224 avdd.n223 0.0154545
R10819 avdd.n244 avdd.n243 0.0154545
R10820 avdd.n8744 avdd.n8743 0.0154545
R10821 avdd.n8704 avdd.n8703 0.0154545
R10822 avdd.n354 avdd.n353 0.0154545
R10823 avdd.n374 avdd.n373 0.0154545
R10824 avdd.n8658 avdd.n8657 0.0154545
R10825 avdd.n8618 avdd.n8617 0.0154545
R10826 avdd.n484 avdd.n483 0.0154545
R10827 avdd.n504 avdd.n503 0.0154545
R10828 avdd.n8572 avdd.n8571 0.0154545
R10829 avdd.n8532 avdd.n8531 0.0154545
R10830 avdd.n614 avdd.n613 0.0154545
R10831 avdd.n634 avdd.n633 0.0154545
R10832 avdd.n8486 avdd.n8485 0.0154545
R10833 avdd.n8446 avdd.n8445 0.0154545
R10834 avdd.n744 avdd.n743 0.0154545
R10835 avdd.n764 avdd.n763 0.0154545
R10836 avdd.n8400 avdd.n8399 0.0154545
R10837 avdd.n8360 avdd.n8359 0.0154545
R10838 avdd.n874 avdd.n873 0.0154545
R10839 avdd.n894 avdd.n893 0.0154545
R10840 avdd.n8314 avdd.n8313 0.0154545
R10841 avdd.n8274 avdd.n8273 0.0154545
R10842 avdd.n1004 avdd.n1003 0.0154545
R10843 avdd.n1024 avdd.n1023 0.0154545
R10844 avdd.n8228 avdd.n8227 0.0154545
R10845 avdd.n8188 avdd.n8187 0.0154545
R10846 avdd.n1134 avdd.n1133 0.0154545
R10847 avdd.n1154 avdd.n1153 0.0154545
R10848 avdd.n8142 avdd.n8141 0.0154545
R10849 avdd.n8102 avdd.n8101 0.0154545
R10850 avdd.n1264 avdd.n1263 0.0154545
R10851 avdd.n1284 avdd.n1283 0.0154545
R10852 avdd.n8056 avdd.n8055 0.0154545
R10853 avdd.n8016 avdd.n8015 0.0154545
R10854 avdd.n1394 avdd.n1393 0.0154545
R10855 avdd.n1414 avdd.n1413 0.0154545
R10856 avdd.n7970 avdd.n7969 0.0154545
R10857 avdd.n7930 avdd.n7929 0.0154545
R10858 avdd.n1524 avdd.n1523 0.0154545
R10859 avdd.n1544 avdd.n1543 0.0154545
R10860 avdd.n7884 avdd.n7883 0.0154545
R10861 avdd.n4640 avdd.n4616 0.0150833
R10862 avdd.n4586 avdd.n4574 0.0150833
R10863 avdd.n4464 avdd 0.0149231
R10864 avdd.n2073 avdd.n1949 0.0147424
R10865 avdd.n2212 avdd.n2210 0.0147424
R10866 avdd.n2427 avdd.n2425 0.0147424
R10867 avdd.n2642 avdd.n2640 0.0147424
R10868 avdd.n2857 avdd.n2855 0.0147424
R10869 avdd.n3072 avdd.n3070 0.0147424
R10870 avdd.n3362 avdd.n3239 0.0147424
R10871 avdd.n3577 avdd.n3454 0.0147424
R10872 avdd.n3792 avdd.n3669 0.0147424
R10873 avdd.n4007 avdd.n3884 0.0147424
R10874 avdd.n4222 avdd.n4099 0.0147424
R10875 avdd.n4437 avdd.n4314 0.0147424
R10876 avdd.n4934 avdd.n4932 0.0147424
R10877 avdd.n5150 avdd.n5148 0.0147424
R10878 avdd.n5366 avdd.n5364 0.0147424
R10879 avdd.n5582 avdd.n5580 0.0147424
R10880 avdd.n5798 avdd.n5796 0.0147424
R10881 avdd.n6014 avdd.n6012 0.0147424
R10882 avdd.n6230 avdd.n6228 0.0147424
R10883 avdd.n6446 avdd.n6444 0.0147424
R10884 avdd.n6662 avdd.n6660 0.0147424
R10885 avdd.n6878 avdd.n6876 0.0147424
R10886 avdd.n7094 avdd.n7092 0.0147424
R10887 avdd.n7310 avdd.n7308 0.0147424
R10888 avdd.n7681 avdd.n7680 0.0147424
R10889 avdd.n10160 avdd.n10159 0.0147424
R10890 avdd.n9944 avdd.n9943 0.0147424
R10891 avdd.n9830 avdd.n9829 0.0147424
R10892 avdd.n9716 avdd.n9715 0.0147424
R10893 avdd.n9603 avdd.n9602 0.0147424
R10894 avdd.n9488 avdd.n9487 0.0147424
R10895 avdd.n9374 avdd.n9373 0.0147424
R10896 avdd.n9260 avdd.n9259 0.0147424
R10897 avdd.n9146 avdd.n9145 0.0147424
R10898 avdd.n9032 avdd.n9031 0.0147424
R10899 avdd.n8918 avdd.n8917 0.0147424
R10900 avdd.n164 avdd.n163 0.0147424
R10901 avdd.n294 avdd.n293 0.0147424
R10902 avdd.n424 avdd.n423 0.0147424
R10903 avdd.n554 avdd.n553 0.0147424
R10904 avdd.n684 avdd.n683 0.0147424
R10905 avdd.n814 avdd.n813 0.0147424
R10906 avdd.n944 avdd.n943 0.0147424
R10907 avdd.n1074 avdd.n1073 0.0147424
R10908 avdd.n1204 avdd.n1203 0.0147424
R10909 avdd.n1334 avdd.n1333 0.0147424
R10910 avdd.n1464 avdd.n1463 0.0147424
R10911 avdd.n1594 avdd.n1593 0.0147424
R10912 avdd.n2045 avdd.n1994 0.0140303
R10913 avdd.n1927 avdd.n1878 0.0140303
R10914 avdd.n2276 avdd.n2271 0.0140303
R10915 avdd.n2195 avdd.n2143 0.0140303
R10916 avdd.n2491 avdd.n2486 0.0140303
R10917 avdd.n2410 avdd.n2358 0.0140303
R10918 avdd.n2706 avdd.n2701 0.0140303
R10919 avdd.n2625 avdd.n2573 0.0140303
R10920 avdd.n2921 avdd.n2916 0.0140303
R10921 avdd.n2840 avdd.n2788 0.0140303
R10922 avdd.n3136 avdd.n3131 0.0140303
R10923 avdd.n3055 avdd.n3003 0.0140303
R10924 avdd.n3334 avdd.n3284 0.0140303
R10925 avdd.n3217 avdd.n3169 0.0140303
R10926 avdd.n3549 avdd.n3499 0.0140303
R10927 avdd.n3432 avdd.n3384 0.0140303
R10928 avdd.n3764 avdd.n3714 0.0140303
R10929 avdd.n3647 avdd.n3599 0.0140303
R10930 avdd.n3979 avdd.n3929 0.0140303
R10931 avdd.n3862 avdd.n3814 0.0140303
R10932 avdd.n4194 avdd.n4144 0.0140303
R10933 avdd.n4077 avdd.n4029 0.0140303
R10934 avdd.n4409 avdd.n4359 0.0140303
R10935 avdd.n4292 avdd.n4244 0.0140303
R10936 avdd.n4995 avdd.n4993 0.0140303
R10937 avdd.n4903 avdd.n4866 0.0140303
R10938 avdd.n5211 avdd.n5209 0.0140303
R10939 avdd.n5119 avdd.n5082 0.0140303
R10940 avdd.n5427 avdd.n5425 0.0140303
R10941 avdd.n5335 avdd.n5298 0.0140303
R10942 avdd.n5643 avdd.n5641 0.0140303
R10943 avdd.n5551 avdd.n5514 0.0140303
R10944 avdd.n5859 avdd.n5857 0.0140303
R10945 avdd.n5767 avdd.n5730 0.0140303
R10946 avdd.n6075 avdd.n6073 0.0140303
R10947 avdd.n5983 avdd.n5946 0.0140303
R10948 avdd.n6291 avdd.n6289 0.0140303
R10949 avdd.n6199 avdd.n6162 0.0140303
R10950 avdd.n6507 avdd.n6505 0.0140303
R10951 avdd.n6415 avdd.n6378 0.0140303
R10952 avdd.n6723 avdd.n6721 0.0140303
R10953 avdd.n6631 avdd.n6594 0.0140303
R10954 avdd.n6939 avdd.n6937 0.0140303
R10955 avdd.n6847 avdd.n6810 0.0140303
R10956 avdd.n7155 avdd.n7153 0.0140303
R10957 avdd.n7063 avdd.n7026 0.0140303
R10958 avdd.n7371 avdd.n7369 0.0140303
R10959 avdd.n7279 avdd.n7242 0.0140303
R10960 avdd.n7779 avdd.n7778 0.0140303
R10961 avdd.n7762 avdd.n7761 0.0140303
R10962 avdd.n10039 avdd.n10038 0.0140303
R10963 avdd.n10241 avdd.n10240 0.0140303
R10964 avdd.n10255 avdd.n10254 0.0140303
R10965 avdd.n10027 avdd.n10005 0.0140303
R10966 avdd.n10357 avdd.n10356 0.0140303
R10967 avdd.n9913 avdd.n9891 0.0140303
R10968 avdd.n10459 avdd.n10458 0.0140303
R10969 avdd.n9799 avdd.n9777 0.0140303
R10970 avdd.n10561 avdd.n10560 0.0140303
R10971 avdd.n9685 avdd.n9664 0.0140303
R10972 avdd.n10663 avdd.n10662 0.0140303
R10973 avdd.n9571 avdd.n9549 0.0140303
R10974 avdd.n10765 avdd.n10764 0.0140303
R10975 avdd.n9457 avdd.n9435 0.0140303
R10976 avdd.n10867 avdd.n10866 0.0140303
R10977 avdd.n9343 avdd.n9321 0.0140303
R10978 avdd.n10969 avdd.n10968 0.0140303
R10979 avdd.n9229 avdd.n9207 0.0140303
R10980 avdd.n11071 avdd.n11070 0.0140303
R10981 avdd.n9115 avdd.n9093 0.0140303
R10982 avdd.n11173 avdd.n11172 0.0140303
R10983 avdd.n9001 avdd.n8979 0.0140303
R10984 avdd.n8882 avdd.n8881 0.0140303
R10985 avdd.n186 avdd.n94 0.0140303
R10986 avdd.n8796 avdd.n8795 0.0140303
R10987 avdd.n316 avdd.n224 0.0140303
R10988 avdd.n8710 avdd.n8709 0.0140303
R10989 avdd.n446 avdd.n354 0.0140303
R10990 avdd.n8624 avdd.n8623 0.0140303
R10991 avdd.n576 avdd.n484 0.0140303
R10992 avdd.n8538 avdd.n8537 0.0140303
R10993 avdd.n706 avdd.n614 0.0140303
R10994 avdd.n8452 avdd.n8451 0.0140303
R10995 avdd.n836 avdd.n744 0.0140303
R10996 avdd.n8366 avdd.n8365 0.0140303
R10997 avdd.n966 avdd.n874 0.0140303
R10998 avdd.n8280 avdd.n8279 0.0140303
R10999 avdd.n1096 avdd.n1004 0.0140303
R11000 avdd.n8194 avdd.n8193 0.0140303
R11001 avdd.n1226 avdd.n1134 0.0140303
R11002 avdd.n8108 avdd.n8107 0.0140303
R11003 avdd.n1356 avdd.n1264 0.0140303
R11004 avdd.n8022 avdd.n8021 0.0140303
R11005 avdd.n1486 avdd.n1394 0.0140303
R11006 avdd.n7936 avdd.n7935 0.0140303
R11007 avdd.n1616 avdd.n1524 0.0140303
R11008 avdd.n2014 avdd.n2012 0.0137576
R11009 avdd.n1983 avdd.n1975 0.0137576
R11010 avdd.n2081 avdd.n1887 0.0137576
R11011 avdd.n1920 avdd.n1893 0.0137576
R11012 avdd.n2287 avdd.n2101 0.0137576
R11013 avdd.n2245 avdd.n2111 0.0137576
R11014 avdd.n2204 avdd.n2130 0.0137576
R11015 avdd.n2174 avdd.n2148 0.0137576
R11016 avdd.n2502 avdd.n2316 0.0137576
R11017 avdd.n2460 avdd.n2326 0.0137576
R11018 avdd.n2419 avdd.n2345 0.0137576
R11019 avdd.n2389 avdd.n2363 0.0137576
R11020 avdd.n2717 avdd.n2531 0.0137576
R11021 avdd.n2675 avdd.n2541 0.0137576
R11022 avdd.n2634 avdd.n2560 0.0137576
R11023 avdd.n2604 avdd.n2578 0.0137576
R11024 avdd.n2932 avdd.n2746 0.0137576
R11025 avdd.n2890 avdd.n2756 0.0137576
R11026 avdd.n2849 avdd.n2775 0.0137576
R11027 avdd.n2819 avdd.n2793 0.0137576
R11028 avdd.n3147 avdd.n2961 0.0137576
R11029 avdd.n3105 avdd.n2971 0.0137576
R11030 avdd.n3064 avdd.n2990 0.0137576
R11031 avdd.n3034 avdd.n3008 0.0137576
R11032 avdd.n3310 avdd.n3307 0.0137576
R11033 avdd.n3273 avdd.n3265 0.0137576
R11034 avdd.n3370 avdd.n3177 0.0137576
R11035 avdd.n3210 avdd.n3183 0.0137576
R11036 avdd.n3525 avdd.n3522 0.0137576
R11037 avdd.n3488 avdd.n3480 0.0137576
R11038 avdd.n3585 avdd.n3392 0.0137576
R11039 avdd.n3425 avdd.n3398 0.0137576
R11040 avdd.n3740 avdd.n3737 0.0137576
R11041 avdd.n3703 avdd.n3695 0.0137576
R11042 avdd.n3800 avdd.n3607 0.0137576
R11043 avdd.n3640 avdd.n3613 0.0137576
R11044 avdd.n3955 avdd.n3952 0.0137576
R11045 avdd.n3918 avdd.n3910 0.0137576
R11046 avdd.n4015 avdd.n3822 0.0137576
R11047 avdd.n3855 avdd.n3828 0.0137576
R11048 avdd.n4170 avdd.n4167 0.0137576
R11049 avdd.n4133 avdd.n4125 0.0137576
R11050 avdd.n4230 avdd.n4037 0.0137576
R11051 avdd.n4070 avdd.n4043 0.0137576
R11052 avdd.n4385 avdd.n4382 0.0137576
R11053 avdd.n4348 avdd.n4340 0.0137576
R11054 avdd.n4445 avdd.n4252 0.0137576
R11055 avdd.n4285 avdd.n4258 0.0137576
R11056 avdd.n4896 avdd.n4870 0.0137576
R11057 avdd.n4926 avdd.n4852 0.0137576
R11058 avdd.n4967 avdd.n4833 0.0137576
R11059 avdd.n5005 avdd.n4822 0.0137576
R11060 avdd.n5112 avdd.n5086 0.0137576
R11061 avdd.n5142 avdd.n5068 0.0137576
R11062 avdd.n5183 avdd.n5049 0.0137576
R11063 avdd.n5221 avdd.n5038 0.0137576
R11064 avdd.n5328 avdd.n5302 0.0137576
R11065 avdd.n5358 avdd.n5284 0.0137576
R11066 avdd.n5399 avdd.n5265 0.0137576
R11067 avdd.n5437 avdd.n5254 0.0137576
R11068 avdd.n5544 avdd.n5518 0.0137576
R11069 avdd.n5574 avdd.n5500 0.0137576
R11070 avdd.n5615 avdd.n5481 0.0137576
R11071 avdd.n5653 avdd.n5470 0.0137576
R11072 avdd.n5760 avdd.n5734 0.0137576
R11073 avdd.n5790 avdd.n5716 0.0137576
R11074 avdd.n5831 avdd.n5697 0.0137576
R11075 avdd.n5869 avdd.n5686 0.0137576
R11076 avdd.n5976 avdd.n5950 0.0137576
R11077 avdd.n6006 avdd.n5932 0.0137576
R11078 avdd.n6047 avdd.n5913 0.0137576
R11079 avdd.n6085 avdd.n5902 0.0137576
R11080 avdd.n6192 avdd.n6166 0.0137576
R11081 avdd.n6222 avdd.n6148 0.0137576
R11082 avdd.n6263 avdd.n6129 0.0137576
R11083 avdd.n6301 avdd.n6118 0.0137576
R11084 avdd.n6408 avdd.n6382 0.0137576
R11085 avdd.n6438 avdd.n6364 0.0137576
R11086 avdd.n6479 avdd.n6345 0.0137576
R11087 avdd.n6517 avdd.n6334 0.0137576
R11088 avdd.n6624 avdd.n6598 0.0137576
R11089 avdd.n6654 avdd.n6580 0.0137576
R11090 avdd.n6695 avdd.n6561 0.0137576
R11091 avdd.n6733 avdd.n6550 0.0137576
R11092 avdd.n6840 avdd.n6814 0.0137576
R11093 avdd.n6870 avdd.n6796 0.0137576
R11094 avdd.n6911 avdd.n6777 0.0137576
R11095 avdd.n6949 avdd.n6766 0.0137576
R11096 avdd.n7056 avdd.n7030 0.0137576
R11097 avdd.n7086 avdd.n7012 0.0137576
R11098 avdd.n7127 avdd.n6993 0.0137576
R11099 avdd.n7165 avdd.n6982 0.0137576
R11100 avdd.n7272 avdd.n7246 0.0137576
R11101 avdd.n7302 avdd.n7228 0.0137576
R11102 avdd.n7343 avdd.n7209 0.0137576
R11103 avdd.n7381 avdd.n7198 0.0137576
R11104 avdd.n7715 avdd.n7714 0.0137576
R11105 avdd.n7695 avdd.n7694 0.0137576
R11106 avdd.n7804 avdd.n7803 0.0137576
R11107 avdd.n7842 avdd.n7841 0.0137576
R11108 avdd.n10194 avdd.n10193 0.0137576
R11109 avdd.n10174 avdd.n10173 0.0137576
R11110 avdd.n10062 avdd.n10061 0.0137576
R11111 avdd.n10100 avdd.n10099 0.0137576
R11112 avdd.n9998 avdd.n9997 0.0137576
R11113 avdd.n9958 avdd.n9957 0.0137576
R11114 avdd.n10294 avdd.n10293 0.0137576
R11115 avdd.n10332 avdd.n10331 0.0137576
R11116 avdd.n9884 avdd.n9883 0.0137576
R11117 avdd.n9844 avdd.n9843 0.0137576
R11118 avdd.n10396 avdd.n10395 0.0137576
R11119 avdd.n10434 avdd.n10433 0.0137576
R11120 avdd.n9770 avdd.n9769 0.0137576
R11121 avdd.n9730 avdd.n9729 0.0137576
R11122 avdd.n10498 avdd.n10497 0.0137576
R11123 avdd.n10536 avdd.n10535 0.0137576
R11124 avdd.n9657 avdd.n9656 0.0137576
R11125 avdd.n9617 avdd.n9616 0.0137576
R11126 avdd.n10600 avdd.n10599 0.0137576
R11127 avdd.n10638 avdd.n10637 0.0137576
R11128 avdd.n9542 avdd.n9541 0.0137576
R11129 avdd.n9502 avdd.n9501 0.0137576
R11130 avdd.n10702 avdd.n10701 0.0137576
R11131 avdd.n10740 avdd.n10739 0.0137576
R11132 avdd.n9428 avdd.n9427 0.0137576
R11133 avdd.n9388 avdd.n9387 0.0137576
R11134 avdd.n10804 avdd.n10803 0.0137576
R11135 avdd.n10842 avdd.n10841 0.0137576
R11136 avdd.n9314 avdd.n9313 0.0137576
R11137 avdd.n9274 avdd.n9273 0.0137576
R11138 avdd.n10906 avdd.n10905 0.0137576
R11139 avdd.n10944 avdd.n10943 0.0137576
R11140 avdd.n9200 avdd.n9199 0.0137576
R11141 avdd.n9160 avdd.n9159 0.0137576
R11142 avdd.n11008 avdd.n11007 0.0137576
R11143 avdd.n11046 avdd.n11045 0.0137576
R11144 avdd.n9086 avdd.n9085 0.0137576
R11145 avdd.n9046 avdd.n9045 0.0137576
R11146 avdd.n11110 avdd.n11109 0.0137576
R11147 avdd.n11148 avdd.n11147 0.0137576
R11148 avdd.n8972 avdd.n8971 0.0137576
R11149 avdd.n8932 avdd.n8931 0.0137576
R11150 avdd.n11212 avdd.n11211 0.0137576
R11151 avdd.n11250 avdd.n11249 0.0137576
R11152 avdd.n8863 avdd.n8862 0.0137576
R11153 avdd.n8825 avdd.n8824 0.0137576
R11154 avdd.n178 avdd.n177 0.0137576
R11155 avdd.n109 avdd.n108 0.0137576
R11156 avdd.n8777 avdd.n8776 0.0137576
R11157 avdd.n8739 avdd.n8738 0.0137576
R11158 avdd.n308 avdd.n307 0.0137576
R11159 avdd.n239 avdd.n238 0.0137576
R11160 avdd.n8691 avdd.n8690 0.0137576
R11161 avdd.n8653 avdd.n8652 0.0137576
R11162 avdd.n438 avdd.n437 0.0137576
R11163 avdd.n369 avdd.n368 0.0137576
R11164 avdd.n8605 avdd.n8604 0.0137576
R11165 avdd.n8567 avdd.n8566 0.0137576
R11166 avdd.n568 avdd.n567 0.0137576
R11167 avdd.n499 avdd.n498 0.0137576
R11168 avdd.n8519 avdd.n8518 0.0137576
R11169 avdd.n8481 avdd.n8480 0.0137576
R11170 avdd.n698 avdd.n697 0.0137576
R11171 avdd.n629 avdd.n628 0.0137576
R11172 avdd.n8433 avdd.n8432 0.0137576
R11173 avdd.n8395 avdd.n8394 0.0137576
R11174 avdd.n828 avdd.n827 0.0137576
R11175 avdd.n759 avdd.n758 0.0137576
R11176 avdd.n8347 avdd.n8346 0.0137576
R11177 avdd.n8309 avdd.n8308 0.0137576
R11178 avdd.n958 avdd.n957 0.0137576
R11179 avdd.n889 avdd.n888 0.0137576
R11180 avdd.n8261 avdd.n8260 0.0137576
R11181 avdd.n8223 avdd.n8222 0.0137576
R11182 avdd.n1088 avdd.n1087 0.0137576
R11183 avdd.n1019 avdd.n1018 0.0137576
R11184 avdd.n8175 avdd.n8174 0.0137576
R11185 avdd.n8137 avdd.n8136 0.0137576
R11186 avdd.n1218 avdd.n1217 0.0137576
R11187 avdd.n1149 avdd.n1148 0.0137576
R11188 avdd.n8089 avdd.n8088 0.0137576
R11189 avdd.n8051 avdd.n8050 0.0137576
R11190 avdd.n1348 avdd.n1347 0.0137576
R11191 avdd.n1279 avdd.n1278 0.0137576
R11192 avdd.n8003 avdd.n8002 0.0137576
R11193 avdd.n7965 avdd.n7964 0.0137576
R11194 avdd.n1478 avdd.n1477 0.0137576
R11195 avdd.n1409 avdd.n1408 0.0137576
R11196 avdd.n7917 avdd.n7916 0.0137576
R11197 avdd.n7879 avdd.n7878 0.0137576
R11198 avdd.n1608 avdd.n1607 0.0137576
R11199 avdd.n1539 avdd.n1538 0.0137576
R11200 avdd.n2086 avdd.n2085 0.0126061
R11201 avdd.n1919 avdd.n1899 0.0126061
R11202 avdd.n2090 avdd.n1880 0.0126061
R11203 avdd.n2063 avdd.n1959 0.0126061
R11204 avdd.n1982 avdd.n1973 0.0126061
R11205 avdd.n2032 avdd.n1996 0.0126061
R11206 avdd.n2024 avdd.n2023 0.0126061
R11207 avdd.n2208 avdd.n2133 0.0126061
R11208 avdd.n2173 avdd.n2153 0.0126061
R11209 avdd.n2198 avdd.n2197 0.0126061
R11210 avdd.n2235 avdd.n2234 0.0126061
R11211 avdd.n2244 avdd.n2116 0.0126061
R11212 avdd.n2278 avdd.n2277 0.0126061
R11213 avdd.n2297 avdd.n2098 0.0126061
R11214 avdd.n2423 avdd.n2348 0.0126061
R11215 avdd.n2388 avdd.n2368 0.0126061
R11216 avdd.n2413 avdd.n2412 0.0126061
R11217 avdd.n2450 avdd.n2449 0.0126061
R11218 avdd.n2459 avdd.n2331 0.0126061
R11219 avdd.n2493 avdd.n2492 0.0126061
R11220 avdd.n2512 avdd.n2313 0.0126061
R11221 avdd.n2638 avdd.n2563 0.0126061
R11222 avdd.n2603 avdd.n2583 0.0126061
R11223 avdd.n2628 avdd.n2627 0.0126061
R11224 avdd.n2665 avdd.n2664 0.0126061
R11225 avdd.n2674 avdd.n2546 0.0126061
R11226 avdd.n2708 avdd.n2707 0.0126061
R11227 avdd.n2727 avdd.n2528 0.0126061
R11228 avdd.n2853 avdd.n2778 0.0126061
R11229 avdd.n2818 avdd.n2798 0.0126061
R11230 avdd.n2843 avdd.n2842 0.0126061
R11231 avdd.n2880 avdd.n2879 0.0126061
R11232 avdd.n2889 avdd.n2761 0.0126061
R11233 avdd.n2923 avdd.n2922 0.0126061
R11234 avdd.n2942 avdd.n2743 0.0126061
R11235 avdd.n3068 avdd.n2993 0.0126061
R11236 avdd.n3033 avdd.n3013 0.0126061
R11237 avdd.n3058 avdd.n3057 0.0126061
R11238 avdd.n3095 avdd.n3094 0.0126061
R11239 avdd.n3104 avdd.n2976 0.0126061
R11240 avdd.n3138 avdd.n3137 0.0126061
R11241 avdd.n3157 avdd.n2958 0.0126061
R11242 avdd.n3375 avdd.n3374 0.0126061
R11243 avdd.n3209 avdd.n3189 0.0126061
R11244 avdd.n3380 avdd.n3171 0.0126061
R11245 avdd.n3352 avdd.n3249 0.0126061
R11246 avdd.n3272 avdd.n3263 0.0126061
R11247 avdd.n3300 avdd.n3286 0.0126061
R11248 avdd.n3318 avdd.n3317 0.0126061
R11249 avdd.n3590 avdd.n3589 0.0126061
R11250 avdd.n3424 avdd.n3404 0.0126061
R11251 avdd.n3595 avdd.n3386 0.0126061
R11252 avdd.n3567 avdd.n3464 0.0126061
R11253 avdd.n3487 avdd.n3478 0.0126061
R11254 avdd.n3515 avdd.n3501 0.0126061
R11255 avdd.n3533 avdd.n3532 0.0126061
R11256 avdd.n3805 avdd.n3804 0.0126061
R11257 avdd.n3639 avdd.n3619 0.0126061
R11258 avdd.n3810 avdd.n3601 0.0126061
R11259 avdd.n3782 avdd.n3679 0.0126061
R11260 avdd.n3702 avdd.n3693 0.0126061
R11261 avdd.n3730 avdd.n3716 0.0126061
R11262 avdd.n3748 avdd.n3747 0.0126061
R11263 avdd.n4020 avdd.n4019 0.0126061
R11264 avdd.n3854 avdd.n3834 0.0126061
R11265 avdd.n4025 avdd.n3816 0.0126061
R11266 avdd.n3997 avdd.n3894 0.0126061
R11267 avdd.n3917 avdd.n3908 0.0126061
R11268 avdd.n3945 avdd.n3931 0.0126061
R11269 avdd.n3963 avdd.n3962 0.0126061
R11270 avdd.n4235 avdd.n4234 0.0126061
R11271 avdd.n4069 avdd.n4049 0.0126061
R11272 avdd.n4240 avdd.n4031 0.0126061
R11273 avdd.n4212 avdd.n4109 0.0126061
R11274 avdd.n4132 avdd.n4123 0.0126061
R11275 avdd.n4160 avdd.n4146 0.0126061
R11276 avdd.n4178 avdd.n4177 0.0126061
R11277 avdd.n4450 avdd.n4449 0.0126061
R11278 avdd.n4284 avdd.n4264 0.0126061
R11279 avdd.n4455 avdd.n4246 0.0126061
R11280 avdd.n4427 avdd.n4324 0.0126061
R11281 avdd.n4347 avdd.n4338 0.0126061
R11282 avdd.n4375 avdd.n4361 0.0126061
R11283 avdd.n4393 avdd.n4392 0.0126061
R11284 avdd.n4930 avdd.n4855 0.0126061
R11285 avdd.n4895 avdd.n4875 0.0126061
R11286 avdd.n4920 avdd.n4919 0.0126061
R11287 avdd.n4957 avdd.n4956 0.0126061
R11288 avdd.n4966 avdd.n4838 0.0126061
R11289 avdd.n4997 avdd.n4996 0.0126061
R11290 avdd.n5016 avdd.n4820 0.0126061
R11291 avdd.n5146 avdd.n5071 0.0126061
R11292 avdd.n5111 avdd.n5091 0.0126061
R11293 avdd.n5136 avdd.n5135 0.0126061
R11294 avdd.n5173 avdd.n5172 0.0126061
R11295 avdd.n5182 avdd.n5054 0.0126061
R11296 avdd.n5213 avdd.n5212 0.0126061
R11297 avdd.n5232 avdd.n5036 0.0126061
R11298 avdd.n5362 avdd.n5287 0.0126061
R11299 avdd.n5327 avdd.n5307 0.0126061
R11300 avdd.n5352 avdd.n5351 0.0126061
R11301 avdd.n5389 avdd.n5388 0.0126061
R11302 avdd.n5398 avdd.n5270 0.0126061
R11303 avdd.n5429 avdd.n5428 0.0126061
R11304 avdd.n5448 avdd.n5252 0.0126061
R11305 avdd.n5578 avdd.n5503 0.0126061
R11306 avdd.n5543 avdd.n5523 0.0126061
R11307 avdd.n5568 avdd.n5567 0.0126061
R11308 avdd.n5605 avdd.n5604 0.0126061
R11309 avdd.n5614 avdd.n5486 0.0126061
R11310 avdd.n5645 avdd.n5644 0.0126061
R11311 avdd.n5664 avdd.n5468 0.0126061
R11312 avdd.n5794 avdd.n5719 0.0126061
R11313 avdd.n5759 avdd.n5739 0.0126061
R11314 avdd.n5784 avdd.n5783 0.0126061
R11315 avdd.n5821 avdd.n5820 0.0126061
R11316 avdd.n5830 avdd.n5702 0.0126061
R11317 avdd.n5861 avdd.n5860 0.0126061
R11318 avdd.n5880 avdd.n5684 0.0126061
R11319 avdd.n6010 avdd.n5935 0.0126061
R11320 avdd.n5975 avdd.n5955 0.0126061
R11321 avdd.n6000 avdd.n5999 0.0126061
R11322 avdd.n6037 avdd.n6036 0.0126061
R11323 avdd.n6046 avdd.n5918 0.0126061
R11324 avdd.n6077 avdd.n6076 0.0126061
R11325 avdd.n6096 avdd.n5900 0.0126061
R11326 avdd.n6226 avdd.n6151 0.0126061
R11327 avdd.n6191 avdd.n6171 0.0126061
R11328 avdd.n6216 avdd.n6215 0.0126061
R11329 avdd.n6253 avdd.n6252 0.0126061
R11330 avdd.n6262 avdd.n6134 0.0126061
R11331 avdd.n6293 avdd.n6292 0.0126061
R11332 avdd.n6312 avdd.n6116 0.0126061
R11333 avdd.n6442 avdd.n6367 0.0126061
R11334 avdd.n6407 avdd.n6387 0.0126061
R11335 avdd.n6432 avdd.n6431 0.0126061
R11336 avdd.n6469 avdd.n6468 0.0126061
R11337 avdd.n6478 avdd.n6350 0.0126061
R11338 avdd.n6509 avdd.n6508 0.0126061
R11339 avdd.n6528 avdd.n6332 0.0126061
R11340 avdd.n6658 avdd.n6583 0.0126061
R11341 avdd.n6623 avdd.n6603 0.0126061
R11342 avdd.n6648 avdd.n6647 0.0126061
R11343 avdd.n6685 avdd.n6684 0.0126061
R11344 avdd.n6694 avdd.n6566 0.0126061
R11345 avdd.n6725 avdd.n6724 0.0126061
R11346 avdd.n6744 avdd.n6548 0.0126061
R11347 avdd.n6874 avdd.n6799 0.0126061
R11348 avdd.n6839 avdd.n6819 0.0126061
R11349 avdd.n6864 avdd.n6863 0.0126061
R11350 avdd.n6901 avdd.n6900 0.0126061
R11351 avdd.n6910 avdd.n6782 0.0126061
R11352 avdd.n6941 avdd.n6940 0.0126061
R11353 avdd.n6960 avdd.n6764 0.0126061
R11354 avdd.n7090 avdd.n7015 0.0126061
R11355 avdd.n7055 avdd.n7035 0.0126061
R11356 avdd.n7080 avdd.n7079 0.0126061
R11357 avdd.n7117 avdd.n7116 0.0126061
R11358 avdd.n7126 avdd.n6998 0.0126061
R11359 avdd.n7157 avdd.n7156 0.0126061
R11360 avdd.n7176 avdd.n6980 0.0126061
R11361 avdd.n7306 avdd.n7231 0.0126061
R11362 avdd.n7271 avdd.n7251 0.0126061
R11363 avdd.n7296 avdd.n7295 0.0126061
R11364 avdd.n7333 avdd.n7332 0.0126061
R11365 avdd.n7342 avdd.n7214 0.0126061
R11366 avdd.n7373 avdd.n7372 0.0126061
R11367 avdd.n7392 avdd.n7196 0.0126061
R11368 avdd.n7651 avdd.n7650 0.0126061
R11369 avdd.n7716 avdd.n7704 0.0126061
R11370 avdd.n7738 avdd.n7737 0.0126061
R11371 avdd.n7663 avdd.n7662 0.0126061
R11372 avdd.n7805 avdd.n7797 0.0126061
R11373 avdd.n7828 avdd.n7827 0.0126061
R11374 avdd.n7790 avdd.n7783 0.0126061
R11375 avdd.n10128 avdd.n10127 0.0126061
R11376 avdd.n10195 avdd.n10183 0.0126061
R11377 avdd.n10217 avdd.n10216 0.0126061
R11378 avdd.n10142 avdd.n10141 0.0126061
R11379 avdd.n10063 avdd.n10056 0.0126061
R11380 avdd.n10086 avdd.n10085 0.0126061
R11381 avdd.n10050 avdd.n10043 0.0126061
R11382 avdd.n9964 avdd.n9928 0.0126061
R11383 avdd.n9999 avdd.n9994 0.0126061
R11384 avdd.n10023 avdd.n10022 0.0126061
R11385 avdd.n10279 avdd.n10272 0.0126061
R11386 avdd.n10295 avdd.n10286 0.0126061
R11387 avdd.n10318 avdd.n10317 0.0126061
R11388 avdd.n10266 avdd.n10259 0.0126061
R11389 avdd.n9850 avdd.n9814 0.0126061
R11390 avdd.n9885 avdd.n9880 0.0126061
R11391 avdd.n9909 avdd.n9908 0.0126061
R11392 avdd.n10381 avdd.n10374 0.0126061
R11393 avdd.n10397 avdd.n10388 0.0126061
R11394 avdd.n10420 avdd.n10419 0.0126061
R11395 avdd.n10368 avdd.n10361 0.0126061
R11396 avdd.n9736 avdd.n9700 0.0126061
R11397 avdd.n9771 avdd.n9766 0.0126061
R11398 avdd.n9795 avdd.n9794 0.0126061
R11399 avdd.n10483 avdd.n10476 0.0126061
R11400 avdd.n10499 avdd.n10490 0.0126061
R11401 avdd.n10522 avdd.n10521 0.0126061
R11402 avdd.n10470 avdd.n10463 0.0126061
R11403 avdd.n9623 avdd.n9586 0.0126061
R11404 avdd.n9658 avdd.n9653 0.0126061
R11405 avdd.n9682 avdd.n9681 0.0126061
R11406 avdd.n10585 avdd.n10578 0.0126061
R11407 avdd.n10601 avdd.n10592 0.0126061
R11408 avdd.n10624 avdd.n10623 0.0126061
R11409 avdd.n10572 avdd.n10565 0.0126061
R11410 avdd.n9508 avdd.n9472 0.0126061
R11411 avdd.n9543 avdd.n9538 0.0126061
R11412 avdd.n9567 avdd.n9566 0.0126061
R11413 avdd.n10687 avdd.n10680 0.0126061
R11414 avdd.n10703 avdd.n10694 0.0126061
R11415 avdd.n10726 avdd.n10725 0.0126061
R11416 avdd.n10674 avdd.n10667 0.0126061
R11417 avdd.n9394 avdd.n9358 0.0126061
R11418 avdd.n9429 avdd.n9424 0.0126061
R11419 avdd.n9453 avdd.n9452 0.0126061
R11420 avdd.n10789 avdd.n10782 0.0126061
R11421 avdd.n10805 avdd.n10796 0.0126061
R11422 avdd.n10828 avdd.n10827 0.0126061
R11423 avdd.n10776 avdd.n10769 0.0126061
R11424 avdd.n9280 avdd.n9244 0.0126061
R11425 avdd.n9315 avdd.n9310 0.0126061
R11426 avdd.n9339 avdd.n9338 0.0126061
R11427 avdd.n10891 avdd.n10884 0.0126061
R11428 avdd.n10907 avdd.n10898 0.0126061
R11429 avdd.n10930 avdd.n10929 0.0126061
R11430 avdd.n10878 avdd.n10871 0.0126061
R11431 avdd.n9166 avdd.n9130 0.0126061
R11432 avdd.n9201 avdd.n9196 0.0126061
R11433 avdd.n9225 avdd.n9224 0.0126061
R11434 avdd.n10993 avdd.n10986 0.0126061
R11435 avdd.n11009 avdd.n11000 0.0126061
R11436 avdd.n11032 avdd.n11031 0.0126061
R11437 avdd.n10980 avdd.n10973 0.0126061
R11438 avdd.n9052 avdd.n9016 0.0126061
R11439 avdd.n9087 avdd.n9082 0.0126061
R11440 avdd.n9111 avdd.n9110 0.0126061
R11441 avdd.n11095 avdd.n11088 0.0126061
R11442 avdd.n11111 avdd.n11102 0.0126061
R11443 avdd.n11134 avdd.n11133 0.0126061
R11444 avdd.n11082 avdd.n11075 0.0126061
R11445 avdd.n8938 avdd.n8902 0.0126061
R11446 avdd.n8973 avdd.n8968 0.0126061
R11447 avdd.n8997 avdd.n8996 0.0126061
R11448 avdd.n11197 avdd.n11190 0.0126061
R11449 avdd.n11213 avdd.n11204 0.0126061
R11450 avdd.n11236 avdd.n11235 0.0126061
R11451 avdd.n11184 avdd.n11177 0.0126061
R11452 avdd.n72 avdd.n71 0.0126061
R11453 avdd.n110 avdd.n98 0.0126061
R11454 avdd.n133 avdd.n132 0.0126061
R11455 avdd.n146 avdd.n145 0.0126061
R11456 avdd.n8826 avdd.n8819 0.0126061
R11457 avdd.n8849 avdd.n8848 0.0126061
R11458 avdd.n8813 avdd.n8806 0.0126061
R11459 avdd.n202 avdd.n201 0.0126061
R11460 avdd.n240 avdd.n228 0.0126061
R11461 avdd.n263 avdd.n262 0.0126061
R11462 avdd.n276 avdd.n275 0.0126061
R11463 avdd.n8740 avdd.n8733 0.0126061
R11464 avdd.n8763 avdd.n8762 0.0126061
R11465 avdd.n8727 avdd.n8720 0.0126061
R11466 avdd.n332 avdd.n331 0.0126061
R11467 avdd.n370 avdd.n358 0.0126061
R11468 avdd.n393 avdd.n392 0.0126061
R11469 avdd.n406 avdd.n405 0.0126061
R11470 avdd.n8654 avdd.n8647 0.0126061
R11471 avdd.n8677 avdd.n8676 0.0126061
R11472 avdd.n8641 avdd.n8634 0.0126061
R11473 avdd.n462 avdd.n461 0.0126061
R11474 avdd.n500 avdd.n488 0.0126061
R11475 avdd.n523 avdd.n522 0.0126061
R11476 avdd.n536 avdd.n535 0.0126061
R11477 avdd.n8568 avdd.n8561 0.0126061
R11478 avdd.n8591 avdd.n8590 0.0126061
R11479 avdd.n8555 avdd.n8548 0.0126061
R11480 avdd.n592 avdd.n591 0.0126061
R11481 avdd.n630 avdd.n618 0.0126061
R11482 avdd.n653 avdd.n652 0.0126061
R11483 avdd.n666 avdd.n665 0.0126061
R11484 avdd.n8482 avdd.n8475 0.0126061
R11485 avdd.n8505 avdd.n8504 0.0126061
R11486 avdd.n8469 avdd.n8462 0.0126061
R11487 avdd.n722 avdd.n721 0.0126061
R11488 avdd.n760 avdd.n748 0.0126061
R11489 avdd.n783 avdd.n782 0.0126061
R11490 avdd.n796 avdd.n795 0.0126061
R11491 avdd.n8396 avdd.n8389 0.0126061
R11492 avdd.n8419 avdd.n8418 0.0126061
R11493 avdd.n8383 avdd.n8376 0.0126061
R11494 avdd.n852 avdd.n851 0.0126061
R11495 avdd.n890 avdd.n878 0.0126061
R11496 avdd.n913 avdd.n912 0.0126061
R11497 avdd.n926 avdd.n925 0.0126061
R11498 avdd.n8310 avdd.n8303 0.0126061
R11499 avdd.n8333 avdd.n8332 0.0126061
R11500 avdd.n8297 avdd.n8290 0.0126061
R11501 avdd.n982 avdd.n981 0.0126061
R11502 avdd.n1020 avdd.n1008 0.0126061
R11503 avdd.n1043 avdd.n1042 0.0126061
R11504 avdd.n1056 avdd.n1055 0.0126061
R11505 avdd.n8224 avdd.n8217 0.0126061
R11506 avdd.n8247 avdd.n8246 0.0126061
R11507 avdd.n8211 avdd.n8204 0.0126061
R11508 avdd.n1112 avdd.n1111 0.0126061
R11509 avdd.n1150 avdd.n1138 0.0126061
R11510 avdd.n1173 avdd.n1172 0.0126061
R11511 avdd.n1186 avdd.n1185 0.0126061
R11512 avdd.n8138 avdd.n8131 0.0126061
R11513 avdd.n8161 avdd.n8160 0.0126061
R11514 avdd.n8125 avdd.n8118 0.0126061
R11515 avdd.n1242 avdd.n1241 0.0126061
R11516 avdd.n1280 avdd.n1268 0.0126061
R11517 avdd.n1303 avdd.n1302 0.0126061
R11518 avdd.n1316 avdd.n1315 0.0126061
R11519 avdd.n8052 avdd.n8045 0.0126061
R11520 avdd.n8075 avdd.n8074 0.0126061
R11521 avdd.n8039 avdd.n8032 0.0126061
R11522 avdd.n1372 avdd.n1371 0.0126061
R11523 avdd.n1410 avdd.n1398 0.0126061
R11524 avdd.n1433 avdd.n1432 0.0126061
R11525 avdd.n1446 avdd.n1445 0.0126061
R11526 avdd.n7966 avdd.n7959 0.0126061
R11527 avdd.n7989 avdd.n7988 0.0126061
R11528 avdd.n7953 avdd.n7946 0.0126061
R11529 avdd.n1502 avdd.n1501 0.0126061
R11530 avdd.n1540 avdd.n1528 0.0126061
R11531 avdd.n1563 avdd.n1562 0.0126061
R11532 avdd.n1576 avdd.n1575 0.0126061
R11533 avdd.n7880 avdd.n7873 0.0126061
R11534 avdd.n7903 avdd.n7902 0.0126061
R11535 avdd.n7867 avdd.n7860 0.0126061
R11536 avdd.n1965 avdd.n1964 0.0126061
R11537 avdd.n2128 avdd.n2124 0.0126061
R11538 avdd.n2343 avdd.n2339 0.0126061
R11539 avdd.n2558 avdd.n2554 0.0126061
R11540 avdd.n2773 avdd.n2769 0.0126061
R11541 avdd.n2988 avdd.n2984 0.0126061
R11542 avdd.n3255 avdd.n3254 0.0126061
R11543 avdd.n3470 avdd.n3469 0.0126061
R11544 avdd.n3685 avdd.n3684 0.0126061
R11545 avdd.n3900 avdd.n3899 0.0126061
R11546 avdd.n4115 avdd.n4114 0.0126061
R11547 avdd.n4330 avdd.n4329 0.0126061
R11548 avdd.n4850 avdd.n4846 0.0126061
R11549 avdd.n5066 avdd.n5062 0.0126061
R11550 avdd.n5282 avdd.n5278 0.0126061
R11551 avdd.n5498 avdd.n5494 0.0126061
R11552 avdd.n5714 avdd.n5710 0.0126061
R11553 avdd.n5930 avdd.n5926 0.0126061
R11554 avdd.n6146 avdd.n6142 0.0126061
R11555 avdd.n6362 avdd.n6358 0.0126061
R11556 avdd.n6578 avdd.n6574 0.0126061
R11557 avdd.n6794 avdd.n6790 0.0126061
R11558 avdd.n7010 avdd.n7006 0.0126061
R11559 avdd.n7226 avdd.n7222 0.0126061
R11560 avdd.n7677 avdd.n7668 0.0126061
R11561 avdd.n10156 avdd.n10147 0.0126061
R11562 avdd.n9940 avdd.n9932 0.0126061
R11563 avdd.n9826 avdd.n9818 0.0126061
R11564 avdd.n9712 avdd.n9704 0.0126061
R11565 avdd.n9599 avdd.n9591 0.0126061
R11566 avdd.n9484 avdd.n9476 0.0126061
R11567 avdd.n9370 avdd.n9362 0.0126061
R11568 avdd.n9256 avdd.n9248 0.0126061
R11569 avdd.n9142 avdd.n9134 0.0126061
R11570 avdd.n9028 avdd.n9020 0.0126061
R11571 avdd.n8914 avdd.n8906 0.0126061
R11572 avdd.n160 avdd.n151 0.0126061
R11573 avdd.n290 avdd.n281 0.0126061
R11574 avdd.n420 avdd.n411 0.0126061
R11575 avdd.n550 avdd.n541 0.0126061
R11576 avdd.n680 avdd.n671 0.0126061
R11577 avdd.n810 avdd.n801 0.0126061
R11578 avdd.n940 avdd.n931 0.0126061
R11579 avdd.n1070 avdd.n1061 0.0126061
R11580 avdd.n1200 avdd.n1191 0.0126061
R11581 avdd.n1330 avdd.n1321 0.0126061
R11582 avdd.n1460 avdd.n1451 0.0126061
R11583 avdd.n1590 avdd.n1581 0.0126061
R11584 avdd.n2018 avdd.n2012 0.0118636
R11585 avdd.n1999 avdd.n1998 0.0118636
R11586 avdd.n1967 avdd.n1966 0.0118636
R11587 avdd.n2077 avdd.n1887 0.0118636
R11588 avdd.n1938 avdd.n1890 0.0118636
R11589 avdd.n2292 avdd.n2101 0.0118636
R11590 avdd.n2266 avdd.n2263 0.0118636
R11591 avdd.n2224 avdd.n2126 0.0118636
R11592 avdd.n2219 avdd.n2130 0.0118636
R11593 avdd.n2190 avdd.n2187 0.0118636
R11594 avdd.n2507 avdd.n2316 0.0118636
R11595 avdd.n2481 avdd.n2478 0.0118636
R11596 avdd.n2439 avdd.n2341 0.0118636
R11597 avdd.n2434 avdd.n2345 0.0118636
R11598 avdd.n2405 avdd.n2402 0.0118636
R11599 avdd.n2722 avdd.n2531 0.0118636
R11600 avdd.n2696 avdd.n2693 0.0118636
R11601 avdd.n2654 avdd.n2556 0.0118636
R11602 avdd.n2649 avdd.n2560 0.0118636
R11603 avdd.n2620 avdd.n2617 0.0118636
R11604 avdd.n2937 avdd.n2746 0.0118636
R11605 avdd.n2911 avdd.n2908 0.0118636
R11606 avdd.n2869 avdd.n2771 0.0118636
R11607 avdd.n2864 avdd.n2775 0.0118636
R11608 avdd.n2835 avdd.n2832 0.0118636
R11609 avdd.n3152 avdd.n2961 0.0118636
R11610 avdd.n3126 avdd.n3123 0.0118636
R11611 avdd.n3084 avdd.n2986 0.0118636
R11612 avdd.n3079 avdd.n2990 0.0118636
R11613 avdd.n3050 avdd.n3047 0.0118636
R11614 avdd.n3311 avdd.n3310 0.0118636
R11615 avdd.n3289 avdd.n3288 0.0118636
R11616 avdd.n3257 avdd.n3256 0.0118636
R11617 avdd.n3366 avdd.n3177 0.0118636
R11618 avdd.n3228 avdd.n3180 0.0118636
R11619 avdd.n3526 avdd.n3525 0.0118636
R11620 avdd.n3504 avdd.n3503 0.0118636
R11621 avdd.n3472 avdd.n3471 0.0118636
R11622 avdd.n3581 avdd.n3392 0.0118636
R11623 avdd.n3443 avdd.n3395 0.0118636
R11624 avdd.n3741 avdd.n3740 0.0118636
R11625 avdd.n3719 avdd.n3718 0.0118636
R11626 avdd.n3687 avdd.n3686 0.0118636
R11627 avdd.n3796 avdd.n3607 0.0118636
R11628 avdd.n3658 avdd.n3610 0.0118636
R11629 avdd.n3956 avdd.n3955 0.0118636
R11630 avdd.n3934 avdd.n3933 0.0118636
R11631 avdd.n3902 avdd.n3901 0.0118636
R11632 avdd.n4011 avdd.n3822 0.0118636
R11633 avdd.n3873 avdd.n3825 0.0118636
R11634 avdd.n4171 avdd.n4170 0.0118636
R11635 avdd.n4149 avdd.n4148 0.0118636
R11636 avdd.n4117 avdd.n4116 0.0118636
R11637 avdd.n4226 avdd.n4037 0.0118636
R11638 avdd.n4088 avdd.n4040 0.0118636
R11639 avdd.n4386 avdd.n4385 0.0118636
R11640 avdd.n4364 avdd.n4363 0.0118636
R11641 avdd.n4332 avdd.n4331 0.0118636
R11642 avdd.n4441 avdd.n4252 0.0118636
R11643 avdd.n4303 avdd.n4255 0.0118636
R11644 avdd.n4913 avdd.n4910 0.0118636
R11645 avdd.n4941 avdd.n4852 0.0118636
R11646 avdd.n4946 avdd.n4848 0.0118636
R11647 avdd.n4988 avdd.n4985 0.0118636
R11648 avdd.n5009 avdd.n4822 0.0118636
R11649 avdd.n5129 avdd.n5126 0.0118636
R11650 avdd.n5157 avdd.n5068 0.0118636
R11651 avdd.n5162 avdd.n5064 0.0118636
R11652 avdd.n5204 avdd.n5201 0.0118636
R11653 avdd.n5225 avdd.n5038 0.0118636
R11654 avdd.n5345 avdd.n5342 0.0118636
R11655 avdd.n5373 avdd.n5284 0.0118636
R11656 avdd.n5378 avdd.n5280 0.0118636
R11657 avdd.n5420 avdd.n5417 0.0118636
R11658 avdd.n5441 avdd.n5254 0.0118636
R11659 avdd.n5561 avdd.n5558 0.0118636
R11660 avdd.n5589 avdd.n5500 0.0118636
R11661 avdd.n5594 avdd.n5496 0.0118636
R11662 avdd.n5636 avdd.n5633 0.0118636
R11663 avdd.n5657 avdd.n5470 0.0118636
R11664 avdd.n5777 avdd.n5774 0.0118636
R11665 avdd.n5805 avdd.n5716 0.0118636
R11666 avdd.n5810 avdd.n5712 0.0118636
R11667 avdd.n5852 avdd.n5849 0.0118636
R11668 avdd.n5873 avdd.n5686 0.0118636
R11669 avdd.n5993 avdd.n5990 0.0118636
R11670 avdd.n6021 avdd.n5932 0.0118636
R11671 avdd.n6026 avdd.n5928 0.0118636
R11672 avdd.n6068 avdd.n6065 0.0118636
R11673 avdd.n6089 avdd.n5902 0.0118636
R11674 avdd.n6209 avdd.n6206 0.0118636
R11675 avdd.n6237 avdd.n6148 0.0118636
R11676 avdd.n6242 avdd.n6144 0.0118636
R11677 avdd.n6284 avdd.n6281 0.0118636
R11678 avdd.n6305 avdd.n6118 0.0118636
R11679 avdd.n6425 avdd.n6422 0.0118636
R11680 avdd.n6453 avdd.n6364 0.0118636
R11681 avdd.n6458 avdd.n6360 0.0118636
R11682 avdd.n6500 avdd.n6497 0.0118636
R11683 avdd.n6521 avdd.n6334 0.0118636
R11684 avdd.n6641 avdd.n6638 0.0118636
R11685 avdd.n6669 avdd.n6580 0.0118636
R11686 avdd.n6674 avdd.n6576 0.0118636
R11687 avdd.n6716 avdd.n6713 0.0118636
R11688 avdd.n6737 avdd.n6550 0.0118636
R11689 avdd.n6857 avdd.n6854 0.0118636
R11690 avdd.n6885 avdd.n6796 0.0118636
R11691 avdd.n6890 avdd.n6792 0.0118636
R11692 avdd.n6932 avdd.n6929 0.0118636
R11693 avdd.n6953 avdd.n6766 0.0118636
R11694 avdd.n7073 avdd.n7070 0.0118636
R11695 avdd.n7101 avdd.n7012 0.0118636
R11696 avdd.n7106 avdd.n7008 0.0118636
R11697 avdd.n7148 avdd.n7145 0.0118636
R11698 avdd.n7169 avdd.n6982 0.0118636
R11699 avdd.n7289 avdd.n7286 0.0118636
R11700 avdd.n7317 avdd.n7228 0.0118636
R11701 avdd.n7322 avdd.n7224 0.0118636
R11702 avdd.n7364 avdd.n7361 0.0118636
R11703 avdd.n7385 avdd.n7198 0.0118636
R11704 avdd.n7734 avdd.n7728 0.0118636
R11705 avdd.n7694 avdd.n7693 0.0118636
R11706 avdd.n7675 avdd.n7674 0.0118636
R11707 avdd.n7824 avdd.n7818 0.0118636
R11708 avdd.n7841 avdd.n7840 0.0118636
R11709 avdd.n10213 avdd.n10207 0.0118636
R11710 avdd.n10173 avdd.n10172 0.0118636
R11711 avdd.n10154 avdd.n10153 0.0118636
R11712 avdd.n10082 avdd.n10076 0.0118636
R11713 avdd.n10099 avdd.n10098 0.0118636
R11714 avdd.n10019 avdd.n10013 0.0118636
R11715 avdd.n9957 avdd.n9956 0.0118636
R11716 avdd.n9938 avdd.n9937 0.0118636
R11717 avdd.n10314 avdd.n10308 0.0118636
R11718 avdd.n10331 avdd.n10330 0.0118636
R11719 avdd.n9905 avdd.n9899 0.0118636
R11720 avdd.n9843 avdd.n9842 0.0118636
R11721 avdd.n9824 avdd.n9823 0.0118636
R11722 avdd.n10416 avdd.n10410 0.0118636
R11723 avdd.n10433 avdd.n10432 0.0118636
R11724 avdd.n9791 avdd.n9785 0.0118636
R11725 avdd.n9729 avdd.n9728 0.0118636
R11726 avdd.n9710 avdd.n9709 0.0118636
R11727 avdd.n10518 avdd.n10512 0.0118636
R11728 avdd.n10535 avdd.n10534 0.0118636
R11729 avdd.n9678 avdd.n9672 0.0118636
R11730 avdd.n9616 avdd.n9615 0.0118636
R11731 avdd.n9597 avdd.n9596 0.0118636
R11732 avdd.n10620 avdd.n10614 0.0118636
R11733 avdd.n10637 avdd.n10636 0.0118636
R11734 avdd.n9563 avdd.n9557 0.0118636
R11735 avdd.n9501 avdd.n9500 0.0118636
R11736 avdd.n9482 avdd.n9481 0.0118636
R11737 avdd.n10722 avdd.n10716 0.0118636
R11738 avdd.n10739 avdd.n10738 0.0118636
R11739 avdd.n9449 avdd.n9443 0.0118636
R11740 avdd.n9387 avdd.n9386 0.0118636
R11741 avdd.n9368 avdd.n9367 0.0118636
R11742 avdd.n10824 avdd.n10818 0.0118636
R11743 avdd.n10841 avdd.n10840 0.0118636
R11744 avdd.n9335 avdd.n9329 0.0118636
R11745 avdd.n9273 avdd.n9272 0.0118636
R11746 avdd.n9254 avdd.n9253 0.0118636
R11747 avdd.n10926 avdd.n10920 0.0118636
R11748 avdd.n10943 avdd.n10942 0.0118636
R11749 avdd.n9221 avdd.n9215 0.0118636
R11750 avdd.n9159 avdd.n9158 0.0118636
R11751 avdd.n9140 avdd.n9139 0.0118636
R11752 avdd.n11028 avdd.n11022 0.0118636
R11753 avdd.n11045 avdd.n11044 0.0118636
R11754 avdd.n9107 avdd.n9101 0.0118636
R11755 avdd.n9045 avdd.n9044 0.0118636
R11756 avdd.n9026 avdd.n9025 0.0118636
R11757 avdd.n11130 avdd.n11124 0.0118636
R11758 avdd.n11147 avdd.n11146 0.0118636
R11759 avdd.n8993 avdd.n8987 0.0118636
R11760 avdd.n8931 avdd.n8930 0.0118636
R11761 avdd.n8912 avdd.n8911 0.0118636
R11762 avdd.n11232 avdd.n11226 0.0118636
R11763 avdd.n11249 avdd.n11248 0.0118636
R11764 avdd.n8862 avdd.n8861 0.0118636
R11765 avdd.n8845 avdd.n8839 0.0118636
R11766 avdd.n158 avdd.n157 0.0118636
R11767 avdd.n177 avdd.n176 0.0118636
R11768 avdd.n129 avdd.n123 0.0118636
R11769 avdd.n8776 avdd.n8775 0.0118636
R11770 avdd.n8759 avdd.n8753 0.0118636
R11771 avdd.n288 avdd.n287 0.0118636
R11772 avdd.n307 avdd.n306 0.0118636
R11773 avdd.n259 avdd.n253 0.0118636
R11774 avdd.n8690 avdd.n8689 0.0118636
R11775 avdd.n8673 avdd.n8667 0.0118636
R11776 avdd.n418 avdd.n417 0.0118636
R11777 avdd.n437 avdd.n436 0.0118636
R11778 avdd.n389 avdd.n383 0.0118636
R11779 avdd.n8604 avdd.n8603 0.0118636
R11780 avdd.n8587 avdd.n8581 0.0118636
R11781 avdd.n548 avdd.n547 0.0118636
R11782 avdd.n567 avdd.n566 0.0118636
R11783 avdd.n519 avdd.n513 0.0118636
R11784 avdd.n8518 avdd.n8517 0.0118636
R11785 avdd.n8501 avdd.n8495 0.0118636
R11786 avdd.n678 avdd.n677 0.0118636
R11787 avdd.n697 avdd.n696 0.0118636
R11788 avdd.n649 avdd.n643 0.0118636
R11789 avdd.n8432 avdd.n8431 0.0118636
R11790 avdd.n8415 avdd.n8409 0.0118636
R11791 avdd.n808 avdd.n807 0.0118636
R11792 avdd.n827 avdd.n826 0.0118636
R11793 avdd.n779 avdd.n773 0.0118636
R11794 avdd.n8346 avdd.n8345 0.0118636
R11795 avdd.n8329 avdd.n8323 0.0118636
R11796 avdd.n938 avdd.n937 0.0118636
R11797 avdd.n957 avdd.n956 0.0118636
R11798 avdd.n909 avdd.n903 0.0118636
R11799 avdd.n8260 avdd.n8259 0.0118636
R11800 avdd.n8243 avdd.n8237 0.0118636
R11801 avdd.n1068 avdd.n1067 0.0118636
R11802 avdd.n1087 avdd.n1086 0.0118636
R11803 avdd.n1039 avdd.n1033 0.0118636
R11804 avdd.n8174 avdd.n8173 0.0118636
R11805 avdd.n8157 avdd.n8151 0.0118636
R11806 avdd.n1198 avdd.n1197 0.0118636
R11807 avdd.n1217 avdd.n1216 0.0118636
R11808 avdd.n1169 avdd.n1163 0.0118636
R11809 avdd.n8088 avdd.n8087 0.0118636
R11810 avdd.n8071 avdd.n8065 0.0118636
R11811 avdd.n1328 avdd.n1327 0.0118636
R11812 avdd.n1347 avdd.n1346 0.0118636
R11813 avdd.n1299 avdd.n1293 0.0118636
R11814 avdd.n8002 avdd.n8001 0.0118636
R11815 avdd.n7985 avdd.n7979 0.0118636
R11816 avdd.n1458 avdd.n1457 0.0118636
R11817 avdd.n1477 avdd.n1476 0.0118636
R11818 avdd.n1429 avdd.n1423 0.0118636
R11819 avdd.n7916 avdd.n7915 0.0118636
R11820 avdd.n7899 avdd.n7893 0.0118636
R11821 avdd.n1588 avdd.n1587 0.0118636
R11822 avdd.n1607 avdd.n1606 0.0118636
R11823 avdd.n1559 avdd.n1553 0.0118636
R11824 avdd.n2087 avdd.n2086 0.0111818
R11825 avdd.n1907 avdd.n1903 0.0111818
R11826 avdd.n1941 avdd.n1940 0.0111818
R11827 avdd.n2088 avdd.n1882 0.0111818
R11828 avdd.n2060 avdd.n1961 0.0111818
R11829 avdd.n2044 avdd.n1995 0.0111818
R11830 avdd.n2142 avdd.n2133 0.0111818
R11831 avdd.n2161 avdd.n2157 0.0111818
R11832 avdd.n2188 avdd.n2138 0.0111818
R11833 avdd.n2141 avdd.n2140 0.0111818
R11834 avdd.n2240 avdd.n2119 0.0111818
R11835 avdd.n2264 avdd.n2105 0.0111818
R11836 avdd.n2357 avdd.n2348 0.0111818
R11837 avdd.n2376 avdd.n2372 0.0111818
R11838 avdd.n2403 avdd.n2353 0.0111818
R11839 avdd.n2356 avdd.n2355 0.0111818
R11840 avdd.n2455 avdd.n2334 0.0111818
R11841 avdd.n2479 avdd.n2320 0.0111818
R11842 avdd.n2572 avdd.n2563 0.0111818
R11843 avdd.n2591 avdd.n2587 0.0111818
R11844 avdd.n2618 avdd.n2568 0.0111818
R11845 avdd.n2571 avdd.n2570 0.0111818
R11846 avdd.n2670 avdd.n2549 0.0111818
R11847 avdd.n2694 avdd.n2535 0.0111818
R11848 avdd.n2787 avdd.n2778 0.0111818
R11849 avdd.n2806 avdd.n2802 0.0111818
R11850 avdd.n2833 avdd.n2783 0.0111818
R11851 avdd.n2786 avdd.n2785 0.0111818
R11852 avdd.n2885 avdd.n2764 0.0111818
R11853 avdd.n2909 avdd.n2750 0.0111818
R11854 avdd.n3002 avdd.n2993 0.0111818
R11855 avdd.n3021 avdd.n3017 0.0111818
R11856 avdd.n3048 avdd.n2998 0.0111818
R11857 avdd.n3001 avdd.n3000 0.0111818
R11858 avdd.n3100 avdd.n2979 0.0111818
R11859 avdd.n3124 avdd.n2965 0.0111818
R11860 avdd.n3376 avdd.n3375 0.0111818
R11861 avdd.n3197 avdd.n3193 0.0111818
R11862 avdd.n3231 avdd.n3230 0.0111818
R11863 avdd.n3377 avdd.n3172 0.0111818
R11864 avdd.n3349 avdd.n3251 0.0111818
R11865 avdd.n3333 avdd.n3285 0.0111818
R11866 avdd.n3591 avdd.n3590 0.0111818
R11867 avdd.n3412 avdd.n3408 0.0111818
R11868 avdd.n3446 avdd.n3445 0.0111818
R11869 avdd.n3592 avdd.n3387 0.0111818
R11870 avdd.n3564 avdd.n3466 0.0111818
R11871 avdd.n3548 avdd.n3500 0.0111818
R11872 avdd.n3806 avdd.n3805 0.0111818
R11873 avdd.n3627 avdd.n3623 0.0111818
R11874 avdd.n3661 avdd.n3660 0.0111818
R11875 avdd.n3807 avdd.n3602 0.0111818
R11876 avdd.n3779 avdd.n3681 0.0111818
R11877 avdd.n3763 avdd.n3715 0.0111818
R11878 avdd.n4021 avdd.n4020 0.0111818
R11879 avdd.n3842 avdd.n3838 0.0111818
R11880 avdd.n3876 avdd.n3875 0.0111818
R11881 avdd.n4022 avdd.n3817 0.0111818
R11882 avdd.n3994 avdd.n3896 0.0111818
R11883 avdd.n3978 avdd.n3930 0.0111818
R11884 avdd.n4236 avdd.n4235 0.0111818
R11885 avdd.n4057 avdd.n4053 0.0111818
R11886 avdd.n4091 avdd.n4090 0.0111818
R11887 avdd.n4237 avdd.n4032 0.0111818
R11888 avdd.n4209 avdd.n4111 0.0111818
R11889 avdd.n4193 avdd.n4145 0.0111818
R11890 avdd.n4451 avdd.n4450 0.0111818
R11891 avdd.n4272 avdd.n4268 0.0111818
R11892 avdd.n4306 avdd.n4305 0.0111818
R11893 avdd.n4452 avdd.n4247 0.0111818
R11894 avdd.n4424 avdd.n4326 0.0111818
R11895 avdd.n4408 avdd.n4360 0.0111818
R11896 avdd.n4865 avdd.n4855 0.0111818
R11897 avdd.n4883 avdd.n4879 0.0111818
R11898 avdd.n4911 avdd.n4860 0.0111818
R11899 avdd.n4864 avdd.n4863 0.0111818
R11900 avdd.n4962 avdd.n4841 0.0111818
R11901 avdd.n4986 avdd.n4826 0.0111818
R11902 avdd.n4816 avdd.n4812 0.0111818
R11903 avdd.n5081 avdd.n5071 0.0111818
R11904 avdd.n5099 avdd.n5095 0.0111818
R11905 avdd.n5127 avdd.n5076 0.0111818
R11906 avdd.n5080 avdd.n5079 0.0111818
R11907 avdd.n5178 avdd.n5057 0.0111818
R11908 avdd.n5202 avdd.n5042 0.0111818
R11909 avdd.n5032 avdd.n5028 0.0111818
R11910 avdd.n5297 avdd.n5287 0.0111818
R11911 avdd.n5315 avdd.n5311 0.0111818
R11912 avdd.n5343 avdd.n5292 0.0111818
R11913 avdd.n5296 avdd.n5295 0.0111818
R11914 avdd.n5394 avdd.n5273 0.0111818
R11915 avdd.n5418 avdd.n5258 0.0111818
R11916 avdd.n5248 avdd.n5244 0.0111818
R11917 avdd.n5513 avdd.n5503 0.0111818
R11918 avdd.n5531 avdd.n5527 0.0111818
R11919 avdd.n5559 avdd.n5508 0.0111818
R11920 avdd.n5512 avdd.n5511 0.0111818
R11921 avdd.n5610 avdd.n5489 0.0111818
R11922 avdd.n5634 avdd.n5474 0.0111818
R11923 avdd.n5464 avdd.n5460 0.0111818
R11924 avdd.n5729 avdd.n5719 0.0111818
R11925 avdd.n5747 avdd.n5743 0.0111818
R11926 avdd.n5775 avdd.n5724 0.0111818
R11927 avdd.n5728 avdd.n5727 0.0111818
R11928 avdd.n5826 avdd.n5705 0.0111818
R11929 avdd.n5850 avdd.n5690 0.0111818
R11930 avdd.n5680 avdd.n5676 0.0111818
R11931 avdd.n5945 avdd.n5935 0.0111818
R11932 avdd.n5963 avdd.n5959 0.0111818
R11933 avdd.n5991 avdd.n5940 0.0111818
R11934 avdd.n5944 avdd.n5943 0.0111818
R11935 avdd.n6042 avdd.n5921 0.0111818
R11936 avdd.n6066 avdd.n5906 0.0111818
R11937 avdd.n5896 avdd.n5892 0.0111818
R11938 avdd.n6161 avdd.n6151 0.0111818
R11939 avdd.n6179 avdd.n6175 0.0111818
R11940 avdd.n6207 avdd.n6156 0.0111818
R11941 avdd.n6160 avdd.n6159 0.0111818
R11942 avdd.n6258 avdd.n6137 0.0111818
R11943 avdd.n6282 avdd.n6122 0.0111818
R11944 avdd.n6112 avdd.n6108 0.0111818
R11945 avdd.n6377 avdd.n6367 0.0111818
R11946 avdd.n6395 avdd.n6391 0.0111818
R11947 avdd.n6423 avdd.n6372 0.0111818
R11948 avdd.n6376 avdd.n6375 0.0111818
R11949 avdd.n6474 avdd.n6353 0.0111818
R11950 avdd.n6498 avdd.n6338 0.0111818
R11951 avdd.n6328 avdd.n6324 0.0111818
R11952 avdd.n6593 avdd.n6583 0.0111818
R11953 avdd.n6611 avdd.n6607 0.0111818
R11954 avdd.n6639 avdd.n6588 0.0111818
R11955 avdd.n6592 avdd.n6591 0.0111818
R11956 avdd.n6690 avdd.n6569 0.0111818
R11957 avdd.n6714 avdd.n6554 0.0111818
R11958 avdd.n6544 avdd.n6540 0.0111818
R11959 avdd.n6809 avdd.n6799 0.0111818
R11960 avdd.n6827 avdd.n6823 0.0111818
R11961 avdd.n6855 avdd.n6804 0.0111818
R11962 avdd.n6808 avdd.n6807 0.0111818
R11963 avdd.n6906 avdd.n6785 0.0111818
R11964 avdd.n6930 avdd.n6770 0.0111818
R11965 avdd.n6760 avdd.n6756 0.0111818
R11966 avdd.n7025 avdd.n7015 0.0111818
R11967 avdd.n7043 avdd.n7039 0.0111818
R11968 avdd.n7071 avdd.n7020 0.0111818
R11969 avdd.n7024 avdd.n7023 0.0111818
R11970 avdd.n7122 avdd.n7001 0.0111818
R11971 avdd.n7146 avdd.n6986 0.0111818
R11972 avdd.n6976 avdd.n6972 0.0111818
R11973 avdd.n7241 avdd.n7231 0.0111818
R11974 avdd.n7259 avdd.n7255 0.0111818
R11975 avdd.n7287 avdd.n7236 0.0111818
R11976 avdd.n7240 avdd.n7239 0.0111818
R11977 avdd.n7338 avdd.n7217 0.0111818
R11978 avdd.n7362 avdd.n7202 0.0111818
R11979 avdd.n7192 avdd.n7188 0.0111818
R11980 avdd.n7652 avdd.n7651 0.0111818
R11981 avdd.n7744 avdd.n7743 0.0111818
R11982 avdd.n7736 avdd.n7735 0.0111818
R11983 avdd.n7701 avdd.n7700 0.0111818
R11984 avdd.n7655 avdd.n7654 0.0111818
R11985 avdd.n7826 avdd.n7825 0.0111818
R11986 avdd.n10129 avdd.n10128 0.0111818
R11987 avdd.n10223 avdd.n10222 0.0111818
R11988 avdd.n10215 avdd.n10214 0.0111818
R11989 avdd.n10180 avdd.n10179 0.0111818
R11990 avdd.n10133 avdd.n10132 0.0111818
R11991 avdd.n10084 avdd.n10083 0.0111818
R11992 avdd.n9965 avdd.n9964 0.0111818
R11993 avdd.n9970 avdd.n9969 0.0111818
R11994 avdd.n10021 avdd.n10020 0.0111818
R11995 avdd.n10281 avdd.n10280 0.0111818
R11996 avdd.n10316 avdd.n10315 0.0111818
R11997 avdd.n10322 avdd.n10321 0.0111818
R11998 avdd.n9851 avdd.n9850 0.0111818
R11999 avdd.n9856 avdd.n9855 0.0111818
R12000 avdd.n9907 avdd.n9906 0.0111818
R12001 avdd.n10383 avdd.n10382 0.0111818
R12002 avdd.n10418 avdd.n10417 0.0111818
R12003 avdd.n10424 avdd.n10423 0.0111818
R12004 avdd.n9737 avdd.n9736 0.0111818
R12005 avdd.n9742 avdd.n9741 0.0111818
R12006 avdd.n9793 avdd.n9792 0.0111818
R12007 avdd.n10485 avdd.n10484 0.0111818
R12008 avdd.n10520 avdd.n10519 0.0111818
R12009 avdd.n10526 avdd.n10525 0.0111818
R12010 avdd.n9624 avdd.n9623 0.0111818
R12011 avdd.n9629 avdd.n9628 0.0111818
R12012 avdd.n9680 avdd.n9679 0.0111818
R12013 avdd.n9622 avdd.n9587 0.0111818
R12014 avdd.n10587 avdd.n10586 0.0111818
R12015 avdd.n10622 avdd.n10621 0.0111818
R12016 avdd.n10628 avdd.n10627 0.0111818
R12017 avdd.n9509 avdd.n9508 0.0111818
R12018 avdd.n9514 avdd.n9513 0.0111818
R12019 avdd.n9565 avdd.n9564 0.0111818
R12020 avdd.n10689 avdd.n10688 0.0111818
R12021 avdd.n10724 avdd.n10723 0.0111818
R12022 avdd.n10730 avdd.n10729 0.0111818
R12023 avdd.n9395 avdd.n9394 0.0111818
R12024 avdd.n9400 avdd.n9399 0.0111818
R12025 avdd.n9451 avdd.n9450 0.0111818
R12026 avdd.n10791 avdd.n10790 0.0111818
R12027 avdd.n10826 avdd.n10825 0.0111818
R12028 avdd.n10832 avdd.n10831 0.0111818
R12029 avdd.n9281 avdd.n9280 0.0111818
R12030 avdd.n9286 avdd.n9285 0.0111818
R12031 avdd.n9337 avdd.n9336 0.0111818
R12032 avdd.n10893 avdd.n10892 0.0111818
R12033 avdd.n10928 avdd.n10927 0.0111818
R12034 avdd.n10934 avdd.n10933 0.0111818
R12035 avdd.n9167 avdd.n9166 0.0111818
R12036 avdd.n9172 avdd.n9171 0.0111818
R12037 avdd.n9223 avdd.n9222 0.0111818
R12038 avdd.n10995 avdd.n10994 0.0111818
R12039 avdd.n11030 avdd.n11029 0.0111818
R12040 avdd.n11036 avdd.n11035 0.0111818
R12041 avdd.n9053 avdd.n9052 0.0111818
R12042 avdd.n9058 avdd.n9057 0.0111818
R12043 avdd.n9109 avdd.n9108 0.0111818
R12044 avdd.n11097 avdd.n11096 0.0111818
R12045 avdd.n11132 avdd.n11131 0.0111818
R12046 avdd.n11138 avdd.n11137 0.0111818
R12047 avdd.n8939 avdd.n8938 0.0111818
R12048 avdd.n8944 avdd.n8943 0.0111818
R12049 avdd.n8995 avdd.n8994 0.0111818
R12050 avdd.n11199 avdd.n11198 0.0111818
R12051 avdd.n11234 avdd.n11233 0.0111818
R12052 avdd.n11240 avdd.n11239 0.0111818
R12053 avdd.n73 avdd.n72 0.0111818
R12054 avdd.n77 avdd.n76 0.0111818
R12055 avdd.n131 avdd.n130 0.0111818
R12056 avdd.n184 avdd.n183 0.0111818
R12057 avdd.n137 avdd.n136 0.0111818
R12058 avdd.n8847 avdd.n8846 0.0111818
R12059 avdd.n203 avdd.n202 0.0111818
R12060 avdd.n207 avdd.n206 0.0111818
R12061 avdd.n261 avdd.n260 0.0111818
R12062 avdd.n314 avdd.n313 0.0111818
R12063 avdd.n267 avdd.n266 0.0111818
R12064 avdd.n8761 avdd.n8760 0.0111818
R12065 avdd.n333 avdd.n332 0.0111818
R12066 avdd.n337 avdd.n336 0.0111818
R12067 avdd.n391 avdd.n390 0.0111818
R12068 avdd.n444 avdd.n443 0.0111818
R12069 avdd.n397 avdd.n396 0.0111818
R12070 avdd.n8675 avdd.n8674 0.0111818
R12071 avdd.n463 avdd.n462 0.0111818
R12072 avdd.n467 avdd.n466 0.0111818
R12073 avdd.n521 avdd.n520 0.0111818
R12074 avdd.n574 avdd.n573 0.0111818
R12075 avdd.n527 avdd.n526 0.0111818
R12076 avdd.n8589 avdd.n8588 0.0111818
R12077 avdd.n593 avdd.n592 0.0111818
R12078 avdd.n597 avdd.n596 0.0111818
R12079 avdd.n651 avdd.n650 0.0111818
R12080 avdd.n704 avdd.n703 0.0111818
R12081 avdd.n657 avdd.n656 0.0111818
R12082 avdd.n8503 avdd.n8502 0.0111818
R12083 avdd.n723 avdd.n722 0.0111818
R12084 avdd.n727 avdd.n726 0.0111818
R12085 avdd.n781 avdd.n780 0.0111818
R12086 avdd.n834 avdd.n833 0.0111818
R12087 avdd.n787 avdd.n786 0.0111818
R12088 avdd.n8417 avdd.n8416 0.0111818
R12089 avdd.n853 avdd.n852 0.0111818
R12090 avdd.n857 avdd.n856 0.0111818
R12091 avdd.n911 avdd.n910 0.0111818
R12092 avdd.n964 avdd.n963 0.0111818
R12093 avdd.n917 avdd.n916 0.0111818
R12094 avdd.n8331 avdd.n8330 0.0111818
R12095 avdd.n983 avdd.n982 0.0111818
R12096 avdd.n987 avdd.n986 0.0111818
R12097 avdd.n1041 avdd.n1040 0.0111818
R12098 avdd.n1094 avdd.n1093 0.0111818
R12099 avdd.n1047 avdd.n1046 0.0111818
R12100 avdd.n8245 avdd.n8244 0.0111818
R12101 avdd.n1113 avdd.n1112 0.0111818
R12102 avdd.n1117 avdd.n1116 0.0111818
R12103 avdd.n1171 avdd.n1170 0.0111818
R12104 avdd.n1224 avdd.n1223 0.0111818
R12105 avdd.n1177 avdd.n1176 0.0111818
R12106 avdd.n8159 avdd.n8158 0.0111818
R12107 avdd.n1243 avdd.n1242 0.0111818
R12108 avdd.n1247 avdd.n1246 0.0111818
R12109 avdd.n1301 avdd.n1300 0.0111818
R12110 avdd.n1354 avdd.n1353 0.0111818
R12111 avdd.n1307 avdd.n1306 0.0111818
R12112 avdd.n8073 avdd.n8072 0.0111818
R12113 avdd.n1373 avdd.n1372 0.0111818
R12114 avdd.n1377 avdd.n1376 0.0111818
R12115 avdd.n1431 avdd.n1430 0.0111818
R12116 avdd.n1484 avdd.n1483 0.0111818
R12117 avdd.n1437 avdd.n1436 0.0111818
R12118 avdd.n7987 avdd.n7986 0.0111818
R12119 avdd.n1503 avdd.n1502 0.0111818
R12120 avdd.n1507 avdd.n1506 0.0111818
R12121 avdd.n1561 avdd.n1560 0.0111818
R12122 avdd.n1614 avdd.n1613 0.0111818
R12123 avdd.n1567 avdd.n1566 0.0111818
R12124 avdd.n7901 avdd.n7900 0.0111818
R12125 avdd.n4627 avdd.n4626 0.0109167
R12126 avdd.n7639 avdd 0.0108238
R12127 avdd.n2017 avdd.n2007 0.0105866
R12128 avdd.n2011 avdd.n2007 0.0105866
R12129 avdd.n2291 avdd.n2290 0.0105866
R12130 avdd.n2290 avdd.n2094 0.0105866
R12131 avdd.n2506 avdd.n2505 0.0105866
R12132 avdd.n2505 avdd.n2309 0.0105866
R12133 avdd.n2721 avdd.n2720 0.0105866
R12134 avdd.n2720 avdd.n2524 0.0105866
R12135 avdd.n2936 avdd.n2935 0.0105866
R12136 avdd.n2935 avdd.n2739 0.0105866
R12137 avdd.n3151 avdd.n3150 0.0105866
R12138 avdd.n3150 avdd.n2954 0.0105866
R12139 avdd.n5008 avdd.n4814 0.0105866
R12140 avdd.n4814 avdd.n4810 0.0105866
R12141 avdd.n5224 avdd.n5030 0.0105866
R12142 avdd.n5030 avdd.n5026 0.0105866
R12143 avdd.n5440 avdd.n5246 0.0105866
R12144 avdd.n5246 avdd.n5242 0.0105866
R12145 avdd.n5656 avdd.n5462 0.0105866
R12146 avdd.n5462 avdd.n5458 0.0105866
R12147 avdd.n5872 avdd.n5678 0.0105866
R12148 avdd.n5678 avdd.n5674 0.0105866
R12149 avdd.n6088 avdd.n5894 0.0105866
R12150 avdd.n5894 avdd.n5890 0.0105866
R12151 avdd.n6304 avdd.n6110 0.0105866
R12152 avdd.n6110 avdd.n6106 0.0105866
R12153 avdd.n6520 avdd.n6326 0.0105866
R12154 avdd.n6326 avdd.n6322 0.0105866
R12155 avdd.n6736 avdd.n6542 0.0105866
R12156 avdd.n6542 avdd.n6538 0.0105866
R12157 avdd.n6952 avdd.n6758 0.0105866
R12158 avdd.n6758 avdd.n6754 0.0105866
R12159 avdd.n7168 avdd.n6974 0.0105866
R12160 avdd.n6974 avdd.n6970 0.0105866
R12161 avdd.n7384 avdd.n7190 0.0105866
R12162 avdd.n7190 avdd.n7186 0.0105866
R12163 avdd.n10338 avdd.n10337 0.0105866
R12164 avdd.n10339 avdd.n10338 0.0105866
R12165 avdd.n10440 avdd.n10439 0.0105866
R12166 avdd.n10441 avdd.n10440 0.0105866
R12167 avdd.n10542 avdd.n10541 0.0105866
R12168 avdd.n10543 avdd.n10542 0.0105866
R12169 avdd.n10644 avdd.n10643 0.0105866
R12170 avdd.n10645 avdd.n10644 0.0105866
R12171 avdd.n10746 avdd.n10745 0.0105866
R12172 avdd.n10747 avdd.n10746 0.0105866
R12173 avdd.n10848 avdd.n10847 0.0105866
R12174 avdd.n10849 avdd.n10848 0.0105866
R12175 avdd.n10950 avdd.n10949 0.0105866
R12176 avdd.n10951 avdd.n10950 0.0105866
R12177 avdd.n11052 avdd.n11051 0.0105866
R12178 avdd.n11053 avdd.n11052 0.0105866
R12179 avdd.n11154 avdd.n11153 0.0105866
R12180 avdd.n11155 avdd.n11154 0.0105866
R12181 avdd.n11256 avdd.n11255 0.0105866
R12182 avdd.n11257 avdd.n11256 0.0105866
R12183 avdd.n8869 avdd.n8868 0.0105866
R12184 avdd.n8870 avdd.n8869 0.0105866
R12185 avdd.n8783 avdd.n8782 0.0105866
R12186 avdd.n8784 avdd.n8783 0.0105866
R12187 avdd.n8697 avdd.n8696 0.0105866
R12188 avdd.n8698 avdd.n8697 0.0105866
R12189 avdd.n8611 avdd.n8610 0.0105866
R12190 avdd.n8612 avdd.n8611 0.0105866
R12191 avdd.n8525 avdd.n8524 0.0105866
R12192 avdd.n8526 avdd.n8525 0.0105866
R12193 avdd.n8439 avdd.n8438 0.0105866
R12194 avdd.n8440 avdd.n8439 0.0105866
R12195 avdd.n8353 avdd.n8352 0.0105866
R12196 avdd.n8354 avdd.n8353 0.0105866
R12197 avdd.n8267 avdd.n8266 0.0105866
R12198 avdd.n8268 avdd.n8267 0.0105866
R12199 avdd.n8181 avdd.n8180 0.0105866
R12200 avdd.n8182 avdd.n8181 0.0105866
R12201 avdd.n8095 avdd.n8094 0.0105866
R12202 avdd.n8096 avdd.n8095 0.0105866
R12203 avdd.n8009 avdd.n8008 0.0105866
R12204 avdd.n8010 avdd.n8009 0.0105866
R12205 avdd.n7923 avdd.n7922 0.0105866
R12206 avdd.n7924 avdd.n7923 0.0105866
R12207 avdd.n1904 avdd.n1903 0.0104697
R12208 avdd.n2060 avdd.n2059 0.0104697
R12209 avdd.n2158 avdd.n2157 0.0104697
R12210 avdd.n2240 avdd.n2239 0.0104697
R12211 avdd.n2373 avdd.n2372 0.0104697
R12212 avdd.n2455 avdd.n2454 0.0104697
R12213 avdd.n2588 avdd.n2587 0.0104697
R12214 avdd.n2670 avdd.n2669 0.0104697
R12215 avdd.n2803 avdd.n2802 0.0104697
R12216 avdd.n2885 avdd.n2884 0.0104697
R12217 avdd.n3018 avdd.n3017 0.0104697
R12218 avdd.n3100 avdd.n3099 0.0104697
R12219 avdd.n3194 avdd.n3193 0.0104697
R12220 avdd.n3349 avdd.n3348 0.0104697
R12221 avdd.n3409 avdd.n3408 0.0104697
R12222 avdd.n3564 avdd.n3563 0.0104697
R12223 avdd.n3624 avdd.n3623 0.0104697
R12224 avdd.n3779 avdd.n3778 0.0104697
R12225 avdd.n3839 avdd.n3838 0.0104697
R12226 avdd.n3994 avdd.n3993 0.0104697
R12227 avdd.n4054 avdd.n4053 0.0104697
R12228 avdd.n4209 avdd.n4208 0.0104697
R12229 avdd.n4269 avdd.n4268 0.0104697
R12230 avdd.n4424 avdd.n4423 0.0104697
R12231 avdd.n4880 avdd.n4879 0.0104697
R12232 avdd.n4962 avdd.n4961 0.0104697
R12233 avdd.n5096 avdd.n5095 0.0104697
R12234 avdd.n5178 avdd.n5177 0.0104697
R12235 avdd.n5312 avdd.n5311 0.0104697
R12236 avdd.n5394 avdd.n5393 0.0104697
R12237 avdd.n5528 avdd.n5527 0.0104697
R12238 avdd.n5610 avdd.n5609 0.0104697
R12239 avdd.n5744 avdd.n5743 0.0104697
R12240 avdd.n5826 avdd.n5825 0.0104697
R12241 avdd.n5960 avdd.n5959 0.0104697
R12242 avdd.n6042 avdd.n6041 0.0104697
R12243 avdd.n6176 avdd.n6175 0.0104697
R12244 avdd.n6258 avdd.n6257 0.0104697
R12245 avdd.n6392 avdd.n6391 0.0104697
R12246 avdd.n6474 avdd.n6473 0.0104697
R12247 avdd.n6608 avdd.n6607 0.0104697
R12248 avdd.n6690 avdd.n6689 0.0104697
R12249 avdd.n6824 avdd.n6823 0.0104697
R12250 avdd.n6906 avdd.n6905 0.0104697
R12251 avdd.n7040 avdd.n7039 0.0104697
R12252 avdd.n7122 avdd.n7121 0.0104697
R12253 avdd.n7256 avdd.n7255 0.0104697
R12254 avdd.n7338 avdd.n7337 0.0104697
R12255 avdd.n7743 avdd.n7742 0.0104697
R12256 avdd.n7654 avdd.n7653 0.0104697
R12257 avdd.n10222 avdd.n10221 0.0104697
R12258 avdd.n10132 avdd.n10131 0.0104697
R12259 avdd.n9969 avdd.n9968 0.0104697
R12260 avdd.n10282 avdd.n10281 0.0104697
R12261 avdd.n9855 avdd.n9854 0.0104697
R12262 avdd.n10384 avdd.n10383 0.0104697
R12263 avdd.n9741 avdd.n9740 0.0104697
R12264 avdd.n10486 avdd.n10485 0.0104697
R12265 avdd.n9628 avdd.n9627 0.0104697
R12266 avdd.n10588 avdd.n10587 0.0104697
R12267 avdd.n9513 avdd.n9512 0.0104697
R12268 avdd.n10690 avdd.n10689 0.0104697
R12269 avdd.n9399 avdd.n9398 0.0104697
R12270 avdd.n10792 avdd.n10791 0.0104697
R12271 avdd.n9285 avdd.n9284 0.0104697
R12272 avdd.n10894 avdd.n10893 0.0104697
R12273 avdd.n9171 avdd.n9170 0.0104697
R12274 avdd.n10996 avdd.n10995 0.0104697
R12275 avdd.n9057 avdd.n9056 0.0104697
R12276 avdd.n11098 avdd.n11097 0.0104697
R12277 avdd.n8943 avdd.n8942 0.0104697
R12278 avdd.n11200 avdd.n11199 0.0104697
R12279 avdd.n76 avdd.n75 0.0104697
R12280 avdd.n136 avdd.n135 0.0104697
R12281 avdd.n206 avdd.n205 0.0104697
R12282 avdd.n266 avdd.n265 0.0104697
R12283 avdd.n336 avdd.n335 0.0104697
R12284 avdd.n396 avdd.n395 0.0104697
R12285 avdd.n466 avdd.n465 0.0104697
R12286 avdd.n526 avdd.n525 0.0104697
R12287 avdd.n596 avdd.n595 0.0104697
R12288 avdd.n656 avdd.n655 0.0104697
R12289 avdd.n726 avdd.n725 0.0104697
R12290 avdd.n786 avdd.n785 0.0104697
R12291 avdd.n856 avdd.n855 0.0104697
R12292 avdd.n916 avdd.n915 0.0104697
R12293 avdd.n986 avdd.n985 0.0104697
R12294 avdd.n1046 avdd.n1045 0.0104697
R12295 avdd.n1116 avdd.n1115 0.0104697
R12296 avdd.n1176 avdd.n1175 0.0104697
R12297 avdd.n1246 avdd.n1245 0.0104697
R12298 avdd.n1306 avdd.n1305 0.0104697
R12299 avdd.n1376 avdd.n1375 0.0104697
R12300 avdd.n1436 avdd.n1435 0.0104697
R12301 avdd.n1506 avdd.n1505 0.0104697
R12302 avdd.n1566 avdd.n1565 0.0104697
R12303 avdd.n1909 avdd.n1908 0.00997968
R12304 avdd.n2163 avdd.n2162 0.00997968
R12305 avdd.n2378 avdd.n2377 0.00997968
R12306 avdd.n2593 avdd.n2592 0.00997968
R12307 avdd.n2808 avdd.n2807 0.00997968
R12308 avdd.n3023 avdd.n3022 0.00997968
R12309 avdd.n3199 avdd.n3198 0.00997968
R12310 avdd.n3414 avdd.n3413 0.00997968
R12311 avdd.n3629 avdd.n3628 0.00997968
R12312 avdd.n3844 avdd.n3843 0.00997968
R12313 avdd.n4059 avdd.n4058 0.00997968
R12314 avdd.n4274 avdd.n4273 0.00997968
R12315 avdd.n4885 avdd.n4884 0.00997968
R12316 avdd.n5101 avdd.n5100 0.00997968
R12317 avdd.n5317 avdd.n5316 0.00997968
R12318 avdd.n5533 avdd.n5532 0.00997968
R12319 avdd.n5749 avdd.n5748 0.00997968
R12320 avdd.n5965 avdd.n5964 0.00997968
R12321 avdd.n6181 avdd.n6180 0.00997968
R12322 avdd.n6397 avdd.n6396 0.00997968
R12323 avdd.n6613 avdd.n6612 0.00997968
R12324 avdd.n6829 avdd.n6828 0.00997968
R12325 avdd.n7045 avdd.n7044 0.00997968
R12326 avdd.n7261 avdd.n7260 0.00997968
R12327 avdd.n7754 avdd.n7753 0.00997968
R12328 avdd.n10233 avdd.n10232 0.00997968
R12329 avdd.n9987 avdd.n9986 0.00997968
R12330 avdd.n9873 avdd.n9872 0.00997968
R12331 avdd.n9759 avdd.n9758 0.00997968
R12332 avdd.n9646 avdd.n9645 0.00997968
R12333 avdd.n9531 avdd.n9530 0.00997968
R12334 avdd.n9417 avdd.n9416 0.00997968
R12335 avdd.n9303 avdd.n9302 0.00997968
R12336 avdd.n9189 avdd.n9188 0.00997968
R12337 avdd.n9075 avdd.n9074 0.00997968
R12338 avdd.n8961 avdd.n8960 0.00997968
R12339 avdd.n87 avdd.n86 0.00997968
R12340 avdd.n217 avdd.n216 0.00997968
R12341 avdd.n347 avdd.n346 0.00997968
R12342 avdd.n477 avdd.n476 0.00997968
R12343 avdd.n607 avdd.n606 0.00997968
R12344 avdd.n737 avdd.n736 0.00997968
R12345 avdd.n867 avdd.n866 0.00997968
R12346 avdd.n997 avdd.n996 0.00997968
R12347 avdd.n1127 avdd.n1126 0.00997968
R12348 avdd.n1257 avdd.n1256 0.00997968
R12349 avdd.n1387 avdd.n1386 0.00997968
R12350 avdd.n1517 avdd.n1516 0.00997968
R12351 avdd.n1963 avdd.n1948 0.0099697
R12352 avdd.n2026 avdd.n2025 0.0099697
R12353 avdd.n2226 avdd.n2225 0.0099697
R12354 avdd.n2300 avdd.n2299 0.0099697
R12355 avdd.n2441 avdd.n2440 0.0099697
R12356 avdd.n2515 avdd.n2514 0.0099697
R12357 avdd.n2656 avdd.n2655 0.0099697
R12358 avdd.n2730 avdd.n2729 0.0099697
R12359 avdd.n2871 avdd.n2870 0.0099697
R12360 avdd.n2945 avdd.n2944 0.0099697
R12361 avdd.n3086 avdd.n3085 0.0099697
R12362 avdd.n3160 avdd.n3159 0.0099697
R12363 avdd.n3253 avdd.n3238 0.0099697
R12364 avdd.n3320 avdd.n3314 0.0099697
R12365 avdd.n3468 avdd.n3453 0.0099697
R12366 avdd.n3535 avdd.n3529 0.0099697
R12367 avdd.n3683 avdd.n3668 0.0099697
R12368 avdd.n3750 avdd.n3744 0.0099697
R12369 avdd.n3898 avdd.n3883 0.0099697
R12370 avdd.n3965 avdd.n3959 0.0099697
R12371 avdd.n4113 avdd.n4098 0.0099697
R12372 avdd.n4180 avdd.n4174 0.0099697
R12373 avdd.n4328 avdd.n4313 0.0099697
R12374 avdd.n4395 avdd.n4389 0.0099697
R12375 avdd.n4948 avdd.n4947 0.0099697
R12376 avdd.n5017 avdd.n5014 0.0099697
R12377 avdd.n5164 avdd.n5163 0.0099697
R12378 avdd.n5233 avdd.n5230 0.0099697
R12379 avdd.n5380 avdd.n5379 0.0099697
R12380 avdd.n5449 avdd.n5446 0.0099697
R12381 avdd.n5596 avdd.n5595 0.0099697
R12382 avdd.n5665 avdd.n5662 0.0099697
R12383 avdd.n5812 avdd.n5811 0.0099697
R12384 avdd.n5881 avdd.n5878 0.0099697
R12385 avdd.n6028 avdd.n6027 0.0099697
R12386 avdd.n6097 avdd.n6094 0.0099697
R12387 avdd.n6244 avdd.n6243 0.0099697
R12388 avdd.n6313 avdd.n6310 0.0099697
R12389 avdd.n6460 avdd.n6459 0.0099697
R12390 avdd.n6529 avdd.n6526 0.0099697
R12391 avdd.n6676 avdd.n6675 0.0099697
R12392 avdd.n6745 avdd.n6742 0.0099697
R12393 avdd.n6892 avdd.n6891 0.0099697
R12394 avdd.n6961 avdd.n6958 0.0099697
R12395 avdd.n7108 avdd.n7107 0.0099697
R12396 avdd.n7177 avdd.n7174 0.0099697
R12397 avdd.n7324 avdd.n7323 0.0099697
R12398 avdd.n7393 avdd.n7390 0.0099697
R12399 avdd.n7676 avdd.n7673 0.0099697
R12400 avdd.n7789 avdd.n7786 0.0099697
R12401 avdd.n10155 avdd.n10152 0.0099697
R12402 avdd.n10049 avdd.n10046 0.0099697
R12403 avdd.n9939 avdd.n9936 0.0099697
R12404 avdd.n10265 avdd.n10262 0.0099697
R12405 avdd.n9825 avdd.n9822 0.0099697
R12406 avdd.n10367 avdd.n10364 0.0099697
R12407 avdd.n9711 avdd.n9708 0.0099697
R12408 avdd.n10469 avdd.n10466 0.0099697
R12409 avdd.n9598 avdd.n9595 0.0099697
R12410 avdd.n10571 avdd.n10568 0.0099697
R12411 avdd.n9483 avdd.n9480 0.0099697
R12412 avdd.n10673 avdd.n10670 0.0099697
R12413 avdd.n9369 avdd.n9366 0.0099697
R12414 avdd.n10775 avdd.n10772 0.0099697
R12415 avdd.n9255 avdd.n9252 0.0099697
R12416 avdd.n10877 avdd.n10874 0.0099697
R12417 avdd.n9141 avdd.n9138 0.0099697
R12418 avdd.n10979 avdd.n10976 0.0099697
R12419 avdd.n9027 avdd.n9024 0.0099697
R12420 avdd.n11081 avdd.n11078 0.0099697
R12421 avdd.n8913 avdd.n8910 0.0099697
R12422 avdd.n11183 avdd.n11180 0.0099697
R12423 avdd.n159 avdd.n156 0.0099697
R12424 avdd.n8812 avdd.n8809 0.0099697
R12425 avdd.n289 avdd.n286 0.0099697
R12426 avdd.n8726 avdd.n8723 0.0099697
R12427 avdd.n419 avdd.n416 0.0099697
R12428 avdd.n8640 avdd.n8637 0.0099697
R12429 avdd.n549 avdd.n546 0.0099697
R12430 avdd.n8554 avdd.n8551 0.0099697
R12431 avdd.n679 avdd.n676 0.0099697
R12432 avdd.n8468 avdd.n8465 0.0099697
R12433 avdd.n809 avdd.n806 0.0099697
R12434 avdd.n8382 avdd.n8379 0.0099697
R12435 avdd.n939 avdd.n936 0.0099697
R12436 avdd.n8296 avdd.n8293 0.0099697
R12437 avdd.n1069 avdd.n1066 0.0099697
R12438 avdd.n8210 avdd.n8207 0.0099697
R12439 avdd.n1199 avdd.n1196 0.0099697
R12440 avdd.n8124 avdd.n8121 0.0099697
R12441 avdd.n1329 avdd.n1326 0.0099697
R12442 avdd.n8038 avdd.n8035 0.0099697
R12443 avdd.n1459 avdd.n1456 0.0099697
R12444 avdd.n7952 avdd.n7949 0.0099697
R12445 avdd.n1589 avdd.n1586 0.0099697
R12446 avdd.n7866 avdd.n7863 0.0099697
R12447 avdd.n1935 avdd.n1934 0.00987834
R12448 avdd.n1934 avdd.n1879 0.00987834
R12449 avdd.n2194 avdd.n2193 0.00987834
R12450 avdd.n2194 avdd.n2145 0.00987834
R12451 avdd.n2409 avdd.n2408 0.00987834
R12452 avdd.n2409 avdd.n2360 0.00987834
R12453 avdd.n2624 avdd.n2623 0.00987834
R12454 avdd.n2624 avdd.n2575 0.00987834
R12455 avdd.n2839 avdd.n2838 0.00987834
R12456 avdd.n2839 avdd.n2790 0.00987834
R12457 avdd.n3054 avdd.n3053 0.00987834
R12458 avdd.n3054 avdd.n3005 0.00987834
R12459 avdd.n118 avdd.n117 0.00987834
R12460 avdd.n117 avdd.n116 0.00987834
R12461 avdd.n248 avdd.n247 0.00987834
R12462 avdd.n247 avdd.n246 0.00987834
R12463 avdd.n378 avdd.n377 0.00987834
R12464 avdd.n377 avdd.n376 0.00987834
R12465 avdd.n508 avdd.n507 0.00987834
R12466 avdd.n507 avdd.n506 0.00987834
R12467 avdd.n638 avdd.n637 0.00987834
R12468 avdd.n637 avdd.n636 0.00987834
R12469 avdd.n768 avdd.n767 0.00987834
R12470 avdd.n767 avdd.n766 0.00987834
R12471 avdd.n898 avdd.n897 0.00987834
R12472 avdd.n897 avdd.n896 0.00987834
R12473 avdd.n1028 avdd.n1027 0.00987834
R12474 avdd.n1027 avdd.n1026 0.00987834
R12475 avdd.n1158 avdd.n1157 0.00987834
R12476 avdd.n1157 avdd.n1156 0.00987834
R12477 avdd.n1288 avdd.n1287 0.00987834
R12478 avdd.n1287 avdd.n1286 0.00987834
R12479 avdd.n1418 avdd.n1417 0.00987834
R12480 avdd.n1417 avdd.n1416 0.00987834
R12481 avdd.n1548 avdd.n1547 0.00987834
R12482 avdd.n1547 avdd.n1546 0.00987834
R12483 avdd.n3225 avdd.n3224 0.00987834
R12484 avdd.n3224 avdd.n3170 0.00987834
R12485 avdd.n3440 avdd.n3439 0.00987834
R12486 avdd.n3439 avdd.n3385 0.00987834
R12487 avdd.n3655 avdd.n3654 0.00987834
R12488 avdd.n3654 avdd.n3600 0.00987834
R12489 avdd.n3870 avdd.n3869 0.00987834
R12490 avdd.n3869 avdd.n3815 0.00987834
R12491 avdd.n4085 avdd.n4084 0.00987834
R12492 avdd.n4084 avdd.n4030 0.00987834
R12493 avdd.n4300 avdd.n4299 0.00987834
R12494 avdd.n4299 avdd.n4245 0.00987834
R12495 avdd.n2031 avdd.n1994 0.00975758
R12496 avdd.n1884 avdd.n1882 0.00975758
R12497 avdd.n2084 avdd.n1885 0.00975758
R12498 avdd.n2033 avdd.n2032 0.00975758
R12499 avdd.n2038 avdd.n2002 0.00975758
R12500 avdd.n2037 avdd.n2003 0.00975758
R12501 avdd.n2276 avdd.n2275 0.00975758
R12502 avdd.n2140 avdd.n2134 0.00975758
R12503 avdd.n2207 avdd.n2135 0.00975758
R12504 avdd.n2277 avdd.n2106 0.00975758
R12505 avdd.n2283 avdd.n2095 0.00975758
R12506 avdd.n2284 avdd.n2102 0.00975758
R12507 avdd.n2491 avdd.n2490 0.00975758
R12508 avdd.n2355 avdd.n2349 0.00975758
R12509 avdd.n2422 avdd.n2350 0.00975758
R12510 avdd.n2492 avdd.n2321 0.00975758
R12511 avdd.n2498 avdd.n2310 0.00975758
R12512 avdd.n2499 avdd.n2317 0.00975758
R12513 avdd.n2706 avdd.n2705 0.00975758
R12514 avdd.n2570 avdd.n2564 0.00975758
R12515 avdd.n2637 avdd.n2565 0.00975758
R12516 avdd.n2707 avdd.n2536 0.00975758
R12517 avdd.n2713 avdd.n2525 0.00975758
R12518 avdd.n2714 avdd.n2532 0.00975758
R12519 avdd.n2921 avdd.n2920 0.00975758
R12520 avdd.n2785 avdd.n2779 0.00975758
R12521 avdd.n2852 avdd.n2780 0.00975758
R12522 avdd.n2922 avdd.n2751 0.00975758
R12523 avdd.n2928 avdd.n2740 0.00975758
R12524 avdd.n2929 avdd.n2747 0.00975758
R12525 avdd.n3136 avdd.n3135 0.00975758
R12526 avdd.n3000 avdd.n2994 0.00975758
R12527 avdd.n3067 avdd.n2995 0.00975758
R12528 avdd.n3137 avdd.n2966 0.00975758
R12529 avdd.n3143 avdd.n2955 0.00975758
R12530 avdd.n3144 avdd.n2962 0.00975758
R12531 avdd.n3301 avdd.n3284 0.00975758
R12532 avdd.n3174 avdd.n3172 0.00975758
R12533 avdd.n3373 avdd.n3175 0.00975758
R12534 avdd.n3302 avdd.n3300 0.00975758
R12535 avdd.n3327 avdd.n3292 0.00975758
R12536 avdd.n3326 avdd.n3293 0.00975758
R12537 avdd.n3516 avdd.n3499 0.00975758
R12538 avdd.n3389 avdd.n3387 0.00975758
R12539 avdd.n3588 avdd.n3390 0.00975758
R12540 avdd.n3517 avdd.n3515 0.00975758
R12541 avdd.n3542 avdd.n3507 0.00975758
R12542 avdd.n3541 avdd.n3508 0.00975758
R12543 avdd.n3731 avdd.n3714 0.00975758
R12544 avdd.n3604 avdd.n3602 0.00975758
R12545 avdd.n3803 avdd.n3605 0.00975758
R12546 avdd.n3732 avdd.n3730 0.00975758
R12547 avdd.n3757 avdd.n3722 0.00975758
R12548 avdd.n3756 avdd.n3723 0.00975758
R12549 avdd.n3946 avdd.n3929 0.00975758
R12550 avdd.n3819 avdd.n3817 0.00975758
R12551 avdd.n4018 avdd.n3820 0.00975758
R12552 avdd.n3947 avdd.n3945 0.00975758
R12553 avdd.n3972 avdd.n3937 0.00975758
R12554 avdd.n3971 avdd.n3938 0.00975758
R12555 avdd.n4161 avdd.n4144 0.00975758
R12556 avdd.n4034 avdd.n4032 0.00975758
R12557 avdd.n4233 avdd.n4035 0.00975758
R12558 avdd.n4162 avdd.n4160 0.00975758
R12559 avdd.n4187 avdd.n4152 0.00975758
R12560 avdd.n4186 avdd.n4153 0.00975758
R12561 avdd.n4376 avdd.n4359 0.00975758
R12562 avdd.n4249 avdd.n4247 0.00975758
R12563 avdd.n4448 avdd.n4250 0.00975758
R12564 avdd.n4377 avdd.n4375 0.00975758
R12565 avdd.n4402 avdd.n4367 0.00975758
R12566 avdd.n4401 avdd.n4368 0.00975758
R12567 avdd.n4995 avdd.n4994 0.00975758
R12568 avdd.n4863 avdd.n4856 0.00975758
R12569 avdd.n4929 avdd.n4857 0.00975758
R12570 avdd.n4996 avdd.n4828 0.00975758
R12571 avdd.n5001 avdd.n4812 0.00975758
R12572 avdd.n4823 avdd.n4815 0.00975758
R12573 avdd.n5211 avdd.n5210 0.00975758
R12574 avdd.n5079 avdd.n5072 0.00975758
R12575 avdd.n5145 avdd.n5073 0.00975758
R12576 avdd.n5212 avdd.n5044 0.00975758
R12577 avdd.n5217 avdd.n5028 0.00975758
R12578 avdd.n5039 avdd.n5031 0.00975758
R12579 avdd.n5427 avdd.n5426 0.00975758
R12580 avdd.n5295 avdd.n5288 0.00975758
R12581 avdd.n5361 avdd.n5289 0.00975758
R12582 avdd.n5428 avdd.n5260 0.00975758
R12583 avdd.n5433 avdd.n5244 0.00975758
R12584 avdd.n5255 avdd.n5247 0.00975758
R12585 avdd.n5643 avdd.n5642 0.00975758
R12586 avdd.n5511 avdd.n5504 0.00975758
R12587 avdd.n5577 avdd.n5505 0.00975758
R12588 avdd.n5644 avdd.n5476 0.00975758
R12589 avdd.n5649 avdd.n5460 0.00975758
R12590 avdd.n5471 avdd.n5463 0.00975758
R12591 avdd.n5859 avdd.n5858 0.00975758
R12592 avdd.n5727 avdd.n5720 0.00975758
R12593 avdd.n5793 avdd.n5721 0.00975758
R12594 avdd.n5860 avdd.n5692 0.00975758
R12595 avdd.n5865 avdd.n5676 0.00975758
R12596 avdd.n5687 avdd.n5679 0.00975758
R12597 avdd.n6075 avdd.n6074 0.00975758
R12598 avdd.n5943 avdd.n5936 0.00975758
R12599 avdd.n6009 avdd.n5937 0.00975758
R12600 avdd.n6076 avdd.n5908 0.00975758
R12601 avdd.n6081 avdd.n5892 0.00975758
R12602 avdd.n5903 avdd.n5895 0.00975758
R12603 avdd.n6291 avdd.n6290 0.00975758
R12604 avdd.n6159 avdd.n6152 0.00975758
R12605 avdd.n6225 avdd.n6153 0.00975758
R12606 avdd.n6292 avdd.n6124 0.00975758
R12607 avdd.n6297 avdd.n6108 0.00975758
R12608 avdd.n6119 avdd.n6111 0.00975758
R12609 avdd.n6507 avdd.n6506 0.00975758
R12610 avdd.n6375 avdd.n6368 0.00975758
R12611 avdd.n6441 avdd.n6369 0.00975758
R12612 avdd.n6508 avdd.n6340 0.00975758
R12613 avdd.n6513 avdd.n6324 0.00975758
R12614 avdd.n6335 avdd.n6327 0.00975758
R12615 avdd.n6723 avdd.n6722 0.00975758
R12616 avdd.n6591 avdd.n6584 0.00975758
R12617 avdd.n6657 avdd.n6585 0.00975758
R12618 avdd.n6724 avdd.n6556 0.00975758
R12619 avdd.n6729 avdd.n6540 0.00975758
R12620 avdd.n6551 avdd.n6543 0.00975758
R12621 avdd.n6939 avdd.n6938 0.00975758
R12622 avdd.n6807 avdd.n6800 0.00975758
R12623 avdd.n6873 avdd.n6801 0.00975758
R12624 avdd.n6940 avdd.n6772 0.00975758
R12625 avdd.n6945 avdd.n6756 0.00975758
R12626 avdd.n6767 avdd.n6759 0.00975758
R12627 avdd.n7155 avdd.n7154 0.00975758
R12628 avdd.n7023 avdd.n7016 0.00975758
R12629 avdd.n7089 avdd.n7017 0.00975758
R12630 avdd.n7156 avdd.n6988 0.00975758
R12631 avdd.n7161 avdd.n6972 0.00975758
R12632 avdd.n6983 avdd.n6975 0.00975758
R12633 avdd.n7371 avdd.n7370 0.00975758
R12634 avdd.n7239 avdd.n7232 0.00975758
R12635 avdd.n7305 avdd.n7233 0.00975758
R12636 avdd.n7372 avdd.n7204 0.00975758
R12637 avdd.n7377 avdd.n7188 0.00975758
R12638 avdd.n7199 avdd.n7191 0.00975758
R12639 avdd.n7780 avdd.n7779 0.00975758
R12640 avdd.n7700 avdd.n7699 0.00975758
R12641 avdd.n7698 avdd.n7697 0.00975758
R12642 avdd.n7829 avdd.n7828 0.00975758
R12643 avdd.n7833 avdd.n7832 0.00975758
R12644 avdd.n7844 avdd.n7834 0.00975758
R12645 avdd.n10040 avdd.n10039 0.00975758
R12646 avdd.n10179 avdd.n10178 0.00975758
R12647 avdd.n10177 avdd.n10176 0.00975758
R12648 avdd.n10087 avdd.n10086 0.00975758
R12649 avdd.n10091 avdd.n10090 0.00975758
R12650 avdd.n10102 avdd.n10092 0.00975758
R12651 avdd.n10256 avdd.n10255 0.00975758
R12652 avdd.n9963 avdd.n9962 0.00975758
R12653 avdd.n9961 avdd.n9960 0.00975758
R12654 avdd.n10319 avdd.n10318 0.00975758
R12655 avdd.n10323 avdd.n10322 0.00975758
R12656 avdd.n10334 avdd.n10324 0.00975758
R12657 avdd.n10358 avdd.n10357 0.00975758
R12658 avdd.n9849 avdd.n9848 0.00975758
R12659 avdd.n9847 avdd.n9846 0.00975758
R12660 avdd.n10421 avdd.n10420 0.00975758
R12661 avdd.n10425 avdd.n10424 0.00975758
R12662 avdd.n10436 avdd.n10426 0.00975758
R12663 avdd.n10460 avdd.n10459 0.00975758
R12664 avdd.n9735 avdd.n9734 0.00975758
R12665 avdd.n9733 avdd.n9732 0.00975758
R12666 avdd.n10523 avdd.n10522 0.00975758
R12667 avdd.n10527 avdd.n10526 0.00975758
R12668 avdd.n10538 avdd.n10528 0.00975758
R12669 avdd.n10562 avdd.n10561 0.00975758
R12670 avdd.n9622 avdd.n9621 0.00975758
R12671 avdd.n9620 avdd.n9619 0.00975758
R12672 avdd.n10625 avdd.n10624 0.00975758
R12673 avdd.n10629 avdd.n10628 0.00975758
R12674 avdd.n10640 avdd.n10630 0.00975758
R12675 avdd.n10664 avdd.n10663 0.00975758
R12676 avdd.n9507 avdd.n9506 0.00975758
R12677 avdd.n9505 avdd.n9504 0.00975758
R12678 avdd.n10727 avdd.n10726 0.00975758
R12679 avdd.n10731 avdd.n10730 0.00975758
R12680 avdd.n10742 avdd.n10732 0.00975758
R12681 avdd.n10766 avdd.n10765 0.00975758
R12682 avdd.n9393 avdd.n9392 0.00975758
R12683 avdd.n9391 avdd.n9390 0.00975758
R12684 avdd.n10829 avdd.n10828 0.00975758
R12685 avdd.n10833 avdd.n10832 0.00975758
R12686 avdd.n10844 avdd.n10834 0.00975758
R12687 avdd.n10868 avdd.n10867 0.00975758
R12688 avdd.n9279 avdd.n9278 0.00975758
R12689 avdd.n9277 avdd.n9276 0.00975758
R12690 avdd.n10931 avdd.n10930 0.00975758
R12691 avdd.n10935 avdd.n10934 0.00975758
R12692 avdd.n10946 avdd.n10936 0.00975758
R12693 avdd.n10970 avdd.n10969 0.00975758
R12694 avdd.n9165 avdd.n9164 0.00975758
R12695 avdd.n9163 avdd.n9162 0.00975758
R12696 avdd.n11033 avdd.n11032 0.00975758
R12697 avdd.n11037 avdd.n11036 0.00975758
R12698 avdd.n11048 avdd.n11038 0.00975758
R12699 avdd.n11072 avdd.n11071 0.00975758
R12700 avdd.n9051 avdd.n9050 0.00975758
R12701 avdd.n9049 avdd.n9048 0.00975758
R12702 avdd.n11135 avdd.n11134 0.00975758
R12703 avdd.n11139 avdd.n11138 0.00975758
R12704 avdd.n11150 avdd.n11140 0.00975758
R12705 avdd.n11174 avdd.n11173 0.00975758
R12706 avdd.n8937 avdd.n8936 0.00975758
R12707 avdd.n8935 avdd.n8934 0.00975758
R12708 avdd.n11237 avdd.n11236 0.00975758
R12709 avdd.n11241 avdd.n11240 0.00975758
R12710 avdd.n11252 avdd.n11242 0.00975758
R12711 avdd.n8883 avdd.n8882 0.00975758
R12712 avdd.n183 avdd.n182 0.00975758
R12713 avdd.n181 avdd.n180 0.00975758
R12714 avdd.n8850 avdd.n8849 0.00975758
R12715 avdd.n8854 avdd.n8853 0.00975758
R12716 avdd.n8865 avdd.n8855 0.00975758
R12717 avdd.n8797 avdd.n8796 0.00975758
R12718 avdd.n313 avdd.n312 0.00975758
R12719 avdd.n311 avdd.n310 0.00975758
R12720 avdd.n8764 avdd.n8763 0.00975758
R12721 avdd.n8768 avdd.n8767 0.00975758
R12722 avdd.n8779 avdd.n8769 0.00975758
R12723 avdd.n8711 avdd.n8710 0.00975758
R12724 avdd.n443 avdd.n442 0.00975758
R12725 avdd.n441 avdd.n440 0.00975758
R12726 avdd.n8678 avdd.n8677 0.00975758
R12727 avdd.n8682 avdd.n8681 0.00975758
R12728 avdd.n8693 avdd.n8683 0.00975758
R12729 avdd.n8625 avdd.n8624 0.00975758
R12730 avdd.n573 avdd.n572 0.00975758
R12731 avdd.n571 avdd.n570 0.00975758
R12732 avdd.n8592 avdd.n8591 0.00975758
R12733 avdd.n8596 avdd.n8595 0.00975758
R12734 avdd.n8607 avdd.n8597 0.00975758
R12735 avdd.n8539 avdd.n8538 0.00975758
R12736 avdd.n703 avdd.n702 0.00975758
R12737 avdd.n701 avdd.n700 0.00975758
R12738 avdd.n8506 avdd.n8505 0.00975758
R12739 avdd.n8510 avdd.n8509 0.00975758
R12740 avdd.n8521 avdd.n8511 0.00975758
R12741 avdd.n8453 avdd.n8452 0.00975758
R12742 avdd.n833 avdd.n832 0.00975758
R12743 avdd.n831 avdd.n830 0.00975758
R12744 avdd.n8420 avdd.n8419 0.00975758
R12745 avdd.n8424 avdd.n8423 0.00975758
R12746 avdd.n8435 avdd.n8425 0.00975758
R12747 avdd.n8367 avdd.n8366 0.00975758
R12748 avdd.n963 avdd.n962 0.00975758
R12749 avdd.n961 avdd.n960 0.00975758
R12750 avdd.n8334 avdd.n8333 0.00975758
R12751 avdd.n8338 avdd.n8337 0.00975758
R12752 avdd.n8349 avdd.n8339 0.00975758
R12753 avdd.n8281 avdd.n8280 0.00975758
R12754 avdd.n1093 avdd.n1092 0.00975758
R12755 avdd.n1091 avdd.n1090 0.00975758
R12756 avdd.n8248 avdd.n8247 0.00975758
R12757 avdd.n8252 avdd.n8251 0.00975758
R12758 avdd.n8263 avdd.n8253 0.00975758
R12759 avdd.n8195 avdd.n8194 0.00975758
R12760 avdd.n1223 avdd.n1222 0.00975758
R12761 avdd.n1221 avdd.n1220 0.00975758
R12762 avdd.n8162 avdd.n8161 0.00975758
R12763 avdd.n8166 avdd.n8165 0.00975758
R12764 avdd.n8177 avdd.n8167 0.00975758
R12765 avdd.n8109 avdd.n8108 0.00975758
R12766 avdd.n1353 avdd.n1352 0.00975758
R12767 avdd.n1351 avdd.n1350 0.00975758
R12768 avdd.n8076 avdd.n8075 0.00975758
R12769 avdd.n8080 avdd.n8079 0.00975758
R12770 avdd.n8091 avdd.n8081 0.00975758
R12771 avdd.n8023 avdd.n8022 0.00975758
R12772 avdd.n1483 avdd.n1482 0.00975758
R12773 avdd.n1481 avdd.n1480 0.00975758
R12774 avdd.n7990 avdd.n7989 0.00975758
R12775 avdd.n7994 avdd.n7993 0.00975758
R12776 avdd.n8005 avdd.n7995 0.00975758
R12777 avdd.n7937 avdd.n7936 0.00975758
R12778 avdd.n1613 avdd.n1612 0.00975758
R12779 avdd.n1611 avdd.n1610 0.00975758
R12780 avdd.n7904 avdd.n7903 0.00975758
R12781 avdd.n7908 avdd.n7907 0.00975758
R12782 avdd.n7919 avdd.n7909 0.00975758
R12783 avdd.n2066 avdd.n1959 0.00904545
R12784 avdd.n2234 avdd.n2232 0.00904545
R12785 avdd.n2449 avdd.n2447 0.00904545
R12786 avdd.n2664 avdd.n2662 0.00904545
R12787 avdd.n2879 avdd.n2877 0.00904545
R12788 avdd.n3094 avdd.n3092 0.00904545
R12789 avdd.n3355 avdd.n3249 0.00904545
R12790 avdd.n3570 avdd.n3464 0.00904545
R12791 avdd.n3785 avdd.n3679 0.00904545
R12792 avdd.n4000 avdd.n3894 0.00904545
R12793 avdd.n4215 avdd.n4109 0.00904545
R12794 avdd.n4430 avdd.n4324 0.00904545
R12795 avdd.n4956 avdd.n4954 0.00904545
R12796 avdd.n5172 avdd.n5170 0.00904545
R12797 avdd.n5388 avdd.n5386 0.00904545
R12798 avdd.n5604 avdd.n5602 0.00904545
R12799 avdd.n5820 avdd.n5818 0.00904545
R12800 avdd.n6036 avdd.n6034 0.00904545
R12801 avdd.n6252 avdd.n6250 0.00904545
R12802 avdd.n6468 avdd.n6466 0.00904545
R12803 avdd.n6684 avdd.n6682 0.00904545
R12804 avdd.n6900 avdd.n6898 0.00904545
R12805 avdd.n7116 avdd.n7114 0.00904545
R12806 avdd.n7332 avdd.n7330 0.00904545
R12807 avdd.n7664 avdd.n7663 0.00904545
R12808 avdd.n10143 avdd.n10142 0.00904545
R12809 avdd.n10272 avdd.n10271 0.00904545
R12810 avdd.n10374 avdd.n10373 0.00904545
R12811 avdd.n10476 avdd.n10475 0.00904545
R12812 avdd.n10578 avdd.n10577 0.00904545
R12813 avdd.n10680 avdd.n10679 0.00904545
R12814 avdd.n10782 avdd.n10781 0.00904545
R12815 avdd.n10884 avdd.n10883 0.00904545
R12816 avdd.n10986 avdd.n10985 0.00904545
R12817 avdd.n11088 avdd.n11087 0.00904545
R12818 avdd.n11190 avdd.n11189 0.00904545
R12819 avdd.n147 avdd.n146 0.00904545
R12820 avdd.n277 avdd.n276 0.00904545
R12821 avdd.n407 avdd.n406 0.00904545
R12822 avdd.n537 avdd.n536 0.00904545
R12823 avdd.n667 avdd.n666 0.00904545
R12824 avdd.n797 avdd.n796 0.00904545
R12825 avdd.n927 avdd.n926 0.00904545
R12826 avdd.n1057 avdd.n1056 0.00904545
R12827 avdd.n1187 avdd.n1186 0.00904545
R12828 avdd.n1317 avdd.n1316 0.00904545
R12829 avdd.n1447 avdd.n1446 0.00904545
R12830 avdd.n1577 avdd.n1576 0.00904545
R12831 avdd.n4594 avdd.n4593 0.00883333
R12832 avdd.n1987 avdd.n1972 0.00833333
R12833 avdd.n1928 avdd.n1926 0.00833333
R12834 avdd.n1997 avdd.n1980 0.00833333
R12835 avdd.n2257 avdd.n2251 0.00833333
R12836 avdd.n2181 avdd.n2180 0.00833333
R12837 avdd.n2265 avdd.n2109 0.00833333
R12838 avdd.n2472 avdd.n2466 0.00833333
R12839 avdd.n2396 avdd.n2395 0.00833333
R12840 avdd.n2480 avdd.n2324 0.00833333
R12841 avdd.n2687 avdd.n2681 0.00833333
R12842 avdd.n2611 avdd.n2610 0.00833333
R12843 avdd.n2695 avdd.n2539 0.00833333
R12844 avdd.n2902 avdd.n2896 0.00833333
R12845 avdd.n2826 avdd.n2825 0.00833333
R12846 avdd.n2910 avdd.n2754 0.00833333
R12847 avdd.n3117 avdd.n3111 0.00833333
R12848 avdd.n3041 avdd.n3040 0.00833333
R12849 avdd.n3125 avdd.n2969 0.00833333
R12850 avdd.n3277 avdd.n3262 0.00833333
R12851 avdd.n3218 avdd.n3216 0.00833333
R12852 avdd.n3287 avdd.n3270 0.00833333
R12853 avdd.n3492 avdd.n3477 0.00833333
R12854 avdd.n3433 avdd.n3431 0.00833333
R12855 avdd.n3502 avdd.n3485 0.00833333
R12856 avdd.n3707 avdd.n3692 0.00833333
R12857 avdd.n3648 avdd.n3646 0.00833333
R12858 avdd.n3717 avdd.n3700 0.00833333
R12859 avdd.n3922 avdd.n3907 0.00833333
R12860 avdd.n3863 avdd.n3861 0.00833333
R12861 avdd.n3932 avdd.n3915 0.00833333
R12862 avdd.n4137 avdd.n4122 0.00833333
R12863 avdd.n4078 avdd.n4076 0.00833333
R12864 avdd.n4147 avdd.n4130 0.00833333
R12865 avdd.n4352 avdd.n4337 0.00833333
R12866 avdd.n4293 avdd.n4291 0.00833333
R12867 avdd.n4362 avdd.n4345 0.00833333
R12868 avdd.n4979 avdd.n4973 0.00833333
R12869 avdd.n4904 avdd.n4902 0.00833333
R12870 avdd.n4987 avdd.n4831 0.00833333
R12871 avdd.n5195 avdd.n5189 0.00833333
R12872 avdd.n5120 avdd.n5118 0.00833333
R12873 avdd.n5203 avdd.n5047 0.00833333
R12874 avdd.n5411 avdd.n5405 0.00833333
R12875 avdd.n5336 avdd.n5334 0.00833333
R12876 avdd.n5419 avdd.n5263 0.00833333
R12877 avdd.n5627 avdd.n5621 0.00833333
R12878 avdd.n5552 avdd.n5550 0.00833333
R12879 avdd.n5635 avdd.n5479 0.00833333
R12880 avdd.n5843 avdd.n5837 0.00833333
R12881 avdd.n5768 avdd.n5766 0.00833333
R12882 avdd.n5851 avdd.n5695 0.00833333
R12883 avdd.n6059 avdd.n6053 0.00833333
R12884 avdd.n5984 avdd.n5982 0.00833333
R12885 avdd.n6067 avdd.n5911 0.00833333
R12886 avdd.n6275 avdd.n6269 0.00833333
R12887 avdd.n6200 avdd.n6198 0.00833333
R12888 avdd.n6283 avdd.n6127 0.00833333
R12889 avdd.n6491 avdd.n6485 0.00833333
R12890 avdd.n6416 avdd.n6414 0.00833333
R12891 avdd.n6499 avdd.n6343 0.00833333
R12892 avdd.n6707 avdd.n6701 0.00833333
R12893 avdd.n6632 avdd.n6630 0.00833333
R12894 avdd.n6715 avdd.n6559 0.00833333
R12895 avdd.n6923 avdd.n6917 0.00833333
R12896 avdd.n6848 avdd.n6846 0.00833333
R12897 avdd.n6931 avdd.n6775 0.00833333
R12898 avdd.n7139 avdd.n7133 0.00833333
R12899 avdd.n7064 avdd.n7062 0.00833333
R12900 avdd.n7147 avdd.n6991 0.00833333
R12901 avdd.n7355 avdd.n7349 0.00833333
R12902 avdd.n7280 avdd.n7278 0.00833333
R12903 avdd.n7363 avdd.n7207 0.00833333
R12904 avdd.n7772 avdd.n7771 0.00833333
R12905 avdd.n7760 avdd.n7759 0.00833333
R12906 avdd.n7815 avdd.n7814 0.00833333
R12907 avdd.n10032 avdd.n10031 0.00833333
R12908 avdd.n10239 avdd.n10238 0.00833333
R12909 avdd.n10073 avdd.n10072 0.00833333
R12910 avdd.n10248 avdd.n10247 0.00833333
R12911 avdd.n10004 avdd.n9992 0.00833333
R12912 avdd.n10305 avdd.n10304 0.00833333
R12913 avdd.n10350 avdd.n10349 0.00833333
R12914 avdd.n9890 avdd.n9878 0.00833333
R12915 avdd.n10407 avdd.n10406 0.00833333
R12916 avdd.n10452 avdd.n10451 0.00833333
R12917 avdd.n9776 avdd.n9764 0.00833333
R12918 avdd.n10509 avdd.n10508 0.00833333
R12919 avdd.n10554 avdd.n10553 0.00833333
R12920 avdd.n9663 avdd.n9651 0.00833333
R12921 avdd.n10611 avdd.n10610 0.00833333
R12922 avdd.n10656 avdd.n10655 0.00833333
R12923 avdd.n9548 avdd.n9536 0.00833333
R12924 avdd.n10713 avdd.n10712 0.00833333
R12925 avdd.n10758 avdd.n10757 0.00833333
R12926 avdd.n9434 avdd.n9422 0.00833333
R12927 avdd.n10815 avdd.n10814 0.00833333
R12928 avdd.n10860 avdd.n10859 0.00833333
R12929 avdd.n9320 avdd.n9308 0.00833333
R12930 avdd.n10917 avdd.n10916 0.00833333
R12931 avdd.n10962 avdd.n10961 0.00833333
R12932 avdd.n9206 avdd.n9194 0.00833333
R12933 avdd.n11019 avdd.n11018 0.00833333
R12934 avdd.n11064 avdd.n11063 0.00833333
R12935 avdd.n9092 avdd.n9080 0.00833333
R12936 avdd.n11121 avdd.n11120 0.00833333
R12937 avdd.n11166 avdd.n11165 0.00833333
R12938 avdd.n8978 avdd.n8966 0.00833333
R12939 avdd.n11223 avdd.n11222 0.00833333
R12940 avdd.n8875 avdd.n8874 0.00833333
R12941 avdd.n93 avdd.n92 0.00833333
R12942 avdd.n8836 avdd.n8835 0.00833333
R12943 avdd.n8789 avdd.n8788 0.00833333
R12944 avdd.n223 avdd.n222 0.00833333
R12945 avdd.n8750 avdd.n8749 0.00833333
R12946 avdd.n8703 avdd.n8702 0.00833333
R12947 avdd.n353 avdd.n352 0.00833333
R12948 avdd.n8664 avdd.n8663 0.00833333
R12949 avdd.n8617 avdd.n8616 0.00833333
R12950 avdd.n483 avdd.n482 0.00833333
R12951 avdd.n8578 avdd.n8577 0.00833333
R12952 avdd.n8531 avdd.n8530 0.00833333
R12953 avdd.n613 avdd.n612 0.00833333
R12954 avdd.n8492 avdd.n8491 0.00833333
R12955 avdd.n8445 avdd.n8444 0.00833333
R12956 avdd.n743 avdd.n742 0.00833333
R12957 avdd.n8406 avdd.n8405 0.00833333
R12958 avdd.n8359 avdd.n8358 0.00833333
R12959 avdd.n873 avdd.n872 0.00833333
R12960 avdd.n8320 avdd.n8319 0.00833333
R12961 avdd.n8273 avdd.n8272 0.00833333
R12962 avdd.n1003 avdd.n1002 0.00833333
R12963 avdd.n8234 avdd.n8233 0.00833333
R12964 avdd.n8187 avdd.n8186 0.00833333
R12965 avdd.n1133 avdd.n1132 0.00833333
R12966 avdd.n8148 avdd.n8147 0.00833333
R12967 avdd.n8101 avdd.n8100 0.00833333
R12968 avdd.n1263 avdd.n1262 0.00833333
R12969 avdd.n8062 avdd.n8061 0.00833333
R12970 avdd.n8015 avdd.n8014 0.00833333
R12971 avdd.n1393 avdd.n1392 0.00833333
R12972 avdd.n7976 avdd.n7975 0.00833333
R12973 avdd.n7929 avdd.n7928 0.00833333
R12974 avdd.n1523 avdd.n1522 0.00833333
R12975 avdd.n7890 avdd.n7889 0.00833333
R12976 avdd.n1939 avdd.n1891 0.00833333
R12977 avdd.n2189 avdd.n2146 0.00833333
R12978 avdd.n2404 avdd.n2361 0.00833333
R12979 avdd.n2619 avdd.n2576 0.00833333
R12980 avdd.n2834 avdd.n2791 0.00833333
R12981 avdd.n3049 avdd.n3006 0.00833333
R12982 avdd.n3229 avdd.n3181 0.00833333
R12983 avdd.n3444 avdd.n3396 0.00833333
R12984 avdd.n3659 avdd.n3611 0.00833333
R12985 avdd.n3874 avdd.n3826 0.00833333
R12986 avdd.n4089 avdd.n4041 0.00833333
R12987 avdd.n4304 avdd.n4256 0.00833333
R12988 avdd.n4912 avdd.n4868 0.00833333
R12989 avdd.n5128 avdd.n5084 0.00833333
R12990 avdd.n5344 avdd.n5300 0.00833333
R12991 avdd.n5560 avdd.n5516 0.00833333
R12992 avdd.n5776 avdd.n5732 0.00833333
R12993 avdd.n5992 avdd.n5948 0.00833333
R12994 avdd.n6208 avdd.n6164 0.00833333
R12995 avdd.n6424 avdd.n6380 0.00833333
R12996 avdd.n6640 avdd.n6596 0.00833333
R12997 avdd.n6856 avdd.n6812 0.00833333
R12998 avdd.n7072 avdd.n7028 0.00833333
R12999 avdd.n7288 avdd.n7244 0.00833333
R13000 avdd.n7725 avdd.n7724 0.00833333
R13001 avdd.n10204 avdd.n10203 0.00833333
R13002 avdd.n10007 avdd.n10006 0.00833333
R13003 avdd.n9893 avdd.n9892 0.00833333
R13004 avdd.n9779 avdd.n9778 0.00833333
R13005 avdd.n9666 avdd.n9665 0.00833333
R13006 avdd.n9551 avdd.n9550 0.00833333
R13007 avdd.n9437 avdd.n9436 0.00833333
R13008 avdd.n9323 avdd.n9322 0.00833333
R13009 avdd.n9209 avdd.n9208 0.00833333
R13010 avdd.n9095 avdd.n9094 0.00833333
R13011 avdd.n8981 avdd.n8980 0.00833333
R13012 avdd.n120 avdd.n119 0.00833333
R13013 avdd.n250 avdd.n249 0.00833333
R13014 avdd.n380 avdd.n379 0.00833333
R13015 avdd.n510 avdd.n509 0.00833333
R13016 avdd.n640 avdd.n639 0.00833333
R13017 avdd.n770 avdd.n769 0.00833333
R13018 avdd.n900 avdd.n899 0.00833333
R13019 avdd.n1030 avdd.n1029 0.00833333
R13020 avdd.n1160 avdd.n1159 0.00833333
R13021 avdd.n1290 avdd.n1289 0.00833333
R13022 avdd.n1420 avdd.n1419 0.00833333
R13023 avdd.n1550 avdd.n1549 0.00833333
R13024 avdd.n2039 avdd.n2001 0.00807576
R13025 avdd.n2048 avdd.n1978 0.00807576
R13026 avdd.n2053 avdd.n2052 0.00807576
R13027 avdd.n2083 avdd.n1886 0.00807576
R13028 avdd.n1937 avdd.n1936 0.00807576
R13029 avdd.n1922 avdd.n1921 0.00807576
R13030 avdd.n2285 avdd.n2282 0.00807576
R13031 avdd.n2268 avdd.n2267 0.00807576
R13032 avdd.n2247 avdd.n2246 0.00807576
R13033 avdd.n2206 avdd.n2202 0.00807576
R13034 avdd.n2192 avdd.n2191 0.00807576
R13035 avdd.n2176 avdd.n2175 0.00807576
R13036 avdd.n2500 avdd.n2497 0.00807576
R13037 avdd.n2483 avdd.n2482 0.00807576
R13038 avdd.n2462 avdd.n2461 0.00807576
R13039 avdd.n2421 avdd.n2417 0.00807576
R13040 avdd.n2407 avdd.n2406 0.00807576
R13041 avdd.n2391 avdd.n2390 0.00807576
R13042 avdd.n2715 avdd.n2712 0.00807576
R13043 avdd.n2698 avdd.n2697 0.00807576
R13044 avdd.n2677 avdd.n2676 0.00807576
R13045 avdd.n2636 avdd.n2632 0.00807576
R13046 avdd.n2622 avdd.n2621 0.00807576
R13047 avdd.n2606 avdd.n2605 0.00807576
R13048 avdd.n2930 avdd.n2927 0.00807576
R13049 avdd.n2913 avdd.n2912 0.00807576
R13050 avdd.n2892 avdd.n2891 0.00807576
R13051 avdd.n2851 avdd.n2847 0.00807576
R13052 avdd.n2837 avdd.n2836 0.00807576
R13053 avdd.n2821 avdd.n2820 0.00807576
R13054 avdd.n3145 avdd.n3142 0.00807576
R13055 avdd.n3128 avdd.n3127 0.00807576
R13056 avdd.n3107 avdd.n3106 0.00807576
R13057 avdd.n3066 avdd.n3062 0.00807576
R13058 avdd.n3052 avdd.n3051 0.00807576
R13059 avdd.n3036 avdd.n3035 0.00807576
R13060 avdd.n3328 avdd.n3291 0.00807576
R13061 avdd.n3337 avdd.n3268 0.00807576
R13062 avdd.n3342 avdd.n3341 0.00807576
R13063 avdd.n3372 avdd.n3176 0.00807576
R13064 avdd.n3227 avdd.n3226 0.00807576
R13065 avdd.n3212 avdd.n3211 0.00807576
R13066 avdd.n3543 avdd.n3506 0.00807576
R13067 avdd.n3552 avdd.n3483 0.00807576
R13068 avdd.n3557 avdd.n3556 0.00807576
R13069 avdd.n3587 avdd.n3391 0.00807576
R13070 avdd.n3442 avdd.n3441 0.00807576
R13071 avdd.n3427 avdd.n3426 0.00807576
R13072 avdd.n3758 avdd.n3721 0.00807576
R13073 avdd.n3767 avdd.n3698 0.00807576
R13074 avdd.n3772 avdd.n3771 0.00807576
R13075 avdd.n3802 avdd.n3606 0.00807576
R13076 avdd.n3657 avdd.n3656 0.00807576
R13077 avdd.n3642 avdd.n3641 0.00807576
R13078 avdd.n3973 avdd.n3936 0.00807576
R13079 avdd.n3982 avdd.n3913 0.00807576
R13080 avdd.n3987 avdd.n3986 0.00807576
R13081 avdd.n4017 avdd.n3821 0.00807576
R13082 avdd.n3872 avdd.n3871 0.00807576
R13083 avdd.n3857 avdd.n3856 0.00807576
R13084 avdd.n4188 avdd.n4151 0.00807576
R13085 avdd.n4197 avdd.n4128 0.00807576
R13086 avdd.n4202 avdd.n4201 0.00807576
R13087 avdd.n4232 avdd.n4036 0.00807576
R13088 avdd.n4087 avdd.n4086 0.00807576
R13089 avdd.n4072 avdd.n4071 0.00807576
R13090 avdd.n4403 avdd.n4366 0.00807576
R13091 avdd.n4412 avdd.n4343 0.00807576
R13092 avdd.n4417 avdd.n4416 0.00807576
R13093 avdd.n4447 avdd.n4251 0.00807576
R13094 avdd.n4302 avdd.n4301 0.00807576
R13095 avdd.n4287 avdd.n4286 0.00807576
R13096 avdd.n4898 avdd.n4897 0.00807576
R13097 avdd.n4915 avdd.n4914 0.00807576
R13098 avdd.n4928 avdd.n4924 0.00807576
R13099 avdd.n4969 avdd.n4968 0.00807576
R13100 avdd.n4990 avdd.n4989 0.00807576
R13101 avdd.n5003 avdd.n5002 0.00807576
R13102 avdd.n5114 avdd.n5113 0.00807576
R13103 avdd.n5131 avdd.n5130 0.00807576
R13104 avdd.n5144 avdd.n5140 0.00807576
R13105 avdd.n5185 avdd.n5184 0.00807576
R13106 avdd.n5206 avdd.n5205 0.00807576
R13107 avdd.n5219 avdd.n5218 0.00807576
R13108 avdd.n5330 avdd.n5329 0.00807576
R13109 avdd.n5347 avdd.n5346 0.00807576
R13110 avdd.n5360 avdd.n5356 0.00807576
R13111 avdd.n5401 avdd.n5400 0.00807576
R13112 avdd.n5422 avdd.n5421 0.00807576
R13113 avdd.n5435 avdd.n5434 0.00807576
R13114 avdd.n5546 avdd.n5545 0.00807576
R13115 avdd.n5563 avdd.n5562 0.00807576
R13116 avdd.n5576 avdd.n5572 0.00807576
R13117 avdd.n5617 avdd.n5616 0.00807576
R13118 avdd.n5638 avdd.n5637 0.00807576
R13119 avdd.n5651 avdd.n5650 0.00807576
R13120 avdd.n5762 avdd.n5761 0.00807576
R13121 avdd.n5779 avdd.n5778 0.00807576
R13122 avdd.n5792 avdd.n5788 0.00807576
R13123 avdd.n5833 avdd.n5832 0.00807576
R13124 avdd.n5854 avdd.n5853 0.00807576
R13125 avdd.n5867 avdd.n5866 0.00807576
R13126 avdd.n5978 avdd.n5977 0.00807576
R13127 avdd.n5995 avdd.n5994 0.00807576
R13128 avdd.n6008 avdd.n6004 0.00807576
R13129 avdd.n6049 avdd.n6048 0.00807576
R13130 avdd.n6070 avdd.n6069 0.00807576
R13131 avdd.n6083 avdd.n6082 0.00807576
R13132 avdd.n6194 avdd.n6193 0.00807576
R13133 avdd.n6211 avdd.n6210 0.00807576
R13134 avdd.n6224 avdd.n6220 0.00807576
R13135 avdd.n6265 avdd.n6264 0.00807576
R13136 avdd.n6286 avdd.n6285 0.00807576
R13137 avdd.n6299 avdd.n6298 0.00807576
R13138 avdd.n6410 avdd.n6409 0.00807576
R13139 avdd.n6427 avdd.n6426 0.00807576
R13140 avdd.n6440 avdd.n6436 0.00807576
R13141 avdd.n6481 avdd.n6480 0.00807576
R13142 avdd.n6502 avdd.n6501 0.00807576
R13143 avdd.n6515 avdd.n6514 0.00807576
R13144 avdd.n6626 avdd.n6625 0.00807576
R13145 avdd.n6643 avdd.n6642 0.00807576
R13146 avdd.n6656 avdd.n6652 0.00807576
R13147 avdd.n6697 avdd.n6696 0.00807576
R13148 avdd.n6718 avdd.n6717 0.00807576
R13149 avdd.n6731 avdd.n6730 0.00807576
R13150 avdd.n6842 avdd.n6841 0.00807576
R13151 avdd.n6859 avdd.n6858 0.00807576
R13152 avdd.n6872 avdd.n6868 0.00807576
R13153 avdd.n6913 avdd.n6912 0.00807576
R13154 avdd.n6934 avdd.n6933 0.00807576
R13155 avdd.n6947 avdd.n6946 0.00807576
R13156 avdd.n7058 avdd.n7057 0.00807576
R13157 avdd.n7075 avdd.n7074 0.00807576
R13158 avdd.n7088 avdd.n7084 0.00807576
R13159 avdd.n7129 avdd.n7128 0.00807576
R13160 avdd.n7150 avdd.n7149 0.00807576
R13161 avdd.n7163 avdd.n7162 0.00807576
R13162 avdd.n7274 avdd.n7273 0.00807576
R13163 avdd.n7291 avdd.n7290 0.00807576
R13164 avdd.n7304 avdd.n7300 0.00807576
R13165 avdd.n7345 avdd.n7344 0.00807576
R13166 avdd.n7366 avdd.n7365 0.00807576
R13167 avdd.n7379 avdd.n7378 0.00807576
R13168 avdd.n7708 avdd.n7707 0.00807576
R13169 avdd.n7727 avdd.n7726 0.00807576
R13170 avdd.n7692 avdd.n7691 0.00807576
R13171 avdd.n7799 avdd.n7798 0.00807576
R13172 avdd.n7817 avdd.n7816 0.00807576
R13173 avdd.n7839 avdd.n7838 0.00807576
R13174 avdd.n10187 avdd.n10186 0.00807576
R13175 avdd.n10206 avdd.n10205 0.00807576
R13176 avdd.n10171 avdd.n10170 0.00807576
R13177 avdd.n10058 avdd.n10057 0.00807576
R13178 avdd.n10075 avdd.n10074 0.00807576
R13179 avdd.n10097 avdd.n10096 0.00807576
R13180 avdd.n9979 avdd.n9978 0.00807576
R13181 avdd.n10012 avdd.n10011 0.00807576
R13182 avdd.n9955 avdd.n9954 0.00807576
R13183 avdd.n10288 avdd.n10287 0.00807576
R13184 avdd.n10307 avdd.n10306 0.00807576
R13185 avdd.n10329 avdd.n10328 0.00807576
R13186 avdd.n9865 avdd.n9864 0.00807576
R13187 avdd.n9898 avdd.n9897 0.00807576
R13188 avdd.n9841 avdd.n9840 0.00807576
R13189 avdd.n10390 avdd.n10389 0.00807576
R13190 avdd.n10409 avdd.n10408 0.00807576
R13191 avdd.n10431 avdd.n10430 0.00807576
R13192 avdd.n9751 avdd.n9750 0.00807576
R13193 avdd.n9784 avdd.n9783 0.00807576
R13194 avdd.n9727 avdd.n9726 0.00807576
R13195 avdd.n10492 avdd.n10491 0.00807576
R13196 avdd.n10511 avdd.n10510 0.00807576
R13197 avdd.n10533 avdd.n10532 0.00807576
R13198 avdd.n9638 avdd.n9637 0.00807576
R13199 avdd.n9671 avdd.n9670 0.00807576
R13200 avdd.n9614 avdd.n9613 0.00807576
R13201 avdd.n10594 avdd.n10593 0.00807576
R13202 avdd.n10613 avdd.n10612 0.00807576
R13203 avdd.n10635 avdd.n10634 0.00807576
R13204 avdd.n9523 avdd.n9522 0.00807576
R13205 avdd.n9556 avdd.n9555 0.00807576
R13206 avdd.n9499 avdd.n9498 0.00807576
R13207 avdd.n10696 avdd.n10695 0.00807576
R13208 avdd.n10715 avdd.n10714 0.00807576
R13209 avdd.n10737 avdd.n10736 0.00807576
R13210 avdd.n9409 avdd.n9408 0.00807576
R13211 avdd.n9442 avdd.n9441 0.00807576
R13212 avdd.n9385 avdd.n9384 0.00807576
R13213 avdd.n10798 avdd.n10797 0.00807576
R13214 avdd.n10817 avdd.n10816 0.00807576
R13215 avdd.n10839 avdd.n10838 0.00807576
R13216 avdd.n9295 avdd.n9294 0.00807576
R13217 avdd.n9328 avdd.n9327 0.00807576
R13218 avdd.n9271 avdd.n9270 0.00807576
R13219 avdd.n10900 avdd.n10899 0.00807576
R13220 avdd.n10919 avdd.n10918 0.00807576
R13221 avdd.n10941 avdd.n10940 0.00807576
R13222 avdd.n9181 avdd.n9180 0.00807576
R13223 avdd.n9214 avdd.n9213 0.00807576
R13224 avdd.n9157 avdd.n9156 0.00807576
R13225 avdd.n11002 avdd.n11001 0.00807576
R13226 avdd.n11021 avdd.n11020 0.00807576
R13227 avdd.n11043 avdd.n11042 0.00807576
R13228 avdd.n9067 avdd.n9066 0.00807576
R13229 avdd.n9100 avdd.n9099 0.00807576
R13230 avdd.n9043 avdd.n9042 0.00807576
R13231 avdd.n11104 avdd.n11103 0.00807576
R13232 avdd.n11123 avdd.n11122 0.00807576
R13233 avdd.n11145 avdd.n11144 0.00807576
R13234 avdd.n8953 avdd.n8952 0.00807576
R13235 avdd.n8986 avdd.n8985 0.00807576
R13236 avdd.n8929 avdd.n8928 0.00807576
R13237 avdd.n11206 avdd.n11205 0.00807576
R13238 avdd.n11225 avdd.n11224 0.00807576
R13239 avdd.n11247 avdd.n11246 0.00807576
R13240 avdd.n8860 avdd.n8859 0.00807576
R13241 avdd.n8838 avdd.n8837 0.00807576
R13242 avdd.n8821 avdd.n8820 0.00807576
R13243 avdd.n175 avdd.n174 0.00807576
R13244 avdd.n122 avdd.n121 0.00807576
R13245 avdd.n102 avdd.n101 0.00807576
R13246 avdd.n8774 avdd.n8773 0.00807576
R13247 avdd.n8752 avdd.n8751 0.00807576
R13248 avdd.n8735 avdd.n8734 0.00807576
R13249 avdd.n305 avdd.n304 0.00807576
R13250 avdd.n252 avdd.n251 0.00807576
R13251 avdd.n232 avdd.n231 0.00807576
R13252 avdd.n8688 avdd.n8687 0.00807576
R13253 avdd.n8666 avdd.n8665 0.00807576
R13254 avdd.n8649 avdd.n8648 0.00807576
R13255 avdd.n435 avdd.n434 0.00807576
R13256 avdd.n382 avdd.n381 0.00807576
R13257 avdd.n362 avdd.n361 0.00807576
R13258 avdd.n8602 avdd.n8601 0.00807576
R13259 avdd.n8580 avdd.n8579 0.00807576
R13260 avdd.n8563 avdd.n8562 0.00807576
R13261 avdd.n565 avdd.n564 0.00807576
R13262 avdd.n512 avdd.n511 0.00807576
R13263 avdd.n492 avdd.n491 0.00807576
R13264 avdd.n8516 avdd.n8515 0.00807576
R13265 avdd.n8494 avdd.n8493 0.00807576
R13266 avdd.n8477 avdd.n8476 0.00807576
R13267 avdd.n695 avdd.n694 0.00807576
R13268 avdd.n642 avdd.n641 0.00807576
R13269 avdd.n622 avdd.n621 0.00807576
R13270 avdd.n8430 avdd.n8429 0.00807576
R13271 avdd.n8408 avdd.n8407 0.00807576
R13272 avdd.n8391 avdd.n8390 0.00807576
R13273 avdd.n825 avdd.n824 0.00807576
R13274 avdd.n772 avdd.n771 0.00807576
R13275 avdd.n752 avdd.n751 0.00807576
R13276 avdd.n8344 avdd.n8343 0.00807576
R13277 avdd.n8322 avdd.n8321 0.00807576
R13278 avdd.n8305 avdd.n8304 0.00807576
R13279 avdd.n955 avdd.n954 0.00807576
R13280 avdd.n902 avdd.n901 0.00807576
R13281 avdd.n882 avdd.n881 0.00807576
R13282 avdd.n8258 avdd.n8257 0.00807576
R13283 avdd.n8236 avdd.n8235 0.00807576
R13284 avdd.n8219 avdd.n8218 0.00807576
R13285 avdd.n1085 avdd.n1084 0.00807576
R13286 avdd.n1032 avdd.n1031 0.00807576
R13287 avdd.n1012 avdd.n1011 0.00807576
R13288 avdd.n8172 avdd.n8171 0.00807576
R13289 avdd.n8150 avdd.n8149 0.00807576
R13290 avdd.n8133 avdd.n8132 0.00807576
R13291 avdd.n1215 avdd.n1214 0.00807576
R13292 avdd.n1162 avdd.n1161 0.00807576
R13293 avdd.n1142 avdd.n1141 0.00807576
R13294 avdd.n8086 avdd.n8085 0.00807576
R13295 avdd.n8064 avdd.n8063 0.00807576
R13296 avdd.n8047 avdd.n8046 0.00807576
R13297 avdd.n1345 avdd.n1344 0.00807576
R13298 avdd.n1292 avdd.n1291 0.00807576
R13299 avdd.n1272 avdd.n1271 0.00807576
R13300 avdd.n8000 avdd.n7999 0.00807576
R13301 avdd.n7978 avdd.n7977 0.00807576
R13302 avdd.n7961 avdd.n7960 0.00807576
R13303 avdd.n1475 avdd.n1474 0.00807576
R13304 avdd.n1422 avdd.n1421 0.00807576
R13305 avdd.n1402 avdd.n1401 0.00807576
R13306 avdd.n7914 avdd.n7913 0.00807576
R13307 avdd.n7892 avdd.n7891 0.00807576
R13308 avdd.n7875 avdd.n7874 0.00807576
R13309 avdd.n1605 avdd.n1604 0.00807576
R13310 avdd.n1552 avdd.n1551 0.00807576
R13311 avdd.n1532 avdd.n1531 0.00807576
R13312 avdd.n1930 avdd.n1894 0.00762121
R13313 avdd.n2080 avdd.n1885 0.00762121
R13314 avdd.n1985 avdd.n1984 0.00762121
R13315 avdd.n2015 avdd.n2003 0.00762121
R13316 avdd.n2183 avdd.n2149 0.00762121
R13317 avdd.n2203 avdd.n2135 0.00762121
R13318 avdd.n2259 avdd.n2112 0.00762121
R13319 avdd.n2288 avdd.n2102 0.00762121
R13320 avdd.n2398 avdd.n2364 0.00762121
R13321 avdd.n2418 avdd.n2350 0.00762121
R13322 avdd.n2474 avdd.n2327 0.00762121
R13323 avdd.n2503 avdd.n2317 0.00762121
R13324 avdd.n2613 avdd.n2579 0.00762121
R13325 avdd.n2633 avdd.n2565 0.00762121
R13326 avdd.n2689 avdd.n2542 0.00762121
R13327 avdd.n2718 avdd.n2532 0.00762121
R13328 avdd.n2828 avdd.n2794 0.00762121
R13329 avdd.n2848 avdd.n2780 0.00762121
R13330 avdd.n2904 avdd.n2757 0.00762121
R13331 avdd.n2933 avdd.n2747 0.00762121
R13332 avdd.n3043 avdd.n3009 0.00762121
R13333 avdd.n3063 avdd.n2995 0.00762121
R13334 avdd.n3119 avdd.n2972 0.00762121
R13335 avdd.n3148 avdd.n2962 0.00762121
R13336 avdd.n3220 avdd.n3184 0.00762121
R13337 avdd.n3369 avdd.n3175 0.00762121
R13338 avdd.n3275 avdd.n3274 0.00762121
R13339 avdd.n3308 avdd.n3293 0.00762121
R13340 avdd.n3435 avdd.n3399 0.00762121
R13341 avdd.n3584 avdd.n3390 0.00762121
R13342 avdd.n3490 avdd.n3489 0.00762121
R13343 avdd.n3523 avdd.n3508 0.00762121
R13344 avdd.n3650 avdd.n3614 0.00762121
R13345 avdd.n3799 avdd.n3605 0.00762121
R13346 avdd.n3705 avdd.n3704 0.00762121
R13347 avdd.n3738 avdd.n3723 0.00762121
R13348 avdd.n3865 avdd.n3829 0.00762121
R13349 avdd.n4014 avdd.n3820 0.00762121
R13350 avdd.n3920 avdd.n3919 0.00762121
R13351 avdd.n3953 avdd.n3938 0.00762121
R13352 avdd.n4080 avdd.n4044 0.00762121
R13353 avdd.n4229 avdd.n4035 0.00762121
R13354 avdd.n4135 avdd.n4134 0.00762121
R13355 avdd.n4168 avdd.n4153 0.00762121
R13356 avdd.n4295 avdd.n4259 0.00762121
R13357 avdd.n4444 avdd.n4250 0.00762121
R13358 avdd.n4350 avdd.n4349 0.00762121
R13359 avdd.n4383 avdd.n4368 0.00762121
R13360 avdd.n4906 avdd.n4871 0.00762121
R13361 avdd.n4925 avdd.n4857 0.00762121
R13362 avdd.n4981 avdd.n4834 0.00762121
R13363 avdd.n5006 avdd.n4823 0.00762121
R13364 avdd.n5122 avdd.n5087 0.00762121
R13365 avdd.n5141 avdd.n5073 0.00762121
R13366 avdd.n5197 avdd.n5050 0.00762121
R13367 avdd.n5222 avdd.n5039 0.00762121
R13368 avdd.n5338 avdd.n5303 0.00762121
R13369 avdd.n5357 avdd.n5289 0.00762121
R13370 avdd.n5413 avdd.n5266 0.00762121
R13371 avdd.n5438 avdd.n5255 0.00762121
R13372 avdd.n5554 avdd.n5519 0.00762121
R13373 avdd.n5573 avdd.n5505 0.00762121
R13374 avdd.n5629 avdd.n5482 0.00762121
R13375 avdd.n5654 avdd.n5471 0.00762121
R13376 avdd.n5770 avdd.n5735 0.00762121
R13377 avdd.n5789 avdd.n5721 0.00762121
R13378 avdd.n5845 avdd.n5698 0.00762121
R13379 avdd.n5870 avdd.n5687 0.00762121
R13380 avdd.n5986 avdd.n5951 0.00762121
R13381 avdd.n6005 avdd.n5937 0.00762121
R13382 avdd.n6061 avdd.n5914 0.00762121
R13383 avdd.n6086 avdd.n5903 0.00762121
R13384 avdd.n6202 avdd.n6167 0.00762121
R13385 avdd.n6221 avdd.n6153 0.00762121
R13386 avdd.n6277 avdd.n6130 0.00762121
R13387 avdd.n6302 avdd.n6119 0.00762121
R13388 avdd.n6418 avdd.n6383 0.00762121
R13389 avdd.n6437 avdd.n6369 0.00762121
R13390 avdd.n6493 avdd.n6346 0.00762121
R13391 avdd.n6518 avdd.n6335 0.00762121
R13392 avdd.n6634 avdd.n6599 0.00762121
R13393 avdd.n6653 avdd.n6585 0.00762121
R13394 avdd.n6709 avdd.n6562 0.00762121
R13395 avdd.n6734 avdd.n6551 0.00762121
R13396 avdd.n6850 avdd.n6815 0.00762121
R13397 avdd.n6869 avdd.n6801 0.00762121
R13398 avdd.n6925 avdd.n6778 0.00762121
R13399 avdd.n6950 avdd.n6767 0.00762121
R13400 avdd.n7066 avdd.n7031 0.00762121
R13401 avdd.n7085 avdd.n7017 0.00762121
R13402 avdd.n7141 avdd.n6994 0.00762121
R13403 avdd.n7166 avdd.n6983 0.00762121
R13404 avdd.n7282 avdd.n7247 0.00762121
R13405 avdd.n7301 avdd.n7233 0.00762121
R13406 avdd.n7357 avdd.n7210 0.00762121
R13407 avdd.n7382 avdd.n7199 0.00762121
R13408 avdd.n7718 avdd.n7717 0.00762121
R13409 avdd.n7697 avdd.n7687 0.00762121
R13410 avdd.n7807 avdd.n7806 0.00762121
R13411 avdd.n7845 avdd.n7844 0.00762121
R13412 avdd.n10197 avdd.n10196 0.00762121
R13413 avdd.n10176 avdd.n10166 0.00762121
R13414 avdd.n10065 avdd.n10064 0.00762121
R13415 avdd.n10103 avdd.n10102 0.00762121
R13416 avdd.n10001 avdd.n10000 0.00762121
R13417 avdd.n9960 avdd.n9950 0.00762121
R13418 avdd.n10297 avdd.n10296 0.00762121
R13419 avdd.n10335 avdd.n10334 0.00762121
R13420 avdd.n9887 avdd.n9886 0.00762121
R13421 avdd.n9846 avdd.n9836 0.00762121
R13422 avdd.n10399 avdd.n10398 0.00762121
R13423 avdd.n10437 avdd.n10436 0.00762121
R13424 avdd.n9773 avdd.n9772 0.00762121
R13425 avdd.n9732 avdd.n9722 0.00762121
R13426 avdd.n10501 avdd.n10500 0.00762121
R13427 avdd.n10539 avdd.n10538 0.00762121
R13428 avdd.n9660 avdd.n9659 0.00762121
R13429 avdd.n9619 avdd.n9609 0.00762121
R13430 avdd.n10603 avdd.n10602 0.00762121
R13431 avdd.n10641 avdd.n10640 0.00762121
R13432 avdd.n9545 avdd.n9544 0.00762121
R13433 avdd.n9504 avdd.n9494 0.00762121
R13434 avdd.n10705 avdd.n10704 0.00762121
R13435 avdd.n10743 avdd.n10742 0.00762121
R13436 avdd.n9431 avdd.n9430 0.00762121
R13437 avdd.n9390 avdd.n9380 0.00762121
R13438 avdd.n10807 avdd.n10806 0.00762121
R13439 avdd.n10845 avdd.n10844 0.00762121
R13440 avdd.n9317 avdd.n9316 0.00762121
R13441 avdd.n9276 avdd.n9266 0.00762121
R13442 avdd.n10909 avdd.n10908 0.00762121
R13443 avdd.n10947 avdd.n10946 0.00762121
R13444 avdd.n9203 avdd.n9202 0.00762121
R13445 avdd.n9162 avdd.n9152 0.00762121
R13446 avdd.n11011 avdd.n11010 0.00762121
R13447 avdd.n11049 avdd.n11048 0.00762121
R13448 avdd.n9089 avdd.n9088 0.00762121
R13449 avdd.n9048 avdd.n9038 0.00762121
R13450 avdd.n11113 avdd.n11112 0.00762121
R13451 avdd.n11151 avdd.n11150 0.00762121
R13452 avdd.n8975 avdd.n8974 0.00762121
R13453 avdd.n8934 avdd.n8924 0.00762121
R13454 avdd.n11215 avdd.n11214 0.00762121
R13455 avdd.n11253 avdd.n11252 0.00762121
R13456 avdd.n112 avdd.n111 0.00762121
R13457 avdd.n180 avdd.n170 0.00762121
R13458 avdd.n8828 avdd.n8827 0.00762121
R13459 avdd.n8866 avdd.n8865 0.00762121
R13460 avdd.n242 avdd.n241 0.00762121
R13461 avdd.n310 avdd.n300 0.00762121
R13462 avdd.n8742 avdd.n8741 0.00762121
R13463 avdd.n8780 avdd.n8779 0.00762121
R13464 avdd.n372 avdd.n371 0.00762121
R13465 avdd.n440 avdd.n430 0.00762121
R13466 avdd.n8656 avdd.n8655 0.00762121
R13467 avdd.n8694 avdd.n8693 0.00762121
R13468 avdd.n502 avdd.n501 0.00762121
R13469 avdd.n570 avdd.n560 0.00762121
R13470 avdd.n8570 avdd.n8569 0.00762121
R13471 avdd.n8608 avdd.n8607 0.00762121
R13472 avdd.n632 avdd.n631 0.00762121
R13473 avdd.n700 avdd.n690 0.00762121
R13474 avdd.n8484 avdd.n8483 0.00762121
R13475 avdd.n8522 avdd.n8521 0.00762121
R13476 avdd.n762 avdd.n761 0.00762121
R13477 avdd.n830 avdd.n820 0.00762121
R13478 avdd.n8398 avdd.n8397 0.00762121
R13479 avdd.n8436 avdd.n8435 0.00762121
R13480 avdd.n892 avdd.n891 0.00762121
R13481 avdd.n960 avdd.n950 0.00762121
R13482 avdd.n8312 avdd.n8311 0.00762121
R13483 avdd.n8350 avdd.n8349 0.00762121
R13484 avdd.n1022 avdd.n1021 0.00762121
R13485 avdd.n1090 avdd.n1080 0.00762121
R13486 avdd.n8226 avdd.n8225 0.00762121
R13487 avdd.n8264 avdd.n8263 0.00762121
R13488 avdd.n1152 avdd.n1151 0.00762121
R13489 avdd.n1220 avdd.n1210 0.00762121
R13490 avdd.n8140 avdd.n8139 0.00762121
R13491 avdd.n8178 avdd.n8177 0.00762121
R13492 avdd.n1282 avdd.n1281 0.00762121
R13493 avdd.n1350 avdd.n1340 0.00762121
R13494 avdd.n8054 avdd.n8053 0.00762121
R13495 avdd.n8092 avdd.n8091 0.00762121
R13496 avdd.n1412 avdd.n1411 0.00762121
R13497 avdd.n1480 avdd.n1470 0.00762121
R13498 avdd.n7968 avdd.n7967 0.00762121
R13499 avdd.n8006 avdd.n8005 0.00762121
R13500 avdd.n1542 avdd.n1541 0.00762121
R13501 avdd.n1610 avdd.n1600 0.00762121
R13502 avdd.n7882 avdd.n7881 0.00762121
R13503 avdd.n7920 avdd.n7919 0.00762121
R13504 avdd.n2071 avdd.n2070 0.00690909
R13505 avdd.n2072 avdd.n1950 0.00690909
R13506 avdd.n2029 avdd.n2009 0.00690909
R13507 avdd.n2228 avdd.n2122 0.00690909
R13508 avdd.n2227 avdd.n2123 0.00690909
R13509 avdd.n2304 avdd.n2301 0.00690909
R13510 avdd.n2443 avdd.n2337 0.00690909
R13511 avdd.n2442 avdd.n2338 0.00690909
R13512 avdd.n2519 avdd.n2516 0.00690909
R13513 avdd.n2658 avdd.n2552 0.00690909
R13514 avdd.n2657 avdd.n2553 0.00690909
R13515 avdd.n2734 avdd.n2731 0.00690909
R13516 avdd.n2873 avdd.n2767 0.00690909
R13517 avdd.n2872 avdd.n2768 0.00690909
R13518 avdd.n2949 avdd.n2946 0.00690909
R13519 avdd.n3088 avdd.n2982 0.00690909
R13520 avdd.n3087 avdd.n2983 0.00690909
R13521 avdd.n3164 avdd.n3161 0.00690909
R13522 avdd.n3360 avdd.n3359 0.00690909
R13523 avdd.n3361 avdd.n3240 0.00690909
R13524 avdd.n3575 avdd.n3574 0.00690909
R13525 avdd.n3576 avdd.n3455 0.00690909
R13526 avdd.n3790 avdd.n3789 0.00690909
R13527 avdd.n3791 avdd.n3670 0.00690909
R13528 avdd.n4005 avdd.n4004 0.00690909
R13529 avdd.n4006 avdd.n3885 0.00690909
R13530 avdd.n4220 avdd.n4219 0.00690909
R13531 avdd.n4221 avdd.n4100 0.00690909
R13532 avdd.n4435 avdd.n4434 0.00690909
R13533 avdd.n4436 avdd.n4315 0.00690909
R13534 avdd.n4950 avdd.n4844 0.00690909
R13535 avdd.n4949 avdd.n4845 0.00690909
R13536 avdd.n5166 avdd.n5060 0.00690909
R13537 avdd.n5165 avdd.n5061 0.00690909
R13538 avdd.n5382 avdd.n5276 0.00690909
R13539 avdd.n5381 avdd.n5277 0.00690909
R13540 avdd.n5598 avdd.n5492 0.00690909
R13541 avdd.n5597 avdd.n5493 0.00690909
R13542 avdd.n5814 avdd.n5708 0.00690909
R13543 avdd.n5813 avdd.n5709 0.00690909
R13544 avdd.n6030 avdd.n5924 0.00690909
R13545 avdd.n6029 avdd.n5925 0.00690909
R13546 avdd.n6246 avdd.n6140 0.00690909
R13547 avdd.n6245 avdd.n6141 0.00690909
R13548 avdd.n6462 avdd.n6356 0.00690909
R13549 avdd.n6461 avdd.n6357 0.00690909
R13550 avdd.n6678 avdd.n6572 0.00690909
R13551 avdd.n6677 avdd.n6573 0.00690909
R13552 avdd.n6894 avdd.n6788 0.00690909
R13553 avdd.n6893 avdd.n6789 0.00690909
R13554 avdd.n7110 avdd.n7004 0.00690909
R13555 avdd.n7109 avdd.n7005 0.00690909
R13556 avdd.n7326 avdd.n7220 0.00690909
R13557 avdd.n7325 avdd.n7221 0.00690909
R13558 avdd.n7644 avdd.n7643 0.00690909
R13559 avdd.n7679 avdd.n7678 0.00690909
R13560 avdd.n7792 avdd.n7791 0.00690909
R13561 avdd.n10121 avdd.n10120 0.00690909
R13562 avdd.n10158 avdd.n10157 0.00690909
R13563 avdd.n10052 avdd.n10051 0.00690909
R13564 avdd.n9922 avdd.n9921 0.00690909
R13565 avdd.n9942 avdd.n9941 0.00690909
R13566 avdd.n9808 avdd.n9807 0.00690909
R13567 avdd.n9828 avdd.n9827 0.00690909
R13568 avdd.n9694 avdd.n9693 0.00690909
R13569 avdd.n9714 avdd.n9713 0.00690909
R13570 avdd.n9580 avdd.n9579 0.00690909
R13571 avdd.n9601 avdd.n9600 0.00690909
R13572 avdd.n9466 avdd.n9465 0.00690909
R13573 avdd.n9486 avdd.n9485 0.00690909
R13574 avdd.n9352 avdd.n9351 0.00690909
R13575 avdd.n9372 avdd.n9371 0.00690909
R13576 avdd.n9238 avdd.n9237 0.00690909
R13577 avdd.n9258 avdd.n9257 0.00690909
R13578 avdd.n9124 avdd.n9123 0.00690909
R13579 avdd.n9144 avdd.n9143 0.00690909
R13580 avdd.n9010 avdd.n9009 0.00690909
R13581 avdd.n9030 avdd.n9029 0.00690909
R13582 avdd.n8896 avdd.n8895 0.00690909
R13583 avdd.n8916 avdd.n8915 0.00690909
R13584 avdd.n65 avdd.n64 0.00690909
R13585 avdd.n162 avdd.n161 0.00690909
R13586 avdd.n8815 avdd.n8814 0.00690909
R13587 avdd.n195 avdd.n194 0.00690909
R13588 avdd.n292 avdd.n291 0.00690909
R13589 avdd.n8729 avdd.n8728 0.00690909
R13590 avdd.n325 avdd.n324 0.00690909
R13591 avdd.n422 avdd.n421 0.00690909
R13592 avdd.n8643 avdd.n8642 0.00690909
R13593 avdd.n455 avdd.n454 0.00690909
R13594 avdd.n552 avdd.n551 0.00690909
R13595 avdd.n8557 avdd.n8556 0.00690909
R13596 avdd.n585 avdd.n584 0.00690909
R13597 avdd.n682 avdd.n681 0.00690909
R13598 avdd.n8471 avdd.n8470 0.00690909
R13599 avdd.n715 avdd.n714 0.00690909
R13600 avdd.n812 avdd.n811 0.00690909
R13601 avdd.n8385 avdd.n8384 0.00690909
R13602 avdd.n845 avdd.n844 0.00690909
R13603 avdd.n942 avdd.n941 0.00690909
R13604 avdd.n8299 avdd.n8298 0.00690909
R13605 avdd.n975 avdd.n974 0.00690909
R13606 avdd.n1072 avdd.n1071 0.00690909
R13607 avdd.n8213 avdd.n8212 0.00690909
R13608 avdd.n1105 avdd.n1104 0.00690909
R13609 avdd.n1202 avdd.n1201 0.00690909
R13610 avdd.n8127 avdd.n8126 0.00690909
R13611 avdd.n1235 avdd.n1234 0.00690909
R13612 avdd.n1332 avdd.n1331 0.00690909
R13613 avdd.n8041 avdd.n8040 0.00690909
R13614 avdd.n1365 avdd.n1364 0.00690909
R13615 avdd.n1462 avdd.n1461 0.00690909
R13616 avdd.n7955 avdd.n7954 0.00690909
R13617 avdd.n1495 avdd.n1494 0.00690909
R13618 avdd.n1592 avdd.n1591 0.00690909
R13619 avdd.n7869 avdd.n7868 0.00690909
R13620 avdd.n2006 avdd.n2002 0.00633256
R13621 avdd.n2272 avdd.n2095 0.00633256
R13622 avdd.n2487 avdd.n2310 0.00633256
R13623 avdd.n2702 avdd.n2525 0.00633256
R13624 avdd.n2917 avdd.n2740 0.00633256
R13625 avdd.n3132 avdd.n2955 0.00633256
R13626 avdd.n3304 avdd.n3292 0.00633256
R13627 avdd.n3519 avdd.n3507 0.00633256
R13628 avdd.n3734 avdd.n3722 0.00633256
R13629 avdd.n3949 avdd.n3937 0.00633256
R13630 avdd.n4164 avdd.n4152 0.00633256
R13631 avdd.n4379 avdd.n4367 0.00633256
R13632 avdd.n7832 avdd.n7831 0.00633256
R13633 avdd.n10090 avdd.n10089 0.00633256
R13634 avdd.n8853 avdd.n8852 0.00633256
R13635 avdd.n8767 avdd.n8766 0.00633256
R13636 avdd.n8681 avdd.n8680 0.00633256
R13637 avdd.n8595 avdd.n8594 0.00633256
R13638 avdd.n8509 avdd.n8508 0.00633256
R13639 avdd.n8423 avdd.n8422 0.00633256
R13640 avdd.n8337 avdd.n8336 0.00633256
R13641 avdd.n8251 avdd.n8250 0.00633256
R13642 avdd.n8165 avdd.n8164 0.00633256
R13643 avdd.n8079 avdd.n8078 0.00633256
R13644 avdd.n7993 avdd.n7992 0.00633256
R13645 avdd.n7907 avdd.n7906 0.00633256
R13646 avdd.n2022 avdd.n2021 0.00585759
R13647 avdd.n2298 avdd.n2295 0.00585759
R13648 avdd.n2513 avdd.n2510 0.00585759
R13649 avdd.n2728 avdd.n2725 0.00585759
R13650 avdd.n2943 avdd.n2940 0.00585759
R13651 avdd.n3158 avdd.n3155 0.00585759
R13652 avdd.n3316 avdd.n3315 0.00585759
R13653 avdd.n3531 avdd.n3530 0.00585759
R13654 avdd.n3746 avdd.n3745 0.00585759
R13655 avdd.n3961 avdd.n3960 0.00585759
R13656 avdd.n4176 avdd.n4175 0.00585759
R13657 avdd.n4391 avdd.n4390 0.00585759
R13658 avdd.n8811 avdd.n8810 0.00585759
R13659 avdd.n8725 avdd.n8724 0.00585759
R13660 avdd.n8639 avdd.n8638 0.00585759
R13661 avdd.n8553 avdd.n8552 0.00585759
R13662 avdd.n8467 avdd.n8466 0.00585759
R13663 avdd.n8381 avdd.n8380 0.00585759
R13664 avdd.n8295 avdd.n8294 0.00585759
R13665 avdd.n8209 avdd.n8208 0.00585759
R13666 avdd.n8123 avdd.n8122 0.00585759
R13667 avdd.n8037 avdd.n8036 0.00585759
R13668 avdd.n7951 avdd.n7950 0.00585759
R13669 avdd.n7865 avdd.n7864 0.00585759
R13670 avdd.n5019 avdd.n5018 0.00585698
R13671 avdd.n5235 avdd.n5234 0.00585698
R13672 avdd.n5451 avdd.n5450 0.00585698
R13673 avdd.n5667 avdd.n5666 0.00585698
R13674 avdd.n5883 avdd.n5882 0.00585698
R13675 avdd.n6099 avdd.n6098 0.00585698
R13676 avdd.n6315 avdd.n6314 0.00585698
R13677 avdd.n6531 avdd.n6530 0.00585698
R13678 avdd.n6747 avdd.n6746 0.00585698
R13679 avdd.n6963 avdd.n6962 0.00585698
R13680 avdd.n7179 avdd.n7178 0.00585698
R13681 avdd.n7395 avdd.n7394 0.00585698
R13682 avdd.n7788 avdd.n7787 0.00585698
R13683 avdd.n10048 avdd.n10047 0.00585698
R13684 avdd.n10264 avdd.n10263 0.00585698
R13685 avdd.n10366 avdd.n10365 0.00585698
R13686 avdd.n10468 avdd.n10467 0.00585698
R13687 avdd.n10570 avdd.n10569 0.00585698
R13688 avdd.n10672 avdd.n10671 0.00585698
R13689 avdd.n10774 avdd.n10773 0.00585698
R13690 avdd.n10876 avdd.n10875 0.00585698
R13691 avdd.n10978 avdd.n10977 0.00585698
R13692 avdd.n11080 avdd.n11079 0.00585698
R13693 avdd.n11182 avdd.n11181 0.00585698
R13694 avdd.n1993 avdd.n1992 0.00548485
R13695 avdd.n1919 avdd.n1894 0.00548485
R13696 avdd.n2080 avdd.n2079 0.00548485
R13697 avdd.n1984 avdd.n1982 0.00548485
R13698 avdd.n1991 avdd.n1979 0.00548485
R13699 avdd.n2016 avdd.n2015 0.00548485
R13700 avdd.n2252 avdd.n2107 0.00548485
R13701 avdd.n2173 avdd.n2149 0.00548485
R13702 avdd.n2203 avdd.n2131 0.00548485
R13703 avdd.n2244 avdd.n2112 0.00548485
R13704 avdd.n2253 avdd.n2108 0.00548485
R13705 avdd.n2289 avdd.n2288 0.00548485
R13706 avdd.n2467 avdd.n2322 0.00548485
R13707 avdd.n2388 avdd.n2364 0.00548485
R13708 avdd.n2418 avdd.n2346 0.00548485
R13709 avdd.n2459 avdd.n2327 0.00548485
R13710 avdd.n2468 avdd.n2323 0.00548485
R13711 avdd.n2504 avdd.n2503 0.00548485
R13712 avdd.n2682 avdd.n2537 0.00548485
R13713 avdd.n2603 avdd.n2579 0.00548485
R13714 avdd.n2633 avdd.n2561 0.00548485
R13715 avdd.n2674 avdd.n2542 0.00548485
R13716 avdd.n2683 avdd.n2538 0.00548485
R13717 avdd.n2719 avdd.n2718 0.00548485
R13718 avdd.n2897 avdd.n2752 0.00548485
R13719 avdd.n2818 avdd.n2794 0.00548485
R13720 avdd.n2848 avdd.n2776 0.00548485
R13721 avdd.n2889 avdd.n2757 0.00548485
R13722 avdd.n2898 avdd.n2753 0.00548485
R13723 avdd.n2934 avdd.n2933 0.00548485
R13724 avdd.n3112 avdd.n2967 0.00548485
R13725 avdd.n3033 avdd.n3009 0.00548485
R13726 avdd.n3063 avdd.n2991 0.00548485
R13727 avdd.n3104 avdd.n2972 0.00548485
R13728 avdd.n3113 avdd.n2968 0.00548485
R13729 avdd.n3149 avdd.n3148 0.00548485
R13730 avdd.n3283 avdd.n3282 0.00548485
R13731 avdd.n3209 avdd.n3184 0.00548485
R13732 avdd.n3369 avdd.n3368 0.00548485
R13733 avdd.n3274 avdd.n3272 0.00548485
R13734 avdd.n3281 avdd.n3269 0.00548485
R13735 avdd.n3309 avdd.n3308 0.00548485
R13736 avdd.n3498 avdd.n3497 0.00548485
R13737 avdd.n3424 avdd.n3399 0.00548485
R13738 avdd.n3584 avdd.n3583 0.00548485
R13739 avdd.n3489 avdd.n3487 0.00548485
R13740 avdd.n3496 avdd.n3484 0.00548485
R13741 avdd.n3524 avdd.n3523 0.00548485
R13742 avdd.n3713 avdd.n3712 0.00548485
R13743 avdd.n3639 avdd.n3614 0.00548485
R13744 avdd.n3799 avdd.n3798 0.00548485
R13745 avdd.n3704 avdd.n3702 0.00548485
R13746 avdd.n3711 avdd.n3699 0.00548485
R13747 avdd.n3739 avdd.n3738 0.00548485
R13748 avdd.n3928 avdd.n3927 0.00548485
R13749 avdd.n3854 avdd.n3829 0.00548485
R13750 avdd.n4014 avdd.n4013 0.00548485
R13751 avdd.n3919 avdd.n3917 0.00548485
R13752 avdd.n3926 avdd.n3914 0.00548485
R13753 avdd.n3954 avdd.n3953 0.00548485
R13754 avdd.n4143 avdd.n4142 0.00548485
R13755 avdd.n4069 avdd.n4044 0.00548485
R13756 avdd.n4229 avdd.n4228 0.00548485
R13757 avdd.n4134 avdd.n4132 0.00548485
R13758 avdd.n4141 avdd.n4129 0.00548485
R13759 avdd.n4169 avdd.n4168 0.00548485
R13760 avdd.n4358 avdd.n4357 0.00548485
R13761 avdd.n4284 avdd.n4259 0.00548485
R13762 avdd.n4444 avdd.n4443 0.00548485
R13763 avdd.n4349 avdd.n4347 0.00548485
R13764 avdd.n4356 avdd.n4344 0.00548485
R13765 avdd.n4384 avdd.n4383 0.00548485
R13766 avdd.n4974 avdd.n4829 0.00548485
R13767 avdd.n4895 avdd.n4871 0.00548485
R13768 avdd.n4925 avdd.n4853 0.00548485
R13769 avdd.n4966 avdd.n4834 0.00548485
R13770 avdd.n4975 avdd.n4830 0.00548485
R13771 avdd.n5007 avdd.n5006 0.00548485
R13772 avdd.n5190 avdd.n5045 0.00548485
R13773 avdd.n5111 avdd.n5087 0.00548485
R13774 avdd.n5141 avdd.n5069 0.00548485
R13775 avdd.n5182 avdd.n5050 0.00548485
R13776 avdd.n5191 avdd.n5046 0.00548485
R13777 avdd.n5223 avdd.n5222 0.00548485
R13778 avdd.n5406 avdd.n5261 0.00548485
R13779 avdd.n5327 avdd.n5303 0.00548485
R13780 avdd.n5357 avdd.n5285 0.00548485
R13781 avdd.n5398 avdd.n5266 0.00548485
R13782 avdd.n5407 avdd.n5262 0.00548485
R13783 avdd.n5439 avdd.n5438 0.00548485
R13784 avdd.n5622 avdd.n5477 0.00548485
R13785 avdd.n5543 avdd.n5519 0.00548485
R13786 avdd.n5573 avdd.n5501 0.00548485
R13787 avdd.n5614 avdd.n5482 0.00548485
R13788 avdd.n5623 avdd.n5478 0.00548485
R13789 avdd.n5655 avdd.n5654 0.00548485
R13790 avdd.n5838 avdd.n5693 0.00548485
R13791 avdd.n5759 avdd.n5735 0.00548485
R13792 avdd.n5789 avdd.n5717 0.00548485
R13793 avdd.n5830 avdd.n5698 0.00548485
R13794 avdd.n5839 avdd.n5694 0.00548485
R13795 avdd.n5871 avdd.n5870 0.00548485
R13796 avdd.n6054 avdd.n5909 0.00548485
R13797 avdd.n5975 avdd.n5951 0.00548485
R13798 avdd.n6005 avdd.n5933 0.00548485
R13799 avdd.n6046 avdd.n5914 0.00548485
R13800 avdd.n6055 avdd.n5910 0.00548485
R13801 avdd.n6087 avdd.n6086 0.00548485
R13802 avdd.n6270 avdd.n6125 0.00548485
R13803 avdd.n6191 avdd.n6167 0.00548485
R13804 avdd.n6221 avdd.n6149 0.00548485
R13805 avdd.n6262 avdd.n6130 0.00548485
R13806 avdd.n6271 avdd.n6126 0.00548485
R13807 avdd.n6303 avdd.n6302 0.00548485
R13808 avdd.n6486 avdd.n6341 0.00548485
R13809 avdd.n6407 avdd.n6383 0.00548485
R13810 avdd.n6437 avdd.n6365 0.00548485
R13811 avdd.n6478 avdd.n6346 0.00548485
R13812 avdd.n6487 avdd.n6342 0.00548485
R13813 avdd.n6519 avdd.n6518 0.00548485
R13814 avdd.n6702 avdd.n6557 0.00548485
R13815 avdd.n6623 avdd.n6599 0.00548485
R13816 avdd.n6653 avdd.n6581 0.00548485
R13817 avdd.n6694 avdd.n6562 0.00548485
R13818 avdd.n6703 avdd.n6558 0.00548485
R13819 avdd.n6735 avdd.n6734 0.00548485
R13820 avdd.n6918 avdd.n6773 0.00548485
R13821 avdd.n6839 avdd.n6815 0.00548485
R13822 avdd.n6869 avdd.n6797 0.00548485
R13823 avdd.n6910 avdd.n6778 0.00548485
R13824 avdd.n6919 avdd.n6774 0.00548485
R13825 avdd.n6951 avdd.n6950 0.00548485
R13826 avdd.n7134 avdd.n6989 0.00548485
R13827 avdd.n7055 avdd.n7031 0.00548485
R13828 avdd.n7085 avdd.n7013 0.00548485
R13829 avdd.n7126 avdd.n6994 0.00548485
R13830 avdd.n7135 avdd.n6990 0.00548485
R13831 avdd.n7167 avdd.n7166 0.00548485
R13832 avdd.n7350 avdd.n7205 0.00548485
R13833 avdd.n7271 avdd.n7247 0.00548485
R13834 avdd.n7301 avdd.n7229 0.00548485
R13835 avdd.n7342 avdd.n7210 0.00548485
R13836 avdd.n7351 avdd.n7206 0.00548485
R13837 avdd.n7383 avdd.n7382 0.00548485
R13838 avdd.n7776 avdd.n7775 0.00548485
R13839 avdd.n7717 avdd.n7716 0.00548485
R13840 avdd.n7687 avdd.n7686 0.00548485
R13841 avdd.n7806 avdd.n7805 0.00548485
R13842 avdd.n7812 avdd.n7811 0.00548485
R13843 avdd.n7846 avdd.n7845 0.00548485
R13844 avdd.n10036 avdd.n10035 0.00548485
R13845 avdd.n10196 avdd.n10195 0.00548485
R13846 avdd.n10166 avdd.n10165 0.00548485
R13847 avdd.n10064 avdd.n10063 0.00548485
R13848 avdd.n10070 avdd.n10069 0.00548485
R13849 avdd.n10104 avdd.n10103 0.00548485
R13850 avdd.n10252 avdd.n10251 0.00548485
R13851 avdd.n10000 avdd.n9999 0.00548485
R13852 avdd.n9950 avdd.n9949 0.00548485
R13853 avdd.n10296 avdd.n10295 0.00548485
R13854 avdd.n10302 avdd.n10301 0.00548485
R13855 avdd.n10336 avdd.n10335 0.00548485
R13856 avdd.n10354 avdd.n10353 0.00548485
R13857 avdd.n9886 avdd.n9885 0.00548485
R13858 avdd.n9836 avdd.n9835 0.00548485
R13859 avdd.n10398 avdd.n10397 0.00548485
R13860 avdd.n10404 avdd.n10403 0.00548485
R13861 avdd.n10438 avdd.n10437 0.00548485
R13862 avdd.n10456 avdd.n10455 0.00548485
R13863 avdd.n9772 avdd.n9771 0.00548485
R13864 avdd.n9722 avdd.n9721 0.00548485
R13865 avdd.n10500 avdd.n10499 0.00548485
R13866 avdd.n10506 avdd.n10505 0.00548485
R13867 avdd.n10540 avdd.n10539 0.00548485
R13868 avdd.n10558 avdd.n10557 0.00548485
R13869 avdd.n9659 avdd.n9658 0.00548485
R13870 avdd.n9609 avdd.n9608 0.00548485
R13871 avdd.n10602 avdd.n10601 0.00548485
R13872 avdd.n10608 avdd.n10607 0.00548485
R13873 avdd.n10642 avdd.n10641 0.00548485
R13874 avdd.n10660 avdd.n10659 0.00548485
R13875 avdd.n9544 avdd.n9543 0.00548485
R13876 avdd.n9494 avdd.n9493 0.00548485
R13877 avdd.n10704 avdd.n10703 0.00548485
R13878 avdd.n10710 avdd.n10709 0.00548485
R13879 avdd.n10744 avdd.n10743 0.00548485
R13880 avdd.n10762 avdd.n10761 0.00548485
R13881 avdd.n9430 avdd.n9429 0.00548485
R13882 avdd.n9380 avdd.n9379 0.00548485
R13883 avdd.n10806 avdd.n10805 0.00548485
R13884 avdd.n10812 avdd.n10811 0.00548485
R13885 avdd.n10846 avdd.n10845 0.00548485
R13886 avdd.n10864 avdd.n10863 0.00548485
R13887 avdd.n9316 avdd.n9315 0.00548485
R13888 avdd.n9266 avdd.n9265 0.00548485
R13889 avdd.n10908 avdd.n10907 0.00548485
R13890 avdd.n10914 avdd.n10913 0.00548485
R13891 avdd.n10948 avdd.n10947 0.00548485
R13892 avdd.n10966 avdd.n10965 0.00548485
R13893 avdd.n9202 avdd.n9201 0.00548485
R13894 avdd.n9152 avdd.n9151 0.00548485
R13895 avdd.n11010 avdd.n11009 0.00548485
R13896 avdd.n11016 avdd.n11015 0.00548485
R13897 avdd.n11050 avdd.n11049 0.00548485
R13898 avdd.n11068 avdd.n11067 0.00548485
R13899 avdd.n9088 avdd.n9087 0.00548485
R13900 avdd.n9038 avdd.n9037 0.00548485
R13901 avdd.n11112 avdd.n11111 0.00548485
R13902 avdd.n11118 avdd.n11117 0.00548485
R13903 avdd.n11152 avdd.n11151 0.00548485
R13904 avdd.n11170 avdd.n11169 0.00548485
R13905 avdd.n8974 avdd.n8973 0.00548485
R13906 avdd.n8924 avdd.n8923 0.00548485
R13907 avdd.n11214 avdd.n11213 0.00548485
R13908 avdd.n11220 avdd.n11219 0.00548485
R13909 avdd.n11254 avdd.n11253 0.00548485
R13910 avdd.n8879 avdd.n8878 0.00548485
R13911 avdd.n111 avdd.n110 0.00548485
R13912 avdd.n170 avdd.n169 0.00548485
R13913 avdd.n8827 avdd.n8826 0.00548485
R13914 avdd.n8833 avdd.n8832 0.00548485
R13915 avdd.n8867 avdd.n8866 0.00548485
R13916 avdd.n8793 avdd.n8792 0.00548485
R13917 avdd.n241 avdd.n240 0.00548485
R13918 avdd.n300 avdd.n299 0.00548485
R13919 avdd.n8741 avdd.n8740 0.00548485
R13920 avdd.n8747 avdd.n8746 0.00548485
R13921 avdd.n8781 avdd.n8780 0.00548485
R13922 avdd.n8707 avdd.n8706 0.00548485
R13923 avdd.n371 avdd.n370 0.00548485
R13924 avdd.n430 avdd.n429 0.00548485
R13925 avdd.n8655 avdd.n8654 0.00548485
R13926 avdd.n8661 avdd.n8660 0.00548485
R13927 avdd.n8695 avdd.n8694 0.00548485
R13928 avdd.n8621 avdd.n8620 0.00548485
R13929 avdd.n501 avdd.n500 0.00548485
R13930 avdd.n560 avdd.n559 0.00548485
R13931 avdd.n8569 avdd.n8568 0.00548485
R13932 avdd.n8575 avdd.n8574 0.00548485
R13933 avdd.n8609 avdd.n8608 0.00548485
R13934 avdd.n8535 avdd.n8534 0.00548485
R13935 avdd.n631 avdd.n630 0.00548485
R13936 avdd.n690 avdd.n689 0.00548485
R13937 avdd.n8483 avdd.n8482 0.00548485
R13938 avdd.n8489 avdd.n8488 0.00548485
R13939 avdd.n8523 avdd.n8522 0.00548485
R13940 avdd.n8449 avdd.n8448 0.00548485
R13941 avdd.n761 avdd.n760 0.00548485
R13942 avdd.n820 avdd.n819 0.00548485
R13943 avdd.n8397 avdd.n8396 0.00548485
R13944 avdd.n8403 avdd.n8402 0.00548485
R13945 avdd.n8437 avdd.n8436 0.00548485
R13946 avdd.n8363 avdd.n8362 0.00548485
R13947 avdd.n891 avdd.n890 0.00548485
R13948 avdd.n950 avdd.n949 0.00548485
R13949 avdd.n8311 avdd.n8310 0.00548485
R13950 avdd.n8317 avdd.n8316 0.00548485
R13951 avdd.n8351 avdd.n8350 0.00548485
R13952 avdd.n8277 avdd.n8276 0.00548485
R13953 avdd.n1021 avdd.n1020 0.00548485
R13954 avdd.n1080 avdd.n1079 0.00548485
R13955 avdd.n8225 avdd.n8224 0.00548485
R13956 avdd.n8231 avdd.n8230 0.00548485
R13957 avdd.n8265 avdd.n8264 0.00548485
R13958 avdd.n8191 avdd.n8190 0.00548485
R13959 avdd.n1151 avdd.n1150 0.00548485
R13960 avdd.n1210 avdd.n1209 0.00548485
R13961 avdd.n8139 avdd.n8138 0.00548485
R13962 avdd.n8145 avdd.n8144 0.00548485
R13963 avdd.n8179 avdd.n8178 0.00548485
R13964 avdd.n8105 avdd.n8104 0.00548485
R13965 avdd.n1281 avdd.n1280 0.00548485
R13966 avdd.n1340 avdd.n1339 0.00548485
R13967 avdd.n8053 avdd.n8052 0.00548485
R13968 avdd.n8059 avdd.n8058 0.00548485
R13969 avdd.n8093 avdd.n8092 0.00548485
R13970 avdd.n8019 avdd.n8018 0.00548485
R13971 avdd.n1411 avdd.n1410 0.00548485
R13972 avdd.n1470 avdd.n1469 0.00548485
R13973 avdd.n7967 avdd.n7966 0.00548485
R13974 avdd.n7973 avdd.n7972 0.00548485
R13975 avdd.n8007 avdd.n8006 0.00548485
R13976 avdd.n7933 avdd.n7932 0.00548485
R13977 avdd.n1541 avdd.n1540 0.00548485
R13978 avdd.n1600 avdd.n1599 0.00548485
R13979 avdd.n7881 avdd.n7880 0.00548485
R13980 avdd.n7887 avdd.n7886 0.00548485
R13981 avdd.n7921 avdd.n7920 0.00548485
R13982 avdd.n2036 avdd.n2030 0.0052
R13983 avdd.n1881 avdd.n1878 0.0052
R13984 avdd.n2091 avdd.n1878 0.0052
R13985 avdd.n2305 avdd.n2093 0.0052
R13986 avdd.n2195 avdd.n2139 0.0052
R13987 avdd.n2195 avdd.n1877 0.0052
R13988 avdd.n2520 avdd.n2308 0.0052
R13989 avdd.n2410 avdd.n2354 0.0052
R13990 avdd.n2410 avdd.n1876 0.0052
R13991 avdd.n2735 avdd.n2523 0.0052
R13992 avdd.n2625 avdd.n2569 0.0052
R13993 avdd.n2625 avdd.n1875 0.0052
R13994 avdd.n2950 avdd.n2738 0.0052
R13995 avdd.n2840 avdd.n2784 0.0052
R13996 avdd.n2840 avdd.n1874 0.0052
R13997 avdd.n3165 avdd.n2953 0.0052
R13998 avdd.n3055 avdd.n2999 0.0052
R13999 avdd.n3055 avdd.n1873 0.0052
R14000 avdd.n3381 avdd.n3169 0.0052
R14001 avdd.n3325 avdd.n3296 0.0052
R14002 avdd.n3325 avdd.n3299 0.0052
R14003 avdd.n3596 avdd.n3384 0.0052
R14004 avdd.n3540 avdd.n3511 0.0052
R14005 avdd.n3540 avdd.n3514 0.0052
R14006 avdd.n3811 avdd.n3599 0.0052
R14007 avdd.n3755 avdd.n3726 0.0052
R14008 avdd.n3755 avdd.n3729 0.0052
R14009 avdd.n4026 avdd.n3814 0.0052
R14010 avdd.n3970 avdd.n3941 0.0052
R14011 avdd.n3970 avdd.n3944 0.0052
R14012 avdd.n4241 avdd.n4029 0.0052
R14013 avdd.n4185 avdd.n4156 0.0052
R14014 avdd.n4185 avdd.n4159 0.0052
R14015 avdd.n4456 avdd.n4244 0.0052
R14016 avdd.n4400 avdd.n4371 0.0052
R14017 avdd.n4400 avdd.n4374 0.0052
R14018 avdd.n5021 avdd.n4819 0.0052
R14019 avdd.n4918 avdd.n4866 0.0052
R14020 avdd.n5237 avdd.n5035 0.0052
R14021 avdd.n5134 avdd.n5082 0.0052
R14022 avdd.n5453 avdd.n5251 0.0052
R14023 avdd.n5350 avdd.n5298 0.0052
R14024 avdd.n5669 avdd.n5467 0.0052
R14025 avdd.n5566 avdd.n5514 0.0052
R14026 avdd.n5885 avdd.n5683 0.0052
R14027 avdd.n5782 avdd.n5730 0.0052
R14028 avdd.n6101 avdd.n5899 0.0052
R14029 avdd.n5998 avdd.n5946 0.0052
R14030 avdd.n6317 avdd.n6115 0.0052
R14031 avdd.n6214 avdd.n6162 0.0052
R14032 avdd.n6533 avdd.n6331 0.0052
R14033 avdd.n6430 avdd.n6378 0.0052
R14034 avdd.n6749 avdd.n6547 0.0052
R14035 avdd.n6646 avdd.n6594 0.0052
R14036 avdd.n6965 avdd.n6763 0.0052
R14037 avdd.n6862 avdd.n6810 0.0052
R14038 avdd.n7181 avdd.n6979 0.0052
R14039 avdd.n7078 avdd.n7026 0.0052
R14040 avdd.n7397 avdd.n7195 0.0052
R14041 avdd.n7294 avdd.n7242 0.0052
R14042 avdd.n7762 avdd.n7740 0.0052
R14043 avdd.n10241 avdd.n10219 0.0052
R14044 avdd.n10342 avdd.n10341 0.0052
R14045 avdd.n10028 avdd.n10027 0.0052
R14046 avdd.n10444 avdd.n10443 0.0052
R14047 avdd.n9914 avdd.n9913 0.0052
R14048 avdd.n10546 avdd.n10545 0.0052
R14049 avdd.n9800 avdd.n9799 0.0052
R14050 avdd.n10648 avdd.n10647 0.0052
R14051 avdd.n9686 avdd.n9685 0.0052
R14052 avdd.n10750 avdd.n10749 0.0052
R14053 avdd.n9572 avdd.n9571 0.0052
R14054 avdd.n10852 avdd.n10851 0.0052
R14055 avdd.n9458 avdd.n9457 0.0052
R14056 avdd.n10954 avdd.n10953 0.0052
R14057 avdd.n9344 avdd.n9343 0.0052
R14058 avdd.n11056 avdd.n11055 0.0052
R14059 avdd.n9230 avdd.n9229 0.0052
R14060 avdd.n11158 avdd.n11157 0.0052
R14061 avdd.n9116 avdd.n9115 0.0052
R14062 avdd.n11260 avdd.n11259 0.0052
R14063 avdd.n9002 avdd.n9001 0.0052
R14064 avdd.n8886 avdd.n8885 0.0052
R14065 avdd.n186 avdd.n95 0.0052
R14066 avdd.n187 avdd.n186 0.0052
R14067 avdd.n8800 avdd.n8799 0.0052
R14068 avdd.n316 avdd.n225 0.0052
R14069 avdd.n317 avdd.n316 0.0052
R14070 avdd.n8714 avdd.n8713 0.0052
R14071 avdd.n446 avdd.n355 0.0052
R14072 avdd.n447 avdd.n446 0.0052
R14073 avdd.n8628 avdd.n8627 0.0052
R14074 avdd.n576 avdd.n485 0.0052
R14075 avdd.n577 avdd.n576 0.0052
R14076 avdd.n8542 avdd.n8541 0.0052
R14077 avdd.n706 avdd.n615 0.0052
R14078 avdd.n707 avdd.n706 0.0052
R14079 avdd.n8456 avdd.n8455 0.0052
R14080 avdd.n836 avdd.n745 0.0052
R14081 avdd.n837 avdd.n836 0.0052
R14082 avdd.n8370 avdd.n8369 0.0052
R14083 avdd.n966 avdd.n875 0.0052
R14084 avdd.n967 avdd.n966 0.0052
R14085 avdd.n8284 avdd.n8283 0.0052
R14086 avdd.n1096 avdd.n1005 0.0052
R14087 avdd.n1097 avdd.n1096 0.0052
R14088 avdd.n8198 avdd.n8197 0.0052
R14089 avdd.n1226 avdd.n1135 0.0052
R14090 avdd.n1227 avdd.n1226 0.0052
R14091 avdd.n8112 avdd.n8111 0.0052
R14092 avdd.n1356 avdd.n1265 0.0052
R14093 avdd.n1357 avdd.n1356 0.0052
R14094 avdd.n8026 avdd.n8025 0.0052
R14095 avdd.n1486 avdd.n1395 0.0052
R14096 avdd.n1487 avdd.n1486 0.0052
R14097 avdd.n7940 avdd.n7939 0.0052
R14098 avdd.n1616 avdd.n1525 0.0052
R14099 avdd.n1617 avdd.n1616 0.0052
R14100 avdd.n7449 avdd.n7448 0.00492753
R14101 avdd.n7488 avdd.n7487 0.00492753
R14102 avdd.n7548 avdd.n7547 0.00492753
R14103 avdd.n7588 avdd.n7587 0.00492753
R14104 avdd.n1811 avdd.n1810 0.00492753
R14105 avdd.n1637 avdd.n1636 0.00492753
R14106 avdd.n1721 avdd.n1720 0.00492753
R14107 avdd.n1673 avdd.n1672 0.00492753
R14108 avdd.n1940 avdd.n1939 0.00477273
R14109 avdd.n2079 avdd.n2078 0.00477273
R14110 avdd.n1965 avdd.n1958 0.00477273
R14111 avdd.n1997 avdd.n1995 0.00477273
R14112 avdd.n2017 avdd.n2016 0.00477273
R14113 avdd.n2023 avdd.n2004 0.00477273
R14114 avdd.n2189 avdd.n2188 0.00477273
R14115 avdd.n2218 avdd.n2131 0.00477273
R14116 avdd.n2128 avdd.n2127 0.00477273
R14117 avdd.n2265 avdd.n2264 0.00477273
R14118 avdd.n2291 avdd.n2289 0.00477273
R14119 avdd.n2297 avdd.n2296 0.00477273
R14120 avdd.n2404 avdd.n2403 0.00477273
R14121 avdd.n2433 avdd.n2346 0.00477273
R14122 avdd.n2343 avdd.n2342 0.00477273
R14123 avdd.n2480 avdd.n2479 0.00477273
R14124 avdd.n2506 avdd.n2504 0.00477273
R14125 avdd.n2512 avdd.n2511 0.00477273
R14126 avdd.n2619 avdd.n2618 0.00477273
R14127 avdd.n2648 avdd.n2561 0.00477273
R14128 avdd.n2558 avdd.n2557 0.00477273
R14129 avdd.n2695 avdd.n2694 0.00477273
R14130 avdd.n2721 avdd.n2719 0.00477273
R14131 avdd.n2727 avdd.n2726 0.00477273
R14132 avdd.n2834 avdd.n2833 0.00477273
R14133 avdd.n2863 avdd.n2776 0.00477273
R14134 avdd.n2773 avdd.n2772 0.00477273
R14135 avdd.n2910 avdd.n2909 0.00477273
R14136 avdd.n2936 avdd.n2934 0.00477273
R14137 avdd.n2942 avdd.n2941 0.00477273
R14138 avdd.n3049 avdd.n3048 0.00477273
R14139 avdd.n3078 avdd.n2991 0.00477273
R14140 avdd.n2988 avdd.n2987 0.00477273
R14141 avdd.n3125 avdd.n3124 0.00477273
R14142 avdd.n3151 avdd.n3149 0.00477273
R14143 avdd.n3157 avdd.n3156 0.00477273
R14144 avdd.n3230 avdd.n3229 0.00477273
R14145 avdd.n3368 avdd.n3367 0.00477273
R14146 avdd.n3255 avdd.n3248 0.00477273
R14147 avdd.n3287 avdd.n3285 0.00477273
R14148 avdd.n3309 avdd.n3297 0.00477273
R14149 avdd.n3317 avdd.n3294 0.00477273
R14150 avdd.n3445 avdd.n3444 0.00477273
R14151 avdd.n3583 avdd.n3582 0.00477273
R14152 avdd.n3470 avdd.n3463 0.00477273
R14153 avdd.n3502 avdd.n3500 0.00477273
R14154 avdd.n3524 avdd.n3512 0.00477273
R14155 avdd.n3532 avdd.n3509 0.00477273
R14156 avdd.n3660 avdd.n3659 0.00477273
R14157 avdd.n3798 avdd.n3797 0.00477273
R14158 avdd.n3685 avdd.n3678 0.00477273
R14159 avdd.n3717 avdd.n3715 0.00477273
R14160 avdd.n3739 avdd.n3727 0.00477273
R14161 avdd.n3747 avdd.n3724 0.00477273
R14162 avdd.n3875 avdd.n3874 0.00477273
R14163 avdd.n4013 avdd.n4012 0.00477273
R14164 avdd.n3900 avdd.n3893 0.00477273
R14165 avdd.n3932 avdd.n3930 0.00477273
R14166 avdd.n3954 avdd.n3942 0.00477273
R14167 avdd.n3962 avdd.n3939 0.00477273
R14168 avdd.n4090 avdd.n4089 0.00477273
R14169 avdd.n4228 avdd.n4227 0.00477273
R14170 avdd.n4115 avdd.n4108 0.00477273
R14171 avdd.n4147 avdd.n4145 0.00477273
R14172 avdd.n4169 avdd.n4157 0.00477273
R14173 avdd.n4177 avdd.n4154 0.00477273
R14174 avdd.n4305 avdd.n4304 0.00477273
R14175 avdd.n4443 avdd.n4442 0.00477273
R14176 avdd.n4330 avdd.n4323 0.00477273
R14177 avdd.n4362 avdd.n4360 0.00477273
R14178 avdd.n4384 avdd.n4372 0.00477273
R14179 avdd.n4392 avdd.n4369 0.00477273
R14180 avdd.n4912 avdd.n4911 0.00477273
R14181 avdd.n4940 avdd.n4853 0.00477273
R14182 avdd.n4850 avdd.n4849 0.00477273
R14183 avdd.n4987 avdd.n4986 0.00477273
R14184 avdd.n5008 avdd.n5007 0.00477273
R14185 avdd.n5020 avdd.n4820 0.00477273
R14186 avdd.n5128 avdd.n5127 0.00477273
R14187 avdd.n5156 avdd.n5069 0.00477273
R14188 avdd.n5066 avdd.n5065 0.00477273
R14189 avdd.n5203 avdd.n5202 0.00477273
R14190 avdd.n5224 avdd.n5223 0.00477273
R14191 avdd.n5236 avdd.n5036 0.00477273
R14192 avdd.n5344 avdd.n5343 0.00477273
R14193 avdd.n5372 avdd.n5285 0.00477273
R14194 avdd.n5282 avdd.n5281 0.00477273
R14195 avdd.n5419 avdd.n5418 0.00477273
R14196 avdd.n5440 avdd.n5439 0.00477273
R14197 avdd.n5452 avdd.n5252 0.00477273
R14198 avdd.n5560 avdd.n5559 0.00477273
R14199 avdd.n5588 avdd.n5501 0.00477273
R14200 avdd.n5498 avdd.n5497 0.00477273
R14201 avdd.n5635 avdd.n5634 0.00477273
R14202 avdd.n5656 avdd.n5655 0.00477273
R14203 avdd.n5668 avdd.n5468 0.00477273
R14204 avdd.n5776 avdd.n5775 0.00477273
R14205 avdd.n5804 avdd.n5717 0.00477273
R14206 avdd.n5714 avdd.n5713 0.00477273
R14207 avdd.n5851 avdd.n5850 0.00477273
R14208 avdd.n5872 avdd.n5871 0.00477273
R14209 avdd.n5884 avdd.n5684 0.00477273
R14210 avdd.n5992 avdd.n5991 0.00477273
R14211 avdd.n6020 avdd.n5933 0.00477273
R14212 avdd.n5930 avdd.n5929 0.00477273
R14213 avdd.n6067 avdd.n6066 0.00477273
R14214 avdd.n6088 avdd.n6087 0.00477273
R14215 avdd.n6100 avdd.n5900 0.00477273
R14216 avdd.n6208 avdd.n6207 0.00477273
R14217 avdd.n6236 avdd.n6149 0.00477273
R14218 avdd.n6146 avdd.n6145 0.00477273
R14219 avdd.n6283 avdd.n6282 0.00477273
R14220 avdd.n6304 avdd.n6303 0.00477273
R14221 avdd.n6316 avdd.n6116 0.00477273
R14222 avdd.n6424 avdd.n6423 0.00477273
R14223 avdd.n6452 avdd.n6365 0.00477273
R14224 avdd.n6362 avdd.n6361 0.00477273
R14225 avdd.n6499 avdd.n6498 0.00477273
R14226 avdd.n6520 avdd.n6519 0.00477273
R14227 avdd.n6532 avdd.n6332 0.00477273
R14228 avdd.n6640 avdd.n6639 0.00477273
R14229 avdd.n6668 avdd.n6581 0.00477273
R14230 avdd.n6578 avdd.n6577 0.00477273
R14231 avdd.n6715 avdd.n6714 0.00477273
R14232 avdd.n6736 avdd.n6735 0.00477273
R14233 avdd.n6748 avdd.n6548 0.00477273
R14234 avdd.n6856 avdd.n6855 0.00477273
R14235 avdd.n6884 avdd.n6797 0.00477273
R14236 avdd.n6794 avdd.n6793 0.00477273
R14237 avdd.n6931 avdd.n6930 0.00477273
R14238 avdd.n6952 avdd.n6951 0.00477273
R14239 avdd.n6964 avdd.n6764 0.00477273
R14240 avdd.n7072 avdd.n7071 0.00477273
R14241 avdd.n7100 avdd.n7013 0.00477273
R14242 avdd.n7010 avdd.n7009 0.00477273
R14243 avdd.n7147 avdd.n7146 0.00477273
R14244 avdd.n7168 avdd.n7167 0.00477273
R14245 avdd.n7180 avdd.n6980 0.00477273
R14246 avdd.n7288 avdd.n7287 0.00477273
R14247 avdd.n7316 avdd.n7229 0.00477273
R14248 avdd.n7226 avdd.n7225 0.00477273
R14249 avdd.n7363 avdd.n7362 0.00477273
R14250 avdd.n7384 avdd.n7383 0.00477273
R14251 avdd.n7396 avdd.n7196 0.00477273
R14252 avdd.n7735 avdd.n7725 0.00477273
R14253 avdd.n7686 avdd.n7685 0.00477273
R14254 avdd.n7668 avdd.n7667 0.00477273
R14255 avdd.n7825 avdd.n7815 0.00477273
R14256 avdd.n7847 avdd.n7846 0.00477273
R14257 avdd.n7783 avdd.n7782 0.00477273
R14258 avdd.n10214 avdd.n10204 0.00477273
R14259 avdd.n10165 avdd.n10164 0.00477273
R14260 avdd.n10147 avdd.n10146 0.00477273
R14261 avdd.n10083 avdd.n10073 0.00477273
R14262 avdd.n10105 avdd.n10104 0.00477273
R14263 avdd.n10043 avdd.n10042 0.00477273
R14264 avdd.n9949 avdd.n9948 0.00477273
R14265 avdd.n9932 avdd.n9931 0.00477273
R14266 avdd.n10315 avdd.n10305 0.00477273
R14267 avdd.n10337 avdd.n10336 0.00477273
R14268 avdd.n10259 avdd.n10258 0.00477273
R14269 avdd.n9835 avdd.n9834 0.00477273
R14270 avdd.n9818 avdd.n9817 0.00477273
R14271 avdd.n10417 avdd.n10407 0.00477273
R14272 avdd.n10439 avdd.n10438 0.00477273
R14273 avdd.n10361 avdd.n10360 0.00477273
R14274 avdd.n9721 avdd.n9720 0.00477273
R14275 avdd.n9704 avdd.n9703 0.00477273
R14276 avdd.n10519 avdd.n10509 0.00477273
R14277 avdd.n10541 avdd.n10540 0.00477273
R14278 avdd.n10463 avdd.n10462 0.00477273
R14279 avdd.n9608 avdd.n9607 0.00477273
R14280 avdd.n9591 avdd.n9590 0.00477273
R14281 avdd.n10621 avdd.n10611 0.00477273
R14282 avdd.n10643 avdd.n10642 0.00477273
R14283 avdd.n10565 avdd.n10564 0.00477273
R14284 avdd.n9493 avdd.n9492 0.00477273
R14285 avdd.n9476 avdd.n9475 0.00477273
R14286 avdd.n10723 avdd.n10713 0.00477273
R14287 avdd.n10745 avdd.n10744 0.00477273
R14288 avdd.n10667 avdd.n10666 0.00477273
R14289 avdd.n9379 avdd.n9378 0.00477273
R14290 avdd.n9362 avdd.n9361 0.00477273
R14291 avdd.n10825 avdd.n10815 0.00477273
R14292 avdd.n10847 avdd.n10846 0.00477273
R14293 avdd.n10769 avdd.n10768 0.00477273
R14294 avdd.n9265 avdd.n9264 0.00477273
R14295 avdd.n9248 avdd.n9247 0.00477273
R14296 avdd.n10927 avdd.n10917 0.00477273
R14297 avdd.n10949 avdd.n10948 0.00477273
R14298 avdd.n10871 avdd.n10870 0.00477273
R14299 avdd.n9151 avdd.n9150 0.00477273
R14300 avdd.n9134 avdd.n9133 0.00477273
R14301 avdd.n11029 avdd.n11019 0.00477273
R14302 avdd.n11051 avdd.n11050 0.00477273
R14303 avdd.n10973 avdd.n10972 0.00477273
R14304 avdd.n9037 avdd.n9036 0.00477273
R14305 avdd.n9020 avdd.n9019 0.00477273
R14306 avdd.n11131 avdd.n11121 0.00477273
R14307 avdd.n11153 avdd.n11152 0.00477273
R14308 avdd.n11075 avdd.n11074 0.00477273
R14309 avdd.n8923 avdd.n8922 0.00477273
R14310 avdd.n8906 avdd.n8905 0.00477273
R14311 avdd.n11233 avdd.n11223 0.00477273
R14312 avdd.n11255 avdd.n11254 0.00477273
R14313 avdd.n11177 avdd.n11176 0.00477273
R14314 avdd.n130 avdd.n120 0.00477273
R14315 avdd.n169 avdd.n168 0.00477273
R14316 avdd.n151 avdd.n150 0.00477273
R14317 avdd.n8846 avdd.n8836 0.00477273
R14318 avdd.n8868 avdd.n8867 0.00477273
R14319 avdd.n8806 avdd.n8805 0.00477273
R14320 avdd.n260 avdd.n250 0.00477273
R14321 avdd.n299 avdd.n298 0.00477273
R14322 avdd.n281 avdd.n280 0.00477273
R14323 avdd.n8760 avdd.n8750 0.00477273
R14324 avdd.n8782 avdd.n8781 0.00477273
R14325 avdd.n8720 avdd.n8719 0.00477273
R14326 avdd.n390 avdd.n380 0.00477273
R14327 avdd.n429 avdd.n428 0.00477273
R14328 avdd.n411 avdd.n410 0.00477273
R14329 avdd.n8674 avdd.n8664 0.00477273
R14330 avdd.n8696 avdd.n8695 0.00477273
R14331 avdd.n8634 avdd.n8633 0.00477273
R14332 avdd.n520 avdd.n510 0.00477273
R14333 avdd.n559 avdd.n558 0.00477273
R14334 avdd.n541 avdd.n540 0.00477273
R14335 avdd.n8588 avdd.n8578 0.00477273
R14336 avdd.n8610 avdd.n8609 0.00477273
R14337 avdd.n8548 avdd.n8547 0.00477273
R14338 avdd.n650 avdd.n640 0.00477273
R14339 avdd.n689 avdd.n688 0.00477273
R14340 avdd.n671 avdd.n670 0.00477273
R14341 avdd.n8502 avdd.n8492 0.00477273
R14342 avdd.n8524 avdd.n8523 0.00477273
R14343 avdd.n8462 avdd.n8461 0.00477273
R14344 avdd.n780 avdd.n770 0.00477273
R14345 avdd.n819 avdd.n818 0.00477273
R14346 avdd.n801 avdd.n800 0.00477273
R14347 avdd.n8416 avdd.n8406 0.00477273
R14348 avdd.n8438 avdd.n8437 0.00477273
R14349 avdd.n8376 avdd.n8375 0.00477273
R14350 avdd.n910 avdd.n900 0.00477273
R14351 avdd.n949 avdd.n948 0.00477273
R14352 avdd.n931 avdd.n930 0.00477273
R14353 avdd.n8330 avdd.n8320 0.00477273
R14354 avdd.n8352 avdd.n8351 0.00477273
R14355 avdd.n8290 avdd.n8289 0.00477273
R14356 avdd.n1040 avdd.n1030 0.00477273
R14357 avdd.n1079 avdd.n1078 0.00477273
R14358 avdd.n1061 avdd.n1060 0.00477273
R14359 avdd.n8244 avdd.n8234 0.00477273
R14360 avdd.n8266 avdd.n8265 0.00477273
R14361 avdd.n8204 avdd.n8203 0.00477273
R14362 avdd.n1170 avdd.n1160 0.00477273
R14363 avdd.n1209 avdd.n1208 0.00477273
R14364 avdd.n1191 avdd.n1190 0.00477273
R14365 avdd.n8158 avdd.n8148 0.00477273
R14366 avdd.n8180 avdd.n8179 0.00477273
R14367 avdd.n8118 avdd.n8117 0.00477273
R14368 avdd.n1300 avdd.n1290 0.00477273
R14369 avdd.n1339 avdd.n1338 0.00477273
R14370 avdd.n1321 avdd.n1320 0.00477273
R14371 avdd.n8072 avdd.n8062 0.00477273
R14372 avdd.n8094 avdd.n8093 0.00477273
R14373 avdd.n8032 avdd.n8031 0.00477273
R14374 avdd.n1430 avdd.n1420 0.00477273
R14375 avdd.n1469 avdd.n1468 0.00477273
R14376 avdd.n1451 avdd.n1450 0.00477273
R14377 avdd.n7986 avdd.n7976 0.00477273
R14378 avdd.n8008 avdd.n8007 0.00477273
R14379 avdd.n7946 avdd.n7945 0.00477273
R14380 avdd.n1560 avdd.n1550 0.00477273
R14381 avdd.n1599 avdd.n1598 0.00477273
R14382 avdd.n1581 avdd.n1580 0.00477273
R14383 avdd.n7900 avdd.n7890 0.00477273
R14384 avdd.n7922 avdd.n7921 0.00477273
R14385 avdd.n7860 avdd.n7859 0.00477273
R14386 avdd.n4607 avdd.n4606 0.00466667
R14387 avdd.n4736 avdd.n4518 0.00466667
R14388 avdd.n2043 avdd.n2042 0.00428788
R14389 avdd.n1943 avdd.n1942 0.00428788
R14390 avdd.n2279 avdd.n2104 0.00428788
R14391 avdd.n2199 avdd.n2137 0.00428788
R14392 avdd.n2494 avdd.n2319 0.00428788
R14393 avdd.n2414 avdd.n2352 0.00428788
R14394 avdd.n2709 avdd.n2534 0.00428788
R14395 avdd.n2629 avdd.n2567 0.00428788
R14396 avdd.n2924 avdd.n2749 0.00428788
R14397 avdd.n2844 avdd.n2782 0.00428788
R14398 avdd.n3139 avdd.n2964 0.00428788
R14399 avdd.n3059 avdd.n2997 0.00428788
R14400 avdd.n3332 avdd.n3331 0.00428788
R14401 avdd.n3233 avdd.n3232 0.00428788
R14402 avdd.n3547 avdd.n3546 0.00428788
R14403 avdd.n3448 avdd.n3447 0.00428788
R14404 avdd.n3762 avdd.n3761 0.00428788
R14405 avdd.n3663 avdd.n3662 0.00428788
R14406 avdd.n3977 avdd.n3976 0.00428788
R14407 avdd.n3878 avdd.n3877 0.00428788
R14408 avdd.n4192 avdd.n4191 0.00428788
R14409 avdd.n4093 avdd.n4092 0.00428788
R14410 avdd.n4407 avdd.n4406 0.00428788
R14411 avdd.n4308 avdd.n4307 0.00428788
R14412 avdd.n4921 avdd.n4859 0.00428788
R14413 avdd.n4998 avdd.n4825 0.00428788
R14414 avdd.n5137 avdd.n5075 0.00428788
R14415 avdd.n5214 avdd.n5041 0.00428788
R14416 avdd.n5353 avdd.n5291 0.00428788
R14417 avdd.n5430 avdd.n5257 0.00428788
R14418 avdd.n5569 avdd.n5507 0.00428788
R14419 avdd.n5646 avdd.n5473 0.00428788
R14420 avdd.n5785 avdd.n5723 0.00428788
R14421 avdd.n5862 avdd.n5689 0.00428788
R14422 avdd.n6001 avdd.n5939 0.00428788
R14423 avdd.n6078 avdd.n5905 0.00428788
R14424 avdd.n6217 avdd.n6155 0.00428788
R14425 avdd.n6294 avdd.n6121 0.00428788
R14426 avdd.n6433 avdd.n6371 0.00428788
R14427 avdd.n6510 avdd.n6337 0.00428788
R14428 avdd.n6649 avdd.n6587 0.00428788
R14429 avdd.n6726 avdd.n6553 0.00428788
R14430 avdd.n6865 avdd.n6803 0.00428788
R14431 avdd.n6942 avdd.n6769 0.00428788
R14432 avdd.n7081 avdd.n7019 0.00428788
R14433 avdd.n7158 avdd.n6985 0.00428788
R14434 avdd.n7297 avdd.n7235 0.00428788
R14435 avdd.n7374 avdd.n7201 0.00428788
R14436 avdd.n7733 avdd.n7732 0.00428788
R14437 avdd.n7823 avdd.n7822 0.00428788
R14438 avdd.n10212 avdd.n10211 0.00428788
R14439 avdd.n10081 avdd.n10080 0.00428788
R14440 avdd.n10018 avdd.n10017 0.00428788
R14441 avdd.n10313 avdd.n10312 0.00428788
R14442 avdd.n9904 avdd.n9903 0.00428788
R14443 avdd.n10415 avdd.n10414 0.00428788
R14444 avdd.n9790 avdd.n9789 0.00428788
R14445 avdd.n10517 avdd.n10516 0.00428788
R14446 avdd.n9677 avdd.n9676 0.00428788
R14447 avdd.n10619 avdd.n10618 0.00428788
R14448 avdd.n9562 avdd.n9561 0.00428788
R14449 avdd.n10721 avdd.n10720 0.00428788
R14450 avdd.n9448 avdd.n9447 0.00428788
R14451 avdd.n10823 avdd.n10822 0.00428788
R14452 avdd.n9334 avdd.n9333 0.00428788
R14453 avdd.n10925 avdd.n10924 0.00428788
R14454 avdd.n9220 avdd.n9219 0.00428788
R14455 avdd.n11027 avdd.n11026 0.00428788
R14456 avdd.n9106 avdd.n9105 0.00428788
R14457 avdd.n11129 avdd.n11128 0.00428788
R14458 avdd.n8992 avdd.n8991 0.00428788
R14459 avdd.n11231 avdd.n11230 0.00428788
R14460 avdd.n8844 avdd.n8843 0.00428788
R14461 avdd.n128 avdd.n127 0.00428788
R14462 avdd.n8758 avdd.n8757 0.00428788
R14463 avdd.n258 avdd.n257 0.00428788
R14464 avdd.n8672 avdd.n8671 0.00428788
R14465 avdd.n388 avdd.n387 0.00428788
R14466 avdd.n8586 avdd.n8585 0.00428788
R14467 avdd.n518 avdd.n517 0.00428788
R14468 avdd.n8500 avdd.n8499 0.00428788
R14469 avdd.n648 avdd.n647 0.00428788
R14470 avdd.n8414 avdd.n8413 0.00428788
R14471 avdd.n778 avdd.n777 0.00428788
R14472 avdd.n8328 avdd.n8327 0.00428788
R14473 avdd.n908 avdd.n907 0.00428788
R14474 avdd.n8242 avdd.n8241 0.00428788
R14475 avdd.n1038 avdd.n1037 0.00428788
R14476 avdd.n8156 avdd.n8155 0.00428788
R14477 avdd.n1168 avdd.n1167 0.00428788
R14478 avdd.n8070 avdd.n8069 0.00428788
R14479 avdd.n1298 avdd.n1297 0.00428788
R14480 avdd.n7984 avdd.n7983 0.00428788
R14481 avdd.n1428 avdd.n1427 0.00428788
R14482 avdd.n7898 avdd.n7897 0.00428788
R14483 avdd.n1558 avdd.n1557 0.00428788
R14484 avdd.n3319 avdd.n3298 0.00420154
R14485 avdd.n3305 avdd.n3298 0.00420154
R14486 avdd.n3534 avdd.n3513 0.00420154
R14487 avdd.n3520 avdd.n3513 0.00420154
R14488 avdd.n3749 avdd.n3728 0.00420154
R14489 avdd.n3735 avdd.n3728 0.00420154
R14490 avdd.n3964 avdd.n3943 0.00420154
R14491 avdd.n3950 avdd.n3943 0.00420154
R14492 avdd.n4179 avdd.n4158 0.00420154
R14493 avdd.n4165 avdd.n4158 0.00420154
R14494 avdd.n4394 avdd.n4373 0.00420154
R14495 avdd.n4380 avdd.n4373 0.00420154
R14496 avdd.n5015 avdd.n4818 0.00420154
R14497 avdd.n4818 avdd.n4811 0.00420154
R14498 avdd.n5231 avdd.n5034 0.00420154
R14499 avdd.n5034 avdd.n5027 0.00420154
R14500 avdd.n5447 avdd.n5250 0.00420154
R14501 avdd.n5250 avdd.n5243 0.00420154
R14502 avdd.n5663 avdd.n5466 0.00420154
R14503 avdd.n5466 avdd.n5459 0.00420154
R14504 avdd.n5879 avdd.n5682 0.00420154
R14505 avdd.n5682 avdd.n5675 0.00420154
R14506 avdd.n6095 avdd.n5898 0.00420154
R14507 avdd.n5898 avdd.n5891 0.00420154
R14508 avdd.n6311 avdd.n6114 0.00420154
R14509 avdd.n6114 avdd.n6107 0.00420154
R14510 avdd.n6527 avdd.n6330 0.00420154
R14511 avdd.n6330 avdd.n6323 0.00420154
R14512 avdd.n6743 avdd.n6546 0.00420154
R14513 avdd.n6546 avdd.n6539 0.00420154
R14514 avdd.n6959 avdd.n6762 0.00420154
R14515 avdd.n6762 avdd.n6755 0.00420154
R14516 avdd.n7175 avdd.n6978 0.00420154
R14517 avdd.n6978 avdd.n6971 0.00420154
R14518 avdd.n7391 avdd.n7194 0.00420154
R14519 avdd.n7194 avdd.n7187 0.00420154
R14520 avdd.n10268 avdd.n10267 0.00420154
R14521 avdd.n10269 avdd.n10268 0.00420154
R14522 avdd.n10370 avdd.n10369 0.00420154
R14523 avdd.n10371 avdd.n10370 0.00420154
R14524 avdd.n10472 avdd.n10471 0.00420154
R14525 avdd.n10473 avdd.n10472 0.00420154
R14526 avdd.n10574 avdd.n10573 0.00420154
R14527 avdd.n10575 avdd.n10574 0.00420154
R14528 avdd.n10676 avdd.n10675 0.00420154
R14529 avdd.n10677 avdd.n10676 0.00420154
R14530 avdd.n10778 avdd.n10777 0.00420154
R14531 avdd.n10779 avdd.n10778 0.00420154
R14532 avdd.n10880 avdd.n10879 0.00420154
R14533 avdd.n10881 avdd.n10880 0.00420154
R14534 avdd.n10982 avdd.n10981 0.00420154
R14535 avdd.n10983 avdd.n10982 0.00420154
R14536 avdd.n11084 avdd.n11083 0.00420154
R14537 avdd.n11085 avdd.n11084 0.00420154
R14538 avdd.n11186 avdd.n11185 0.00420154
R14539 avdd.n11187 avdd.n11186 0.00420154
R14540 avdd.n1952 avdd.n1951 0.00406061
R14541 avdd.n1953 avdd.n1888 0.00406061
R14542 avdd.n1964 avdd.n1950 0.00406061
R14543 avdd.n2024 avdd.n2009 0.00406061
R14544 avdd.n2216 avdd.n2215 0.00406061
R14545 avdd.n2214 avdd.n2132 0.00406061
R14546 avdd.n2227 avdd.n2124 0.00406061
R14547 avdd.n2301 avdd.n2098 0.00406061
R14548 avdd.n2431 avdd.n2430 0.00406061
R14549 avdd.n2429 avdd.n2347 0.00406061
R14550 avdd.n2442 avdd.n2339 0.00406061
R14551 avdd.n2516 avdd.n2313 0.00406061
R14552 avdd.n2646 avdd.n2645 0.00406061
R14553 avdd.n2644 avdd.n2562 0.00406061
R14554 avdd.n2657 avdd.n2554 0.00406061
R14555 avdd.n2731 avdd.n2528 0.00406061
R14556 avdd.n2861 avdd.n2860 0.00406061
R14557 avdd.n2859 avdd.n2777 0.00406061
R14558 avdd.n2872 avdd.n2769 0.00406061
R14559 avdd.n2946 avdd.n2743 0.00406061
R14560 avdd.n3076 avdd.n3075 0.00406061
R14561 avdd.n3074 avdd.n2992 0.00406061
R14562 avdd.n3087 avdd.n2984 0.00406061
R14563 avdd.n3161 avdd.n2958 0.00406061
R14564 avdd.n3242 avdd.n3241 0.00406061
R14565 avdd.n3243 avdd.n3178 0.00406061
R14566 avdd.n3254 avdd.n3240 0.00406061
R14567 avdd.n3319 avdd.n3318 0.00406061
R14568 avdd.n3457 avdd.n3456 0.00406061
R14569 avdd.n3458 avdd.n3393 0.00406061
R14570 avdd.n3469 avdd.n3455 0.00406061
R14571 avdd.n3534 avdd.n3533 0.00406061
R14572 avdd.n3672 avdd.n3671 0.00406061
R14573 avdd.n3673 avdd.n3608 0.00406061
R14574 avdd.n3684 avdd.n3670 0.00406061
R14575 avdd.n3749 avdd.n3748 0.00406061
R14576 avdd.n3887 avdd.n3886 0.00406061
R14577 avdd.n3888 avdd.n3823 0.00406061
R14578 avdd.n3899 avdd.n3885 0.00406061
R14579 avdd.n3964 avdd.n3963 0.00406061
R14580 avdd.n4102 avdd.n4101 0.00406061
R14581 avdd.n4103 avdd.n4038 0.00406061
R14582 avdd.n4114 avdd.n4100 0.00406061
R14583 avdd.n4179 avdd.n4178 0.00406061
R14584 avdd.n4317 avdd.n4316 0.00406061
R14585 avdd.n4318 avdd.n4253 0.00406061
R14586 avdd.n4329 avdd.n4315 0.00406061
R14587 avdd.n4394 avdd.n4393 0.00406061
R14588 avdd.n4938 avdd.n4937 0.00406061
R14589 avdd.n4936 avdd.n4854 0.00406061
R14590 avdd.n4949 avdd.n4846 0.00406061
R14591 avdd.n5016 avdd.n5015 0.00406061
R14592 avdd.n5154 avdd.n5153 0.00406061
R14593 avdd.n5152 avdd.n5070 0.00406061
R14594 avdd.n5165 avdd.n5062 0.00406061
R14595 avdd.n5232 avdd.n5231 0.00406061
R14596 avdd.n5370 avdd.n5369 0.00406061
R14597 avdd.n5368 avdd.n5286 0.00406061
R14598 avdd.n5381 avdd.n5278 0.00406061
R14599 avdd.n5448 avdd.n5447 0.00406061
R14600 avdd.n5586 avdd.n5585 0.00406061
R14601 avdd.n5584 avdd.n5502 0.00406061
R14602 avdd.n5597 avdd.n5494 0.00406061
R14603 avdd.n5664 avdd.n5663 0.00406061
R14604 avdd.n5802 avdd.n5801 0.00406061
R14605 avdd.n5800 avdd.n5718 0.00406061
R14606 avdd.n5813 avdd.n5710 0.00406061
R14607 avdd.n5880 avdd.n5879 0.00406061
R14608 avdd.n6018 avdd.n6017 0.00406061
R14609 avdd.n6016 avdd.n5934 0.00406061
R14610 avdd.n6029 avdd.n5926 0.00406061
R14611 avdd.n6096 avdd.n6095 0.00406061
R14612 avdd.n6234 avdd.n6233 0.00406061
R14613 avdd.n6232 avdd.n6150 0.00406061
R14614 avdd.n6245 avdd.n6142 0.00406061
R14615 avdd.n6312 avdd.n6311 0.00406061
R14616 avdd.n6450 avdd.n6449 0.00406061
R14617 avdd.n6448 avdd.n6366 0.00406061
R14618 avdd.n6461 avdd.n6358 0.00406061
R14619 avdd.n6528 avdd.n6527 0.00406061
R14620 avdd.n6666 avdd.n6665 0.00406061
R14621 avdd.n6664 avdd.n6582 0.00406061
R14622 avdd.n6677 avdd.n6574 0.00406061
R14623 avdd.n6744 avdd.n6743 0.00406061
R14624 avdd.n6882 avdd.n6881 0.00406061
R14625 avdd.n6880 avdd.n6798 0.00406061
R14626 avdd.n6893 avdd.n6790 0.00406061
R14627 avdd.n6960 avdd.n6959 0.00406061
R14628 avdd.n7098 avdd.n7097 0.00406061
R14629 avdd.n7096 avdd.n7014 0.00406061
R14630 avdd.n7109 avdd.n7006 0.00406061
R14631 avdd.n7176 avdd.n7175 0.00406061
R14632 avdd.n7314 avdd.n7313 0.00406061
R14633 avdd.n7312 avdd.n7230 0.00406061
R14634 avdd.n7325 avdd.n7222 0.00406061
R14635 avdd.n7392 avdd.n7391 0.00406061
R14636 avdd.n7648 avdd.n7647 0.00406061
R14637 avdd.n7684 avdd.n7683 0.00406061
R14638 avdd.n7678 avdd.n7677 0.00406061
R14639 avdd.n7791 avdd.n7790 0.00406061
R14640 avdd.n10125 avdd.n10124 0.00406061
R14641 avdd.n10163 avdd.n10162 0.00406061
R14642 avdd.n10157 avdd.n10156 0.00406061
R14643 avdd.n10051 avdd.n10050 0.00406061
R14644 avdd.n9926 avdd.n9925 0.00406061
R14645 avdd.n9947 avdd.n9946 0.00406061
R14646 avdd.n9941 avdd.n9940 0.00406061
R14647 avdd.n10267 avdd.n10266 0.00406061
R14648 avdd.n9812 avdd.n9811 0.00406061
R14649 avdd.n9833 avdd.n9832 0.00406061
R14650 avdd.n9827 avdd.n9826 0.00406061
R14651 avdd.n10369 avdd.n10368 0.00406061
R14652 avdd.n9698 avdd.n9697 0.00406061
R14653 avdd.n9719 avdd.n9718 0.00406061
R14654 avdd.n9713 avdd.n9712 0.00406061
R14655 avdd.n10471 avdd.n10470 0.00406061
R14656 avdd.n9584 avdd.n9583 0.00406061
R14657 avdd.n9606 avdd.n9605 0.00406061
R14658 avdd.n9600 avdd.n9599 0.00406061
R14659 avdd.n10573 avdd.n10572 0.00406061
R14660 avdd.n9470 avdd.n9469 0.00406061
R14661 avdd.n9491 avdd.n9490 0.00406061
R14662 avdd.n9485 avdd.n9484 0.00406061
R14663 avdd.n10675 avdd.n10674 0.00406061
R14664 avdd.n9356 avdd.n9355 0.00406061
R14665 avdd.n9377 avdd.n9376 0.00406061
R14666 avdd.n9371 avdd.n9370 0.00406061
R14667 avdd.n10777 avdd.n10776 0.00406061
R14668 avdd.n9242 avdd.n9241 0.00406061
R14669 avdd.n9263 avdd.n9262 0.00406061
R14670 avdd.n9257 avdd.n9256 0.00406061
R14671 avdd.n10879 avdd.n10878 0.00406061
R14672 avdd.n9128 avdd.n9127 0.00406061
R14673 avdd.n9149 avdd.n9148 0.00406061
R14674 avdd.n9143 avdd.n9142 0.00406061
R14675 avdd.n10981 avdd.n10980 0.00406061
R14676 avdd.n9014 avdd.n9013 0.00406061
R14677 avdd.n9035 avdd.n9034 0.00406061
R14678 avdd.n9029 avdd.n9028 0.00406061
R14679 avdd.n11083 avdd.n11082 0.00406061
R14680 avdd.n8900 avdd.n8899 0.00406061
R14681 avdd.n8921 avdd.n8920 0.00406061
R14682 avdd.n8915 avdd.n8914 0.00406061
R14683 avdd.n11185 avdd.n11184 0.00406061
R14684 avdd.n69 avdd.n68 0.00406061
R14685 avdd.n167 avdd.n166 0.00406061
R14686 avdd.n161 avdd.n160 0.00406061
R14687 avdd.n8814 avdd.n8813 0.00406061
R14688 avdd.n199 avdd.n198 0.00406061
R14689 avdd.n297 avdd.n296 0.00406061
R14690 avdd.n291 avdd.n290 0.00406061
R14691 avdd.n8728 avdd.n8727 0.00406061
R14692 avdd.n329 avdd.n328 0.00406061
R14693 avdd.n427 avdd.n426 0.00406061
R14694 avdd.n421 avdd.n420 0.00406061
R14695 avdd.n8642 avdd.n8641 0.00406061
R14696 avdd.n459 avdd.n458 0.00406061
R14697 avdd.n557 avdd.n556 0.00406061
R14698 avdd.n551 avdd.n550 0.00406061
R14699 avdd.n8556 avdd.n8555 0.00406061
R14700 avdd.n589 avdd.n588 0.00406061
R14701 avdd.n687 avdd.n686 0.00406061
R14702 avdd.n681 avdd.n680 0.00406061
R14703 avdd.n8470 avdd.n8469 0.00406061
R14704 avdd.n719 avdd.n718 0.00406061
R14705 avdd.n817 avdd.n816 0.00406061
R14706 avdd.n811 avdd.n810 0.00406061
R14707 avdd.n8384 avdd.n8383 0.00406061
R14708 avdd.n849 avdd.n848 0.00406061
R14709 avdd.n947 avdd.n946 0.00406061
R14710 avdd.n941 avdd.n940 0.00406061
R14711 avdd.n8298 avdd.n8297 0.00406061
R14712 avdd.n979 avdd.n978 0.00406061
R14713 avdd.n1077 avdd.n1076 0.00406061
R14714 avdd.n1071 avdd.n1070 0.00406061
R14715 avdd.n8212 avdd.n8211 0.00406061
R14716 avdd.n1109 avdd.n1108 0.00406061
R14717 avdd.n1207 avdd.n1206 0.00406061
R14718 avdd.n1201 avdd.n1200 0.00406061
R14719 avdd.n8126 avdd.n8125 0.00406061
R14720 avdd.n1239 avdd.n1238 0.00406061
R14721 avdd.n1337 avdd.n1336 0.00406061
R14722 avdd.n1331 avdd.n1330 0.00406061
R14723 avdd.n8040 avdd.n8039 0.00406061
R14724 avdd.n1369 avdd.n1368 0.00406061
R14725 avdd.n1467 avdd.n1466 0.00406061
R14726 avdd.n1461 avdd.n1460 0.00406061
R14727 avdd.n7954 avdd.n7953 0.00406061
R14728 avdd.n1499 avdd.n1498 0.00406061
R14729 avdd.n1597 avdd.n1596 0.00406061
R14730 avdd.n1591 avdd.n1590 0.00406061
R14731 avdd.n7868 avdd.n7867 0.00406061
R14732 avdd.n1923 avdd.n1899 0.00334848
R14733 avdd.n1935 avdd.n1891 0.00334848
R14734 avdd.n2084 avdd.n1884 0.00334848
R14735 avdd.n2054 avdd.n1973 0.00334848
R14736 avdd.n2047 avdd.n1980 0.00334848
R14737 avdd.n2038 avdd.n2037 0.00334848
R14738 avdd.n2177 avdd.n2153 0.00334848
R14739 avdd.n2193 avdd.n2146 0.00334848
R14740 avdd.n2207 avdd.n2134 0.00334848
R14741 avdd.n2248 avdd.n2116 0.00334848
R14742 avdd.n2269 avdd.n2109 0.00334848
R14743 avdd.n2284 avdd.n2283 0.00334848
R14744 avdd.n2392 avdd.n2368 0.00334848
R14745 avdd.n2408 avdd.n2361 0.00334848
R14746 avdd.n2422 avdd.n2349 0.00334848
R14747 avdd.n2463 avdd.n2331 0.00334848
R14748 avdd.n2484 avdd.n2324 0.00334848
R14749 avdd.n2499 avdd.n2498 0.00334848
R14750 avdd.n2607 avdd.n2583 0.00334848
R14751 avdd.n2623 avdd.n2576 0.00334848
R14752 avdd.n2637 avdd.n2564 0.00334848
R14753 avdd.n2678 avdd.n2546 0.00334848
R14754 avdd.n2699 avdd.n2539 0.00334848
R14755 avdd.n2714 avdd.n2713 0.00334848
R14756 avdd.n2822 avdd.n2798 0.00334848
R14757 avdd.n2838 avdd.n2791 0.00334848
R14758 avdd.n2852 avdd.n2779 0.00334848
R14759 avdd.n2893 avdd.n2761 0.00334848
R14760 avdd.n2914 avdd.n2754 0.00334848
R14761 avdd.n2929 avdd.n2928 0.00334848
R14762 avdd.n3037 avdd.n3013 0.00334848
R14763 avdd.n3053 avdd.n3006 0.00334848
R14764 avdd.n3067 avdd.n2994 0.00334848
R14765 avdd.n3108 avdd.n2976 0.00334848
R14766 avdd.n3129 avdd.n2969 0.00334848
R14767 avdd.n3144 avdd.n3143 0.00334848
R14768 avdd.n3213 avdd.n3189 0.00334848
R14769 avdd.n3225 avdd.n3181 0.00334848
R14770 avdd.n3373 avdd.n3174 0.00334848
R14771 avdd.n3343 avdd.n3263 0.00334848
R14772 avdd.n3336 avdd.n3270 0.00334848
R14773 avdd.n3327 avdd.n3326 0.00334848
R14774 avdd.n3428 avdd.n3404 0.00334848
R14775 avdd.n3440 avdd.n3396 0.00334848
R14776 avdd.n3588 avdd.n3389 0.00334848
R14777 avdd.n3558 avdd.n3478 0.00334848
R14778 avdd.n3551 avdd.n3485 0.00334848
R14779 avdd.n3542 avdd.n3541 0.00334848
R14780 avdd.n3643 avdd.n3619 0.00334848
R14781 avdd.n3655 avdd.n3611 0.00334848
R14782 avdd.n3803 avdd.n3604 0.00334848
R14783 avdd.n3773 avdd.n3693 0.00334848
R14784 avdd.n3766 avdd.n3700 0.00334848
R14785 avdd.n3757 avdd.n3756 0.00334848
R14786 avdd.n3858 avdd.n3834 0.00334848
R14787 avdd.n3870 avdd.n3826 0.00334848
R14788 avdd.n4018 avdd.n3819 0.00334848
R14789 avdd.n3988 avdd.n3908 0.00334848
R14790 avdd.n3981 avdd.n3915 0.00334848
R14791 avdd.n3972 avdd.n3971 0.00334848
R14792 avdd.n4073 avdd.n4049 0.00334848
R14793 avdd.n4085 avdd.n4041 0.00334848
R14794 avdd.n4233 avdd.n4034 0.00334848
R14795 avdd.n4203 avdd.n4123 0.00334848
R14796 avdd.n4196 avdd.n4130 0.00334848
R14797 avdd.n4187 avdd.n4186 0.00334848
R14798 avdd.n4288 avdd.n4264 0.00334848
R14799 avdd.n4300 avdd.n4256 0.00334848
R14800 avdd.n4448 avdd.n4249 0.00334848
R14801 avdd.n4418 avdd.n4338 0.00334848
R14802 avdd.n4411 avdd.n4345 0.00334848
R14803 avdd.n4402 avdd.n4401 0.00334848
R14804 avdd.n4899 avdd.n4875 0.00334848
R14805 avdd.n4916 avdd.n4868 0.00334848
R14806 avdd.n4929 avdd.n4856 0.00334848
R14807 avdd.n4970 avdd.n4838 0.00334848
R14808 avdd.n4991 avdd.n4831 0.00334848
R14809 avdd.n5001 avdd.n4815 0.00334848
R14810 avdd.n5115 avdd.n5091 0.00334848
R14811 avdd.n5132 avdd.n5084 0.00334848
R14812 avdd.n5145 avdd.n5072 0.00334848
R14813 avdd.n5186 avdd.n5054 0.00334848
R14814 avdd.n5207 avdd.n5047 0.00334848
R14815 avdd.n5217 avdd.n5031 0.00334848
R14816 avdd.n5331 avdd.n5307 0.00334848
R14817 avdd.n5348 avdd.n5300 0.00334848
R14818 avdd.n5361 avdd.n5288 0.00334848
R14819 avdd.n5402 avdd.n5270 0.00334848
R14820 avdd.n5423 avdd.n5263 0.00334848
R14821 avdd.n5433 avdd.n5247 0.00334848
R14822 avdd.n5547 avdd.n5523 0.00334848
R14823 avdd.n5564 avdd.n5516 0.00334848
R14824 avdd.n5577 avdd.n5504 0.00334848
R14825 avdd.n5618 avdd.n5486 0.00334848
R14826 avdd.n5639 avdd.n5479 0.00334848
R14827 avdd.n5649 avdd.n5463 0.00334848
R14828 avdd.n5763 avdd.n5739 0.00334848
R14829 avdd.n5780 avdd.n5732 0.00334848
R14830 avdd.n5793 avdd.n5720 0.00334848
R14831 avdd.n5834 avdd.n5702 0.00334848
R14832 avdd.n5855 avdd.n5695 0.00334848
R14833 avdd.n5865 avdd.n5679 0.00334848
R14834 avdd.n5979 avdd.n5955 0.00334848
R14835 avdd.n5996 avdd.n5948 0.00334848
R14836 avdd.n6009 avdd.n5936 0.00334848
R14837 avdd.n6050 avdd.n5918 0.00334848
R14838 avdd.n6071 avdd.n5911 0.00334848
R14839 avdd.n6081 avdd.n5895 0.00334848
R14840 avdd.n6195 avdd.n6171 0.00334848
R14841 avdd.n6212 avdd.n6164 0.00334848
R14842 avdd.n6225 avdd.n6152 0.00334848
R14843 avdd.n6266 avdd.n6134 0.00334848
R14844 avdd.n6287 avdd.n6127 0.00334848
R14845 avdd.n6297 avdd.n6111 0.00334848
R14846 avdd.n6411 avdd.n6387 0.00334848
R14847 avdd.n6428 avdd.n6380 0.00334848
R14848 avdd.n6441 avdd.n6368 0.00334848
R14849 avdd.n6482 avdd.n6350 0.00334848
R14850 avdd.n6503 avdd.n6343 0.00334848
R14851 avdd.n6513 avdd.n6327 0.00334848
R14852 avdd.n6627 avdd.n6603 0.00334848
R14853 avdd.n6644 avdd.n6596 0.00334848
R14854 avdd.n6657 avdd.n6584 0.00334848
R14855 avdd.n6698 avdd.n6566 0.00334848
R14856 avdd.n6719 avdd.n6559 0.00334848
R14857 avdd.n6729 avdd.n6543 0.00334848
R14858 avdd.n6843 avdd.n6819 0.00334848
R14859 avdd.n6860 avdd.n6812 0.00334848
R14860 avdd.n6873 avdd.n6800 0.00334848
R14861 avdd.n6914 avdd.n6782 0.00334848
R14862 avdd.n6935 avdd.n6775 0.00334848
R14863 avdd.n6945 avdd.n6759 0.00334848
R14864 avdd.n7059 avdd.n7035 0.00334848
R14865 avdd.n7076 avdd.n7028 0.00334848
R14866 avdd.n7089 avdd.n7016 0.00334848
R14867 avdd.n7130 avdd.n6998 0.00334848
R14868 avdd.n7151 avdd.n6991 0.00334848
R14869 avdd.n7161 avdd.n6975 0.00334848
R14870 avdd.n7275 avdd.n7251 0.00334848
R14871 avdd.n7292 avdd.n7244 0.00334848
R14872 avdd.n7305 avdd.n7232 0.00334848
R14873 avdd.n7346 avdd.n7214 0.00334848
R14874 avdd.n7367 avdd.n7207 0.00334848
R14875 avdd.n7377 avdd.n7191 0.00334848
R14876 avdd.n7704 avdd.n7703 0.00334848
R14877 avdd.n7724 avdd.n7723 0.00334848
R14878 avdd.n7699 avdd.n7698 0.00334848
R14879 avdd.n7797 avdd.n7796 0.00334848
R14880 avdd.n7814 avdd.n7813 0.00334848
R14881 avdd.n7834 avdd.n7833 0.00334848
R14882 avdd.n10183 avdd.n10182 0.00334848
R14883 avdd.n10203 avdd.n10202 0.00334848
R14884 avdd.n10178 avdd.n10177 0.00334848
R14885 avdd.n10056 avdd.n10055 0.00334848
R14886 avdd.n10072 avdd.n10071 0.00334848
R14887 avdd.n10092 avdd.n10091 0.00334848
R14888 avdd.n9994 avdd.n9993 0.00334848
R14889 avdd.n10008 avdd.n10007 0.00334848
R14890 avdd.n9962 avdd.n9961 0.00334848
R14891 avdd.n10286 avdd.n10285 0.00334848
R14892 avdd.n10304 avdd.n10303 0.00334848
R14893 avdd.n10324 avdd.n10323 0.00334848
R14894 avdd.n9880 avdd.n9879 0.00334848
R14895 avdd.n9894 avdd.n9893 0.00334848
R14896 avdd.n9848 avdd.n9847 0.00334848
R14897 avdd.n10388 avdd.n10387 0.00334848
R14898 avdd.n10406 avdd.n10405 0.00334848
R14899 avdd.n10426 avdd.n10425 0.00334848
R14900 avdd.n9766 avdd.n9765 0.00334848
R14901 avdd.n9780 avdd.n9779 0.00334848
R14902 avdd.n9734 avdd.n9733 0.00334848
R14903 avdd.n10490 avdd.n10489 0.00334848
R14904 avdd.n10508 avdd.n10507 0.00334848
R14905 avdd.n10528 avdd.n10527 0.00334848
R14906 avdd.n9653 avdd.n9652 0.00334848
R14907 avdd.n9667 avdd.n9666 0.00334848
R14908 avdd.n9621 avdd.n9620 0.00334848
R14909 avdd.n10592 avdd.n10591 0.00334848
R14910 avdd.n10610 avdd.n10609 0.00334848
R14911 avdd.n10630 avdd.n10629 0.00334848
R14912 avdd.n9538 avdd.n9537 0.00334848
R14913 avdd.n9552 avdd.n9551 0.00334848
R14914 avdd.n9506 avdd.n9505 0.00334848
R14915 avdd.n10694 avdd.n10693 0.00334848
R14916 avdd.n10712 avdd.n10711 0.00334848
R14917 avdd.n10732 avdd.n10731 0.00334848
R14918 avdd.n9424 avdd.n9423 0.00334848
R14919 avdd.n9438 avdd.n9437 0.00334848
R14920 avdd.n9392 avdd.n9391 0.00334848
R14921 avdd.n10796 avdd.n10795 0.00334848
R14922 avdd.n10814 avdd.n10813 0.00334848
R14923 avdd.n10834 avdd.n10833 0.00334848
R14924 avdd.n9310 avdd.n9309 0.00334848
R14925 avdd.n9324 avdd.n9323 0.00334848
R14926 avdd.n9278 avdd.n9277 0.00334848
R14927 avdd.n10898 avdd.n10897 0.00334848
R14928 avdd.n10916 avdd.n10915 0.00334848
R14929 avdd.n10936 avdd.n10935 0.00334848
R14930 avdd.n9196 avdd.n9195 0.00334848
R14931 avdd.n9210 avdd.n9209 0.00334848
R14932 avdd.n9164 avdd.n9163 0.00334848
R14933 avdd.n11000 avdd.n10999 0.00334848
R14934 avdd.n11018 avdd.n11017 0.00334848
R14935 avdd.n11038 avdd.n11037 0.00334848
R14936 avdd.n9082 avdd.n9081 0.00334848
R14937 avdd.n9096 avdd.n9095 0.00334848
R14938 avdd.n9050 avdd.n9049 0.00334848
R14939 avdd.n11102 avdd.n11101 0.00334848
R14940 avdd.n11120 avdd.n11119 0.00334848
R14941 avdd.n11140 avdd.n11139 0.00334848
R14942 avdd.n8968 avdd.n8967 0.00334848
R14943 avdd.n8982 avdd.n8981 0.00334848
R14944 avdd.n8936 avdd.n8935 0.00334848
R14945 avdd.n11204 avdd.n11203 0.00334848
R14946 avdd.n11222 avdd.n11221 0.00334848
R14947 avdd.n11242 avdd.n11241 0.00334848
R14948 avdd.n98 avdd.n97 0.00334848
R14949 avdd.n119 avdd.n118 0.00334848
R14950 avdd.n182 avdd.n181 0.00334848
R14951 avdd.n8819 avdd.n8818 0.00334848
R14952 avdd.n8835 avdd.n8834 0.00334848
R14953 avdd.n8855 avdd.n8854 0.00334848
R14954 avdd.n228 avdd.n227 0.00334848
R14955 avdd.n249 avdd.n248 0.00334848
R14956 avdd.n312 avdd.n311 0.00334848
R14957 avdd.n8733 avdd.n8732 0.00334848
R14958 avdd.n8749 avdd.n8748 0.00334848
R14959 avdd.n8769 avdd.n8768 0.00334848
R14960 avdd.n358 avdd.n357 0.00334848
R14961 avdd.n379 avdd.n378 0.00334848
R14962 avdd.n442 avdd.n441 0.00334848
R14963 avdd.n8647 avdd.n8646 0.00334848
R14964 avdd.n8663 avdd.n8662 0.00334848
R14965 avdd.n8683 avdd.n8682 0.00334848
R14966 avdd.n488 avdd.n487 0.00334848
R14967 avdd.n509 avdd.n508 0.00334848
R14968 avdd.n572 avdd.n571 0.00334848
R14969 avdd.n8561 avdd.n8560 0.00334848
R14970 avdd.n8577 avdd.n8576 0.00334848
R14971 avdd.n8597 avdd.n8596 0.00334848
R14972 avdd.n618 avdd.n617 0.00334848
R14973 avdd.n639 avdd.n638 0.00334848
R14974 avdd.n702 avdd.n701 0.00334848
R14975 avdd.n8475 avdd.n8474 0.00334848
R14976 avdd.n8491 avdd.n8490 0.00334848
R14977 avdd.n8511 avdd.n8510 0.00334848
R14978 avdd.n748 avdd.n747 0.00334848
R14979 avdd.n769 avdd.n768 0.00334848
R14980 avdd.n832 avdd.n831 0.00334848
R14981 avdd.n8389 avdd.n8388 0.00334848
R14982 avdd.n8405 avdd.n8404 0.00334848
R14983 avdd.n8425 avdd.n8424 0.00334848
R14984 avdd.n878 avdd.n877 0.00334848
R14985 avdd.n899 avdd.n898 0.00334848
R14986 avdd.n962 avdd.n961 0.00334848
R14987 avdd.n8303 avdd.n8302 0.00334848
R14988 avdd.n8319 avdd.n8318 0.00334848
R14989 avdd.n8339 avdd.n8338 0.00334848
R14990 avdd.n1008 avdd.n1007 0.00334848
R14991 avdd.n1029 avdd.n1028 0.00334848
R14992 avdd.n1092 avdd.n1091 0.00334848
R14993 avdd.n8217 avdd.n8216 0.00334848
R14994 avdd.n8233 avdd.n8232 0.00334848
R14995 avdd.n8253 avdd.n8252 0.00334848
R14996 avdd.n1138 avdd.n1137 0.00334848
R14997 avdd.n1159 avdd.n1158 0.00334848
R14998 avdd.n1222 avdd.n1221 0.00334848
R14999 avdd.n8131 avdd.n8130 0.00334848
R15000 avdd.n8147 avdd.n8146 0.00334848
R15001 avdd.n8167 avdd.n8166 0.00334848
R15002 avdd.n1268 avdd.n1267 0.00334848
R15003 avdd.n1289 avdd.n1288 0.00334848
R15004 avdd.n1352 avdd.n1351 0.00334848
R15005 avdd.n8045 avdd.n8044 0.00334848
R15006 avdd.n8061 avdd.n8060 0.00334848
R15007 avdd.n8081 avdd.n8080 0.00334848
R15008 avdd.n1398 avdd.n1397 0.00334848
R15009 avdd.n1419 avdd.n1418 0.00334848
R15010 avdd.n1482 avdd.n1481 0.00334848
R15011 avdd.n7959 avdd.n7958 0.00334848
R15012 avdd.n7975 avdd.n7974 0.00334848
R15013 avdd.n7995 avdd.n7994 0.00334848
R15014 avdd.n1528 avdd.n1527 0.00334848
R15015 avdd.n1549 avdd.n1548 0.00334848
R15016 avdd.n1612 avdd.n1611 0.00334848
R15017 avdd.n7873 avdd.n7872 0.00334848
R15018 avdd.n7889 avdd.n7888 0.00334848
R15019 avdd.n7909 avdd.n7908 0.00334848
R15020 avdd.n2036 avdd.n2005 0.00334838
R15021 avdd.n2010 avdd.n2005 0.00334838
R15022 avdd.n2303 avdd.n2093 0.00334838
R15023 avdd.n2303 avdd.n2302 0.00334838
R15024 avdd.n2518 avdd.n2308 0.00334838
R15025 avdd.n2518 avdd.n2517 0.00334838
R15026 avdd.n2733 avdd.n2523 0.00334838
R15027 avdd.n2733 avdd.n2732 0.00334838
R15028 avdd.n2948 avdd.n2738 0.00334838
R15029 avdd.n2948 avdd.n2947 0.00334838
R15030 avdd.n3163 avdd.n2953 0.00334838
R15031 avdd.n3163 avdd.n3162 0.00334838
R15032 avdd.n3379 avdd.n3169 0.00334838
R15033 avdd.n3594 avdd.n3384 0.00334838
R15034 avdd.n3809 avdd.n3599 0.00334838
R15035 avdd.n4024 avdd.n3814 0.00334838
R15036 avdd.n4239 avdd.n4029 0.00334838
R15037 avdd.n4454 avdd.n4244 0.00334838
R15038 avdd.n5022 avdd.n5021 0.00334838
R15039 avdd.n5023 avdd.n5022 0.00334838
R15040 avdd.n5238 avdd.n5237 0.00334838
R15041 avdd.n5239 avdd.n5238 0.00334838
R15042 avdd.n5454 avdd.n5453 0.00334838
R15043 avdd.n5455 avdd.n5454 0.00334838
R15044 avdd.n5670 avdd.n5669 0.00334838
R15045 avdd.n5671 avdd.n5670 0.00334838
R15046 avdd.n5886 avdd.n5885 0.00334838
R15047 avdd.n5887 avdd.n5886 0.00334838
R15048 avdd.n6102 avdd.n6101 0.00334838
R15049 avdd.n6103 avdd.n6102 0.00334838
R15050 avdd.n6318 avdd.n6317 0.00334838
R15051 avdd.n6319 avdd.n6318 0.00334838
R15052 avdd.n6534 avdd.n6533 0.00334838
R15053 avdd.n6535 avdd.n6534 0.00334838
R15054 avdd.n6750 avdd.n6749 0.00334838
R15055 avdd.n6751 avdd.n6750 0.00334838
R15056 avdd.n6966 avdd.n6965 0.00334838
R15057 avdd.n6967 avdd.n6966 0.00334838
R15058 avdd.n7182 avdd.n7181 0.00334838
R15059 avdd.n7183 avdd.n7182 0.00334838
R15060 avdd.n7398 avdd.n7397 0.00334838
R15061 avdd.n7399 avdd.n7398 0.00334838
R15062 avdd.n7763 avdd.n7762 0.00334838
R15063 avdd.n7764 avdd.n7763 0.00334838
R15064 avdd.n7854 avdd.n7853 0.00334838
R15065 avdd.n7851 avdd.n7850 0.00334838
R15066 avdd.n7853 avdd.n7852 0.00334838
R15067 avdd.n7852 avdd.n7851 0.00334838
R15068 avdd.n10242 avdd.n10241 0.00334838
R15069 avdd.n10243 avdd.n10242 0.00334838
R15070 avdd.n10112 avdd.n10111 0.00334838
R15071 avdd.n10109 avdd.n10108 0.00334838
R15072 avdd.n10111 avdd.n10110 0.00334838
R15073 avdd.n10110 avdd.n10109 0.00334838
R15074 avdd.n10343 avdd.n10342 0.00334838
R15075 avdd.n10344 avdd.n10343 0.00334838
R15076 avdd.n10445 avdd.n10444 0.00334838
R15077 avdd.n10446 avdd.n10445 0.00334838
R15078 avdd.n10547 avdd.n10546 0.00334838
R15079 avdd.n10548 avdd.n10547 0.00334838
R15080 avdd.n10649 avdd.n10648 0.00334838
R15081 avdd.n10650 avdd.n10649 0.00334838
R15082 avdd.n10751 avdd.n10750 0.00334838
R15083 avdd.n10752 avdd.n10751 0.00334838
R15084 avdd.n10853 avdd.n10852 0.00334838
R15085 avdd.n10854 avdd.n10853 0.00334838
R15086 avdd.n10955 avdd.n10954 0.00334838
R15087 avdd.n10956 avdd.n10955 0.00334838
R15088 avdd.n11057 avdd.n11056 0.00334838
R15089 avdd.n11058 avdd.n11057 0.00334838
R15090 avdd.n11159 avdd.n11158 0.00334838
R15091 avdd.n11160 avdd.n11159 0.00334838
R15092 avdd.n11261 avdd.n11260 0.00334838
R15093 avdd.n11262 avdd.n11261 0.00334838
R15094 avdd.n8885 avdd.n8804 0.00334838
R15095 avdd.n8804 avdd.n8803 0.00334838
R15096 avdd.n8799 avdd.n8718 0.00334838
R15097 avdd.n8718 avdd.n8717 0.00334838
R15098 avdd.n8713 avdd.n8632 0.00334838
R15099 avdd.n8632 avdd.n8631 0.00334838
R15100 avdd.n8627 avdd.n8546 0.00334838
R15101 avdd.n8546 avdd.n8545 0.00334838
R15102 avdd.n8541 avdd.n8460 0.00334838
R15103 avdd.n8460 avdd.n8459 0.00334838
R15104 avdd.n8455 avdd.n8374 0.00334838
R15105 avdd.n8374 avdd.n8373 0.00334838
R15106 avdd.n8369 avdd.n8288 0.00334838
R15107 avdd.n8288 avdd.n8287 0.00334838
R15108 avdd.n8283 avdd.n8202 0.00334838
R15109 avdd.n8202 avdd.n8201 0.00334838
R15110 avdd.n8197 avdd.n8116 0.00334838
R15111 avdd.n8116 avdd.n8115 0.00334838
R15112 avdd.n8111 avdd.n8030 0.00334838
R15113 avdd.n8030 avdd.n8029 0.00334838
R15114 avdd.n8025 avdd.n7944 0.00334838
R15115 avdd.n7944 avdd.n7943 0.00334838
R15116 avdd.n7939 avdd.n7858 0.00334838
R15117 avdd.n7858 avdd.n7857 0.00334838
R15118 avdd.n7455 avdd.n7454 0.00310417
R15119 avdd.n7493 avdd.n7477 0.00310417
R15120 avdd.n7554 avdd.n7553 0.00310417
R15121 avdd.n7593 avdd.n7577 0.00310417
R15122 avdd.n1691 avdd.n1690 0.00310417
R15123 avdd.n1730 avdd.n1713 0.00310417
R15124 avdd.n1781 avdd.n1780 0.00310417
R15125 avdd.n1820 avdd.n1803 0.00310417
R15126 avdd.n2073 avdd.n2072 0.00263636
R15127 avdd.n2029 avdd.n2028 0.00263636
R15128 avdd.n2210 avdd.n2123 0.00263636
R15129 avdd.n2304 avdd.n2097 0.00263636
R15130 avdd.n2425 avdd.n2338 0.00263636
R15131 avdd.n2519 avdd.n2312 0.00263636
R15132 avdd.n2640 avdd.n2553 0.00263636
R15133 avdd.n2734 avdd.n2527 0.00263636
R15134 avdd.n2855 avdd.n2768 0.00263636
R15135 avdd.n2949 avdd.n2742 0.00263636
R15136 avdd.n3070 avdd.n2983 0.00263636
R15137 avdd.n3164 avdd.n2957 0.00263636
R15138 avdd.n3362 avdd.n3361 0.00263636
R15139 avdd.n3322 avdd.n3305 0.00263636
R15140 avdd.n3577 avdd.n3576 0.00263636
R15141 avdd.n3537 avdd.n3520 0.00263636
R15142 avdd.n3792 avdd.n3791 0.00263636
R15143 avdd.n3752 avdd.n3735 0.00263636
R15144 avdd.n4007 avdd.n4006 0.00263636
R15145 avdd.n3967 avdd.n3950 0.00263636
R15146 avdd.n4222 avdd.n4221 0.00263636
R15147 avdd.n4182 avdd.n4165 0.00263636
R15148 avdd.n4437 avdd.n4436 0.00263636
R15149 avdd.n4397 avdd.n4380 0.00263636
R15150 avdd.n4932 avdd.n4845 0.00263636
R15151 avdd.n5012 avdd.n4811 0.00263636
R15152 avdd.n5148 avdd.n5061 0.00263636
R15153 avdd.n5228 avdd.n5027 0.00263636
R15154 avdd.n5364 avdd.n5277 0.00263636
R15155 avdd.n5444 avdd.n5243 0.00263636
R15156 avdd.n5580 avdd.n5493 0.00263636
R15157 avdd.n5660 avdd.n5459 0.00263636
R15158 avdd.n5796 avdd.n5709 0.00263636
R15159 avdd.n5876 avdd.n5675 0.00263636
R15160 avdd.n6012 avdd.n5925 0.00263636
R15161 avdd.n6092 avdd.n5891 0.00263636
R15162 avdd.n6228 avdd.n6141 0.00263636
R15163 avdd.n6308 avdd.n6107 0.00263636
R15164 avdd.n6444 avdd.n6357 0.00263636
R15165 avdd.n6524 avdd.n6323 0.00263636
R15166 avdd.n6660 avdd.n6573 0.00263636
R15167 avdd.n6740 avdd.n6539 0.00263636
R15168 avdd.n6876 avdd.n6789 0.00263636
R15169 avdd.n6956 avdd.n6755 0.00263636
R15170 avdd.n7092 avdd.n7005 0.00263636
R15171 avdd.n7172 avdd.n6971 0.00263636
R15172 avdd.n7308 avdd.n7221 0.00263636
R15173 avdd.n7388 avdd.n7187 0.00263636
R15174 avdd.n7680 avdd.n7679 0.00263636
R15175 avdd.n7793 avdd.n7792 0.00263636
R15176 avdd.n10159 avdd.n10158 0.00263636
R15177 avdd.n10053 avdd.n10052 0.00263636
R15178 avdd.n9943 avdd.n9942 0.00263636
R15179 avdd.n10270 avdd.n10269 0.00263636
R15180 avdd.n9829 avdd.n9828 0.00263636
R15181 avdd.n10372 avdd.n10371 0.00263636
R15182 avdd.n9715 avdd.n9714 0.00263636
R15183 avdd.n10474 avdd.n10473 0.00263636
R15184 avdd.n9602 avdd.n9601 0.00263636
R15185 avdd.n10576 avdd.n10575 0.00263636
R15186 avdd.n9487 avdd.n9486 0.00263636
R15187 avdd.n10678 avdd.n10677 0.00263636
R15188 avdd.n9373 avdd.n9372 0.00263636
R15189 avdd.n10780 avdd.n10779 0.00263636
R15190 avdd.n9259 avdd.n9258 0.00263636
R15191 avdd.n10882 avdd.n10881 0.00263636
R15192 avdd.n9145 avdd.n9144 0.00263636
R15193 avdd.n10984 avdd.n10983 0.00263636
R15194 avdd.n9031 avdd.n9030 0.00263636
R15195 avdd.n11086 avdd.n11085 0.00263636
R15196 avdd.n8917 avdd.n8916 0.00263636
R15197 avdd.n11188 avdd.n11187 0.00263636
R15198 avdd.n163 avdd.n162 0.00263636
R15199 avdd.n8816 avdd.n8815 0.00263636
R15200 avdd.n293 avdd.n292 0.00263636
R15201 avdd.n8730 avdd.n8729 0.00263636
R15202 avdd.n423 avdd.n422 0.00263636
R15203 avdd.n8644 avdd.n8643 0.00263636
R15204 avdd.n553 avdd.n552 0.00263636
R15205 avdd.n8558 avdd.n8557 0.00263636
R15206 avdd.n683 avdd.n682 0.00263636
R15207 avdd.n8472 avdd.n8471 0.00263636
R15208 avdd.n813 avdd.n812 0.00263636
R15209 avdd.n8386 avdd.n8385 0.00263636
R15210 avdd.n943 avdd.n942 0.00263636
R15211 avdd.n8300 avdd.n8299 0.00263636
R15212 avdd.n1073 avdd.n1072 0.00263636
R15213 avdd.n8214 avdd.n8213 0.00263636
R15214 avdd.n1203 avdd.n1202 0.00263636
R15215 avdd.n8128 avdd.n8127 0.00263636
R15216 avdd.n1333 avdd.n1332 0.00263636
R15217 avdd.n8042 avdd.n8041 0.00263636
R15218 avdd.n1463 avdd.n1462 0.00263636
R15219 avdd.n7956 avdd.n7955 0.00263636
R15220 avdd.n1593 avdd.n1592 0.00263636
R15221 avdd.n7870 avdd.n7869 0.00263636
R15222 avdd.n4866 avdd.n4861 0.002423
R15223 avdd.n5082 avdd.n5077 0.002423
R15224 avdd.n5298 avdd.n5293 0.002423
R15225 avdd.n5514 avdd.n5509 0.002423
R15226 avdd.n5730 avdd.n5725 0.002423
R15227 avdd.n5946 avdd.n5941 0.002423
R15228 avdd.n6162 avdd.n6157 0.002423
R15229 avdd.n6378 avdd.n6373 0.002423
R15230 avdd.n6594 avdd.n6589 0.002423
R15231 avdd.n6810 avdd.n6805 0.002423
R15232 avdd.n7026 avdd.n7021 0.002423
R15233 avdd.n7242 avdd.n7237 0.002423
R15234 avdd.n10027 avdd.n10026 0.002423
R15235 avdd.n9913 avdd.n9912 0.002423
R15236 avdd.n9799 avdd.n9798 0.002423
R15237 avdd.n9685 avdd.n9684 0.002423
R15238 avdd.n9571 avdd.n9570 0.002423
R15239 avdd.n9457 avdd.n9456 0.002423
R15240 avdd.n9343 avdd.n9342 0.002423
R15241 avdd.n9229 avdd.n9228 0.002423
R15242 avdd.n9115 avdd.n9114 0.002423
R15243 avdd.n9001 avdd.n9000 0.002423
R15244 avdd.n2064 avdd.n1960 0.00192424
R15245 avdd.n1908 avdd.n1907 0.00192424
R15246 avdd.n1941 avdd.n1880 0.00192424
R15247 avdd.n2063 avdd.n1961 0.00192424
R15248 avdd.n2044 avdd.n1996 0.00192424
R15249 avdd.n2237 avdd.n2236 0.00192424
R15250 avdd.n2162 avdd.n2161 0.00192424
R15251 avdd.n2198 avdd.n2138 0.00192424
R15252 avdd.n2235 avdd.n2119 0.00192424
R15253 avdd.n2278 avdd.n2105 0.00192424
R15254 avdd.n2452 avdd.n2451 0.00192424
R15255 avdd.n2377 avdd.n2376 0.00192424
R15256 avdd.n2413 avdd.n2353 0.00192424
R15257 avdd.n2450 avdd.n2334 0.00192424
R15258 avdd.n2493 avdd.n2320 0.00192424
R15259 avdd.n2667 avdd.n2666 0.00192424
R15260 avdd.n2592 avdd.n2591 0.00192424
R15261 avdd.n2628 avdd.n2568 0.00192424
R15262 avdd.n2665 avdd.n2549 0.00192424
R15263 avdd.n2708 avdd.n2535 0.00192424
R15264 avdd.n2882 avdd.n2881 0.00192424
R15265 avdd.n2807 avdd.n2806 0.00192424
R15266 avdd.n2843 avdd.n2783 0.00192424
R15267 avdd.n2880 avdd.n2764 0.00192424
R15268 avdd.n2923 avdd.n2750 0.00192424
R15269 avdd.n3097 avdd.n3096 0.00192424
R15270 avdd.n3022 avdd.n3021 0.00192424
R15271 avdd.n3058 avdd.n2998 0.00192424
R15272 avdd.n3095 avdd.n2979 0.00192424
R15273 avdd.n3138 avdd.n2965 0.00192424
R15274 avdd.n3353 avdd.n3250 0.00192424
R15275 avdd.n3198 avdd.n3197 0.00192424
R15276 avdd.n3231 avdd.n3171 0.00192424
R15277 avdd.n3352 avdd.n3251 0.00192424
R15278 avdd.n3333 avdd.n3286 0.00192424
R15279 avdd.n3568 avdd.n3465 0.00192424
R15280 avdd.n3413 avdd.n3412 0.00192424
R15281 avdd.n3446 avdd.n3386 0.00192424
R15282 avdd.n3567 avdd.n3466 0.00192424
R15283 avdd.n3548 avdd.n3501 0.00192424
R15284 avdd.n3783 avdd.n3680 0.00192424
R15285 avdd.n3628 avdd.n3627 0.00192424
R15286 avdd.n3661 avdd.n3601 0.00192424
R15287 avdd.n3782 avdd.n3681 0.00192424
R15288 avdd.n3763 avdd.n3716 0.00192424
R15289 avdd.n3998 avdd.n3895 0.00192424
R15290 avdd.n3843 avdd.n3842 0.00192424
R15291 avdd.n3876 avdd.n3816 0.00192424
R15292 avdd.n3997 avdd.n3896 0.00192424
R15293 avdd.n3978 avdd.n3931 0.00192424
R15294 avdd.n4213 avdd.n4110 0.00192424
R15295 avdd.n4058 avdd.n4057 0.00192424
R15296 avdd.n4091 avdd.n4031 0.00192424
R15297 avdd.n4212 avdd.n4111 0.00192424
R15298 avdd.n4193 avdd.n4146 0.00192424
R15299 avdd.n4428 avdd.n4325 0.00192424
R15300 avdd.n4273 avdd.n4272 0.00192424
R15301 avdd.n4306 avdd.n4246 0.00192424
R15302 avdd.n4427 avdd.n4326 0.00192424
R15303 avdd.n4408 avdd.n4361 0.00192424
R15304 avdd.n4959 avdd.n4958 0.00192424
R15305 avdd.n4884 avdd.n4883 0.00192424
R15306 avdd.n4920 avdd.n4860 0.00192424
R15307 avdd.n4957 avdd.n4841 0.00192424
R15308 avdd.n4997 avdd.n4826 0.00192424
R15309 avdd.n5175 avdd.n5174 0.00192424
R15310 avdd.n5100 avdd.n5099 0.00192424
R15311 avdd.n5136 avdd.n5076 0.00192424
R15312 avdd.n5173 avdd.n5057 0.00192424
R15313 avdd.n5213 avdd.n5042 0.00192424
R15314 avdd.n5391 avdd.n5390 0.00192424
R15315 avdd.n5316 avdd.n5315 0.00192424
R15316 avdd.n5352 avdd.n5292 0.00192424
R15317 avdd.n5389 avdd.n5273 0.00192424
R15318 avdd.n5429 avdd.n5258 0.00192424
R15319 avdd.n5607 avdd.n5606 0.00192424
R15320 avdd.n5532 avdd.n5531 0.00192424
R15321 avdd.n5568 avdd.n5508 0.00192424
R15322 avdd.n5605 avdd.n5489 0.00192424
R15323 avdd.n5645 avdd.n5474 0.00192424
R15324 avdd.n5823 avdd.n5822 0.00192424
R15325 avdd.n5748 avdd.n5747 0.00192424
R15326 avdd.n5784 avdd.n5724 0.00192424
R15327 avdd.n5821 avdd.n5705 0.00192424
R15328 avdd.n5861 avdd.n5690 0.00192424
R15329 avdd.n6039 avdd.n6038 0.00192424
R15330 avdd.n5964 avdd.n5963 0.00192424
R15331 avdd.n6000 avdd.n5940 0.00192424
R15332 avdd.n6037 avdd.n5921 0.00192424
R15333 avdd.n6077 avdd.n5906 0.00192424
R15334 avdd.n6255 avdd.n6254 0.00192424
R15335 avdd.n6180 avdd.n6179 0.00192424
R15336 avdd.n6216 avdd.n6156 0.00192424
R15337 avdd.n6253 avdd.n6137 0.00192424
R15338 avdd.n6293 avdd.n6122 0.00192424
R15339 avdd.n6471 avdd.n6470 0.00192424
R15340 avdd.n6396 avdd.n6395 0.00192424
R15341 avdd.n6432 avdd.n6372 0.00192424
R15342 avdd.n6469 avdd.n6353 0.00192424
R15343 avdd.n6509 avdd.n6338 0.00192424
R15344 avdd.n6687 avdd.n6686 0.00192424
R15345 avdd.n6612 avdd.n6611 0.00192424
R15346 avdd.n6648 avdd.n6588 0.00192424
R15347 avdd.n6685 avdd.n6569 0.00192424
R15348 avdd.n6725 avdd.n6554 0.00192424
R15349 avdd.n6903 avdd.n6902 0.00192424
R15350 avdd.n6828 avdd.n6827 0.00192424
R15351 avdd.n6864 avdd.n6804 0.00192424
R15352 avdd.n6901 avdd.n6785 0.00192424
R15353 avdd.n6941 avdd.n6770 0.00192424
R15354 avdd.n7119 avdd.n7118 0.00192424
R15355 avdd.n7044 avdd.n7043 0.00192424
R15356 avdd.n7080 avdd.n7020 0.00192424
R15357 avdd.n7117 avdd.n7001 0.00192424
R15358 avdd.n7157 avdd.n6986 0.00192424
R15359 avdd.n7335 avdd.n7334 0.00192424
R15360 avdd.n7260 avdd.n7259 0.00192424
R15361 avdd.n7296 avdd.n7236 0.00192424
R15362 avdd.n7333 avdd.n7217 0.00192424
R15363 avdd.n7373 avdd.n7202 0.00192424
R15364 avdd.n7767 avdd.n7766 0.00192424
R15365 avdd.n7753 avdd.n7744 0.00192424
R15366 avdd.n7737 avdd.n7736 0.00192424
R15367 avdd.n7662 avdd.n7655 0.00192424
R15368 avdd.n7827 avdd.n7826 0.00192424
R15369 avdd.n10116 avdd.n10115 0.00192424
R15370 avdd.n10232 avdd.n10223 0.00192424
R15371 avdd.n10216 avdd.n10215 0.00192424
R15372 avdd.n10141 avdd.n10133 0.00192424
R15373 avdd.n10085 avdd.n10084 0.00192424
R15374 avdd.n9917 avdd.n9916 0.00192424
R15375 avdd.n9986 avdd.n9970 0.00192424
R15376 avdd.n10022 avdd.n10021 0.00192424
R15377 avdd.n10280 avdd.n10279 0.00192424
R15378 avdd.n10317 avdd.n10316 0.00192424
R15379 avdd.n9803 avdd.n9802 0.00192424
R15380 avdd.n9872 avdd.n9856 0.00192424
R15381 avdd.n9908 avdd.n9907 0.00192424
R15382 avdd.n10382 avdd.n10381 0.00192424
R15383 avdd.n10419 avdd.n10418 0.00192424
R15384 avdd.n9689 avdd.n9688 0.00192424
R15385 avdd.n9758 avdd.n9742 0.00192424
R15386 avdd.n9794 avdd.n9793 0.00192424
R15387 avdd.n10484 avdd.n10483 0.00192424
R15388 avdd.n10521 avdd.n10520 0.00192424
R15389 avdd.n9575 avdd.n9574 0.00192424
R15390 avdd.n9645 avdd.n9629 0.00192424
R15391 avdd.n9681 avdd.n9680 0.00192424
R15392 avdd.n10586 avdd.n10585 0.00192424
R15393 avdd.n10623 avdd.n10622 0.00192424
R15394 avdd.n9461 avdd.n9460 0.00192424
R15395 avdd.n9530 avdd.n9514 0.00192424
R15396 avdd.n9566 avdd.n9565 0.00192424
R15397 avdd.n10688 avdd.n10687 0.00192424
R15398 avdd.n10725 avdd.n10724 0.00192424
R15399 avdd.n9347 avdd.n9346 0.00192424
R15400 avdd.n9416 avdd.n9400 0.00192424
R15401 avdd.n9452 avdd.n9451 0.00192424
R15402 avdd.n10790 avdd.n10789 0.00192424
R15403 avdd.n10827 avdd.n10826 0.00192424
R15404 avdd.n9233 avdd.n9232 0.00192424
R15405 avdd.n9302 avdd.n9286 0.00192424
R15406 avdd.n9338 avdd.n9337 0.00192424
R15407 avdd.n10892 avdd.n10891 0.00192424
R15408 avdd.n10929 avdd.n10928 0.00192424
R15409 avdd.n9119 avdd.n9118 0.00192424
R15410 avdd.n9188 avdd.n9172 0.00192424
R15411 avdd.n9224 avdd.n9223 0.00192424
R15412 avdd.n10994 avdd.n10993 0.00192424
R15413 avdd.n11031 avdd.n11030 0.00192424
R15414 avdd.n9005 avdd.n9004 0.00192424
R15415 avdd.n9074 avdd.n9058 0.00192424
R15416 avdd.n9110 avdd.n9109 0.00192424
R15417 avdd.n11096 avdd.n11095 0.00192424
R15418 avdd.n11133 avdd.n11132 0.00192424
R15419 avdd.n8891 avdd.n8890 0.00192424
R15420 avdd.n8960 avdd.n8944 0.00192424
R15421 avdd.n8996 avdd.n8995 0.00192424
R15422 avdd.n11198 avdd.n11197 0.00192424
R15423 avdd.n11235 avdd.n11234 0.00192424
R15424 avdd.n60 avdd.n59 0.00192424
R15425 avdd.n86 avdd.n77 0.00192424
R15426 avdd.n132 avdd.n131 0.00192424
R15427 avdd.n145 avdd.n137 0.00192424
R15428 avdd.n8848 avdd.n8847 0.00192424
R15429 avdd.n190 avdd.n189 0.00192424
R15430 avdd.n216 avdd.n207 0.00192424
R15431 avdd.n262 avdd.n261 0.00192424
R15432 avdd.n275 avdd.n267 0.00192424
R15433 avdd.n8762 avdd.n8761 0.00192424
R15434 avdd.n320 avdd.n319 0.00192424
R15435 avdd.n346 avdd.n337 0.00192424
R15436 avdd.n392 avdd.n391 0.00192424
R15437 avdd.n405 avdd.n397 0.00192424
R15438 avdd.n8676 avdd.n8675 0.00192424
R15439 avdd.n450 avdd.n449 0.00192424
R15440 avdd.n476 avdd.n467 0.00192424
R15441 avdd.n522 avdd.n521 0.00192424
R15442 avdd.n535 avdd.n527 0.00192424
R15443 avdd.n8590 avdd.n8589 0.00192424
R15444 avdd.n580 avdd.n579 0.00192424
R15445 avdd.n606 avdd.n597 0.00192424
R15446 avdd.n652 avdd.n651 0.00192424
R15447 avdd.n665 avdd.n657 0.00192424
R15448 avdd.n8504 avdd.n8503 0.00192424
R15449 avdd.n710 avdd.n709 0.00192424
R15450 avdd.n736 avdd.n727 0.00192424
R15451 avdd.n782 avdd.n781 0.00192424
R15452 avdd.n795 avdd.n787 0.00192424
R15453 avdd.n8418 avdd.n8417 0.00192424
R15454 avdd.n840 avdd.n839 0.00192424
R15455 avdd.n866 avdd.n857 0.00192424
R15456 avdd.n912 avdd.n911 0.00192424
R15457 avdd.n925 avdd.n917 0.00192424
R15458 avdd.n8332 avdd.n8331 0.00192424
R15459 avdd.n970 avdd.n969 0.00192424
R15460 avdd.n996 avdd.n987 0.00192424
R15461 avdd.n1042 avdd.n1041 0.00192424
R15462 avdd.n1055 avdd.n1047 0.00192424
R15463 avdd.n8246 avdd.n8245 0.00192424
R15464 avdd.n1100 avdd.n1099 0.00192424
R15465 avdd.n1126 avdd.n1117 0.00192424
R15466 avdd.n1172 avdd.n1171 0.00192424
R15467 avdd.n1185 avdd.n1177 0.00192424
R15468 avdd.n8160 avdd.n8159 0.00192424
R15469 avdd.n1230 avdd.n1229 0.00192424
R15470 avdd.n1256 avdd.n1247 0.00192424
R15471 avdd.n1302 avdd.n1301 0.00192424
R15472 avdd.n1315 avdd.n1307 0.00192424
R15473 avdd.n8074 avdd.n8073 0.00192424
R15474 avdd.n1360 avdd.n1359 0.00192424
R15475 avdd.n1386 avdd.n1377 0.00192424
R15476 avdd.n1432 avdd.n1431 0.00192424
R15477 avdd.n1445 avdd.n1437 0.00192424
R15478 avdd.n7988 avdd.n7987 0.00192424
R15479 avdd.n1490 avdd.n1489 0.00192424
R15480 avdd.n1516 avdd.n1507 0.00192424
R15481 avdd.n1562 avdd.n1561 0.00192424
R15482 avdd.n1575 avdd.n1567 0.00192424
R15483 avdd.n7902 avdd.n7901 0.00192424
R15484 avdd.n1930 avdd.n1929 0.00121212
R15485 avdd.n1986 avdd.n1985 0.00121212
R15486 avdd.n2183 avdd.n2182 0.00121212
R15487 avdd.n2259 avdd.n2258 0.00121212
R15488 avdd.n2398 avdd.n2397 0.00121212
R15489 avdd.n2474 avdd.n2473 0.00121212
R15490 avdd.n2613 avdd.n2612 0.00121212
R15491 avdd.n2689 avdd.n2688 0.00121212
R15492 avdd.n2828 avdd.n2827 0.00121212
R15493 avdd.n2904 avdd.n2903 0.00121212
R15494 avdd.n3043 avdd.n3042 0.00121212
R15495 avdd.n3119 avdd.n3118 0.00121212
R15496 avdd.n3220 avdd.n3219 0.00121212
R15497 avdd.n3276 avdd.n3275 0.00121212
R15498 avdd.n3435 avdd.n3434 0.00121212
R15499 avdd.n3491 avdd.n3490 0.00121212
R15500 avdd.n3650 avdd.n3649 0.00121212
R15501 avdd.n3706 avdd.n3705 0.00121212
R15502 avdd.n3865 avdd.n3864 0.00121212
R15503 avdd.n3921 avdd.n3920 0.00121212
R15504 avdd.n4080 avdd.n4079 0.00121212
R15505 avdd.n4136 avdd.n4135 0.00121212
R15506 avdd.n4295 avdd.n4294 0.00121212
R15507 avdd.n4351 avdd.n4350 0.00121212
R15508 avdd.n4906 avdd.n4905 0.00121212
R15509 avdd.n4981 avdd.n4980 0.00121212
R15510 avdd.n5122 avdd.n5121 0.00121212
R15511 avdd.n5197 avdd.n5196 0.00121212
R15512 avdd.n5338 avdd.n5337 0.00121212
R15513 avdd.n5413 avdd.n5412 0.00121212
R15514 avdd.n5554 avdd.n5553 0.00121212
R15515 avdd.n5629 avdd.n5628 0.00121212
R15516 avdd.n5770 avdd.n5769 0.00121212
R15517 avdd.n5845 avdd.n5844 0.00121212
R15518 avdd.n5986 avdd.n5985 0.00121212
R15519 avdd.n6061 avdd.n6060 0.00121212
R15520 avdd.n6202 avdd.n6201 0.00121212
R15521 avdd.n6277 avdd.n6276 0.00121212
R15522 avdd.n6418 avdd.n6417 0.00121212
R15523 avdd.n6493 avdd.n6492 0.00121212
R15524 avdd.n6634 avdd.n6633 0.00121212
R15525 avdd.n6709 avdd.n6708 0.00121212
R15526 avdd.n6850 avdd.n6849 0.00121212
R15527 avdd.n6925 avdd.n6924 0.00121212
R15528 avdd.n7066 avdd.n7065 0.00121212
R15529 avdd.n7141 avdd.n7140 0.00121212
R15530 avdd.n7282 avdd.n7281 0.00121212
R15531 avdd.n7357 avdd.n7356 0.00121212
R15532 avdd.n7719 avdd.n7718 0.00121212
R15533 avdd.n7808 avdd.n7807 0.00121212
R15534 avdd.n10198 avdd.n10197 0.00121212
R15535 avdd.n10066 avdd.n10065 0.00121212
R15536 avdd.n10003 avdd.n10001 0.00121212
R15537 avdd.n10298 avdd.n10297 0.00121212
R15538 avdd.n9889 avdd.n9887 0.00121212
R15539 avdd.n10400 avdd.n10399 0.00121212
R15540 avdd.n9775 avdd.n9773 0.00121212
R15541 avdd.n10502 avdd.n10501 0.00121212
R15542 avdd.n9662 avdd.n9660 0.00121212
R15543 avdd.n10604 avdd.n10603 0.00121212
R15544 avdd.n9547 avdd.n9545 0.00121212
R15545 avdd.n10706 avdd.n10705 0.00121212
R15546 avdd.n9433 avdd.n9431 0.00121212
R15547 avdd.n10808 avdd.n10807 0.00121212
R15548 avdd.n9319 avdd.n9317 0.00121212
R15549 avdd.n10910 avdd.n10909 0.00121212
R15550 avdd.n9205 avdd.n9203 0.00121212
R15551 avdd.n11012 avdd.n11011 0.00121212
R15552 avdd.n9091 avdd.n9089 0.00121212
R15553 avdd.n11114 avdd.n11113 0.00121212
R15554 avdd.n8977 avdd.n8975 0.00121212
R15555 avdd.n11216 avdd.n11215 0.00121212
R15556 avdd.n113 avdd.n112 0.00121212
R15557 avdd.n8829 avdd.n8828 0.00121212
R15558 avdd.n243 avdd.n242 0.00121212
R15559 avdd.n8743 avdd.n8742 0.00121212
R15560 avdd.n373 avdd.n372 0.00121212
R15561 avdd.n8657 avdd.n8656 0.00121212
R15562 avdd.n503 avdd.n502 0.00121212
R15563 avdd.n8571 avdd.n8570 0.00121212
R15564 avdd.n633 avdd.n632 0.00121212
R15565 avdd.n8485 avdd.n8484 0.00121212
R15566 avdd.n763 avdd.n762 0.00121212
R15567 avdd.n8399 avdd.n8398 0.00121212
R15568 avdd.n893 avdd.n892 0.00121212
R15569 avdd.n8313 avdd.n8312 0.00121212
R15570 avdd.n1023 avdd.n1022 0.00121212
R15571 avdd.n8227 avdd.n8226 0.00121212
R15572 avdd.n1153 avdd.n1152 0.00121212
R15573 avdd.n8141 avdd.n8140 0.00121212
R15574 avdd.n1283 avdd.n1282 0.00121212
R15575 avdd.n8055 avdd.n8054 0.00121212
R15576 avdd.n1413 avdd.n1412 0.00121212
R15577 avdd.n7969 avdd.n7968 0.00121212
R15578 avdd.n1543 avdd.n1542 0.00121212
R15579 avdd.n7883 avdd.n7882 0.00121212
R15580 avdd.n1815 avdd.n1814 0.00101841
R15581 avdd.n1641 avdd.n1640 0.00101841
R15582 avdd.n1725 avdd.n1724 0.00101841
R15583 avdd.n1677 avdd.n1676 0.00101841
R15584 avdd.n4762 avdd.n4759 0.000773431
R15585 trim4.n7 trim4.n6 280.8
R15586 trim4.n0 trim4.t2 135.841
R15587 trim4.n2 trim4.t7 135.841
R15588 trim4.n2 trim4.t6 135.52
R15589 trim4.n3 trim4.t3 135.52
R15590 trim4.n4 trim4.t0 135.52
R15591 trim4.n5 trim4.t4 135.52
R15592 trim4.n1 trim4.t1 135.52
R15593 trim4.n0 trim4.t5 135.52
R15594 trim4.n7 trim4 0.593172
R15595 trim4.n1 trim4.n0 0.321152
R15596 trim4.n5 trim4.n4 0.321152
R15597 trim4.n4 trim4.n3 0.321152
R15598 trim4.n3 trim4.n2 0.321152
R15599 trim4 trim4.n7 0.188
R15600 trim4.n6 trim4.n1 0.163543
R15601 trim4.n6 trim4.n5 0.158109
R15602 avss.n3491 avss.n3182 234681
R15603 avss.n3144 avss.n2621 49090.1
R15604 avss.n3144 avss.n2620 49075.8
R15605 avss.n2804 avss.n2803 9913.74
R15606 avss.n2915 avss.n2627 9913.74
R15607 avss.n2652 avss.n2651 9913.74
R15608 avss.n2677 avss.n2676 9913.74
R15609 avss.n2921 avss.n2920 9907.94
R15610 avss.n2971 avss.n2970 9907.94
R15611 avss.n3028 avss.n3023 9907.94
R15612 avss.n3620 avss.n2614 9907.94
R15613 avss.n3143 avss.n2622 6110.51
R15614 avss.n3142 avss.n2917 6110.51
R15615 avss.n3142 avss.n3141 6110.51
R15616 avss.n3143 avss.n2623 6110.51
R15617 avss.n2618 avss.n2615 6110.51
R15618 avss.n2801 avss.n2618 6110.51
R15619 avss.n2924 avss.n2921 5290.03
R15620 avss.n2970 avss.n2967 5290.03
R15621 avss.n3025 avss.n3023 5290.03
R15622 avss.n3617 avss.n2614 5290.03
R15623 avss.n2803 avss.n2797 5290.03
R15624 avss.n2798 avss.n2627 5290.03
R15625 avss.n2651 avss.n2649 5290.03
R15626 avss.n2680 avss.n2677 5290.03
R15627 avss.n3139 avss.n2924 5162.56
R15628 avss.n2967 avss.n2966 5162.56
R15629 avss.n3026 avss.n3025 5162.56
R15630 avss.n3618 avss.n3617 5162.56
R15631 avss.n2806 avss.n2797 5156.76
R15632 avss.n2798 avss.n2626 5156.76
R15633 avss.n2654 avss.n2649 5156.76
R15634 avss.n2681 avss.n2680 5156.76
R15635 avss.n3614 avss.n2616 4871.71
R15636 avss.n3615 avss.n3614 4871.71
R15637 avss.n3614 avss.n2618 2462.31
R15638 avss.n3332 avss.n3331 2404.56
R15639 avss.n3493 avss.n3181 2404.56
R15640 avss.n3498 avss.n3497 2219.15
R15641 avss.n3327 avss.n3300 2195.97
R15642 avss.n2653 avss.n2622 2038.64
R15643 avss.n2917 avss.n2916 2038.64
R15644 avss.n2805 avss.n2801 2038.64
R15645 avss.n3027 avss.n2623 2038.64
R15646 avss.n3141 avss.n3140 2038.64
R15647 avss.n3619 avss.n2615 2038.64
R15648 avss.n2678 avss.n2622 2015.03
R15649 avss.n2917 avss.n2624 2015.03
R15650 avss.n2801 avss.n2800 2015.03
R15651 avss.n2969 avss.n2623 2015.03
R15652 avss.n3141 avss.n2918 2015.03
R15653 avss.n2922 avss.n2615 2015.03
R15654 avss.n3614 avss.n2617 1893.81
R15655 avss.n3614 avss.n3613 1879.36
R15656 avss.n3248 avss.n2619 1734.87
R15657 avss.n3143 avss.n3142 1653.87
R15658 avss.n3142 avss.n2618 1653.87
R15659 avss.n3144 avss.n3143 1478.42
R15660 avss.t204 avss.n2621 1361.72
R15661 avss.t211 avss.n2678 1361.72
R15662 avss.n2653 avss.t274 1361.72
R15663 avss.t266 avss.n2624 1361.72
R15664 avss.n2916 avss.t253 1361.72
R15665 avss.n2800 avss.t249 1361.72
R15666 avss.n2805 avss.t76 1361.72
R15667 avss.t83 avss.n2616 1361.72
R15668 avss.t150 avss.n2620 1361.72
R15669 avss.n2969 avss.t157 1361.72
R15670 avss.n3027 avss.t357 1361.72
R15671 avss.t349 avss.n2918 1361.72
R15672 avss.n3140 avss.t327 1361.72
R15673 avss.t323 avss.n2922 1361.72
R15674 avss.n3619 avss.t140 1361.72
R15675 avss.t147 avss.n3615 1361.72
R15676 avss.t205 avss.t204 928.802
R15677 avss.t209 avss.t205 928.802
R15678 avss.t206 avss.t209 928.802
R15679 avss.t210 avss.t206 928.802
R15680 avss.t207 avss.t202 928.802
R15681 avss.t202 avss.t208 928.802
R15682 avss.t208 avss.t203 928.802
R15683 avss.t203 avss.t211 928.802
R15684 avss.t274 avss.t270 928.802
R15685 avss.t270 avss.t267 928.802
R15686 avss.t267 avss.t272 928.802
R15687 avss.t272 avss.t268 928.802
R15688 avss.t265 avss.t273 928.802
R15689 avss.t273 avss.t269 928.802
R15690 avss.t269 avss.t271 928.802
R15691 avss.t271 avss.t266 928.802
R15692 avss.t247 avss.t253 928.802
R15693 avss.t248 avss.t247 928.802
R15694 avss.t254 avss.t248 928.802
R15695 avss.t250 avss.t254 928.802
R15696 avss.t251 avss.t255 928.802
R15697 avss.t256 avss.t251 928.802
R15698 avss.t252 avss.t256 928.802
R15699 avss.t249 avss.t252 928.802
R15700 avss.t76 avss.t81 928.802
R15701 avss.t81 avss.t77 928.802
R15702 avss.t77 avss.t78 928.802
R15703 avss.t78 avss.t74 928.802
R15704 avss.t79 avss.t82 928.802
R15705 avss.t82 avss.t80 928.802
R15706 avss.t80 avss.t75 928.802
R15707 avss.t75 avss.t83 928.802
R15708 avss.t151 avss.t150 928.802
R15709 avss.t155 avss.t151 928.802
R15710 avss.t152 avss.t155 928.802
R15711 avss.t156 avss.t152 928.802
R15712 avss.t158 avss.t153 928.802
R15713 avss.t154 avss.t158 928.802
R15714 avss.t149 avss.t154 928.802
R15715 avss.t157 avss.t149 928.802
R15716 avss.t353 avss.t357 928.802
R15717 avss.t350 avss.t353 928.802
R15718 avss.t355 avss.t350 928.802
R15719 avss.t351 avss.t355 928.802
R15720 avss.t358 avss.t356 928.802
R15721 avss.t356 avss.t352 928.802
R15722 avss.t352 avss.t354 928.802
R15723 avss.t354 avss.t349 928.802
R15724 avss.t331 avss.t327 928.802
R15725 avss.t332 avss.t331 928.802
R15726 avss.t328 avss.t332 928.802
R15727 avss.t324 avss.t328 928.802
R15728 avss.t329 avss.t325 928.802
R15729 avss.t325 avss.t330 928.802
R15730 avss.t330 avss.t326 928.802
R15731 avss.t326 avss.t323 928.802
R15732 avss.t145 avss.t140 928.802
R15733 avss.t141 avss.t145 928.802
R15734 avss.t142 avss.t141 928.802
R15735 avss.t148 avss.t142 928.802
R15736 avss.t143 avss.t146 928.802
R15737 avss.t146 avss.t144 928.802
R15738 avss.t144 avss.t139 928.802
R15739 avss.t139 avss.t147 928.802
R15740 avss.n3245 avss.t228 803.125
R15741 avss.n3608 avss.n3148 705.89
R15742 avss.n3609 avss.n3608 705.876
R15743 avss avss.n3600 649.827
R15744 avss.n2676 avss.n2621 585
R15745 avss.n2653 avss.n2652 585
R15746 avss.n2916 avss.n2915 585
R15747 avss.n2805 avss.n2804 585
R15748 avss.n3620 avss.n3619 585
R15749 avss.n3028 avss.n3027 585
R15750 avss.n2971 avss.n2620 585
R15751 avss.n3140 avss.n2920 585
R15752 avss.n3213 avss.n3209 585
R15753 avss.n3209 avss.n3207 585
R15754 avss.n3244 avss.n3243 585
R15755 avss.n3400 avss.n3244 585
R15756 avss.n3403 avss.n3402 585
R15757 avss.n3402 avss.n3401 585
R15758 avss.n3419 avss.n3237 585
R15759 avss.n3237 avss.n3235 585
R15760 avss.n3421 avss.n3420 585
R15761 avss.n3422 avss.n3421 585
R15762 avss.n3410 avss.n3227 585
R15763 avss.n3429 avss.n3227 585
R15764 avss.n3241 avss.n3230 585
R15765 avss.n3428 avss.n3230 585
R15766 avss.n3228 avss.n3226 585
R15767 avss.n3430 avss.n3228 585
R15768 avss.n3222 avss.n3221 585
R15769 avss.n3221 avss.n3220 585
R15770 avss.n3212 avss.n3211 585
R15771 avss.n3211 avss.n3205 585
R15772 avss.n3203 avss.n3201 585
R15773 avss.n3448 avss.n3203 585
R15774 avss.n3215 avss.n3214 585
R15775 avss.n3216 avss.n3215 585
R15776 avss.n3474 avss.n3192 585
R15777 avss.n3192 avss.n3190 585
R15778 avss.n3473 avss.n3472 585
R15779 avss.n3472 avss.n3471 585
R15780 avss.n3520 avss.n3519 585
R15781 avss.n3521 avss.n3520 585
R15782 avss.n3518 avss.n3170 585
R15783 avss.n3282 avss.n3281 585
R15784 avss.n3359 avss.n3288 585
R15785 avss.n3376 avss.n3375 585
R15786 avss.n3374 avss.n3279 585
R15787 avss.n3374 avss.n3275 585
R15788 avss.n3384 avss.n3274 585
R15789 avss.n3387 avss.n3386 585
R15790 avss.n3356 avss.n3355 585
R15791 avss.n3290 avss.n3289 585
R15792 avss.n3289 avss.n3275 585
R15793 avss avss.n3602 547.423
R15794 avss.n3611 avss.n3610 516.596
R15795 avss.n3147 avss.n3146 495.408
R15796 avss.n2679 avss.t210 464.401
R15797 avss.n2679 avss.t207 464.401
R15798 avss.t268 avss.n2650 464.401
R15799 avss.n2650 avss.t265 464.401
R15800 avss.n2799 avss.t250 464.401
R15801 avss.t255 avss.n2799 464.401
R15802 avss.t74 avss.n2802 464.401
R15803 avss.n2802 avss.t79 464.401
R15804 avss.n2968 avss.t156 464.401
R15805 avss.t153 avss.n2968 464.401
R15806 avss.n3024 avss.t351 464.401
R15807 avss.n3024 avss.t358 464.401
R15808 avss.n2923 avss.t324 464.401
R15809 avss.n2923 avss.t329 464.401
R15810 avss.n3616 avss.t148 464.401
R15811 avss.n3616 avss.t143 464.401
R15812 avss.n3177 avss.n3162 427.507
R15813 avss.n3327 avss.n3298 394
R15814 avss.n3331 avss.n3298 394
R15815 avss.n3322 avss.n3321 394
R15816 avss.n3319 avss.n3303 394
R15817 avss.n3315 avss.n3314 394
R15818 avss.n3312 avss.n3306 394
R15819 avss.n3308 avss.n3233 394
R15820 avss.n3423 avss.n3233 394
R15821 avss.n3423 avss.n3231 394
R15822 avss.n3427 avss.n3231 394
R15823 avss.n3427 avss.n3219 394
R15824 avss.n3442 avss.n3219 394
R15825 avss.n3442 avss.n3206 394
R15826 avss.n3447 avss.n3206 394
R15827 avss.n3447 avss.n3217 394
R15828 avss.n3217 avss.n3188 394
R15829 avss.n3478 avss.n3188 394
R15830 avss.n3478 avss.n3186 394
R15831 avss.n3489 avss.n3186 394
R15832 avss.n3485 avss.n3185 394
R15833 avss.n3483 avss.n3482 394
R15834 avss.n3493 avss.n3179 394
R15835 avss.n3497 avss.n3179 394
R15836 avss.n3440 avss.n3202 394
R15837 avss.n3476 avss.n3191 394
R15838 avss.n3504 avss.n3167 394
R15839 avss.n3502 avss.n3501 394
R15840 avss.n3440 avss.n3221 370.825
R15841 avss.n3211 avss.n3209 370.825
R15842 avss.n3476 avss.n3192 370.825
R15843 avss.n3417 avss.n3237 359.236
R15844 avss.n3386 avss.n3269 347.647
R15845 avss.n3371 avss.n3281 336.06
R15846 avss.n3254 avss.n3252 325.935
R15847 avss.n3535 avss.n3534 325.935
R15848 avss.n3602 avss.n3601 321.488
R15849 avss.n3398 avss.n3269 318.676
R15850 avss.n3601 avss.n3539 309.844
R15851 avss.n3402 avss.n3236 307.089
R15852 avss.n3417 avss.n3415 307.089
R15853 avss.n3432 avss.n3227 307.089
R15854 avss.n3450 avss.n3202 307.089
R15855 avss.n3210 avss.n3191 307.089
R15856 avss.n3520 avss.n3169 307.089
R15857 avss.n3516 avss.n3167 307.089
R15858 avss.n3602 avss 306.606
R15859 avss.n3604 avss.n3603 293.966
R15860 avss.n3418 avss.n3417 292.5
R15861 avss.n3417 avss.n3416 292.5
R15862 avss.n3440 avss.n3439 292.5
R15863 avss.n3441 avss.n3440 292.5
R15864 avss.n3223 avss.n3202 292.5
R15865 avss.n3204 avss.n3202 292.5
R15866 avss.n3459 avss.n3191 292.5
R15867 avss.n3191 avss.n3189 292.5
R15868 avss.n3476 avss.n3475 292.5
R15869 avss.n3477 avss.n3476 292.5
R15870 avss.n3233 avss.n3232 292.5
R15871 avss.n3400 avss.n3233 292.5
R15872 avss.n3424 avss.n3423 292.5
R15873 avss.n3423 avss.n3422 292.5
R15874 avss.n3425 avss.n3231 292.5
R15875 avss.n3416 avss.n3231 292.5
R15876 avss.n3427 avss.n3426 292.5
R15877 avss.n3428 avss.n3427 292.5
R15878 avss.n3219 avss.n3218 292.5
R15879 avss.n3430 avss.n3219 292.5
R15880 avss.n3443 avss.n3442 292.5
R15881 avss.n3442 avss.n3441 292.5
R15882 avss.n3444 avss.n3206 292.5
R15883 avss.n3206 avss.n3204 292.5
R15884 avss.n3447 avss.n3446 292.5
R15885 avss.n3448 avss.n3447 292.5
R15886 avss.n3445 avss.n3217 292.5
R15887 avss.n3217 avss.n3216 292.5
R15888 avss.n3188 avss.n3187 292.5
R15889 avss.n3189 avss.n3188 292.5
R15890 avss.n3479 avss.n3478 292.5
R15891 avss.n3478 avss.n3477 292.5
R15892 avss.n3480 avss.n3186 292.5
R15893 avss.n3471 avss.n3186 292.5
R15894 avss.n3499 avss.n3498 292.5
R15895 avss.n3501 avss.n3500 292.5
R15896 avss.n3503 avss.n3502 292.5
R15897 avss.n3505 avss.n3504 292.5
R15898 avss.n3521 avss.n3167 292.5
R15899 avss.n3506 avss.n3167 292.5
R15900 avss.n3489 avss.n3488 292.5
R15901 avss.n3487 avss.n3185 292.5
R15902 avss.n3486 avss.n3485 292.5
R15903 avss.n3484 avss.n3483 292.5
R15904 avss.n3482 avss.n3481 292.5
R15905 avss.n3181 avss.n3180 292.5
R15906 avss.n3494 avss.n3493 292.5
R15907 avss.n3493 avss.n3492 292.5
R15908 avss.n3495 avss.n3179 292.5
R15909 avss.n3179 avss.n3178 292.5
R15910 avss.n3497 avss.n3496 292.5
R15911 avss.n3497 avss.n3164 292.5
R15912 avss.n3371 avss.n3370 292.5
R15913 avss.n3388 avss.n3269 292.5
R15914 avss.n3275 avss.n3269 292.5
R15915 avss.n3342 avss.n3341 292.5
R15916 avss.n3335 avss.n3334 292.5
R15917 avss.n3332 avss.n3297 292.5
R15918 avss.n3331 avss.n3299 292.5
R15919 avss.n3331 avss.n3330 292.5
R15920 avss.n3325 avss.n3298 292.5
R15921 avss.n3329 avss.n3298 292.5
R15922 avss.n3327 avss.n3326 292.5
R15923 avss.n3328 avss.n3327 292.5
R15924 avss.n3324 avss.n3300 292.5
R15925 avss.n3323 avss.n3322 292.5
R15926 avss.n3321 avss.n3301 292.5
R15927 avss.n3319 avss.n3318 292.5
R15928 avss.n3317 avss.n3303 292.5
R15929 avss.n3316 avss.n3315 292.5
R15930 avss.n3314 avss.n3304 292.5
R15931 avss.n3312 avss.n3311 292.5
R15932 avss.n3310 avss.n3306 292.5
R15933 avss.n3309 avss.n3308 292.5
R15934 avss.n3148 avss 292.175
R15935 avss.n3147 avss 292.175
R15936 avss.n3610 avss 290.204
R15937 avss.n3609 avss 290.204
R15938 avss.n3613 avss 283.469
R15939 avss.n3612 avss 283.469
R15940 avss.n2617 avss 283.204
R15941 avss.n3145 avss 283.204
R15942 avss.n3608 avss.t307 283.147
R15943 avss.n3385 avss.n3275 281.354
R15944 avss.n3358 avss.n3275 278.7
R15945 avss.n3263 avss.n3262 271.844
R15946 avss.n3264 avss.n3257 267.671
R15947 avss.n3530 avss.n3160 267.671
R15948 avss.t188 avss.t259 237.5
R15949 avss.t200 avss.t129 235.494
R15950 avss avss.t54 220.53
R15951 avss avss.t51 220.53
R15952 avss avss.t11 220.53
R15953 avss avss.t31 220.53
R15954 avss.n3296 avss.n3275 218.815
R15955 avss.t17 avss 215.286
R15956 avss.t37 avss 215.286
R15957 avss.t40 avss 215.286
R15958 avss.t14 avss 215.286
R15959 avss.n3343 avss.n3342 213.625
R15960 avss.n11630 avss.t420 212.081
R15961 avss.n11629 avss.t413 212.081
R15962 avss.n3611 avss.n2619 205.958
R15963 avss.n3146 avss.n2619 205.736
R15964 avss.n3529 avss.n3162 200.185
R15965 avss.n3375 avss.n3276 199.3
R15966 avss.n3357 avss.n3356 199.3
R15967 avss.n2991 avss.t106 193.933
R15968 avss.n2950 avss.t114 193.933
R15969 avss.n3048 avss.t278 193.933
R15970 avss.n2934 avss.t215 193.933
R15971 avss.n3120 avss.t312 193.933
R15972 avss.n3113 avss.t126 193.933
R15973 avss.n3640 avss.t346 193.933
R15974 avss.n2600 avss.t408 193.933
R15975 avss.n2703 avss.t136 193.933
R15976 avss.n2663 avss.t124 193.933
R15977 avss.n2748 avss.t221 193.933
R15978 avss.n2636 avss.t290 193.933
R15979 avss.n2894 avss.t102 193.933
R15980 avss.n2887 avss.t406 193.933
R15981 avss.n2854 avss.t386 193.933
R15982 avss.n2847 avss.t195 193.933
R15983 avss.n2985 avss.t108 192.982
R15984 avss.n2953 avss.t217 192.982
R15985 avss.n3042 avss.t276 192.982
R15986 avss.n2937 avss.t197 192.982
R15987 avss.n3126 avss.t316 192.982
R15988 avss.n3119 avss.t336 192.982
R15989 avss.n3634 avss.t344 192.982
R15990 avss.n2603 avss.t69 192.982
R15991 avss.n2697 avss.t132 192.982
R15992 avss.n2666 avss.t402 192.982
R15993 avss.n2742 avss.t225 192.982
R15994 avss.n2639 avss.t162 192.982
R15995 avss.n2900 avss.t100 192.982
R15996 avss.n2893 avss.t116 192.982
R15997 avss.n2860 avss.t384 192.982
R15998 avss.n2853 avss.t334 192.982
R15999 avss.t54 avss 189.266
R16000 avss.t51 avss 189.266
R16001 avss.t11 avss 189.266
R16002 avss.t31 avss 189.266
R16003 avss avss.t17 184.764
R16004 avss avss.t37 184.764
R16005 avss avss.t40 184.764
R16006 avss avss.t14 184.764
R16007 avss.n2980 avss.t425 183.082
R16008 avss.n3037 avss.t412 183.082
R16009 avss.n3078 avss.t418 183.082
R16010 avss.n3629 avss.t419 183.082
R16011 avss.n2692 avss.t411 183.082
R16012 avss.n2737 avss.t417 183.082
R16013 avss.n2776 avss.t423 183.082
R16014 avss.n2812 avss.t424 183.082
R16015 avss.n3334 avss.n3333 181.275
R16016 avss.n3441 avss.n3204 170.387
R16017 avss.n3477 avss.n3189 170.387
R16018 avss.t187 avss.n3248 165.109
R16019 avss.n3441 avss.n3220 160.364
R16020 avss.n3477 avss.n3190 160.364
R16021 avss.n3299 avss.n3297 156.236
R16022 avss.n3494 avss.n3180 156.236
R16023 avss.n3416 avss.n3235 155.353
R16024 avss.n3372 avss.n3371 152.838
R16025 avss.n3342 avss.n3296 147.374
R16026 avss.n3334 avss.n3296 147.374
R16027 avss.n3326 avss.n3324 142.683
R16028 avss.n11630 avss.t239 139.78
R16029 avss.n11629 avss.t242 139.78
R16030 avss.t173 avss.n3525 137.88
R16031 avss.n3267 avss.t395 136.714
R16032 avss.n3249 avss.n3247 136.405
R16033 avss.n3333 avss.n3275 134.577
R16034 avss.n3264 avss.n3263 134.4
R16035 avss.n3530 avss.n3529 134.4
R16036 avss.n3416 avss.n3229 132.803
R16037 avss.n3431 avss.n3429 132.803
R16038 avss.n3449 avss.n3204 132.803
R16039 avss.n3208 avss.n3189 132.803
R16040 avss.n3145 avss.t8 126.748
R16041 avss.n3526 avss.t64 126.136
R16042 avss.n3207 avss.t179 125.285
R16043 avss.n3266 avss.t119 125.07
R16044 avss.n3662 avss.n3661 124.692
R16045 avss.n3101 avss.n3100 124.692
R16046 avss.n3071 avss.n3069 124.692
R16047 avss.n3013 avss.n3012 124.692
R16048 avss.n2835 avss.n2834 124.692
R16049 avss.n2875 avss.n2874 124.692
R16050 avss.n2770 avss.n2769 124.692
R16051 avss.n2725 avss.n2724 124.692
R16052 avss.t57 avss.n3612 123.77
R16053 avss.n2595 avss.t16 121.956
R16054 avss.n3651 avss.t15 121.956
R16055 avss.n2609 avss.t46 121.956
R16056 avss.n2607 avss.t47 121.956
R16057 avss.n3099 avss.t42 121.956
R16058 avss.n3088 avss.t41 121.956
R16059 avss.n3077 avss.t21 121.956
R16060 avss.n3079 avss.t22 121.956
R16061 avss.n3070 avss.t39 121.956
R16062 avss.n3059 avss.t38 121.956
R16063 avss.n2943 avss.t35 121.956
R16064 avss.n2941 avss.t36 121.956
R16065 avss.n2945 avss.t19 121.956
R16066 avss.n3002 avss.t18 121.956
R16067 avss.n2959 avss.t58 121.956
R16068 avss.n2957 avss.t59 121.956
R16069 avss.n2833 avss.t33 121.956
R16070 avss.n2822 avss.t32 121.956
R16071 avss.n2813 avss.t27 121.956
R16072 avss.n2811 avss.t26 121.956
R16073 avss.n2873 avss.t13 121.956
R16074 avss.n2786 avss.t12 121.956
R16075 avss.n2777 avss.t30 121.956
R16076 avss.n2907 avss.t29 121.956
R16077 avss.n2631 avss.t53 121.956
R16078 avss.n2759 avss.t52 121.956
R16079 avss.n2643 avss.t50 121.956
R16080 avss.n2645 avss.t49 121.956
R16081 avss.n2658 avss.t56 121.956
R16082 avss.n2714 avss.t55 121.956
R16083 avss.n2670 avss.t10 121.956
R16084 avss.n2672 avss.t9 121.956
R16085 avss.n3490 avss.n3489 117.719
R16086 avss.n3302 avss.n3300 117.719
R16087 avss.n3490 avss.n3185 117.719
R16088 avss.n3322 avss.n3302 117.719
R16089 avss.n3320 avss.n3319 117.719
R16090 avss.n3315 avss.n3305 117.719
R16091 avss.n3313 avss.n3312 117.719
R16092 avss.n3308 avss.n3307 117.719
R16093 avss.n3483 avss.n3184 117.719
R16094 avss.n3183 avss.n3181 117.719
R16095 avss.n3502 avss.n3166 117.719
R16096 avss.n3498 avss.n3165 117.719
R16097 avss.n3501 avss.n3165 117.719
R16098 avss.n3504 avss.n3166 117.719
R16099 avss.n3485 avss.n3184 117.719
R16100 avss.n3482 avss.n3183 117.719
R16101 avss.n3321 avss.n3320 117.719
R16102 avss.n3305 avss.n3303 117.719
R16103 avss.n3314 avss.n3313 117.719
R16104 avss.n3307 avss.n3306 117.719
R16105 avss.n4695 avss.t230 116.115
R16106 avss.n4691 avss.t73 116.115
R16107 avss.n4703 avss.t398 116.115
R16108 avss.n4687 avss.t284 116.115
R16109 avss.n4711 avss.t176 116.115
R16110 avss.n4683 avss.t376 116.115
R16111 avss.n4719 avss.t338 116.115
R16112 avss.n4679 avss.t164 116.115
R16113 avss.n4727 avss.t24 116.115
R16114 avss.n3540 avss.t63 116.115
R16115 avss.n3593 avss.t170 116.115
R16116 avss.n3544 avss.t118 116.115
R16117 avss.n3585 avss.t227 116.115
R16118 avss.n3548 avss.t340 116.115
R16119 avss.n3577 avss.t213 116.115
R16120 avss.n3552 avss.t71 116.115
R16121 avss.n3569 avss.t186 116.115
R16122 avss.n3556 avss.t244 116.115
R16123 avss.n3645 avss.n2602 114.713
R16124 avss.n3638 avss.n2605 114.713
R16125 avss.n3086 avss.n3085 114.713
R16126 avss.n3082 avss.n3081 114.713
R16127 avss.n3053 avss.n2936 114.713
R16128 avss.n3046 avss.n2939 114.713
R16129 avss.n2996 avss.n2952 114.713
R16130 avss.n2989 avss.n2955 114.713
R16131 avss.n2701 avss.n2668 114.713
R16132 avss.n2708 avss.n2665 114.713
R16133 avss.n2746 avss.n2641 114.713
R16134 avss.n2753 avss.n2638 114.713
R16135 avss.n2780 avss.n2779 114.713
R16136 avss.n2784 avss.n2783 114.713
R16137 avss.n2816 avss.n2815 114.713
R16138 avss.n2820 avss.n2819 114.713
R16139 avss.n3660 avss.n3659 114.398
R16140 avss.n3094 avss.n3092 114.398
R16141 avss.n3068 avss.n3067 114.398
R16142 avss.n3011 avss.n3010 114.398
R16143 avss.n2828 avss.n2826 114.398
R16144 avss.n2792 avss.n2790 114.398
R16145 avss.n2768 avss.n2767 114.398
R16146 avss.n2723 avss.n2722 114.398
R16147 avss.n4692 avss.t112 113.677
R16148 avss.n4702 avss.t296 113.677
R16149 avss.n4688 avss.t246 113.677
R16150 avss.n4710 avss.t238 113.677
R16151 avss.n4684 avss.t264 113.677
R16152 avss.n4718 avss.t168 113.677
R16153 avss.n4680 avss.t378 113.677
R16154 avss.n4726 avss.t5 113.677
R16155 avss.n3594 avss.t310 113.677
R16156 avss.n3543 avss.t172 113.677
R16157 avss.n3586 avss.t61 113.677
R16158 avss.n3547 avss.t199 113.677
R16159 avss.n3578 avss.t7 113.677
R16160 avss.n3551 avss.t178 113.677
R16161 avss.n3570 avss.t294 113.677
R16162 avss.n3555 avss.t166 113.677
R16163 avss.n3562 avss.t241 113.677
R16164 avss.n4676 avss.t44 113.677
R16165 avss.n3621 avss.n3620 108.785
R16166 avss.n2972 avss.n2971 108.785
R16167 avss.n3029 avss.n3028 108.785
R16168 avss.n2925 avss.n2920 108.785
R16169 avss.n3608 avss.n3144 106.424
R16170 avss.n2804 avss.n2795 104.882
R16171 avss.n2915 avss.n2914 104.882
R16172 avss.n2652 avss.n2647 104.882
R16173 avss.n2676 avss.n2674 104.882
R16174 avss.t86 avss.n3249 98.1277
R16175 avss avss.t48 93.2374
R16176 avss avss.t28 93.2374
R16177 avss avss.t25 93.2374
R16178 avss.t379 avss.n3234 92.7112
R16179 avss.t34 avss 91.0199
R16180 avss.t20 avss 91.0199
R16181 avss.t45 avss 91.0199
R16182 avss.n3333 avss.n3332 90.6382
R16183 avss.n3492 avss.n3491 87.8793
R16184 avss.n3491 avss.n3490 87.3927
R16185 avss.n3302 avss.n3182 87.3927
R16186 avss.n3521 avss.n3165 87.3925
R16187 avss.n3521 avss.n3166 87.3925
R16188 avss.n3491 avss.n3184 87.3925
R16189 avss.n3491 avss.n3183 87.3925
R16190 avss.n3320 avss.n3182 87.3925
R16191 avss.n3305 avss.n3182 87.3925
R16192 avss.n3313 avss.n3182 87.3925
R16193 avss.n3307 avss.n3182 87.3925
R16194 avss.n3499 avss.n3177 87.3417
R16195 avss.n3328 avss.n3182 87.1366
R16196 avss.n3415 avss.n3230 86.9123
R16197 avss.n3450 avss.n3203 86.9123
R16198 avss.n3215 avss.n3210 86.9123
R16199 avss.n3522 avss.n3521 84.4702
R16200 avss.n3275 avss.n3268 83.7564
R16201 avss.n3012 avss.n2947 76.0005
R16202 avss.n3069 avss.n2931 76.0005
R16203 avss.n3102 avss.n3101 76.0005
R16204 avss.n3661 avss.n2597 76.0005
R16205 avss.n2724 avss.n2660 76.0005
R16206 avss.n2769 avss.n2633 76.0005
R16207 avss.n2876 avss.n2875 76.0005
R16208 avss.n2836 avss.n2835 76.0005
R16209 avss.n3521 avss.n3164 75.7581
R16210 avss.n3398 avss.n3244 75.324
R16211 avss.n3432 avss.n3228 75.324
R16212 avss.n3472 avss.n3169 75.324
R16213 avss.n3522 avss.n3163 75.1713
R16214 avss.n3330 avss.n3275 75.1179
R16215 avss.n3170 avss.n3168 74.6377
R16216 avss avss.t131 74.255
R16217 avss avss.t224 74.255
R16218 avss avss.t99 74.255
R16219 avss avss.t383 74.255
R16220 avss.n3525 avss.t257 73.8641
R16221 avss.n3526 avss.t173 73.8641
R16222 avss.n3252 avss.n3151 73.4481
R16223 avss.n3536 avss.n3535 73.4481
R16224 avss.t159 avss.n3267 73.2399
R16225 avss.t395 avss.n3266 73.2399
R16226 avss.t107 avss 72.489
R16227 avss.t275 avss 72.489
R16228 avss.t315 avss 72.489
R16229 avss.t343 avss 72.489
R16230 avss.n3146 avss.n3145 70.8187
R16231 avss.n3260 avss.n3259 70.7972
R16232 avss.n3528 avss.n3527 70.7972
R16233 avss avss.t401 70.3469
R16234 avss avss.t161 70.3469
R16235 avss avss.t115 70.3469
R16236 avss avss.t333 70.3469
R16237 avss.n3534 avss.n3158 69.3723
R16238 avss.n3160 avss.n3159 69.3467
R16239 avss.n3530 avss.n3161 69.3126
R16240 avss.n3254 avss.n3253 69.2957
R16241 avss.n3257 avss.n3256 69.2702
R16242 avss.n3264 avss.n3258 69.2363
R16243 avss.n3612 avss.n3611 69.1715
R16244 avss.t127 avss.t91 68.7958
R16245 avss.t234 avss.t363 68.7958
R16246 avss.t232 avss.t365 68.7958
R16247 avss.t367 avss.t183 68.7958
R16248 avss.t361 avss.t285 68.7958
R16249 avss.t359 avss.t181 68.7958
R16250 avss.t216 avss 68.6739
R16251 avss.t196 avss 68.6739
R16252 avss.t335 avss 68.6739
R16253 avss.t68 avss 68.6739
R16254 avss.n3399 avss.n3268 67.6543
R16255 avss.n3605 avss.n3604 67.4138
R16256 avss.n3539 avss.n3538 67.4138
R16257 avss avss.n2617 65.7939
R16258 avss.n3262 avss.n3261 64.3972
R16259 avss.n3524 avss.n3523 64.3972
R16260 avss.n3613 avss 64.2662
R16261 avss.n3374 avss.n3373 63.7358
R16262 avss.n3421 avss.n3236 63.7358
R16263 avss.n3268 avss.t159 63.4747
R16264 avss.n3245 avss.t67 63.4022
R16265 avss.n3524 avss.n3162 62.5269
R16266 avss.t305 avss.t66 61.5542
R16267 avss.n3263 avss.n3260 61.3652
R16268 avss.n3529 avss.n3528 61.3652
R16269 avss.n11630 avss.n11629 61.346
R16270 avss.t8 avss 60.8557
R16271 avss.t48 avss 60.8557
R16272 avss.t28 avss 60.8557
R16273 avss.t25 avss 60.8557
R16274 avss.n3536 avss.n3156 60.4824
R16275 avss.n3151 avss.n3150 60.4093
R16276 avss.n3539 avss.n3154 60.3406
R16277 avss.n3604 avss.n3153 60.2615
R16278 avss.n3535 avss.n3157 60.0765
R16279 avss.n3252 avss.n3251 60.0059
R16280 avss.n3538 avss.n3155 59.8927
R16281 avss.n3605 avss.n3152 59.8165
R16282 avss avss.t57 59.4084
R16283 avss avss.t34 59.4084
R16284 avss avss.t20 59.4084
R16285 avss avss.t45 59.4084
R16286 avss.n3496 avss.n3177 56.8476
R16287 avss.t257 avss.n3522 55.3035
R16288 avss.n3344 avss.n3289 52.1476
R16289 avss.n3384 avss.n3383 52.1476
R16290 avss.n3246 avss 50.9028
R16291 avss.n3247 avss.n3246 50.6052
R16292 avss.t131 avss.t133 46.8981
R16293 avss.t133 avss.t137 46.8981
R16294 avss.t137 avss.t135 46.8981
R16295 avss.t401 avss.t389 46.8981
R16296 avss.t389 avss.t403 46.8981
R16297 avss.t403 avss.t123 46.8981
R16298 avss.t224 avss.t218 46.8981
R16299 avss.t218 avss.t222 46.8981
R16300 avss.t222 avss.t220 46.8981
R16301 avss.t161 avss.t393 46.8981
R16302 avss.t393 avss.t190 46.8981
R16303 avss.t190 avss.t289 46.8981
R16304 avss.t99 avss.t95 46.8981
R16305 avss.t95 avss.t97 46.8981
R16306 avss.t97 avss.t101 46.8981
R16307 avss.t115 avss.t2 46.8981
R16308 avss.t2 avss.t391 46.8981
R16309 avss.t391 avss.t405 46.8981
R16310 avss.t383 avss.t387 46.8981
R16311 avss.t387 avss.t381 46.8981
R16312 avss.t381 avss.t385 46.8981
R16313 avss.t333 avss.t301 46.8981
R16314 avss.t301 avss.t399 46.8981
R16315 avss.t399 avss.t194 46.8981
R16316 avss.n3356 avss.n3289 46.3534
R16317 avss.t103 avss.t107 45.7827
R16318 avss.t109 avss.t103 45.7827
R16319 avss.t105 avss.t109 45.7827
R16320 avss.t0 avss.t216 45.7827
R16321 avss.t291 avss.t0 45.7827
R16322 avss.t113 avss.t291 45.7827
R16323 avss.t281 avss.t275 45.7827
R16324 avss.t279 avss.t281 45.7827
R16325 avss.t277 avss.t279 45.7827
R16326 avss.t303 avss.t196 45.7827
R16327 avss.t192 avss.t303 45.7827
R16328 avss.t214 avss.t192 45.7827
R16329 avss.t313 avss.t315 45.7827
R16330 avss.t317 avss.t313 45.7827
R16331 avss.t311 avss.t317 45.7827
R16332 avss.t319 avss.t335 45.7827
R16333 avss.t121 avss.t319 45.7827
R16334 avss.t125 avss.t121 45.7827
R16335 avss.t341 avss.t343 45.7827
R16336 avss.t347 avss.t341 45.7827
R16337 avss.t345 avss.t347 45.7827
R16338 avss.t261 avss.t68 45.7827
R16339 avss.t321 avss.t261 45.7827
R16340 avss.t407 avss.t321 45.7827
R16341 avss.t87 avss.t188 44.6975
R16342 avss.t129 avss.t299 44.3197
R16343 avss.t135 avss 41.8734
R16344 avss.t123 avss 41.8734
R16345 avss.t220 avss 41.8734
R16346 avss.t289 avss 41.8734
R16347 avss.t101 avss 41.8734
R16348 avss.t405 avss 41.8734
R16349 avss.t385 avss 41.8734
R16350 avss.t194 avss 41.8734
R16351 avss.t297 avss.t86 41.2777
R16352 avss.t229 avss.n3609 40.9322
R16353 avss.n3148 avss.t62 40.919
R16354 avss avss.t105 40.8775
R16355 avss avss.t113 40.8775
R16356 avss avss.t277 40.8775
R16357 avss avss.t214 40.8775
R16358 avss avss.t311 40.8775
R16359 avss avss.t125 40.8775
R16360 avss avss.t345 40.8775
R16361 avss avss.t407 40.8775
R16362 avss.n3360 avss.n3359 40.5593
R16363 avss.n3401 avss.t379 40.0916
R16364 avss.n4733 avss.n4732 39.2858
R16365 avss.n3561 avss.n3558 39.2858
R16366 avss.n11632 avss.n11630 38.5418
R16367 avss.n3255 avss.n3254 38.024
R16368 avss.n3534 avss.n3533 38.024
R16369 avss.n3257 avss.n3255 37.6476
R16370 avss.n3533 avss.n3160 37.6476
R16371 avss.n3428 avss.n3229 37.5859
R16372 avss.n3449 avss.n3448 37.5859
R16373 avss.n3216 avss.n3208 37.5859
R16374 avss.n3522 avss.t84 37.5859
R16375 avss.t375 avss 35.4412
R16376 avss.n3606 avss.n3151 35.3529
R16377 avss.n3537 avss.n3536 35.3529
R16378 avss.n3606 avss.n3605 35.3122
R16379 avss.n3538 avss.n3537 35.3122
R16380 avss.t23 avss 35.2183
R16381 avss.t337 avss 35.2183
R16382 avss.t175 avss 35.2183
R16383 avss.t283 avss 35.2183
R16384 avss.t72 avss 35.2183
R16385 avss.t179 avss.n3205 35.0802
R16386 avss.t163 avss 34.9954
R16387 avss.t397 avss 34.9954
R16388 avss.n3375 avss.n3374 34.7652
R16389 avss.n3421 avss.n3237 34.7652
R16390 avss.n2989 avss.n2956 34.6358
R16391 avss.n2990 avss.n2989 34.6358
R16392 avss.n2996 avss.n2995 34.6358
R16393 avss.n2997 avss.n2996 34.6358
R16394 avss.n3046 avss.n2940 34.6358
R16395 avss.n3047 avss.n3046 34.6358
R16396 avss.n3053 avss.n3052 34.6358
R16397 avss.n3054 avss.n3053 34.6358
R16398 avss.n3125 avss.n3082 34.6358
R16399 avss.n3121 avss.n3082 34.6358
R16400 avss.n3118 avss.n3086 34.6358
R16401 avss.n3114 avss.n3086 34.6358
R16402 avss.n3638 avss.n2606 34.6358
R16403 avss.n3639 avss.n3638 34.6358
R16404 avss.n3645 avss.n3644 34.6358
R16405 avss.n3646 avss.n3645 34.6358
R16406 avss.n2701 avss.n2669 34.6358
R16407 avss.n2702 avss.n2701 34.6358
R16408 avss.n2708 avss.n2707 34.6358
R16409 avss.n2709 avss.n2708 34.6358
R16410 avss.n2746 avss.n2642 34.6358
R16411 avss.n2747 avss.n2746 34.6358
R16412 avss.n2753 avss.n2752 34.6358
R16413 avss.n2754 avss.n2753 34.6358
R16414 avss.n2899 avss.n2780 34.6358
R16415 avss.n2895 avss.n2780 34.6358
R16416 avss.n2892 avss.n2784 34.6358
R16417 avss.n2888 avss.n2784 34.6358
R16418 avss.n2859 avss.n2816 34.6358
R16419 avss.n2855 avss.n2816 34.6358
R16420 avss.n2852 avss.n2820 34.6358
R16421 avss.n2848 avss.n2820 34.6358
R16422 avss.n3660 avss.t414 34.2973
R16423 avss.n3094 avss.t422 34.2973
R16424 avss.n3068 avss.t410 34.2973
R16425 avss.n3011 avss.t409 34.2973
R16426 avss.n2828 avss.t421 34.2973
R16427 avss.n2792 avss.t426 34.2973
R16428 avss.n2768 avss.t416 34.2973
R16429 avss.n2723 avss.t415 34.2973
R16430 avss.n3610 avss 33.6175
R16431 avss.n2973 avss.n2964 33.1064
R16432 avss.n3030 avss.n3021 33.1064
R16433 avss.n3138 avss.n3137 33.1064
R16434 avss.n3622 avss.n2612 33.1064
R16435 avss.n2808 avss.n2807 33.1064
R16436 avss.n2913 avss.n2628 33.1064
R16437 avss.n2656 avss.n2655 33.1064
R16438 avss.n2683 avss.n2682 33.1064
R16439 avss.n3400 avss.n3399 32.5745
R16440 avss.n3431 avss.n3430 32.5745
R16441 avss.n3471 avss.n3163 32.5745
R16442 avss.n4695 avss.n4694 31.2534
R16443 avss.n2685 avss 29.9309
R16444 avss.n2961 avss 29.9299
R16445 avss.n3667 avss.n3666 29.1367
R16446 avss.n2832 avss.n2829 29.1367
R16447 avss avss.t212 27.8627
R16448 avss.n3600 avss.n3599 27.8593
R16449 avss avss.t169 27.6398
R16450 avss avss.t226 27.6398
R16451 avss avss.t339 27.6398
R16452 avss avss.t70 27.6398
R16453 avss avss.t243 27.6398
R16454 avss.n3358 avss.n3281 27.6046
R16455 avss.n3359 avss.n3358 27.6046
R16456 avss.n3422 avss.n3234 27.5631
R16457 avss avss.t117 27.4169
R16458 avss avss.t185 27.4169
R16459 avss.n3599 avss.n3540 27.1064
R16460 avss.n3246 avss.n3245 27.0889
R16461 avss.n3250 avss.t89 26.0703
R16462 avss.t287 avss.n3149 26.0703
R16463 avss.t373 avss.n3607 26.0703
R16464 avss avss.n3147 26.0522
R16465 avss.n3178 avss.n3164 25.7581
R16466 avss.n4732 avss.n4676 25.6005
R16467 avss.n3326 avss.n3325 25.6005
R16468 avss.n3325 avss.n3299 25.6005
R16469 avss.n3324 avss.n3323 25.6005
R16470 avss.n3323 avss.n3301 25.6005
R16471 avss.n3318 avss.n3301 25.6005
R16472 avss.n3318 avss.n3317 25.6005
R16473 avss.n3317 avss.n3316 25.6005
R16474 avss.n3316 avss.n3304 25.6005
R16475 avss.n3311 avss.n3304 25.6005
R16476 avss.n3311 avss.n3310 25.6005
R16477 avss.n3310 avss.n3309 25.6005
R16478 avss.n3309 avss.n3232 25.6005
R16479 avss.n3424 avss.n3232 25.6005
R16480 avss.n3425 avss.n3424 25.6005
R16481 avss.n3426 avss.n3425 25.6005
R16482 avss.n3426 avss.n3218 25.6005
R16483 avss.n3443 avss.n3218 25.6005
R16484 avss.n3444 avss.n3443 25.6005
R16485 avss.n3446 avss.n3444 25.6005
R16486 avss.n3446 avss.n3445 25.6005
R16487 avss.n3445 avss.n3187 25.6005
R16488 avss.n3479 avss.n3187 25.6005
R16489 avss.n3480 avss.n3479 25.6005
R16490 avss.n3488 avss.n3480 25.6005
R16491 avss.n3488 avss.n3487 25.6005
R16492 avss.n3487 avss.n3486 25.6005
R16493 avss.n3486 avss.n3484 25.6005
R16494 avss.n3484 avss.n3481 25.6005
R16495 avss.n3481 avss.n3180 25.6005
R16496 avss.n3495 avss.n3494 25.6005
R16497 avss.n3496 avss.n3495 25.6005
R16498 avss.n3335 avss.n3297 25.6005
R16499 avss.n3341 avss.n3335 25.6005
R16500 avss.n3506 avss.n3505 25.6005
R16501 avss.n3505 avss.n3503 25.6005
R16502 avss.n3503 avss.n3500 25.6005
R16503 avss.n3500 avss.n3499 25.6005
R16504 avss.n3562 avss.n3561 25.6005
R16505 avss.n3330 avss.n3329 25.5404
R16506 avss.n4696 avss.n4692 25.224
R16507 avss.n4696 avss.n4695 25.224
R16508 avss.n4702 avss.n4690 25.224
R16509 avss.n4691 avss.n4690 25.224
R16510 avss.n4704 avss.n4688 25.224
R16511 avss.n4704 avss.n4703 25.224
R16512 avss.n4710 avss.n4686 25.224
R16513 avss.n4687 avss.n4686 25.224
R16514 avss.n4712 avss.n4684 25.224
R16515 avss.n4712 avss.n4711 25.224
R16516 avss.n4718 avss.n4682 25.224
R16517 avss.n4683 avss.n4682 25.224
R16518 avss.n4720 avss.n4680 25.224
R16519 avss.n4720 avss.n4719 25.224
R16520 avss.n4726 avss.n4678 25.224
R16521 avss.n4679 avss.n4678 25.224
R16522 avss.n4728 avss.n4676 25.224
R16523 avss.n4728 avss.n4727 25.224
R16524 avss.n3595 avss.n3540 25.224
R16525 avss.n3595 avss.n3594 25.224
R16526 avss.n3593 avss.n3592 25.224
R16527 avss.n3592 avss.n3543 25.224
R16528 avss.n3587 avss.n3544 25.224
R16529 avss.n3587 avss.n3586 25.224
R16530 avss.n3585 avss.n3584 25.224
R16531 avss.n3584 avss.n3547 25.224
R16532 avss.n3579 avss.n3548 25.224
R16533 avss.n3579 avss.n3578 25.224
R16534 avss.n3577 avss.n3576 25.224
R16535 avss.n3576 avss.n3551 25.224
R16536 avss.n3571 avss.n3552 25.224
R16537 avss.n3571 avss.n3570 25.224
R16538 avss.n3569 avss.n3568 25.224
R16539 avss.n3568 avss.n3555 25.224
R16540 avss.n3563 avss.n3556 25.224
R16541 avss.n3563 avss.n3562 25.224
R16542 avss.n2602 avss.t262 24.9236
R16543 avss.n2602 avss.t322 24.9236
R16544 avss.n2605 avss.t342 24.9236
R16545 avss.n2605 avss.t348 24.9236
R16546 avss.n3085 avss.t320 24.9236
R16547 avss.n3085 avss.t122 24.9236
R16548 avss.n3081 avss.t314 24.9236
R16549 avss.n3081 avss.t318 24.9236
R16550 avss.n2936 avss.t304 24.9236
R16551 avss.n2936 avss.t193 24.9236
R16552 avss.n2939 avss.t282 24.9236
R16553 avss.n2939 avss.t280 24.9236
R16554 avss.n2952 avss.t1 24.9236
R16555 avss.n2952 avss.t292 24.9236
R16556 avss.n2955 avss.t104 24.9236
R16557 avss.n2955 avss.t110 24.9236
R16558 avss.n2668 avss.t134 24.9236
R16559 avss.n2668 avss.t138 24.9236
R16560 avss.n2665 avss.t390 24.9236
R16561 avss.n2665 avss.t404 24.9236
R16562 avss.n2641 avss.t219 24.9236
R16563 avss.n2641 avss.t223 24.9236
R16564 avss.n2638 avss.t394 24.9236
R16565 avss.n2638 avss.t191 24.9236
R16566 avss.n2779 avss.t96 24.9236
R16567 avss.n2779 avss.t98 24.9236
R16568 avss.n2783 avss.t3 24.9236
R16569 avss.n2783 avss.t392 24.9236
R16570 avss.n2815 avss.t388 24.9236
R16571 avss.n2815 avss.t382 24.9236
R16572 avss.n2819 avss.t302 24.9236
R16573 avss.n2819 avss.t400 24.9236
R16574 avss.n3176 avss.t85 24.7704
R16575 avss.n3273 avss.t380 24.5445
R16576 avss.n3455 avss.t180 24.5445
R16577 avss.n3509 avss.t236 24.5445
R16578 avss.n3286 avss.t231 24.5442
R16579 avss.n3336 avss.t94 24.5442
R16580 avss.n3439 avss.n3222 24.0946
R16581 avss.n3213 avss.n3212 24.0946
R16582 avss.n3475 avss.n3474 24.0946
R16583 avss.n3419 avss.n3418 23.3417
R16584 avss.n3402 avss.n3244 23.177
R16585 avss.n3228 avss.n3221 23.177
R16586 avss.n3472 avss.n3192 23.177
R16587 avss.n3388 avss.n3387 22.5887
R16588 avss.n3531 avss.t64 22.349
R16589 avss.t259 avss.n3531 22.349
R16590 avss.n3532 avss.t87 22.349
R16591 avss.n3385 avss.n3384 22.2943
R16592 avss.n3386 avss.n3385 22.2943
R16593 avss.n2985 avss.n2956 22.2123
R16594 avss.n2991 avss.n2990 22.2123
R16595 avss.n2995 avss.n2953 22.2123
R16596 avss.n2997 avss.n2950 22.2123
R16597 avss.n3042 avss.n2940 22.2123
R16598 avss.n3048 avss.n3047 22.2123
R16599 avss.n3052 avss.n2937 22.2123
R16600 avss.n3054 avss.n2934 22.2123
R16601 avss.n3126 avss.n3125 22.2123
R16602 avss.n3121 avss.n3120 22.2123
R16603 avss.n3119 avss.n3118 22.2123
R16604 avss.n3114 avss.n3113 22.2123
R16605 avss.n3634 avss.n2606 22.2123
R16606 avss.n3640 avss.n3639 22.2123
R16607 avss.n3644 avss.n2603 22.2123
R16608 avss.n3646 avss.n2600 22.2123
R16609 avss.n2697 avss.n2669 22.2123
R16610 avss.n2703 avss.n2702 22.2123
R16611 avss.n2707 avss.n2666 22.2123
R16612 avss.n2709 avss.n2663 22.2123
R16613 avss.n2742 avss.n2642 22.2123
R16614 avss.n2748 avss.n2747 22.2123
R16615 avss.n2752 avss.n2639 22.2123
R16616 avss.n2754 avss.n2636 22.2123
R16617 avss.n2900 avss.n2899 22.2123
R16618 avss.n2895 avss.n2894 22.2123
R16619 avss.n2893 avss.n2892 22.2123
R16620 avss.n2888 avss.n2887 22.2123
R16621 avss.n2860 avss.n2859 22.2123
R16622 avss.n2855 avss.n2854 22.2123
R16623 avss.n2853 avss.n2852 22.2123
R16624 avss.n2848 avss.n2847 22.2123
R16625 avss.t119 avss.n3265 22.1601
R16626 avss.n3265 avss.t200 22.1601
R16627 avss.n3370 avss.n3282 21.8358
R16628 avss.t299 avss.n2619 21.409
R16629 avss.n3262 avss 21.0506
R16630 avss avss.n3524 21.0506
R16631 avss.n4684 avss.n4683 20.3299
R16632 avss.n3578 avss.n3577 20.3299
R16633 avss.n4692 avss.n4691 19.9534
R16634 avss.n4688 avss.n4687 19.9534
R16635 avss.n4711 avss.n4710 19.9534
R16636 avss.n4719 avss.n4718 19.9534
R16637 avss.n4727 avss.n4726 19.9534
R16638 avss.n3594 avss.n3593 19.9534
R16639 avss.n3586 avss.n3585 19.9534
R16640 avss.n3548 avss.n3547 19.9534
R16641 avss.n3552 avss.n3551 19.9534
R16642 avss.n3556 avss.n3555 19.9534
R16643 avss.n4703 avss.n4702 19.577
R16644 avss.n4680 avss.n4679 19.577
R16645 avss.n3544 avss.n3543 19.577
R16646 avss.n3570 avss.n3569 19.577
R16647 avss.n2985 avss.n2984 19.3355
R16648 avss.n3042 avss.n3041 19.3355
R16649 avss.n3127 avss.n3126 19.3355
R16650 avss.n3634 avss.n3633 19.3355
R16651 avss.n2697 avss.n2696 19.3355
R16652 avss.n2742 avss.n2741 19.3355
R16653 avss.n2901 avss.n2900 19.3355
R16654 avss.n2861 avss.n2860 19.3355
R16655 avss.t43 avss.t23 18.7239
R16656 avss.t4 avss.t163 18.7239
R16657 avss.t377 avss.t337 18.7239
R16658 avss.t167 avss.t375 18.7239
R16659 avss.t263 avss.t175 18.7239
R16660 avss.t237 avss.t283 18.7239
R16661 avss.t245 avss.t397 18.7239
R16662 avss.t295 avss.t72 18.7239
R16663 avss.t111 avss.t229 18.7239
R16664 avss.t62 avss.t309 18.7239
R16665 avss.t169 avss.t171 18.7239
R16666 avss.t117 avss.t60 18.7239
R16667 avss.t226 avss.t198 18.7239
R16668 avss.t339 avss.t6 18.7239
R16669 avss.t212 avss.t177 18.7239
R16670 avss.t70 avss.t293 18.7239
R16671 avss.t185 avss.t165 18.7239
R16672 avss.t243 avss.t240 18.7239
R16673 avss.n2991 avss.n2953 18.0711
R16674 avss.n3048 avss.n2937 18.0711
R16675 avss.n3120 avss.n3119 18.0711
R16676 avss.n3640 avss.n2603 18.0711
R16677 avss.n2703 avss.n2666 18.0711
R16678 avss.n2748 avss.n2639 18.0711
R16679 avss.n2894 avss.n2893 18.0711
R16680 avss.n2854 avss.n2853 18.0711
R16681 avss.n3001 avss.n2950 17.4103
R16682 avss.n3058 avss.n2934 17.4103
R16683 avss.n3113 avss.n3112 17.4103
R16684 avss.n3650 avss.n2600 17.4103
R16685 avss.n2713 avss.n2663 17.4103
R16686 avss.n2758 avss.n2636 17.4103
R16687 avss.n2887 avss.n2886 17.4103
R16688 avss.n2847 avss.n2846 17.4103
R16689 avss.n3261 avss.t160 17.4059
R16690 avss.n3259 avss.t396 17.4059
R16691 avss.n3527 avss.t174 17.4059
R16692 avss.n3523 avss.t258 17.4059
R16693 avss.n3152 avss.t184 17.4005
R16694 avss.n3152 avss.t286 17.4005
R16695 avss.n3153 avss.t182 17.4005
R16696 avss.n3153 avss.t308 17.4005
R16697 avss.n3251 avss.t235 17.4005
R16698 avss.n3251 avss.t306 17.4005
R16699 avss.n3150 avss.t233 17.4005
R16700 avss.n3150 avss.t288 17.4005
R16701 avss.n3253 avss.t128 17.4005
R16702 avss.n3253 avss.t298 17.4005
R16703 avss.n3256 avss.t130 17.4005
R16704 avss.n3256 avss.t300 17.4005
R16705 avss.n3258 avss.t120 17.4005
R16706 avss.n3258 avss.t201 17.4005
R16707 avss.n3154 avss.t362 17.4005
R16708 avss.n3154 avss.t360 17.4005
R16709 avss.n3155 avss.t374 17.4005
R16710 avss.n3155 avss.t368 17.4005
R16711 avss.n3156 avss.t372 17.4005
R16712 avss.n3156 avss.t366 17.4005
R16713 avss.n3157 avss.t370 17.4005
R16714 avss.n3157 avss.t364 17.4005
R16715 avss.n3158 avss.t90 17.4005
R16716 avss.n3158 avss.t92 17.4005
R16717 avss.n3159 avss.t189 17.4005
R16718 avss.n3159 avss.t88 17.4005
R16719 avss.n3161 avss.t65 17.4005
R16720 avss.n3161 avss.t260 17.4005
R16721 avss.n3178 avss.t84 17.046
R16722 avss.n3329 avss.t93 16.9019
R16723 avss.t89 avss.t127 16.6562
R16724 avss.t91 avss.t297 16.6562
R16725 avss.t369 avss.t234 16.6562
R16726 avss.t363 avss.t305 16.6562
R16727 avss.t371 avss.t232 16.6562
R16728 avss.t365 avss.t287 16.6562
R16729 avss.n3607 avss.n3149 16.6562
R16730 avss.t183 avss.t373 16.6562
R16731 avss.t285 avss.t367 16.6562
R16732 avss.t181 avss.t361 16.6562
R16733 avss.t307 avss.t359 16.6562
R16734 avss.n3018 avss.n3017 16.0891
R16735 avss.n3076 avss.n2929 16.0891
R16736 avss.n3098 avss.n3095 16.0891
R16737 avss.n2730 avss.n2729 16.0891
R16738 avss.n2908 avss.n2774 16.0891
R16739 avss.n2872 avss.n2793 16.0891
R16740 avss.n3341 avss.n3340 15.8123
R16741 avss.n3260 avss 15.0593
R16742 avss.n3528 avss 15.0593
R16743 avss.n3370 avss.n3369 15.0593
R16744 avss.n3422 avss.n3235 15.0347
R16745 avss.t309 avss 14.9346
R16746 avss.t171 avss 14.9346
R16747 avss.t60 avss 14.9346
R16748 avss.t198 avss 14.9346
R16749 avss.t6 avss 14.9346
R16750 avss.t177 avss 14.9346
R16751 avss.t293 avss 14.9346
R16752 avss.t165 avss 14.9346
R16753 avss.t240 avss 14.9346
R16754 avss.n3389 avss.n3388 14.3064
R16755 avss.n3377 avss.n3376 13.5534
R16756 avss.n3404 avss.n3403 13.5534
R16757 avss.n3418 avss.n3239 13.5534
R16758 avss.n3411 avss.n3410 13.5534
R16759 avss.n3435 avss.n3223 13.5534
R16760 avss.n3519 avss.n3171 13.5534
R16761 avss.n3507 avss.n3506 13.5534
R16762 avss.n3439 avss.n3438 12.8005
R16763 avss.n3438 avss.n3223 12.8005
R16764 avss.n3459 avss.n3193 12.8005
R16765 avss.n3475 avss.n3193 12.8005
R16766 avss.n3460 avss.n3459 12.424
R16767 avss.n3230 avss.n3227 11.5887
R16768 avss.n3211 avss.n3203 11.5887
R16769 avss.n3215 avss.n3209 11.5887
R16770 avss.n3520 avss.n3170 11.5887
R16771 avss.n3355 avss.n3354 11.2946
R16772 avss.n3401 avss.n3400 10.0233
R16773 avss.n3430 avss.n3220 10.0233
R16774 avss.n3471 avss.n3190 10.0233
R16775 avss.n11632 avss.n11627 9.3147
R16776 avss.n11633 avss.n11632 9.3005
R16777 avss.n3631 avss.n3630 9.3005
R16778 avss.n2982 avss.n2981 9.3005
R16779 avss.n2979 avss.n2958 9.3005
R16780 avss.n3036 avss.n2942 9.3005
R16781 avss.n3039 avss.n3038 9.3005
R16782 avss.n3130 avss.n3129 9.3005
R16783 avss.n3131 avss.n2928 9.3005
R16784 avss.n3628 avss.n2608 9.3005
R16785 avss.n2864 avss.n2863 9.3005
R16786 avss.n2903 avss.n2775 9.3005
R16787 avss.n2739 avss.n2738 9.3005
R16788 avss.n2694 avss.n2693 9.3005
R16789 avss.n2865 avss.n2810 9.3005
R16790 avss.n2905 avss.n2904 9.3005
R16791 avss.n2736 avss.n2644 9.3005
R16792 avss.n2691 avss.n2671 9.3005
R16793 avss.n3340 avss.n3339 9.3005
R16794 avss.n3367 avss.n3283 9.3005
R16795 avss.n3379 avss.n3277 9.3005
R16796 avss.n3406 avss.n3405 9.3005
R16797 avss.n3409 avss.n3240 9.3005
R16798 avss.n3225 avss.n3224 9.3005
R16799 avss.n3200 avss.n3199 9.3005
R16800 avss.n3468 avss.n3194 9.3005
R16801 avss.n3369 avss.n3368 9.3005
R16802 avss.n3378 avss.n3377 9.3005
R16803 avss.n3390 avss.n3389 9.3005
R16804 avss.n3404 avss.n3242 9.3005
R16805 avss.n3408 avss.n3239 9.3005
R16806 avss.n3412 avss.n3411 9.3005
R16807 avss.n3436 avss.n3435 9.3005
R16808 avss.n3457 avss.n3456 9.3005
R16809 avss.n3458 avss.n3197 9.3005
R16810 avss.n3467 avss.n3171 9.3005
R16811 avss.n3508 avss.n3507 9.3005
R16812 avss.n3338 avss.n3295 9.3005
R16813 avss.n3287 avss.n3286 9.3005
R16814 avss.n3352 avss.n3291 9.3005
R16815 avss.n3434 avss.n3433 9.3005
R16816 avss.n3433 avss.n3432 9.3005
R16817 avss.n3432 avss.n3431 9.3005
R16818 avss.n3397 avss.n3396 9.3005
R16819 avss.n3398 avss.n3397 9.3005
R16820 avss.n3399 avss.n3398 9.3005
R16821 avss.n3407 avss.n3238 9.3005
R16822 avss.n3238 avss.n3236 9.3005
R16823 avss.n3236 avss.n3234 9.3005
R16824 avss.n3414 avss.n3413 9.3005
R16825 avss.n3415 avss.n3414 9.3005
R16826 avss.n3415 avss.n3229 9.3005
R16827 avss.n3452 avss.n3451 9.3005
R16828 avss.n3451 avss.n3450 9.3005
R16829 avss.n3450 avss.n3449 9.3005
R16830 avss.n3454 avss.n3198 9.3005
R16831 avss.n3210 avss.n3198 9.3005
R16832 avss.n3210 avss.n3208 9.3005
R16833 avss.n3470 avss.n3469 9.3005
R16834 avss.n3470 avss.n3169 9.3005
R16835 avss.n3169 avss.n3163 9.3005
R16836 avss.n3517 avss.n3515 9.3005
R16837 avss.n3517 avss.n3516 9.3005
R16838 avss.n3345 avss.n3294 9.3005
R16839 avss.n3345 avss.n3344 9.3005
R16840 avss.n3361 avss.n3360 9.3005
R16841 avss.n3382 avss.n3381 9.3005
R16842 avss.n3383 avss.n3382 9.3005
R16843 avss.n3280 avss.n3278 9.3005
R16844 avss.n3373 avss.n3280 9.3005
R16845 avss.n11634 avss.n11633 9.01808
R16846 avss.n2975 avss.n2960 9.0005
R16847 avss.n3032 avss.n2944 9.0005
R16848 avss.n3135 avss.n3134 9.0005
R16849 avss.n3034 avss.n3033 9.0005
R16850 avss.n3035 avss.n3034 9.0005
R16851 avss.n2977 avss.n2976 9.0005
R16852 avss.n2978 avss.n2977 9.0005
R16853 avss.n3133 avss.n2926 9.0005
R16854 avss.n3133 avss.n3132 9.0005
R16855 avss.n3624 avss.n2610 9.0005
R16856 avss.n3626 avss.n3625 9.0005
R16857 avss.n3627 avss.n3626 9.0005
R16858 avss.n2868 avss.n2867 9.0005
R16859 avss.n2867 avss.n2866 9.0005
R16860 avss.n2869 avss.n2868 9.0005
R16861 avss.n2911 avss.n2630 9.0005
R16862 avss.n2906 avss.n2630 9.0005
R16863 avss.n2911 avss.n2910 9.0005
R16864 avss.n2734 avss.n2733 9.0005
R16865 avss.n2735 avss.n2734 9.0005
R16866 avss.n2733 avss.n2732 9.0005
R16867 avss.n2689 avss.n2688 9.0005
R16868 avss.n2690 avss.n2689 9.0005
R16869 avss.n2688 avss.n2687 9.0005
R16870 avss.n3366 avss.n3365 9.0005
R16871 avss.n3395 avss.n3394 9.0005
R16872 avss.n3465 avss.n3464 9.0005
R16873 avss.n3175 avss.n3173 9.0005
R16874 avss.n3511 avss.n3510 9.0005
R16875 avss.n3514 avss.n3513 9.0005
R16876 avss.n3463 avss.n3195 9.0005
R16877 avss.n3393 avss.n3271 9.0005
R16878 avss.n3364 avss.n3284 9.0005
R16879 avss.n3349 avss.n3292 9.0005
R16880 avss.n3351 avss.n3350 9.0005
R16881 avss.n3354 avss.n3353 9.0005
R16882 avss.n3391 avss.n3270 9.0005
R16883 avss.n3461 avss.n3460 9.0005
R16884 avss.n3174 avss.n3172 9.0005
R16885 avss.n3347 avss.n3346 9.0005
R16886 avss.n3492 avss.t84 8.71262
R16887 avss.t93 avss.n3328 8.639
R16888 avss.n2807 avss.n2806 8.19978
R16889 avss.n2628 avss.n2626 8.19978
R16890 avss.n2655 avss.n2654 8.19978
R16891 avss.n2682 avss.n2681 8.19978
R16892 avss.n3521 avss.n3168 7.9875
R16893 avss.n3532 avss.n2619 7.95505
R16894 avss.n3139 avss.n3138 7.84627
R16895 avss.n2966 avss.n2964 7.84627
R16896 avss.n3026 avss.n3021 7.84627
R16897 avss.n3618 avss.n2612 7.84627
R16898 avss.n3603 avss 7.52991
R16899 avss.n11636 avss.n11635 7.40831
R16900 avss avss.t43 7.35612
R16901 avss avss.t4 7.35612
R16902 avss avss.t377 7.35612
R16903 avss avss.t167 7.35612
R16904 avss avss.t263 7.35612
R16905 avss avss.t237 7.35612
R16906 avss avss.t245 7.35612
R16907 avss avss.t295 7.35612
R16908 avss avss.t111 7.35612
R16909 avss.t66 avss.t371 7.24211
R16910 avss.n3004 avss.n3003 6.26433
R16911 avss.n3004 avss.n2948 6.26433
R16912 avss.n3061 avss.n3060 6.26433
R16913 avss.n3061 avss.n2932 6.26433
R16914 avss.n3109 avss.n3108 6.26433
R16915 avss.n3108 avss.n3107 6.26433
R16916 avss.n3653 avss.n3652 6.26433
R16917 avss.n3653 avss.n2598 6.26433
R16918 avss.n2716 avss.n2715 6.26433
R16919 avss.n2716 avss.n2661 6.26433
R16920 avss.n2761 avss.n2760 6.26433
R16921 avss.n2761 avss.n2634 6.26433
R16922 avss.n2883 avss.n2882 6.26433
R16923 avss.n2882 avss.n2881 6.26433
R16924 avss.n2843 avss.n2842 6.26433
R16925 avss.n2842 avss.n2841 6.26433
R16926 avss.n3357 avss.n3275 6.03669
R16927 avss.n3276 avss.n3275 6.03669
R16928 avss.n3361 avss.n3287 6.02403
R16929 avss.n3601 avss 5.90819
R16930 avss.n3003 avss.n3002 5.85582
R16931 avss.n3060 avss.n3059 5.85582
R16932 avss.n3109 avss.n3088 5.85582
R16933 avss.n3652 avss.n3651 5.85582
R16934 avss.n2715 avss.n2714 5.85582
R16935 avss.n2760 avss.n2759 5.85582
R16936 avss.n2883 avss.n2786 5.85582
R16937 avss.n2843 avss.n2822 5.85582
R16938 avss.n3343 avss.n3275 5.81255
R16939 avss.n3008 avss.n2948 5.65809
R16940 avss.n3065 avss.n2932 5.65809
R16941 avss.n3107 avss.n3090 5.65809
R16942 avss.n3657 avss.n2598 5.65809
R16943 avss.n2720 avss.n2661 5.65809
R16944 avss.n2765 avss.n2634 5.65809
R16945 avss.n2881 avss.n2788 5.65809
R16946 avss.n2841 avss.n2824 5.65809
R16947 avss.n3345 avss.n3295 5.64756
R16948 avss.n3414 avss.n3240 5.64756
R16949 avss.n3414 avss.n3241 5.64756
R16950 avss.n3451 avss.n3200 5.64756
R16951 avss.n3451 avss.n3201 5.64756
R16952 avss.n3214 avss.n3198 5.64756
R16953 avss.n3518 avss.n3517 5.64756
R16954 avss.n3517 avss.n3172 5.64756
R16955 avss.n4952 avss.n4734 5.28703
R16956 avss.n3458 avss.n3457 5.27109
R16957 avss.n3603 avss 5.06097
R16958 avss.n3429 avss.n3428 5.01189
R16959 avss.n3448 avss.n3205 5.01189
R16960 avss.n3216 avss.n3207 5.01189
R16961 avss.n2978 avss.n2959 5.0092
R16962 avss.n3035 avss.n2943 5.0092
R16963 avss.n3132 avss.n3077 5.0092
R16964 avss.n3627 avss.n2609 5.0092
R16965 avss.n2690 avss.n2672 5.0092
R16966 avss.n2735 avss.n2645 5.0092
R16967 avss.n2907 avss.n2906 5.0092
R16968 avss.n2866 avss.n2811 5.0092
R16969 avss.n3397 avss.n3270 4.89462
R16970 avss.n3397 avss.n3243 4.89462
R16971 avss.n3433 avss.n3225 4.89462
R16972 avss.n3433 avss.n3226 4.89462
R16973 avss.n3473 avss.n3470 4.89462
R16974 avss.n3470 avss.n3194 4.89462
R16975 avss.n3373 avss.n3372 4.86041
R16976 avss.n3661 avss.n3660 4.85762
R16977 avss.n3101 avss.n3094 4.85762
R16978 avss.n3069 avss.n3068 4.85762
R16979 avss.n3012 avss.n3011 4.85762
R16980 avss.n2835 avss.n2828 4.85762
R16981 avss.n2875 avss.n2792 4.85762
R16982 avss.n2769 avss.n2768 4.85762
R16983 avss.n2724 avss.n2723 4.85762
R16984 avss.n3600 avss 4.67784
R16985 avss.n4732 avss.n4731 4.6505
R16986 avss.n4727 avss.n4677 4.6505
R16987 avss.n4726 avss.n4725 4.6505
R16988 avss.n4723 avss.n4679 4.6505
R16989 avss.n4722 avss.n4680 4.6505
R16990 avss.n4719 avss.n4681 4.6505
R16991 avss.n4718 avss.n4717 4.6505
R16992 avss.n4715 avss.n4683 4.6505
R16993 avss.n4714 avss.n4684 4.6505
R16994 avss.n4711 avss.n4685 4.6505
R16995 avss.n4710 avss.n4709 4.6505
R16996 avss.n4707 avss.n4687 4.6505
R16997 avss.n4706 avss.n4688 4.6505
R16998 avss.n4703 avss.n4689 4.6505
R16999 avss.n4702 avss.n4701 4.6505
R17000 avss.n4699 avss.n4691 4.6505
R17001 avss.n4698 avss.n4692 4.6505
R17002 avss.n4695 avss.n4693 4.6505
R17003 avss.n4729 avss.n4728 4.6505
R17004 avss.n4724 avss.n4678 4.6505
R17005 avss.n4721 avss.n4720 4.6505
R17006 avss.n4716 avss.n4682 4.6505
R17007 avss.n4713 avss.n4712 4.6505
R17008 avss.n4708 avss.n4686 4.6505
R17009 avss.n4705 avss.n4704 4.6505
R17010 avss.n4700 avss.n4690 4.6505
R17011 avss.n4697 avss.n4696 4.6505
R17012 avss.n4730 avss.n4676 4.6505
R17013 avss.n3635 avss.n3634 4.6505
R17014 avss.n3641 avss.n3640 4.6505
R17015 avss.n3642 avss.n2603 4.6505
R17016 avss.n3648 avss.n2600 4.6505
R17017 avss.n2962 avss.n2961 4.6505
R17018 avss.n2984 avss.n2983 4.6505
R17019 avss.n2986 avss.n2985 4.6505
R17020 avss.n2987 avss.n2956 4.6505
R17021 avss.n2989 avss.n2988 4.6505
R17022 avss.n2990 avss.n2954 4.6505
R17023 avss.n2992 avss.n2991 4.6505
R17024 avss.n2993 avss.n2953 4.6505
R17025 avss.n2995 avss.n2994 4.6505
R17026 avss.n2996 avss.n2951 4.6505
R17027 avss.n2998 avss.n2997 4.6505
R17028 avss.n2999 avss.n2950 4.6505
R17029 avss.n3001 avss.n3000 4.6505
R17030 avss.n3003 avss.n2949 4.6505
R17031 avss.n3005 avss.n3004 4.6505
R17032 avss.n3006 avss.n2948 4.6505
R17033 avss.n3008 avss.n3007 4.6505
R17034 avss.n3009 avss.n2946 4.6505
R17035 avss.n3015 avss.n3014 4.6505
R17036 avss.n3017 avss.n3016 4.6505
R17037 avss.n3019 avss.n3018 4.6505
R17038 avss.n3041 avss.n3040 4.6505
R17039 avss.n3043 avss.n3042 4.6505
R17040 avss.n3044 avss.n2940 4.6505
R17041 avss.n3046 avss.n3045 4.6505
R17042 avss.n3047 avss.n2938 4.6505
R17043 avss.n3049 avss.n3048 4.6505
R17044 avss.n3050 avss.n2937 4.6505
R17045 avss.n3052 avss.n3051 4.6505
R17046 avss.n3053 avss.n2935 4.6505
R17047 avss.n3055 avss.n3054 4.6505
R17048 avss.n3056 avss.n2934 4.6505
R17049 avss.n3058 avss.n3057 4.6505
R17050 avss.n3060 avss.n2933 4.6505
R17051 avss.n3062 avss.n3061 4.6505
R17052 avss.n3063 avss.n2932 4.6505
R17053 avss.n3065 avss.n3064 4.6505
R17054 avss.n3066 avss.n2930 4.6505
R17055 avss.n3073 avss.n3072 4.6505
R17056 avss.n3074 avss.n2929 4.6505
R17057 avss.n3076 avss.n3075 4.6505
R17058 avss.n3128 avss.n3127 4.6505
R17059 avss.n3126 avss.n3080 4.6505
R17060 avss.n3125 avss.n3124 4.6505
R17061 avss.n3123 avss.n3082 4.6505
R17062 avss.n3122 avss.n3121 4.6505
R17063 avss.n3120 avss.n3083 4.6505
R17064 avss.n3119 avss.n3084 4.6505
R17065 avss.n3118 avss.n3117 4.6505
R17066 avss.n3116 avss.n3086 4.6505
R17067 avss.n3115 avss.n3114 4.6505
R17068 avss.n3113 avss.n3087 4.6505
R17069 avss.n3112 avss.n3111 4.6505
R17070 avss.n3110 avss.n3109 4.6505
R17071 avss.n3108 avss.n3089 4.6505
R17072 avss.n3107 avss.n3106 4.6505
R17073 avss.n3105 avss.n3090 4.6505
R17074 avss.n3104 avss.n3103 4.6505
R17075 avss.n3093 avss.n3091 4.6505
R17076 avss.n3098 avss.n3097 4.6505
R17077 avss.n3096 avss.n3095 4.6505
R17078 avss.n3633 avss.n3632 4.6505
R17079 avss.n3636 avss.n2606 4.6505
R17080 avss.n3638 avss.n3637 4.6505
R17081 avss.n3639 avss.n2604 4.6505
R17082 avss.n3644 avss.n3643 4.6505
R17083 avss.n3645 avss.n2601 4.6505
R17084 avss.n3647 avss.n3646 4.6505
R17085 avss.n3650 avss.n3649 4.6505
R17086 avss.n3652 avss.n2599 4.6505
R17087 avss.n3654 avss.n3653 4.6505
R17088 avss.n3655 avss.n2598 4.6505
R17089 avss.n3657 avss.n3656 4.6505
R17090 avss.n3658 avss.n2596 4.6505
R17091 avss.n3664 avss.n3663 4.6505
R17092 avss.n3666 avss.n3665 4.6505
R17093 avss.n2860 avss.n2814 4.6505
R17094 avss.n2854 avss.n2817 4.6505
R17095 avss.n2853 avss.n2818 4.6505
R17096 avss.n2847 avss.n2821 4.6505
R17097 avss.n2887 avss.n2785 4.6505
R17098 avss.n2893 avss.n2782 4.6505
R17099 avss.n2894 avss.n2781 4.6505
R17100 avss.n2900 avss.n2778 4.6505
R17101 avss.n2756 avss.n2636 4.6505
R17102 avss.n2750 avss.n2639 4.6505
R17103 avss.n2749 avss.n2748 4.6505
R17104 avss.n2743 avss.n2742 4.6505
R17105 avss.n2711 avss.n2663 4.6505
R17106 avss.n2705 avss.n2666 4.6505
R17107 avss.n2704 avss.n2703 4.6505
R17108 avss.n2698 avss.n2697 4.6505
R17109 avss.n2832 avss.n2831 4.6505
R17110 avss.n2827 avss.n2825 4.6505
R17111 avss.n2838 avss.n2837 4.6505
R17112 avss.n2839 avss.n2824 4.6505
R17113 avss.n2841 avss.n2840 4.6505
R17114 avss.n2842 avss.n2823 4.6505
R17115 avss.n2844 avss.n2843 4.6505
R17116 avss.n2846 avss.n2845 4.6505
R17117 avss.n2849 avss.n2848 4.6505
R17118 avss.n2850 avss.n2820 4.6505
R17119 avss.n2852 avss.n2851 4.6505
R17120 avss.n2856 avss.n2855 4.6505
R17121 avss.n2857 avss.n2816 4.6505
R17122 avss.n2859 avss.n2858 4.6505
R17123 avss.n2862 avss.n2861 4.6505
R17124 avss.n2870 avss.n2793 4.6505
R17125 avss.n2872 avss.n2871 4.6505
R17126 avss.n2791 avss.n2789 4.6505
R17127 avss.n2878 avss.n2877 4.6505
R17128 avss.n2879 avss.n2788 4.6505
R17129 avss.n2881 avss.n2880 4.6505
R17130 avss.n2882 avss.n2787 4.6505
R17131 avss.n2884 avss.n2883 4.6505
R17132 avss.n2886 avss.n2885 4.6505
R17133 avss.n2889 avss.n2888 4.6505
R17134 avss.n2890 avss.n2784 4.6505
R17135 avss.n2892 avss.n2891 4.6505
R17136 avss.n2896 avss.n2895 4.6505
R17137 avss.n2897 avss.n2780 4.6505
R17138 avss.n2899 avss.n2898 4.6505
R17139 avss.n2902 avss.n2901 4.6505
R17140 avss.n2909 avss.n2908 4.6505
R17141 avss.n2774 avss.n2773 4.6505
R17142 avss.n2772 avss.n2771 4.6505
R17143 avss.n2766 avss.n2632 4.6505
R17144 avss.n2765 avss.n2764 4.6505
R17145 avss.n2763 avss.n2634 4.6505
R17146 avss.n2762 avss.n2761 4.6505
R17147 avss.n2760 avss.n2635 4.6505
R17148 avss.n2758 avss.n2757 4.6505
R17149 avss.n2755 avss.n2754 4.6505
R17150 avss.n2753 avss.n2637 4.6505
R17151 avss.n2752 avss.n2751 4.6505
R17152 avss.n2747 avss.n2640 4.6505
R17153 avss.n2746 avss.n2745 4.6505
R17154 avss.n2744 avss.n2642 4.6505
R17155 avss.n2741 avss.n2740 4.6505
R17156 avss.n2731 avss.n2730 4.6505
R17157 avss.n2729 avss.n2728 4.6505
R17158 avss.n2727 avss.n2726 4.6505
R17159 avss.n2721 avss.n2659 4.6505
R17160 avss.n2720 avss.n2719 4.6505
R17161 avss.n2718 avss.n2661 4.6505
R17162 avss.n2717 avss.n2716 4.6505
R17163 avss.n2715 avss.n2662 4.6505
R17164 avss.n2713 avss.n2712 4.6505
R17165 avss.n2710 avss.n2709 4.6505
R17166 avss.n2708 avss.n2664 4.6505
R17167 avss.n2707 avss.n2706 4.6505
R17168 avss.n2702 avss.n2667 4.6505
R17169 avss.n2701 avss.n2700 4.6505
R17170 avss.n2699 avss.n2669 4.6505
R17171 avss.n2696 avss.n2695 4.6505
R17172 avss.n2686 avss.n2685 4.6505
R17173 avss.n3466 avss.n3193 4.6505
R17174 avss.n3438 avss.n3437 4.6505
R17175 avss.n3561 avss.n3560 4.6505
R17176 avss.n3562 avss.n3557 4.6505
R17177 avss.n3565 avss.n3556 4.6505
R17178 avss.n3566 avss.n3555 4.6505
R17179 avss.n3569 avss.n3554 4.6505
R17180 avss.n3570 avss.n3553 4.6505
R17181 avss.n3573 avss.n3552 4.6505
R17182 avss.n3574 avss.n3551 4.6505
R17183 avss.n3577 avss.n3550 4.6505
R17184 avss.n3578 avss.n3549 4.6505
R17185 avss.n3581 avss.n3548 4.6505
R17186 avss.n3582 avss.n3547 4.6505
R17187 avss.n3585 avss.n3546 4.6505
R17188 avss.n3586 avss.n3545 4.6505
R17189 avss.n3589 avss.n3544 4.6505
R17190 avss.n3590 avss.n3543 4.6505
R17191 avss.n3593 avss.n3542 4.6505
R17192 avss.n3594 avss.n3541 4.6505
R17193 avss.n3597 avss.n3540 4.6505
R17194 avss.n3564 avss.n3563 4.6505
R17195 avss.n3568 avss.n3567 4.6505
R17196 avss.n3572 avss.n3571 4.6505
R17197 avss.n3576 avss.n3575 4.6505
R17198 avss.n3580 avss.n3579 4.6505
R17199 avss.n3584 avss.n3583 4.6505
R17200 avss.n3588 avss.n3587 4.6505
R17201 avss.n3592 avss.n3591 4.6505
R17202 avss.n3596 avss.n3595 4.6505
R17203 avss.n3599 avss.n3598 4.6505
R17204 avss.n2981 avss.n2980 4.5918
R17205 avss.n3038 avss.n3037 4.5918
R17206 avss.n3130 avss.n3078 4.5918
R17207 avss.n3630 avss.n3629 4.5918
R17208 avss.n2693 avss.n2692 4.5918
R17209 avss.n2738 avss.n2737 4.5918
R17210 avss.n2776 avss.n2775 4.5918
R17211 avss.n2864 avss.n2812 4.5918
R17212 avss.n3336 avss 4.5906
R17213 avss.n3362 avss.n3361 4.57427
R17214 avss.n8762 avss.n8761 4.53698
R17215 avss.n8963 avss.n8952 4.53698
R17216 avss.n8409 avss.n8408 4.53698
R17217 avss.n8610 avss.n8599 4.53698
R17218 avss.n8056 avss.n8055 4.53698
R17219 avss.n8257 avss.n8246 4.53698
R17220 avss.n7703 avss.n7702 4.53698
R17221 avss.n7904 avss.n7893 4.53698
R17222 avss.n7350 avss.n7349 4.53698
R17223 avss.n7551 avss.n7540 4.53698
R17224 avss.n6997 avss.n6996 4.53698
R17225 avss.n7198 avss.n7187 4.53698
R17226 avss.n6644 avss.n6643 4.53698
R17227 avss.n6845 avss.n6834 4.53698
R17228 avss.n6291 avss.n6290 4.53698
R17229 avss.n6492 avss.n6481 4.53698
R17230 avss.n5938 avss.n5937 4.53698
R17231 avss.n6139 avss.n6128 4.53698
R17232 avss.n5585 avss.n5584 4.53698
R17233 avss.n5786 avss.n5775 4.53698
R17234 avss.n5244 avss.n5243 4.53698
R17235 avss.n5433 avss.n5422 4.53698
R17236 avss.n4890 avss.n4889 4.53698
R17237 avss.n5079 avss.n5068 4.53698
R17238 avss.n8783 avss.n8718 4.52562
R17239 avss.n8823 avss.n8647 4.52562
R17240 avss.n8847 avss.n8846 4.52562
R17241 avss.n8931 avss.n8930 4.52562
R17242 avss.n8430 avss.n8365 4.52562
R17243 avss.n8470 avss.n8294 4.52562
R17244 avss.n8494 avss.n8493 4.52562
R17245 avss.n8578 avss.n8577 4.52562
R17246 avss.n8077 avss.n8012 4.52562
R17247 avss.n8117 avss.n7941 4.52562
R17248 avss.n8141 avss.n8140 4.52562
R17249 avss.n8225 avss.n8224 4.52562
R17250 avss.n7724 avss.n7659 4.52562
R17251 avss.n7764 avss.n7588 4.52562
R17252 avss.n7788 avss.n7787 4.52562
R17253 avss.n7872 avss.n7871 4.52562
R17254 avss.n7371 avss.n7306 4.52562
R17255 avss.n7411 avss.n7235 4.52562
R17256 avss.n7435 avss.n7434 4.52562
R17257 avss.n7519 avss.n7518 4.52562
R17258 avss.n7018 avss.n6953 4.52562
R17259 avss.n7058 avss.n6882 4.52562
R17260 avss.n7082 avss.n7081 4.52562
R17261 avss.n7166 avss.n7165 4.52562
R17262 avss.n6665 avss.n6600 4.52562
R17263 avss.n6705 avss.n6529 4.52562
R17264 avss.n6729 avss.n6728 4.52562
R17265 avss.n6813 avss.n6812 4.52562
R17266 avss.n6312 avss.n6247 4.52562
R17267 avss.n6352 avss.n6176 4.52562
R17268 avss.n6376 avss.n6375 4.52562
R17269 avss.n6460 avss.n6459 4.52562
R17270 avss.n5959 avss.n5894 4.52562
R17271 avss.n5999 avss.n5823 4.52562
R17272 avss.n6023 avss.n6022 4.52562
R17273 avss.n6107 avss.n6106 4.52562
R17274 avss.n5606 avss.n5541 4.52562
R17275 avss.n5646 avss.n5470 4.52562
R17276 avss.n5670 avss.n5669 4.52562
R17277 avss.n5754 avss.n5753 4.52562
R17278 avss.n5261 avss.n5195 4.52562
R17279 avss.n5130 avss.n5129 4.52562
R17280 avss.n5317 avss.n5316 4.52562
R17281 avss.n5401 avss.n5400 4.52562
R17282 avss.n4907 avss.n4841 4.52562
R17283 avss.n4776 avss.n4775 4.52562
R17284 avss.n4963 avss.n4962 4.52562
R17285 avss.n5047 avss.n5046 4.52562
R17286 avss.n8799 avss.n8798 4.51426
R17287 avss.n8803 avss.n8678 4.51426
R17288 avss.n8880 avss.n3705 4.51426
R17289 avss.n8901 avss.n8895 4.51426
R17290 avss.n8446 avss.n8445 4.51426
R17291 avss.n8450 avss.n8325 4.51426
R17292 avss.n8527 avss.n3789 4.51426
R17293 avss.n8548 avss.n8542 4.51426
R17294 avss.n8093 avss.n8092 4.51426
R17295 avss.n8097 avss.n7972 4.51426
R17296 avss.n8174 avss.n3873 4.51426
R17297 avss.n8195 avss.n8189 4.51426
R17298 avss.n7740 avss.n7739 4.51426
R17299 avss.n7744 avss.n7619 4.51426
R17300 avss.n7821 avss.n3957 4.51426
R17301 avss.n7842 avss.n7836 4.51426
R17302 avss.n7387 avss.n7386 4.51426
R17303 avss.n7391 avss.n7266 4.51426
R17304 avss.n7468 avss.n4041 4.51426
R17305 avss.n7489 avss.n7483 4.51426
R17306 avss.n7034 avss.n7033 4.51426
R17307 avss.n7038 avss.n6913 4.51426
R17308 avss.n7115 avss.n4125 4.51426
R17309 avss.n7136 avss.n7130 4.51426
R17310 avss.n6681 avss.n6680 4.51426
R17311 avss.n6685 avss.n6560 4.51426
R17312 avss.n6762 avss.n4209 4.51426
R17313 avss.n6783 avss.n6777 4.51426
R17314 avss.n6328 avss.n6327 4.51426
R17315 avss.n6332 avss.n6207 4.51426
R17316 avss.n6409 avss.n4293 4.51426
R17317 avss.n6430 avss.n6424 4.51426
R17318 avss.n5975 avss.n5974 4.51426
R17319 avss.n5979 avss.n5854 4.51426
R17320 avss.n6056 avss.n4377 4.51426
R17321 avss.n6077 avss.n6071 4.51426
R17322 avss.n5622 avss.n5621 4.51426
R17323 avss.n5626 avss.n5501 4.51426
R17324 avss.n5703 avss.n4461 4.51426
R17325 avss.n5724 avss.n5718 4.51426
R17326 avss.n5277 avss.n5276 4.51426
R17327 avss.n5281 avss.n5155 4.51426
R17328 avss.n5350 avss.n4545 4.51426
R17329 avss.n5371 avss.n5365 4.51426
R17330 avss.n4923 avss.n4922 4.51426
R17331 avss.n4927 avss.n4801 4.51426
R17332 avss.n4996 avss.n4629 4.51426
R17333 avss.n5017 avss.n5011 4.51426
R17334 avss.n8764 avss.n8763 4.51047
R17335 avss.n8742 avss.n8741 4.51047
R17336 avss.n8677 avss.n8676 4.51047
R17337 avss.n8815 avss.n8814 4.51047
R17338 avss.n8867 avss.n8866 4.51047
R17339 avss.n8869 avss.n3711 4.51047
R17340 avss.n8942 avss.n8941 4.51047
R17341 avss.n8951 avss.n8950 4.51047
R17342 avss.n8411 avss.n8410 4.51047
R17343 avss.n8389 avss.n8388 4.51047
R17344 avss.n8324 avss.n8323 4.51047
R17345 avss.n8462 avss.n8461 4.51047
R17346 avss.n8514 avss.n8513 4.51047
R17347 avss.n8516 avss.n3795 4.51047
R17348 avss.n8589 avss.n8588 4.51047
R17349 avss.n8598 avss.n8597 4.51047
R17350 avss.n8058 avss.n8057 4.51047
R17351 avss.n8036 avss.n8035 4.51047
R17352 avss.n7971 avss.n7970 4.51047
R17353 avss.n8109 avss.n8108 4.51047
R17354 avss.n8161 avss.n8160 4.51047
R17355 avss.n8163 avss.n3879 4.51047
R17356 avss.n8236 avss.n8235 4.51047
R17357 avss.n8245 avss.n8244 4.51047
R17358 avss.n7705 avss.n7704 4.51047
R17359 avss.n7683 avss.n7682 4.51047
R17360 avss.n7618 avss.n7617 4.51047
R17361 avss.n7756 avss.n7755 4.51047
R17362 avss.n7808 avss.n7807 4.51047
R17363 avss.n7810 avss.n3963 4.51047
R17364 avss.n7883 avss.n7882 4.51047
R17365 avss.n7892 avss.n7891 4.51047
R17366 avss.n7352 avss.n7351 4.51047
R17367 avss.n7330 avss.n7329 4.51047
R17368 avss.n7265 avss.n7264 4.51047
R17369 avss.n7403 avss.n7402 4.51047
R17370 avss.n7455 avss.n7454 4.51047
R17371 avss.n7457 avss.n4047 4.51047
R17372 avss.n7530 avss.n7529 4.51047
R17373 avss.n7539 avss.n7538 4.51047
R17374 avss.n6999 avss.n6998 4.51047
R17375 avss.n6977 avss.n6976 4.51047
R17376 avss.n6912 avss.n6911 4.51047
R17377 avss.n7050 avss.n7049 4.51047
R17378 avss.n7102 avss.n7101 4.51047
R17379 avss.n7104 avss.n4131 4.51047
R17380 avss.n7177 avss.n7176 4.51047
R17381 avss.n7186 avss.n7185 4.51047
R17382 avss.n6646 avss.n6645 4.51047
R17383 avss.n6624 avss.n6623 4.51047
R17384 avss.n6559 avss.n6558 4.51047
R17385 avss.n6697 avss.n6696 4.51047
R17386 avss.n6749 avss.n6748 4.51047
R17387 avss.n6751 avss.n4215 4.51047
R17388 avss.n6824 avss.n6823 4.51047
R17389 avss.n6833 avss.n6832 4.51047
R17390 avss.n6293 avss.n6292 4.51047
R17391 avss.n6271 avss.n6270 4.51047
R17392 avss.n6206 avss.n6205 4.51047
R17393 avss.n6344 avss.n6343 4.51047
R17394 avss.n6396 avss.n6395 4.51047
R17395 avss.n6398 avss.n4299 4.51047
R17396 avss.n6471 avss.n6470 4.51047
R17397 avss.n6480 avss.n6479 4.51047
R17398 avss.n5940 avss.n5939 4.51047
R17399 avss.n5918 avss.n5917 4.51047
R17400 avss.n5853 avss.n5852 4.51047
R17401 avss.n5991 avss.n5990 4.51047
R17402 avss.n6043 avss.n6042 4.51047
R17403 avss.n6045 avss.n4383 4.51047
R17404 avss.n6118 avss.n6117 4.51047
R17405 avss.n6127 avss.n6126 4.51047
R17406 avss.n5587 avss.n5586 4.51047
R17407 avss.n5565 avss.n5564 4.51047
R17408 avss.n5500 avss.n5499 4.51047
R17409 avss.n5638 avss.n5637 4.51047
R17410 avss.n5690 avss.n5689 4.51047
R17411 avss.n5692 avss.n4467 4.51047
R17412 avss.n5765 avss.n5764 4.51047
R17413 avss.n5774 avss.n5773 4.51047
R17414 avss.n5245 avss.n5210 4.51047
R17415 avss.n5225 avss.n5224 4.51047
R17416 avss.n5154 avss.n5153 4.51047
R17417 avss.n5292 avss.n5132 4.51047
R17418 avss.n5337 avss.n5336 4.51047
R17419 avss.n5339 avss.n4551 4.51047
R17420 avss.n5412 avss.n5411 4.51047
R17421 avss.n5421 avss.n5420 4.51047
R17422 avss.n4891 avss.n4856 4.51047
R17423 avss.n4871 avss.n4870 4.51047
R17424 avss.n4800 avss.n4799 4.51047
R17425 avss.n4938 avss.n4778 4.51047
R17426 avss.n4983 avss.n4982 4.51047
R17427 avss.n4985 avss.n4635 4.51047
R17428 avss.n5058 avss.n5057 4.51047
R17429 avss.n5067 avss.n5066 4.51047
R17430 avss.n3453 avss.n3196 4.5005
R17431 avss.n3380 avss.n3272 4.5005
R17432 avss.n3337 avss.n3293 4.5005
R17433 avss.n3372 avss.n3275 4.30475
R17434 avss.n11636 avss.n11626 4.30135
R17435 avss.n3283 avss.n3280 4.14168
R17436 avss.n3280 avss.n3279 4.14168
R17437 avss.n3405 avss.n3238 4.14168
R17438 avss.n3420 avss.n3238 4.14168
R17439 avss.n3288 avss.n3282 3.76521
R17440 avss.n2809 avss 3.61567
R17441 avss avss.n2912 3.61567
R17442 avss.n2657 avss 3.61567
R17443 avss.n2684 avss 3.61567
R17444 avss.n2975 avss.n2974 3.60668
R17445 avss.n3032 avss.n3031 3.60668
R17446 avss.n3136 avss.n3135 3.60668
R17447 avss.n3624 avss.n3623 3.60668
R17448 avss.n3010 avss.n3009 3.50735
R17449 avss.n3067 avss.n3066 3.50735
R17450 avss.n3103 avss.n3092 3.50735
R17451 avss.n3659 avss.n3658 3.50735
R17452 avss.n2722 avss.n2721 3.50735
R17453 avss.n2767 avss.n2766 3.50735
R17454 avss.n2877 avss.n2790 3.50735
R17455 avss.n2837 avss.n2826 3.50735
R17456 avss.n8639 avss.n8629 3.41965
R17457 avss.n8286 avss.n8276 3.41965
R17458 avss.n7933 avss.n7923 3.41965
R17459 avss.n7580 avss.n7570 3.41965
R17460 avss.n7227 avss.n7217 3.41965
R17461 avss.n6874 avss.n6864 3.41965
R17462 avss.n6521 avss.n6511 3.41965
R17463 avss.n6168 avss.n6158 3.41965
R17464 avss.n5815 avss.n5805 3.41965
R17465 avss.n5462 avss.n5452 3.41965
R17466 avss.n5114 avss.n5103 3.41965
R17467 avss.n4760 avss.n4749 3.41965
R17468 avss.n3739 avss.n3729 3.41965
R17469 avss.n3823 avss.n3813 3.41965
R17470 avss.n3907 avss.n3897 3.41965
R17471 avss.n3991 avss.n3981 3.41965
R17472 avss.n4075 avss.n4065 3.41965
R17473 avss.n4159 avss.n4149 3.41965
R17474 avss.n4243 avss.n4233 3.41965
R17475 avss.n4327 avss.n4317 3.41965
R17476 avss.n4411 avss.n4401 3.41965
R17477 avss.n4495 avss.n4485 3.41965
R17478 avss.n4579 avss.n4569 3.41965
R17479 avss.n4663 avss.n4653 3.41965
R17480 avss.n8753 avss.n8751 3.41468
R17481 avss.n8400 avss.n8398 3.41468
R17482 avss.n8047 avss.n8045 3.41468
R17483 avss.n7694 avss.n7692 3.41468
R17484 avss.n7341 avss.n7339 3.41468
R17485 avss.n6988 avss.n6986 3.41468
R17486 avss.n6635 avss.n6633 3.41468
R17487 avss.n6282 avss.n6280 3.41468
R17488 avss.n5929 avss.n5927 3.41468
R17489 avss.n5576 avss.n5574 3.41468
R17490 avss.n5235 avss.n5233 3.41468
R17491 avss.n4881 avss.n4879 3.41468
R17492 avss.n8728 avss.n8723 3.41335
R17493 avss.n8375 avss.n8370 3.41335
R17494 avss.n8022 avss.n8017 3.41335
R17495 avss.n7669 avss.n7664 3.41335
R17496 avss.n7316 avss.n7311 3.41335
R17497 avss.n6963 avss.n6958 3.41335
R17498 avss.n6610 avss.n6605 3.41335
R17499 avss.n6257 avss.n6252 3.41335
R17500 avss.n5904 avss.n5899 3.41335
R17501 avss.n5551 avss.n5546 3.41335
R17502 avss.n5303 avss.n5090 3.41335
R17503 avss.n4949 avss.n4736 3.41335
R17504 avss.n8960 avss.n8959 3.41317
R17505 avss.n8607 avss.n8606 3.41317
R17506 avss.n8254 avss.n8253 3.41317
R17507 avss.n7901 avss.n7900 3.41317
R17508 avss.n7548 avss.n7547 3.41317
R17509 avss.n7195 avss.n7194 3.41317
R17510 avss.n6842 avss.n6841 3.41317
R17511 avss.n6489 avss.n6488 3.41317
R17512 avss.n6136 avss.n6135 3.41317
R17513 avss.n5783 avss.n5782 3.41317
R17514 avss.n5430 avss.n5429 3.41317
R17515 avss.n5076 avss.n5075 3.41317
R17516 avss.n8755 avss.n8754 3.4105
R17517 avss.n8761 avss.n8760 3.4105
R17518 avss.n8765 avss.n8764 3.4105
R17519 avss.n8774 avss.n8727 3.4105
R17520 avss.n8769 avss.n8727 3.4105
R17521 avss.n8741 avss.n8740 3.4105
R17522 avss.n8739 avss.n8730 3.4105
R17523 avss.n8776 avss.n8775 3.4105
R17524 avss.n8774 avss.n8724 3.4105
R17525 avss.n8735 avss.n8724 3.4105
R17526 avss.n8779 avss.n8778 3.4105
R17527 avss.n8782 avss.n8781 3.4105
R17528 avss.n8783 avss.n8782 3.4105
R17529 avss.n8786 avss.n8785 3.4105
R17530 avss.n8714 avss.n8713 3.4105
R17531 avss.n8788 avss.n8716 3.4105
R17532 avss.n8711 avss.n8710 3.4105
R17533 avss.n8795 avss.n8794 3.4105
R17534 avss.n8794 avss.n8793 3.4105
R17535 avss.n8703 avss.n8702 3.4105
R17536 avss.n8697 avss.n8696 3.4105
R17537 avss.n8797 avss.n8796 3.4105
R17538 avss.n8798 avss.n8797 3.4105
R17539 avss.n8694 avss.n8693 3.4105
R17540 avss.n8690 avss.n8687 3.4105
R17541 avss.n8690 avss.n8689 3.4105
R17542 avss.n8804 avss.n8803 3.4105
R17543 avss.n8676 avss.n8670 3.4105
R17544 avss.n8668 avss.n8662 3.4105
R17545 avss.n8808 avss.n8663 3.4105
R17546 avss.n8663 avss.n8661 3.4105
R17547 avss.n8665 avss.n8664 3.4105
R17548 avss.n8817 avss.n8816 3.4105
R17549 avss.n8816 avss.n8815 3.4105
R17550 avss.n8659 avss.n8654 3.4105
R17551 avss.n8624 avss.n8623 3.4105
R17552 avss.n8819 avss.n8818 3.4105
R17553 avss.n8819 avss.n8649 3.4105
R17554 avss.n8828 avss.n8827 3.4105
R17555 avss.n8632 avss.n8625 3.4105
R17556 avss.n8640 avss.n8631 3.4105
R17557 avss.n8631 avss.n8630 3.4105
R17558 avss.n8636 avss.n8633 3.4105
R17559 avss.n8638 avss.n8637 3.4105
R17560 avss.n8644 avss.n8643 3.4105
R17561 avss.n8826 avss.n8825 3.4105
R17562 avss.n8825 avss.n8824 3.4105
R17563 avss.n8821 avss.n8820 3.4105
R17564 avss.n8658 avss.n8657 3.4105
R17565 avss.n8658 avss.n8648 3.4105
R17566 avss.n8812 avss.n8811 3.4105
R17567 avss.n8675 avss.n8674 3.4105
R17568 avss.n8675 avss.n8660 3.4105
R17569 avss.n8802 avss.n8671 3.4105
R17570 avss.n8802 avss.n8801 3.4105
R17571 avss.n8686 avss.n8680 3.4105
R17572 avss.n8684 avss.n8682 3.4105
R17573 avss.n8682 avss.n8681 3.4105
R17574 avss.n8792 avss.n8701 3.4105
R17575 avss.n8784 avss.n8717 3.4105
R17576 avss.n8784 avss.n8705 3.4105
R17577 avss.n8734 avss.n8733 3.4105
R17578 avss.n8738 avss.n8737 3.4105
R17579 avss.n8737 avss.n8729 3.4105
R17580 avss.n8771 avss.n8770 3.4105
R17581 avss.n8766 avss.n8744 3.4105
R17582 avss.n8746 avss.n8744 3.4105
R17583 avss.n8759 avss.n8748 3.4105
R17584 avss.n8748 avss.n8747 3.4105
R17585 avss.n8758 avss.n8757 3.4105
R17586 avss.n8773 avss.n8728 3.4105
R17587 avss.n8773 avss.n8772 3.4105
R17588 avss.n8834 avss.n8622 3.4105
R17589 avss.n8832 avss.n8621 3.4105
R17590 avss.n8647 avss.n8621 3.4105
R17591 avss.n8832 avss.n8831 3.4105
R17592 avss.n8627 avss.n8622 3.4105
R17593 avss.n8835 avss.n8834 3.4105
R17594 avss.n3677 avss.n3671 3.4105
R17595 avss.n8970 avss.n3671 3.4105
R17596 avss.n8964 avss.n8963 3.4105
R17597 avss.n8962 avss.n3681 3.4105
R17598 avss.n8962 avss.n8961 3.4105
R17599 avss.n8955 avss.n8953 3.4105
R17600 avss.n3738 avss.n3737 3.4105
R17601 avss.n3732 avss.n3724 3.4105
R17602 avss.n3736 avss.n3733 3.4105
R17603 avss.n3740 avss.n3731 3.4105
R17604 avss.n3731 avss.n3730 3.4105
R17605 avss.n3744 avss.n3743 3.4105
R17606 avss.n3748 avss.n3747 3.4105
R17607 avss.n3722 avss.n3721 3.4105
R17608 avss.n3721 avss.n3720 3.4105
R17609 avss.n8849 avss.n3718 3.4105
R17610 avss.n8862 avss.n8861 3.4105
R17611 avss.n8842 avss.n8841 3.4105
R17612 avss.n8855 avss.n8854 3.4105
R17613 avss.n8854 avss.n8853 3.4105
R17614 avss.n3715 avss.n3714 3.4105
R17615 avss.n8865 avss.n8864 3.4105
R17616 avss.n8866 avss.n8865 3.4105
R17617 avss.n8851 avss.n8850 3.4105
R17618 avss.n8851 avss.n3713 3.4105
R17619 avss.n8857 avss.n3710 3.4105
R17620 avss.n8859 avss.n8858 3.4105
R17621 avss.n8875 avss.n8874 3.4105
R17622 avss.n8874 avss.n8873 3.4105
R17623 avss.n3711 avss.n3706 3.4105
R17624 avss.n8871 avss.n3712 3.4105
R17625 avss.n8871 avss.n8870 3.4105
R17626 avss.n8881 avss.n3704 3.4105
R17627 avss.n8881 avss.n3699 3.4105
R17628 avss.n8891 avss.n8890 3.4105
R17629 avss.n8880 avss.n8879 3.4105
R17630 avss.n8885 avss.n8884 3.4105
R17631 avss.n8884 avss.n3700 3.4105
R17632 avss.n8893 avss.n8892 3.4105
R17633 avss.n8900 avss.n3698 3.4105
R17634 avss.n8900 avss.n3692 3.4105
R17635 avss.n8909 avss.n3695 3.4105
R17636 avss.n8888 avss.n8887 3.4105
R17637 avss.n8903 avss.n8902 3.4105
R17638 avss.n8902 avss.n8901 3.4105
R17639 avss.n8899 avss.n8898 3.4105
R17640 avss.n8904 avss.n3694 3.4105
R17641 avss.n3694 avss.n3693 3.4105
R17642 avss.n8913 avss.n8912 3.4105
R17643 avss.n8926 avss.n8925 3.4105
R17644 avss.n8906 avss.n8905 3.4105
R17645 avss.n8921 avss.n8920 3.4105
R17646 avss.n8917 avss.n8916 3.4105
R17647 avss.n8929 avss.n8928 3.4105
R17648 avss.n8930 avss.n8929 3.4105
R17649 avss.n3687 avss.n3686 3.4105
R17650 avss.n3686 avss.n3685 3.4105
R17651 avss.n8934 avss.n8933 3.4105
R17652 avss.n8923 avss.n3673 3.4105
R17653 avss.n8968 avss.n3676 3.4105
R17654 avss.n8935 avss.n3676 3.4105
R17655 avss.n8940 avss.n8939 3.4105
R17656 avss.n8968 avss.n3675 3.4105
R17657 avss.n8941 avss.n3675 3.4105
R17658 avss.n8938 avss.n3684 3.4105
R17659 avss.n3684 avss.n3683 3.4105
R17660 avss.n8944 avss.n3670 3.4105
R17661 avss.n8971 avss.n8970 3.4105
R17662 avss.n8945 avss.n3672 3.4105
R17663 avss.n8950 avss.n3680 3.4105
R17664 avss.n8949 avss.n8948 3.4105
R17665 avss.n8949 avss.n3682 3.4105
R17666 avss.n8958 avss.n8954 3.4105
R17667 avss.n8838 avss.n3726 3.4105
R17668 avss.n3726 avss.n3723 3.4105
R17669 avss.n8839 avss.n3723 3.4105
R17670 avss.n8839 avss.n8838 3.4105
R17671 avss.n8843 avss.n3751 3.4105
R17672 avss.n8846 avss.n8845 3.4105
R17673 avss.n8402 avss.n8401 3.4105
R17674 avss.n8408 avss.n8407 3.4105
R17675 avss.n8412 avss.n8411 3.4105
R17676 avss.n8421 avss.n8374 3.4105
R17677 avss.n8416 avss.n8374 3.4105
R17678 avss.n8388 avss.n8387 3.4105
R17679 avss.n8386 avss.n8377 3.4105
R17680 avss.n8423 avss.n8422 3.4105
R17681 avss.n8421 avss.n8371 3.4105
R17682 avss.n8382 avss.n8371 3.4105
R17683 avss.n8426 avss.n8425 3.4105
R17684 avss.n8429 avss.n8428 3.4105
R17685 avss.n8430 avss.n8429 3.4105
R17686 avss.n8433 avss.n8432 3.4105
R17687 avss.n8361 avss.n8360 3.4105
R17688 avss.n8435 avss.n8363 3.4105
R17689 avss.n8358 avss.n8357 3.4105
R17690 avss.n8442 avss.n8441 3.4105
R17691 avss.n8441 avss.n8440 3.4105
R17692 avss.n8350 avss.n8349 3.4105
R17693 avss.n8344 avss.n8343 3.4105
R17694 avss.n8444 avss.n8443 3.4105
R17695 avss.n8445 avss.n8444 3.4105
R17696 avss.n8341 avss.n8340 3.4105
R17697 avss.n8337 avss.n8334 3.4105
R17698 avss.n8337 avss.n8336 3.4105
R17699 avss.n8451 avss.n8450 3.4105
R17700 avss.n8323 avss.n8317 3.4105
R17701 avss.n8315 avss.n8309 3.4105
R17702 avss.n8455 avss.n8310 3.4105
R17703 avss.n8310 avss.n8308 3.4105
R17704 avss.n8312 avss.n8311 3.4105
R17705 avss.n8464 avss.n8463 3.4105
R17706 avss.n8463 avss.n8462 3.4105
R17707 avss.n8306 avss.n8301 3.4105
R17708 avss.n8271 avss.n8270 3.4105
R17709 avss.n8466 avss.n8465 3.4105
R17710 avss.n8466 avss.n8296 3.4105
R17711 avss.n8475 avss.n8474 3.4105
R17712 avss.n8279 avss.n8272 3.4105
R17713 avss.n8287 avss.n8278 3.4105
R17714 avss.n8278 avss.n8277 3.4105
R17715 avss.n8283 avss.n8280 3.4105
R17716 avss.n8285 avss.n8284 3.4105
R17717 avss.n8291 avss.n8290 3.4105
R17718 avss.n8473 avss.n8472 3.4105
R17719 avss.n8472 avss.n8471 3.4105
R17720 avss.n8468 avss.n8467 3.4105
R17721 avss.n8305 avss.n8304 3.4105
R17722 avss.n8305 avss.n8295 3.4105
R17723 avss.n8459 avss.n8458 3.4105
R17724 avss.n8322 avss.n8321 3.4105
R17725 avss.n8322 avss.n8307 3.4105
R17726 avss.n8449 avss.n8318 3.4105
R17727 avss.n8449 avss.n8448 3.4105
R17728 avss.n8333 avss.n8327 3.4105
R17729 avss.n8331 avss.n8329 3.4105
R17730 avss.n8329 avss.n8328 3.4105
R17731 avss.n8439 avss.n8348 3.4105
R17732 avss.n8431 avss.n8364 3.4105
R17733 avss.n8431 avss.n8352 3.4105
R17734 avss.n8381 avss.n8380 3.4105
R17735 avss.n8385 avss.n8384 3.4105
R17736 avss.n8384 avss.n8376 3.4105
R17737 avss.n8418 avss.n8417 3.4105
R17738 avss.n8413 avss.n8391 3.4105
R17739 avss.n8393 avss.n8391 3.4105
R17740 avss.n8406 avss.n8395 3.4105
R17741 avss.n8395 avss.n8394 3.4105
R17742 avss.n8405 avss.n8404 3.4105
R17743 avss.n8420 avss.n8375 3.4105
R17744 avss.n8420 avss.n8419 3.4105
R17745 avss.n8481 avss.n8269 3.4105
R17746 avss.n8479 avss.n8268 3.4105
R17747 avss.n8294 avss.n8268 3.4105
R17748 avss.n8479 avss.n8478 3.4105
R17749 avss.n8274 avss.n8269 3.4105
R17750 avss.n8482 avss.n8481 3.4105
R17751 avss.n3761 avss.n3755 3.4105
R17752 avss.n8617 avss.n3755 3.4105
R17753 avss.n8611 avss.n8610 3.4105
R17754 avss.n8609 avss.n3765 3.4105
R17755 avss.n8609 avss.n8608 3.4105
R17756 avss.n8602 avss.n8600 3.4105
R17757 avss.n3822 avss.n3821 3.4105
R17758 avss.n3816 avss.n3808 3.4105
R17759 avss.n3820 avss.n3817 3.4105
R17760 avss.n3824 avss.n3815 3.4105
R17761 avss.n3815 avss.n3814 3.4105
R17762 avss.n3828 avss.n3827 3.4105
R17763 avss.n3832 avss.n3831 3.4105
R17764 avss.n3806 avss.n3805 3.4105
R17765 avss.n3805 avss.n3804 3.4105
R17766 avss.n8496 avss.n3802 3.4105
R17767 avss.n8509 avss.n8508 3.4105
R17768 avss.n8489 avss.n8488 3.4105
R17769 avss.n8502 avss.n8501 3.4105
R17770 avss.n8501 avss.n8500 3.4105
R17771 avss.n3799 avss.n3798 3.4105
R17772 avss.n8512 avss.n8511 3.4105
R17773 avss.n8513 avss.n8512 3.4105
R17774 avss.n8498 avss.n8497 3.4105
R17775 avss.n8498 avss.n3797 3.4105
R17776 avss.n8504 avss.n3794 3.4105
R17777 avss.n8506 avss.n8505 3.4105
R17778 avss.n8522 avss.n8521 3.4105
R17779 avss.n8521 avss.n8520 3.4105
R17780 avss.n3795 avss.n3790 3.4105
R17781 avss.n8518 avss.n3796 3.4105
R17782 avss.n8518 avss.n8517 3.4105
R17783 avss.n8528 avss.n3788 3.4105
R17784 avss.n8528 avss.n3783 3.4105
R17785 avss.n8538 avss.n8537 3.4105
R17786 avss.n8527 avss.n8526 3.4105
R17787 avss.n8532 avss.n8531 3.4105
R17788 avss.n8531 avss.n3784 3.4105
R17789 avss.n8540 avss.n8539 3.4105
R17790 avss.n8547 avss.n3782 3.4105
R17791 avss.n8547 avss.n3776 3.4105
R17792 avss.n8556 avss.n3779 3.4105
R17793 avss.n8535 avss.n8534 3.4105
R17794 avss.n8550 avss.n8549 3.4105
R17795 avss.n8549 avss.n8548 3.4105
R17796 avss.n8546 avss.n8545 3.4105
R17797 avss.n8551 avss.n3778 3.4105
R17798 avss.n3778 avss.n3777 3.4105
R17799 avss.n8560 avss.n8559 3.4105
R17800 avss.n8573 avss.n8572 3.4105
R17801 avss.n8553 avss.n8552 3.4105
R17802 avss.n8568 avss.n8567 3.4105
R17803 avss.n8564 avss.n8563 3.4105
R17804 avss.n8576 avss.n8575 3.4105
R17805 avss.n8577 avss.n8576 3.4105
R17806 avss.n3771 avss.n3770 3.4105
R17807 avss.n3770 avss.n3769 3.4105
R17808 avss.n8581 avss.n8580 3.4105
R17809 avss.n8570 avss.n3757 3.4105
R17810 avss.n8615 avss.n3760 3.4105
R17811 avss.n8582 avss.n3760 3.4105
R17812 avss.n8587 avss.n8586 3.4105
R17813 avss.n8615 avss.n3759 3.4105
R17814 avss.n8588 avss.n3759 3.4105
R17815 avss.n8585 avss.n3768 3.4105
R17816 avss.n3768 avss.n3767 3.4105
R17817 avss.n8591 avss.n3754 3.4105
R17818 avss.n8618 avss.n8617 3.4105
R17819 avss.n8592 avss.n3756 3.4105
R17820 avss.n8597 avss.n3764 3.4105
R17821 avss.n8596 avss.n8595 3.4105
R17822 avss.n8596 avss.n3766 3.4105
R17823 avss.n8605 avss.n8601 3.4105
R17824 avss.n8485 avss.n3810 3.4105
R17825 avss.n3810 avss.n3807 3.4105
R17826 avss.n8486 avss.n3807 3.4105
R17827 avss.n8486 avss.n8485 3.4105
R17828 avss.n8490 avss.n3835 3.4105
R17829 avss.n8493 avss.n8492 3.4105
R17830 avss.n8049 avss.n8048 3.4105
R17831 avss.n8055 avss.n8054 3.4105
R17832 avss.n8059 avss.n8058 3.4105
R17833 avss.n8068 avss.n8021 3.4105
R17834 avss.n8063 avss.n8021 3.4105
R17835 avss.n8035 avss.n8034 3.4105
R17836 avss.n8033 avss.n8024 3.4105
R17837 avss.n8070 avss.n8069 3.4105
R17838 avss.n8068 avss.n8018 3.4105
R17839 avss.n8029 avss.n8018 3.4105
R17840 avss.n8073 avss.n8072 3.4105
R17841 avss.n8076 avss.n8075 3.4105
R17842 avss.n8077 avss.n8076 3.4105
R17843 avss.n8080 avss.n8079 3.4105
R17844 avss.n8008 avss.n8007 3.4105
R17845 avss.n8082 avss.n8010 3.4105
R17846 avss.n8005 avss.n8004 3.4105
R17847 avss.n8089 avss.n8088 3.4105
R17848 avss.n8088 avss.n8087 3.4105
R17849 avss.n7997 avss.n7996 3.4105
R17850 avss.n7991 avss.n7990 3.4105
R17851 avss.n8091 avss.n8090 3.4105
R17852 avss.n8092 avss.n8091 3.4105
R17853 avss.n7988 avss.n7987 3.4105
R17854 avss.n7984 avss.n7981 3.4105
R17855 avss.n7984 avss.n7983 3.4105
R17856 avss.n8098 avss.n8097 3.4105
R17857 avss.n7970 avss.n7964 3.4105
R17858 avss.n7962 avss.n7956 3.4105
R17859 avss.n8102 avss.n7957 3.4105
R17860 avss.n7957 avss.n7955 3.4105
R17861 avss.n7959 avss.n7958 3.4105
R17862 avss.n8111 avss.n8110 3.4105
R17863 avss.n8110 avss.n8109 3.4105
R17864 avss.n7953 avss.n7948 3.4105
R17865 avss.n7918 avss.n7917 3.4105
R17866 avss.n8113 avss.n8112 3.4105
R17867 avss.n8113 avss.n7943 3.4105
R17868 avss.n8122 avss.n8121 3.4105
R17869 avss.n7926 avss.n7919 3.4105
R17870 avss.n7934 avss.n7925 3.4105
R17871 avss.n7925 avss.n7924 3.4105
R17872 avss.n7930 avss.n7927 3.4105
R17873 avss.n7932 avss.n7931 3.4105
R17874 avss.n7938 avss.n7937 3.4105
R17875 avss.n8120 avss.n8119 3.4105
R17876 avss.n8119 avss.n8118 3.4105
R17877 avss.n8115 avss.n8114 3.4105
R17878 avss.n7952 avss.n7951 3.4105
R17879 avss.n7952 avss.n7942 3.4105
R17880 avss.n8106 avss.n8105 3.4105
R17881 avss.n7969 avss.n7968 3.4105
R17882 avss.n7969 avss.n7954 3.4105
R17883 avss.n8096 avss.n7965 3.4105
R17884 avss.n8096 avss.n8095 3.4105
R17885 avss.n7980 avss.n7974 3.4105
R17886 avss.n7978 avss.n7976 3.4105
R17887 avss.n7976 avss.n7975 3.4105
R17888 avss.n8086 avss.n7995 3.4105
R17889 avss.n8078 avss.n8011 3.4105
R17890 avss.n8078 avss.n7999 3.4105
R17891 avss.n8028 avss.n8027 3.4105
R17892 avss.n8032 avss.n8031 3.4105
R17893 avss.n8031 avss.n8023 3.4105
R17894 avss.n8065 avss.n8064 3.4105
R17895 avss.n8060 avss.n8038 3.4105
R17896 avss.n8040 avss.n8038 3.4105
R17897 avss.n8053 avss.n8042 3.4105
R17898 avss.n8042 avss.n8041 3.4105
R17899 avss.n8052 avss.n8051 3.4105
R17900 avss.n8067 avss.n8022 3.4105
R17901 avss.n8067 avss.n8066 3.4105
R17902 avss.n8128 avss.n7916 3.4105
R17903 avss.n8126 avss.n7915 3.4105
R17904 avss.n7941 avss.n7915 3.4105
R17905 avss.n8126 avss.n8125 3.4105
R17906 avss.n7921 avss.n7916 3.4105
R17907 avss.n8129 avss.n8128 3.4105
R17908 avss.n3845 avss.n3839 3.4105
R17909 avss.n8264 avss.n3839 3.4105
R17910 avss.n8258 avss.n8257 3.4105
R17911 avss.n8256 avss.n3849 3.4105
R17912 avss.n8256 avss.n8255 3.4105
R17913 avss.n8249 avss.n8247 3.4105
R17914 avss.n3906 avss.n3905 3.4105
R17915 avss.n3900 avss.n3892 3.4105
R17916 avss.n3904 avss.n3901 3.4105
R17917 avss.n3908 avss.n3899 3.4105
R17918 avss.n3899 avss.n3898 3.4105
R17919 avss.n3912 avss.n3911 3.4105
R17920 avss.n3916 avss.n3915 3.4105
R17921 avss.n3890 avss.n3889 3.4105
R17922 avss.n3889 avss.n3888 3.4105
R17923 avss.n8143 avss.n3886 3.4105
R17924 avss.n8156 avss.n8155 3.4105
R17925 avss.n8136 avss.n8135 3.4105
R17926 avss.n8149 avss.n8148 3.4105
R17927 avss.n8148 avss.n8147 3.4105
R17928 avss.n3883 avss.n3882 3.4105
R17929 avss.n8159 avss.n8158 3.4105
R17930 avss.n8160 avss.n8159 3.4105
R17931 avss.n8145 avss.n8144 3.4105
R17932 avss.n8145 avss.n3881 3.4105
R17933 avss.n8151 avss.n3878 3.4105
R17934 avss.n8153 avss.n8152 3.4105
R17935 avss.n8169 avss.n8168 3.4105
R17936 avss.n8168 avss.n8167 3.4105
R17937 avss.n3879 avss.n3874 3.4105
R17938 avss.n8165 avss.n3880 3.4105
R17939 avss.n8165 avss.n8164 3.4105
R17940 avss.n8175 avss.n3872 3.4105
R17941 avss.n8175 avss.n3867 3.4105
R17942 avss.n8185 avss.n8184 3.4105
R17943 avss.n8174 avss.n8173 3.4105
R17944 avss.n8179 avss.n8178 3.4105
R17945 avss.n8178 avss.n3868 3.4105
R17946 avss.n8187 avss.n8186 3.4105
R17947 avss.n8194 avss.n3866 3.4105
R17948 avss.n8194 avss.n3860 3.4105
R17949 avss.n8203 avss.n3863 3.4105
R17950 avss.n8182 avss.n8181 3.4105
R17951 avss.n8197 avss.n8196 3.4105
R17952 avss.n8196 avss.n8195 3.4105
R17953 avss.n8193 avss.n8192 3.4105
R17954 avss.n8198 avss.n3862 3.4105
R17955 avss.n3862 avss.n3861 3.4105
R17956 avss.n8207 avss.n8206 3.4105
R17957 avss.n8220 avss.n8219 3.4105
R17958 avss.n8200 avss.n8199 3.4105
R17959 avss.n8215 avss.n8214 3.4105
R17960 avss.n8211 avss.n8210 3.4105
R17961 avss.n8223 avss.n8222 3.4105
R17962 avss.n8224 avss.n8223 3.4105
R17963 avss.n3855 avss.n3854 3.4105
R17964 avss.n3854 avss.n3853 3.4105
R17965 avss.n8228 avss.n8227 3.4105
R17966 avss.n8217 avss.n3841 3.4105
R17967 avss.n8262 avss.n3844 3.4105
R17968 avss.n8229 avss.n3844 3.4105
R17969 avss.n8234 avss.n8233 3.4105
R17970 avss.n8262 avss.n3843 3.4105
R17971 avss.n8235 avss.n3843 3.4105
R17972 avss.n8232 avss.n3852 3.4105
R17973 avss.n3852 avss.n3851 3.4105
R17974 avss.n8238 avss.n3838 3.4105
R17975 avss.n8265 avss.n8264 3.4105
R17976 avss.n8239 avss.n3840 3.4105
R17977 avss.n8244 avss.n3848 3.4105
R17978 avss.n8243 avss.n8242 3.4105
R17979 avss.n8243 avss.n3850 3.4105
R17980 avss.n8252 avss.n8248 3.4105
R17981 avss.n8132 avss.n3894 3.4105
R17982 avss.n3894 avss.n3891 3.4105
R17983 avss.n8133 avss.n3891 3.4105
R17984 avss.n8133 avss.n8132 3.4105
R17985 avss.n8137 avss.n3919 3.4105
R17986 avss.n8140 avss.n8139 3.4105
R17987 avss.n7696 avss.n7695 3.4105
R17988 avss.n7702 avss.n7701 3.4105
R17989 avss.n7706 avss.n7705 3.4105
R17990 avss.n7715 avss.n7668 3.4105
R17991 avss.n7710 avss.n7668 3.4105
R17992 avss.n7682 avss.n7681 3.4105
R17993 avss.n7680 avss.n7671 3.4105
R17994 avss.n7717 avss.n7716 3.4105
R17995 avss.n7715 avss.n7665 3.4105
R17996 avss.n7676 avss.n7665 3.4105
R17997 avss.n7720 avss.n7719 3.4105
R17998 avss.n7723 avss.n7722 3.4105
R17999 avss.n7724 avss.n7723 3.4105
R18000 avss.n7727 avss.n7726 3.4105
R18001 avss.n7655 avss.n7654 3.4105
R18002 avss.n7729 avss.n7657 3.4105
R18003 avss.n7652 avss.n7651 3.4105
R18004 avss.n7736 avss.n7735 3.4105
R18005 avss.n7735 avss.n7734 3.4105
R18006 avss.n7644 avss.n7643 3.4105
R18007 avss.n7638 avss.n7637 3.4105
R18008 avss.n7738 avss.n7737 3.4105
R18009 avss.n7739 avss.n7738 3.4105
R18010 avss.n7635 avss.n7634 3.4105
R18011 avss.n7631 avss.n7628 3.4105
R18012 avss.n7631 avss.n7630 3.4105
R18013 avss.n7745 avss.n7744 3.4105
R18014 avss.n7617 avss.n7611 3.4105
R18015 avss.n7609 avss.n7603 3.4105
R18016 avss.n7749 avss.n7604 3.4105
R18017 avss.n7604 avss.n7602 3.4105
R18018 avss.n7606 avss.n7605 3.4105
R18019 avss.n7758 avss.n7757 3.4105
R18020 avss.n7757 avss.n7756 3.4105
R18021 avss.n7600 avss.n7595 3.4105
R18022 avss.n7565 avss.n7564 3.4105
R18023 avss.n7760 avss.n7759 3.4105
R18024 avss.n7760 avss.n7590 3.4105
R18025 avss.n7769 avss.n7768 3.4105
R18026 avss.n7573 avss.n7566 3.4105
R18027 avss.n7581 avss.n7572 3.4105
R18028 avss.n7572 avss.n7571 3.4105
R18029 avss.n7577 avss.n7574 3.4105
R18030 avss.n7579 avss.n7578 3.4105
R18031 avss.n7585 avss.n7584 3.4105
R18032 avss.n7767 avss.n7766 3.4105
R18033 avss.n7766 avss.n7765 3.4105
R18034 avss.n7762 avss.n7761 3.4105
R18035 avss.n7599 avss.n7598 3.4105
R18036 avss.n7599 avss.n7589 3.4105
R18037 avss.n7753 avss.n7752 3.4105
R18038 avss.n7616 avss.n7615 3.4105
R18039 avss.n7616 avss.n7601 3.4105
R18040 avss.n7743 avss.n7612 3.4105
R18041 avss.n7743 avss.n7742 3.4105
R18042 avss.n7627 avss.n7621 3.4105
R18043 avss.n7625 avss.n7623 3.4105
R18044 avss.n7623 avss.n7622 3.4105
R18045 avss.n7733 avss.n7642 3.4105
R18046 avss.n7725 avss.n7658 3.4105
R18047 avss.n7725 avss.n7646 3.4105
R18048 avss.n7675 avss.n7674 3.4105
R18049 avss.n7679 avss.n7678 3.4105
R18050 avss.n7678 avss.n7670 3.4105
R18051 avss.n7712 avss.n7711 3.4105
R18052 avss.n7707 avss.n7685 3.4105
R18053 avss.n7687 avss.n7685 3.4105
R18054 avss.n7700 avss.n7689 3.4105
R18055 avss.n7689 avss.n7688 3.4105
R18056 avss.n7699 avss.n7698 3.4105
R18057 avss.n7714 avss.n7669 3.4105
R18058 avss.n7714 avss.n7713 3.4105
R18059 avss.n7775 avss.n7563 3.4105
R18060 avss.n7773 avss.n7562 3.4105
R18061 avss.n7588 avss.n7562 3.4105
R18062 avss.n7773 avss.n7772 3.4105
R18063 avss.n7568 avss.n7563 3.4105
R18064 avss.n7776 avss.n7775 3.4105
R18065 avss.n3929 avss.n3923 3.4105
R18066 avss.n7911 avss.n3923 3.4105
R18067 avss.n7905 avss.n7904 3.4105
R18068 avss.n7903 avss.n3933 3.4105
R18069 avss.n7903 avss.n7902 3.4105
R18070 avss.n7896 avss.n7894 3.4105
R18071 avss.n3990 avss.n3989 3.4105
R18072 avss.n3984 avss.n3976 3.4105
R18073 avss.n3988 avss.n3985 3.4105
R18074 avss.n3992 avss.n3983 3.4105
R18075 avss.n3983 avss.n3982 3.4105
R18076 avss.n3996 avss.n3995 3.4105
R18077 avss.n4000 avss.n3999 3.4105
R18078 avss.n3974 avss.n3973 3.4105
R18079 avss.n3973 avss.n3972 3.4105
R18080 avss.n7790 avss.n3970 3.4105
R18081 avss.n7803 avss.n7802 3.4105
R18082 avss.n7783 avss.n7782 3.4105
R18083 avss.n7796 avss.n7795 3.4105
R18084 avss.n7795 avss.n7794 3.4105
R18085 avss.n3967 avss.n3966 3.4105
R18086 avss.n7806 avss.n7805 3.4105
R18087 avss.n7807 avss.n7806 3.4105
R18088 avss.n7792 avss.n7791 3.4105
R18089 avss.n7792 avss.n3965 3.4105
R18090 avss.n7798 avss.n3962 3.4105
R18091 avss.n7800 avss.n7799 3.4105
R18092 avss.n7816 avss.n7815 3.4105
R18093 avss.n7815 avss.n7814 3.4105
R18094 avss.n3963 avss.n3958 3.4105
R18095 avss.n7812 avss.n3964 3.4105
R18096 avss.n7812 avss.n7811 3.4105
R18097 avss.n7822 avss.n3956 3.4105
R18098 avss.n7822 avss.n3951 3.4105
R18099 avss.n7832 avss.n7831 3.4105
R18100 avss.n7821 avss.n7820 3.4105
R18101 avss.n7826 avss.n7825 3.4105
R18102 avss.n7825 avss.n3952 3.4105
R18103 avss.n7834 avss.n7833 3.4105
R18104 avss.n7841 avss.n3950 3.4105
R18105 avss.n7841 avss.n3944 3.4105
R18106 avss.n7850 avss.n3947 3.4105
R18107 avss.n7829 avss.n7828 3.4105
R18108 avss.n7844 avss.n7843 3.4105
R18109 avss.n7843 avss.n7842 3.4105
R18110 avss.n7840 avss.n7839 3.4105
R18111 avss.n7845 avss.n3946 3.4105
R18112 avss.n3946 avss.n3945 3.4105
R18113 avss.n7854 avss.n7853 3.4105
R18114 avss.n7867 avss.n7866 3.4105
R18115 avss.n7847 avss.n7846 3.4105
R18116 avss.n7862 avss.n7861 3.4105
R18117 avss.n7858 avss.n7857 3.4105
R18118 avss.n7870 avss.n7869 3.4105
R18119 avss.n7871 avss.n7870 3.4105
R18120 avss.n3939 avss.n3938 3.4105
R18121 avss.n3938 avss.n3937 3.4105
R18122 avss.n7875 avss.n7874 3.4105
R18123 avss.n7864 avss.n3925 3.4105
R18124 avss.n7909 avss.n3928 3.4105
R18125 avss.n7876 avss.n3928 3.4105
R18126 avss.n7881 avss.n7880 3.4105
R18127 avss.n7909 avss.n3927 3.4105
R18128 avss.n7882 avss.n3927 3.4105
R18129 avss.n7879 avss.n3936 3.4105
R18130 avss.n3936 avss.n3935 3.4105
R18131 avss.n7885 avss.n3922 3.4105
R18132 avss.n7912 avss.n7911 3.4105
R18133 avss.n7886 avss.n3924 3.4105
R18134 avss.n7891 avss.n3932 3.4105
R18135 avss.n7890 avss.n7889 3.4105
R18136 avss.n7890 avss.n3934 3.4105
R18137 avss.n7899 avss.n7895 3.4105
R18138 avss.n7779 avss.n3978 3.4105
R18139 avss.n3978 avss.n3975 3.4105
R18140 avss.n7780 avss.n3975 3.4105
R18141 avss.n7780 avss.n7779 3.4105
R18142 avss.n7784 avss.n4003 3.4105
R18143 avss.n7787 avss.n7786 3.4105
R18144 avss.n7343 avss.n7342 3.4105
R18145 avss.n7349 avss.n7348 3.4105
R18146 avss.n7353 avss.n7352 3.4105
R18147 avss.n7362 avss.n7315 3.4105
R18148 avss.n7357 avss.n7315 3.4105
R18149 avss.n7329 avss.n7328 3.4105
R18150 avss.n7327 avss.n7318 3.4105
R18151 avss.n7364 avss.n7363 3.4105
R18152 avss.n7362 avss.n7312 3.4105
R18153 avss.n7323 avss.n7312 3.4105
R18154 avss.n7367 avss.n7366 3.4105
R18155 avss.n7370 avss.n7369 3.4105
R18156 avss.n7371 avss.n7370 3.4105
R18157 avss.n7374 avss.n7373 3.4105
R18158 avss.n7302 avss.n7301 3.4105
R18159 avss.n7376 avss.n7304 3.4105
R18160 avss.n7299 avss.n7298 3.4105
R18161 avss.n7383 avss.n7382 3.4105
R18162 avss.n7382 avss.n7381 3.4105
R18163 avss.n7291 avss.n7290 3.4105
R18164 avss.n7285 avss.n7284 3.4105
R18165 avss.n7385 avss.n7384 3.4105
R18166 avss.n7386 avss.n7385 3.4105
R18167 avss.n7282 avss.n7281 3.4105
R18168 avss.n7278 avss.n7275 3.4105
R18169 avss.n7278 avss.n7277 3.4105
R18170 avss.n7392 avss.n7391 3.4105
R18171 avss.n7264 avss.n7258 3.4105
R18172 avss.n7256 avss.n7250 3.4105
R18173 avss.n7396 avss.n7251 3.4105
R18174 avss.n7251 avss.n7249 3.4105
R18175 avss.n7253 avss.n7252 3.4105
R18176 avss.n7405 avss.n7404 3.4105
R18177 avss.n7404 avss.n7403 3.4105
R18178 avss.n7247 avss.n7242 3.4105
R18179 avss.n7212 avss.n7211 3.4105
R18180 avss.n7407 avss.n7406 3.4105
R18181 avss.n7407 avss.n7237 3.4105
R18182 avss.n7416 avss.n7415 3.4105
R18183 avss.n7220 avss.n7213 3.4105
R18184 avss.n7228 avss.n7219 3.4105
R18185 avss.n7219 avss.n7218 3.4105
R18186 avss.n7224 avss.n7221 3.4105
R18187 avss.n7226 avss.n7225 3.4105
R18188 avss.n7232 avss.n7231 3.4105
R18189 avss.n7414 avss.n7413 3.4105
R18190 avss.n7413 avss.n7412 3.4105
R18191 avss.n7409 avss.n7408 3.4105
R18192 avss.n7246 avss.n7245 3.4105
R18193 avss.n7246 avss.n7236 3.4105
R18194 avss.n7400 avss.n7399 3.4105
R18195 avss.n7263 avss.n7262 3.4105
R18196 avss.n7263 avss.n7248 3.4105
R18197 avss.n7390 avss.n7259 3.4105
R18198 avss.n7390 avss.n7389 3.4105
R18199 avss.n7274 avss.n7268 3.4105
R18200 avss.n7272 avss.n7270 3.4105
R18201 avss.n7270 avss.n7269 3.4105
R18202 avss.n7380 avss.n7289 3.4105
R18203 avss.n7372 avss.n7305 3.4105
R18204 avss.n7372 avss.n7293 3.4105
R18205 avss.n7322 avss.n7321 3.4105
R18206 avss.n7326 avss.n7325 3.4105
R18207 avss.n7325 avss.n7317 3.4105
R18208 avss.n7359 avss.n7358 3.4105
R18209 avss.n7354 avss.n7332 3.4105
R18210 avss.n7334 avss.n7332 3.4105
R18211 avss.n7347 avss.n7336 3.4105
R18212 avss.n7336 avss.n7335 3.4105
R18213 avss.n7346 avss.n7345 3.4105
R18214 avss.n7361 avss.n7316 3.4105
R18215 avss.n7361 avss.n7360 3.4105
R18216 avss.n7422 avss.n7210 3.4105
R18217 avss.n7420 avss.n7209 3.4105
R18218 avss.n7235 avss.n7209 3.4105
R18219 avss.n7420 avss.n7419 3.4105
R18220 avss.n7215 avss.n7210 3.4105
R18221 avss.n7423 avss.n7422 3.4105
R18222 avss.n4013 avss.n4007 3.4105
R18223 avss.n7558 avss.n4007 3.4105
R18224 avss.n7552 avss.n7551 3.4105
R18225 avss.n7550 avss.n4017 3.4105
R18226 avss.n7550 avss.n7549 3.4105
R18227 avss.n7543 avss.n7541 3.4105
R18228 avss.n4074 avss.n4073 3.4105
R18229 avss.n4068 avss.n4060 3.4105
R18230 avss.n4072 avss.n4069 3.4105
R18231 avss.n4076 avss.n4067 3.4105
R18232 avss.n4067 avss.n4066 3.4105
R18233 avss.n4080 avss.n4079 3.4105
R18234 avss.n4084 avss.n4083 3.4105
R18235 avss.n4058 avss.n4057 3.4105
R18236 avss.n4057 avss.n4056 3.4105
R18237 avss.n7437 avss.n4054 3.4105
R18238 avss.n7450 avss.n7449 3.4105
R18239 avss.n7430 avss.n7429 3.4105
R18240 avss.n7443 avss.n7442 3.4105
R18241 avss.n7442 avss.n7441 3.4105
R18242 avss.n4051 avss.n4050 3.4105
R18243 avss.n7453 avss.n7452 3.4105
R18244 avss.n7454 avss.n7453 3.4105
R18245 avss.n7439 avss.n7438 3.4105
R18246 avss.n7439 avss.n4049 3.4105
R18247 avss.n7445 avss.n4046 3.4105
R18248 avss.n7447 avss.n7446 3.4105
R18249 avss.n7463 avss.n7462 3.4105
R18250 avss.n7462 avss.n7461 3.4105
R18251 avss.n4047 avss.n4042 3.4105
R18252 avss.n7459 avss.n4048 3.4105
R18253 avss.n7459 avss.n7458 3.4105
R18254 avss.n7469 avss.n4040 3.4105
R18255 avss.n7469 avss.n4035 3.4105
R18256 avss.n7479 avss.n7478 3.4105
R18257 avss.n7468 avss.n7467 3.4105
R18258 avss.n7473 avss.n7472 3.4105
R18259 avss.n7472 avss.n4036 3.4105
R18260 avss.n7481 avss.n7480 3.4105
R18261 avss.n7488 avss.n4034 3.4105
R18262 avss.n7488 avss.n4028 3.4105
R18263 avss.n7497 avss.n4031 3.4105
R18264 avss.n7476 avss.n7475 3.4105
R18265 avss.n7491 avss.n7490 3.4105
R18266 avss.n7490 avss.n7489 3.4105
R18267 avss.n7487 avss.n7486 3.4105
R18268 avss.n7492 avss.n4030 3.4105
R18269 avss.n4030 avss.n4029 3.4105
R18270 avss.n7501 avss.n7500 3.4105
R18271 avss.n7514 avss.n7513 3.4105
R18272 avss.n7494 avss.n7493 3.4105
R18273 avss.n7509 avss.n7508 3.4105
R18274 avss.n7505 avss.n7504 3.4105
R18275 avss.n7517 avss.n7516 3.4105
R18276 avss.n7518 avss.n7517 3.4105
R18277 avss.n4023 avss.n4022 3.4105
R18278 avss.n4022 avss.n4021 3.4105
R18279 avss.n7522 avss.n7521 3.4105
R18280 avss.n7511 avss.n4009 3.4105
R18281 avss.n7556 avss.n4012 3.4105
R18282 avss.n7523 avss.n4012 3.4105
R18283 avss.n7528 avss.n7527 3.4105
R18284 avss.n7556 avss.n4011 3.4105
R18285 avss.n7529 avss.n4011 3.4105
R18286 avss.n7526 avss.n4020 3.4105
R18287 avss.n4020 avss.n4019 3.4105
R18288 avss.n7532 avss.n4006 3.4105
R18289 avss.n7559 avss.n7558 3.4105
R18290 avss.n7533 avss.n4008 3.4105
R18291 avss.n7538 avss.n4016 3.4105
R18292 avss.n7537 avss.n7536 3.4105
R18293 avss.n7537 avss.n4018 3.4105
R18294 avss.n7546 avss.n7542 3.4105
R18295 avss.n7426 avss.n4062 3.4105
R18296 avss.n4062 avss.n4059 3.4105
R18297 avss.n7427 avss.n4059 3.4105
R18298 avss.n7427 avss.n7426 3.4105
R18299 avss.n7431 avss.n4087 3.4105
R18300 avss.n7434 avss.n7433 3.4105
R18301 avss.n6990 avss.n6989 3.4105
R18302 avss.n6996 avss.n6995 3.4105
R18303 avss.n7000 avss.n6999 3.4105
R18304 avss.n7009 avss.n6962 3.4105
R18305 avss.n7004 avss.n6962 3.4105
R18306 avss.n6976 avss.n6975 3.4105
R18307 avss.n6974 avss.n6965 3.4105
R18308 avss.n7011 avss.n7010 3.4105
R18309 avss.n7009 avss.n6959 3.4105
R18310 avss.n6970 avss.n6959 3.4105
R18311 avss.n7014 avss.n7013 3.4105
R18312 avss.n7017 avss.n7016 3.4105
R18313 avss.n7018 avss.n7017 3.4105
R18314 avss.n7021 avss.n7020 3.4105
R18315 avss.n6949 avss.n6948 3.4105
R18316 avss.n7023 avss.n6951 3.4105
R18317 avss.n6946 avss.n6945 3.4105
R18318 avss.n7030 avss.n7029 3.4105
R18319 avss.n7029 avss.n7028 3.4105
R18320 avss.n6938 avss.n6937 3.4105
R18321 avss.n6932 avss.n6931 3.4105
R18322 avss.n7032 avss.n7031 3.4105
R18323 avss.n7033 avss.n7032 3.4105
R18324 avss.n6929 avss.n6928 3.4105
R18325 avss.n6925 avss.n6922 3.4105
R18326 avss.n6925 avss.n6924 3.4105
R18327 avss.n7039 avss.n7038 3.4105
R18328 avss.n6911 avss.n6905 3.4105
R18329 avss.n6903 avss.n6897 3.4105
R18330 avss.n7043 avss.n6898 3.4105
R18331 avss.n6898 avss.n6896 3.4105
R18332 avss.n6900 avss.n6899 3.4105
R18333 avss.n7052 avss.n7051 3.4105
R18334 avss.n7051 avss.n7050 3.4105
R18335 avss.n6894 avss.n6889 3.4105
R18336 avss.n6859 avss.n6858 3.4105
R18337 avss.n7054 avss.n7053 3.4105
R18338 avss.n7054 avss.n6884 3.4105
R18339 avss.n7063 avss.n7062 3.4105
R18340 avss.n6867 avss.n6860 3.4105
R18341 avss.n6875 avss.n6866 3.4105
R18342 avss.n6866 avss.n6865 3.4105
R18343 avss.n6871 avss.n6868 3.4105
R18344 avss.n6873 avss.n6872 3.4105
R18345 avss.n6879 avss.n6878 3.4105
R18346 avss.n7061 avss.n7060 3.4105
R18347 avss.n7060 avss.n7059 3.4105
R18348 avss.n7056 avss.n7055 3.4105
R18349 avss.n6893 avss.n6892 3.4105
R18350 avss.n6893 avss.n6883 3.4105
R18351 avss.n7047 avss.n7046 3.4105
R18352 avss.n6910 avss.n6909 3.4105
R18353 avss.n6910 avss.n6895 3.4105
R18354 avss.n7037 avss.n6906 3.4105
R18355 avss.n7037 avss.n7036 3.4105
R18356 avss.n6921 avss.n6915 3.4105
R18357 avss.n6919 avss.n6917 3.4105
R18358 avss.n6917 avss.n6916 3.4105
R18359 avss.n7027 avss.n6936 3.4105
R18360 avss.n7019 avss.n6952 3.4105
R18361 avss.n7019 avss.n6940 3.4105
R18362 avss.n6969 avss.n6968 3.4105
R18363 avss.n6973 avss.n6972 3.4105
R18364 avss.n6972 avss.n6964 3.4105
R18365 avss.n7006 avss.n7005 3.4105
R18366 avss.n7001 avss.n6979 3.4105
R18367 avss.n6981 avss.n6979 3.4105
R18368 avss.n6994 avss.n6983 3.4105
R18369 avss.n6983 avss.n6982 3.4105
R18370 avss.n6993 avss.n6992 3.4105
R18371 avss.n7008 avss.n6963 3.4105
R18372 avss.n7008 avss.n7007 3.4105
R18373 avss.n7069 avss.n6857 3.4105
R18374 avss.n7067 avss.n6856 3.4105
R18375 avss.n6882 avss.n6856 3.4105
R18376 avss.n7067 avss.n7066 3.4105
R18377 avss.n6862 avss.n6857 3.4105
R18378 avss.n7070 avss.n7069 3.4105
R18379 avss.n4097 avss.n4091 3.4105
R18380 avss.n7205 avss.n4091 3.4105
R18381 avss.n7199 avss.n7198 3.4105
R18382 avss.n7197 avss.n4101 3.4105
R18383 avss.n7197 avss.n7196 3.4105
R18384 avss.n7190 avss.n7188 3.4105
R18385 avss.n4158 avss.n4157 3.4105
R18386 avss.n4152 avss.n4144 3.4105
R18387 avss.n4156 avss.n4153 3.4105
R18388 avss.n4160 avss.n4151 3.4105
R18389 avss.n4151 avss.n4150 3.4105
R18390 avss.n4164 avss.n4163 3.4105
R18391 avss.n4168 avss.n4167 3.4105
R18392 avss.n4142 avss.n4141 3.4105
R18393 avss.n4141 avss.n4140 3.4105
R18394 avss.n7084 avss.n4138 3.4105
R18395 avss.n7097 avss.n7096 3.4105
R18396 avss.n7077 avss.n7076 3.4105
R18397 avss.n7090 avss.n7089 3.4105
R18398 avss.n7089 avss.n7088 3.4105
R18399 avss.n4135 avss.n4134 3.4105
R18400 avss.n7100 avss.n7099 3.4105
R18401 avss.n7101 avss.n7100 3.4105
R18402 avss.n7086 avss.n7085 3.4105
R18403 avss.n7086 avss.n4133 3.4105
R18404 avss.n7092 avss.n4130 3.4105
R18405 avss.n7094 avss.n7093 3.4105
R18406 avss.n7110 avss.n7109 3.4105
R18407 avss.n7109 avss.n7108 3.4105
R18408 avss.n4131 avss.n4126 3.4105
R18409 avss.n7106 avss.n4132 3.4105
R18410 avss.n7106 avss.n7105 3.4105
R18411 avss.n7116 avss.n4124 3.4105
R18412 avss.n7116 avss.n4119 3.4105
R18413 avss.n7126 avss.n7125 3.4105
R18414 avss.n7115 avss.n7114 3.4105
R18415 avss.n7120 avss.n7119 3.4105
R18416 avss.n7119 avss.n4120 3.4105
R18417 avss.n7128 avss.n7127 3.4105
R18418 avss.n7135 avss.n4118 3.4105
R18419 avss.n7135 avss.n4112 3.4105
R18420 avss.n7144 avss.n4115 3.4105
R18421 avss.n7123 avss.n7122 3.4105
R18422 avss.n7138 avss.n7137 3.4105
R18423 avss.n7137 avss.n7136 3.4105
R18424 avss.n7134 avss.n7133 3.4105
R18425 avss.n7139 avss.n4114 3.4105
R18426 avss.n4114 avss.n4113 3.4105
R18427 avss.n7148 avss.n7147 3.4105
R18428 avss.n7161 avss.n7160 3.4105
R18429 avss.n7141 avss.n7140 3.4105
R18430 avss.n7156 avss.n7155 3.4105
R18431 avss.n7152 avss.n7151 3.4105
R18432 avss.n7164 avss.n7163 3.4105
R18433 avss.n7165 avss.n7164 3.4105
R18434 avss.n4107 avss.n4106 3.4105
R18435 avss.n4106 avss.n4105 3.4105
R18436 avss.n7169 avss.n7168 3.4105
R18437 avss.n7158 avss.n4093 3.4105
R18438 avss.n7203 avss.n4096 3.4105
R18439 avss.n7170 avss.n4096 3.4105
R18440 avss.n7175 avss.n7174 3.4105
R18441 avss.n7203 avss.n4095 3.4105
R18442 avss.n7176 avss.n4095 3.4105
R18443 avss.n7173 avss.n4104 3.4105
R18444 avss.n4104 avss.n4103 3.4105
R18445 avss.n7179 avss.n4090 3.4105
R18446 avss.n7206 avss.n7205 3.4105
R18447 avss.n7180 avss.n4092 3.4105
R18448 avss.n7185 avss.n4100 3.4105
R18449 avss.n7184 avss.n7183 3.4105
R18450 avss.n7184 avss.n4102 3.4105
R18451 avss.n7193 avss.n7189 3.4105
R18452 avss.n7073 avss.n4146 3.4105
R18453 avss.n4146 avss.n4143 3.4105
R18454 avss.n7074 avss.n4143 3.4105
R18455 avss.n7074 avss.n7073 3.4105
R18456 avss.n7078 avss.n4171 3.4105
R18457 avss.n7081 avss.n7080 3.4105
R18458 avss.n6637 avss.n6636 3.4105
R18459 avss.n6643 avss.n6642 3.4105
R18460 avss.n6647 avss.n6646 3.4105
R18461 avss.n6656 avss.n6609 3.4105
R18462 avss.n6651 avss.n6609 3.4105
R18463 avss.n6623 avss.n6622 3.4105
R18464 avss.n6621 avss.n6612 3.4105
R18465 avss.n6658 avss.n6657 3.4105
R18466 avss.n6656 avss.n6606 3.4105
R18467 avss.n6617 avss.n6606 3.4105
R18468 avss.n6661 avss.n6660 3.4105
R18469 avss.n6664 avss.n6663 3.4105
R18470 avss.n6665 avss.n6664 3.4105
R18471 avss.n6668 avss.n6667 3.4105
R18472 avss.n6596 avss.n6595 3.4105
R18473 avss.n6670 avss.n6598 3.4105
R18474 avss.n6593 avss.n6592 3.4105
R18475 avss.n6677 avss.n6676 3.4105
R18476 avss.n6676 avss.n6675 3.4105
R18477 avss.n6585 avss.n6584 3.4105
R18478 avss.n6579 avss.n6578 3.4105
R18479 avss.n6679 avss.n6678 3.4105
R18480 avss.n6680 avss.n6679 3.4105
R18481 avss.n6576 avss.n6575 3.4105
R18482 avss.n6572 avss.n6569 3.4105
R18483 avss.n6572 avss.n6571 3.4105
R18484 avss.n6686 avss.n6685 3.4105
R18485 avss.n6558 avss.n6552 3.4105
R18486 avss.n6550 avss.n6544 3.4105
R18487 avss.n6690 avss.n6545 3.4105
R18488 avss.n6545 avss.n6543 3.4105
R18489 avss.n6547 avss.n6546 3.4105
R18490 avss.n6699 avss.n6698 3.4105
R18491 avss.n6698 avss.n6697 3.4105
R18492 avss.n6541 avss.n6536 3.4105
R18493 avss.n6506 avss.n6505 3.4105
R18494 avss.n6701 avss.n6700 3.4105
R18495 avss.n6701 avss.n6531 3.4105
R18496 avss.n6710 avss.n6709 3.4105
R18497 avss.n6514 avss.n6507 3.4105
R18498 avss.n6522 avss.n6513 3.4105
R18499 avss.n6513 avss.n6512 3.4105
R18500 avss.n6518 avss.n6515 3.4105
R18501 avss.n6520 avss.n6519 3.4105
R18502 avss.n6526 avss.n6525 3.4105
R18503 avss.n6708 avss.n6707 3.4105
R18504 avss.n6707 avss.n6706 3.4105
R18505 avss.n6703 avss.n6702 3.4105
R18506 avss.n6540 avss.n6539 3.4105
R18507 avss.n6540 avss.n6530 3.4105
R18508 avss.n6694 avss.n6693 3.4105
R18509 avss.n6557 avss.n6556 3.4105
R18510 avss.n6557 avss.n6542 3.4105
R18511 avss.n6684 avss.n6553 3.4105
R18512 avss.n6684 avss.n6683 3.4105
R18513 avss.n6568 avss.n6562 3.4105
R18514 avss.n6566 avss.n6564 3.4105
R18515 avss.n6564 avss.n6563 3.4105
R18516 avss.n6674 avss.n6583 3.4105
R18517 avss.n6666 avss.n6599 3.4105
R18518 avss.n6666 avss.n6587 3.4105
R18519 avss.n6616 avss.n6615 3.4105
R18520 avss.n6620 avss.n6619 3.4105
R18521 avss.n6619 avss.n6611 3.4105
R18522 avss.n6653 avss.n6652 3.4105
R18523 avss.n6648 avss.n6626 3.4105
R18524 avss.n6628 avss.n6626 3.4105
R18525 avss.n6641 avss.n6630 3.4105
R18526 avss.n6630 avss.n6629 3.4105
R18527 avss.n6640 avss.n6639 3.4105
R18528 avss.n6655 avss.n6610 3.4105
R18529 avss.n6655 avss.n6654 3.4105
R18530 avss.n6716 avss.n6504 3.4105
R18531 avss.n6714 avss.n6503 3.4105
R18532 avss.n6529 avss.n6503 3.4105
R18533 avss.n6714 avss.n6713 3.4105
R18534 avss.n6509 avss.n6504 3.4105
R18535 avss.n6717 avss.n6716 3.4105
R18536 avss.n4181 avss.n4175 3.4105
R18537 avss.n6852 avss.n4175 3.4105
R18538 avss.n6846 avss.n6845 3.4105
R18539 avss.n6844 avss.n4185 3.4105
R18540 avss.n6844 avss.n6843 3.4105
R18541 avss.n6837 avss.n6835 3.4105
R18542 avss.n4242 avss.n4241 3.4105
R18543 avss.n4236 avss.n4228 3.4105
R18544 avss.n4240 avss.n4237 3.4105
R18545 avss.n4244 avss.n4235 3.4105
R18546 avss.n4235 avss.n4234 3.4105
R18547 avss.n4248 avss.n4247 3.4105
R18548 avss.n4252 avss.n4251 3.4105
R18549 avss.n4226 avss.n4225 3.4105
R18550 avss.n4225 avss.n4224 3.4105
R18551 avss.n6731 avss.n4222 3.4105
R18552 avss.n6744 avss.n6743 3.4105
R18553 avss.n6724 avss.n6723 3.4105
R18554 avss.n6737 avss.n6736 3.4105
R18555 avss.n6736 avss.n6735 3.4105
R18556 avss.n4219 avss.n4218 3.4105
R18557 avss.n6747 avss.n6746 3.4105
R18558 avss.n6748 avss.n6747 3.4105
R18559 avss.n6733 avss.n6732 3.4105
R18560 avss.n6733 avss.n4217 3.4105
R18561 avss.n6739 avss.n4214 3.4105
R18562 avss.n6741 avss.n6740 3.4105
R18563 avss.n6757 avss.n6756 3.4105
R18564 avss.n6756 avss.n6755 3.4105
R18565 avss.n4215 avss.n4210 3.4105
R18566 avss.n6753 avss.n4216 3.4105
R18567 avss.n6753 avss.n6752 3.4105
R18568 avss.n6763 avss.n4208 3.4105
R18569 avss.n6763 avss.n4203 3.4105
R18570 avss.n6773 avss.n6772 3.4105
R18571 avss.n6762 avss.n6761 3.4105
R18572 avss.n6767 avss.n6766 3.4105
R18573 avss.n6766 avss.n4204 3.4105
R18574 avss.n6775 avss.n6774 3.4105
R18575 avss.n6782 avss.n4202 3.4105
R18576 avss.n6782 avss.n4196 3.4105
R18577 avss.n6791 avss.n4199 3.4105
R18578 avss.n6770 avss.n6769 3.4105
R18579 avss.n6785 avss.n6784 3.4105
R18580 avss.n6784 avss.n6783 3.4105
R18581 avss.n6781 avss.n6780 3.4105
R18582 avss.n6786 avss.n4198 3.4105
R18583 avss.n4198 avss.n4197 3.4105
R18584 avss.n6795 avss.n6794 3.4105
R18585 avss.n6808 avss.n6807 3.4105
R18586 avss.n6788 avss.n6787 3.4105
R18587 avss.n6803 avss.n6802 3.4105
R18588 avss.n6799 avss.n6798 3.4105
R18589 avss.n6811 avss.n6810 3.4105
R18590 avss.n6812 avss.n6811 3.4105
R18591 avss.n4191 avss.n4190 3.4105
R18592 avss.n4190 avss.n4189 3.4105
R18593 avss.n6816 avss.n6815 3.4105
R18594 avss.n6805 avss.n4177 3.4105
R18595 avss.n6850 avss.n4180 3.4105
R18596 avss.n6817 avss.n4180 3.4105
R18597 avss.n6822 avss.n6821 3.4105
R18598 avss.n6850 avss.n4179 3.4105
R18599 avss.n6823 avss.n4179 3.4105
R18600 avss.n6820 avss.n4188 3.4105
R18601 avss.n4188 avss.n4187 3.4105
R18602 avss.n6826 avss.n4174 3.4105
R18603 avss.n6853 avss.n6852 3.4105
R18604 avss.n6827 avss.n4176 3.4105
R18605 avss.n6832 avss.n4184 3.4105
R18606 avss.n6831 avss.n6830 3.4105
R18607 avss.n6831 avss.n4186 3.4105
R18608 avss.n6840 avss.n6836 3.4105
R18609 avss.n6720 avss.n4230 3.4105
R18610 avss.n4230 avss.n4227 3.4105
R18611 avss.n6721 avss.n4227 3.4105
R18612 avss.n6721 avss.n6720 3.4105
R18613 avss.n6725 avss.n4255 3.4105
R18614 avss.n6728 avss.n6727 3.4105
R18615 avss.n6284 avss.n6283 3.4105
R18616 avss.n6290 avss.n6289 3.4105
R18617 avss.n6294 avss.n6293 3.4105
R18618 avss.n6303 avss.n6256 3.4105
R18619 avss.n6298 avss.n6256 3.4105
R18620 avss.n6270 avss.n6269 3.4105
R18621 avss.n6268 avss.n6259 3.4105
R18622 avss.n6305 avss.n6304 3.4105
R18623 avss.n6303 avss.n6253 3.4105
R18624 avss.n6264 avss.n6253 3.4105
R18625 avss.n6308 avss.n6307 3.4105
R18626 avss.n6311 avss.n6310 3.4105
R18627 avss.n6312 avss.n6311 3.4105
R18628 avss.n6315 avss.n6314 3.4105
R18629 avss.n6243 avss.n6242 3.4105
R18630 avss.n6317 avss.n6245 3.4105
R18631 avss.n6240 avss.n6239 3.4105
R18632 avss.n6324 avss.n6323 3.4105
R18633 avss.n6323 avss.n6322 3.4105
R18634 avss.n6232 avss.n6231 3.4105
R18635 avss.n6226 avss.n6225 3.4105
R18636 avss.n6326 avss.n6325 3.4105
R18637 avss.n6327 avss.n6326 3.4105
R18638 avss.n6223 avss.n6222 3.4105
R18639 avss.n6219 avss.n6216 3.4105
R18640 avss.n6219 avss.n6218 3.4105
R18641 avss.n6333 avss.n6332 3.4105
R18642 avss.n6205 avss.n6199 3.4105
R18643 avss.n6197 avss.n6191 3.4105
R18644 avss.n6337 avss.n6192 3.4105
R18645 avss.n6192 avss.n6190 3.4105
R18646 avss.n6194 avss.n6193 3.4105
R18647 avss.n6346 avss.n6345 3.4105
R18648 avss.n6345 avss.n6344 3.4105
R18649 avss.n6188 avss.n6183 3.4105
R18650 avss.n6153 avss.n6152 3.4105
R18651 avss.n6348 avss.n6347 3.4105
R18652 avss.n6348 avss.n6178 3.4105
R18653 avss.n6357 avss.n6356 3.4105
R18654 avss.n6161 avss.n6154 3.4105
R18655 avss.n6169 avss.n6160 3.4105
R18656 avss.n6160 avss.n6159 3.4105
R18657 avss.n6165 avss.n6162 3.4105
R18658 avss.n6167 avss.n6166 3.4105
R18659 avss.n6173 avss.n6172 3.4105
R18660 avss.n6355 avss.n6354 3.4105
R18661 avss.n6354 avss.n6353 3.4105
R18662 avss.n6350 avss.n6349 3.4105
R18663 avss.n6187 avss.n6186 3.4105
R18664 avss.n6187 avss.n6177 3.4105
R18665 avss.n6341 avss.n6340 3.4105
R18666 avss.n6204 avss.n6203 3.4105
R18667 avss.n6204 avss.n6189 3.4105
R18668 avss.n6331 avss.n6200 3.4105
R18669 avss.n6331 avss.n6330 3.4105
R18670 avss.n6215 avss.n6209 3.4105
R18671 avss.n6213 avss.n6211 3.4105
R18672 avss.n6211 avss.n6210 3.4105
R18673 avss.n6321 avss.n6230 3.4105
R18674 avss.n6313 avss.n6246 3.4105
R18675 avss.n6313 avss.n6234 3.4105
R18676 avss.n6263 avss.n6262 3.4105
R18677 avss.n6267 avss.n6266 3.4105
R18678 avss.n6266 avss.n6258 3.4105
R18679 avss.n6300 avss.n6299 3.4105
R18680 avss.n6295 avss.n6273 3.4105
R18681 avss.n6275 avss.n6273 3.4105
R18682 avss.n6288 avss.n6277 3.4105
R18683 avss.n6277 avss.n6276 3.4105
R18684 avss.n6287 avss.n6286 3.4105
R18685 avss.n6302 avss.n6257 3.4105
R18686 avss.n6302 avss.n6301 3.4105
R18687 avss.n6363 avss.n6151 3.4105
R18688 avss.n6361 avss.n6150 3.4105
R18689 avss.n6176 avss.n6150 3.4105
R18690 avss.n6361 avss.n6360 3.4105
R18691 avss.n6156 avss.n6151 3.4105
R18692 avss.n6364 avss.n6363 3.4105
R18693 avss.n4265 avss.n4259 3.4105
R18694 avss.n6499 avss.n4259 3.4105
R18695 avss.n6493 avss.n6492 3.4105
R18696 avss.n6491 avss.n4269 3.4105
R18697 avss.n6491 avss.n6490 3.4105
R18698 avss.n6484 avss.n6482 3.4105
R18699 avss.n4326 avss.n4325 3.4105
R18700 avss.n4320 avss.n4312 3.4105
R18701 avss.n4324 avss.n4321 3.4105
R18702 avss.n4328 avss.n4319 3.4105
R18703 avss.n4319 avss.n4318 3.4105
R18704 avss.n4332 avss.n4331 3.4105
R18705 avss.n4336 avss.n4335 3.4105
R18706 avss.n4310 avss.n4309 3.4105
R18707 avss.n4309 avss.n4308 3.4105
R18708 avss.n6378 avss.n4306 3.4105
R18709 avss.n6391 avss.n6390 3.4105
R18710 avss.n6371 avss.n6370 3.4105
R18711 avss.n6384 avss.n6383 3.4105
R18712 avss.n6383 avss.n6382 3.4105
R18713 avss.n4303 avss.n4302 3.4105
R18714 avss.n6394 avss.n6393 3.4105
R18715 avss.n6395 avss.n6394 3.4105
R18716 avss.n6380 avss.n6379 3.4105
R18717 avss.n6380 avss.n4301 3.4105
R18718 avss.n6386 avss.n4298 3.4105
R18719 avss.n6388 avss.n6387 3.4105
R18720 avss.n6404 avss.n6403 3.4105
R18721 avss.n6403 avss.n6402 3.4105
R18722 avss.n4299 avss.n4294 3.4105
R18723 avss.n6400 avss.n4300 3.4105
R18724 avss.n6400 avss.n6399 3.4105
R18725 avss.n6410 avss.n4292 3.4105
R18726 avss.n6410 avss.n4287 3.4105
R18727 avss.n6420 avss.n6419 3.4105
R18728 avss.n6409 avss.n6408 3.4105
R18729 avss.n6414 avss.n6413 3.4105
R18730 avss.n6413 avss.n4288 3.4105
R18731 avss.n6422 avss.n6421 3.4105
R18732 avss.n6429 avss.n4286 3.4105
R18733 avss.n6429 avss.n4280 3.4105
R18734 avss.n6438 avss.n4283 3.4105
R18735 avss.n6417 avss.n6416 3.4105
R18736 avss.n6432 avss.n6431 3.4105
R18737 avss.n6431 avss.n6430 3.4105
R18738 avss.n6428 avss.n6427 3.4105
R18739 avss.n6433 avss.n4282 3.4105
R18740 avss.n4282 avss.n4281 3.4105
R18741 avss.n6442 avss.n6441 3.4105
R18742 avss.n6455 avss.n6454 3.4105
R18743 avss.n6435 avss.n6434 3.4105
R18744 avss.n6450 avss.n6449 3.4105
R18745 avss.n6446 avss.n6445 3.4105
R18746 avss.n6458 avss.n6457 3.4105
R18747 avss.n6459 avss.n6458 3.4105
R18748 avss.n4275 avss.n4274 3.4105
R18749 avss.n4274 avss.n4273 3.4105
R18750 avss.n6463 avss.n6462 3.4105
R18751 avss.n6452 avss.n4261 3.4105
R18752 avss.n6497 avss.n4264 3.4105
R18753 avss.n6464 avss.n4264 3.4105
R18754 avss.n6469 avss.n6468 3.4105
R18755 avss.n6497 avss.n4263 3.4105
R18756 avss.n6470 avss.n4263 3.4105
R18757 avss.n6467 avss.n4272 3.4105
R18758 avss.n4272 avss.n4271 3.4105
R18759 avss.n6473 avss.n4258 3.4105
R18760 avss.n6500 avss.n6499 3.4105
R18761 avss.n6474 avss.n4260 3.4105
R18762 avss.n6479 avss.n4268 3.4105
R18763 avss.n6478 avss.n6477 3.4105
R18764 avss.n6478 avss.n4270 3.4105
R18765 avss.n6487 avss.n6483 3.4105
R18766 avss.n6367 avss.n4314 3.4105
R18767 avss.n4314 avss.n4311 3.4105
R18768 avss.n6368 avss.n4311 3.4105
R18769 avss.n6368 avss.n6367 3.4105
R18770 avss.n6372 avss.n4339 3.4105
R18771 avss.n6375 avss.n6374 3.4105
R18772 avss.n5931 avss.n5930 3.4105
R18773 avss.n5937 avss.n5936 3.4105
R18774 avss.n5941 avss.n5940 3.4105
R18775 avss.n5950 avss.n5903 3.4105
R18776 avss.n5945 avss.n5903 3.4105
R18777 avss.n5917 avss.n5916 3.4105
R18778 avss.n5915 avss.n5906 3.4105
R18779 avss.n5952 avss.n5951 3.4105
R18780 avss.n5950 avss.n5900 3.4105
R18781 avss.n5911 avss.n5900 3.4105
R18782 avss.n5955 avss.n5954 3.4105
R18783 avss.n5958 avss.n5957 3.4105
R18784 avss.n5959 avss.n5958 3.4105
R18785 avss.n5962 avss.n5961 3.4105
R18786 avss.n5890 avss.n5889 3.4105
R18787 avss.n5964 avss.n5892 3.4105
R18788 avss.n5887 avss.n5886 3.4105
R18789 avss.n5971 avss.n5970 3.4105
R18790 avss.n5970 avss.n5969 3.4105
R18791 avss.n5879 avss.n5878 3.4105
R18792 avss.n5873 avss.n5872 3.4105
R18793 avss.n5973 avss.n5972 3.4105
R18794 avss.n5974 avss.n5973 3.4105
R18795 avss.n5870 avss.n5869 3.4105
R18796 avss.n5866 avss.n5863 3.4105
R18797 avss.n5866 avss.n5865 3.4105
R18798 avss.n5980 avss.n5979 3.4105
R18799 avss.n5852 avss.n5846 3.4105
R18800 avss.n5844 avss.n5838 3.4105
R18801 avss.n5984 avss.n5839 3.4105
R18802 avss.n5839 avss.n5837 3.4105
R18803 avss.n5841 avss.n5840 3.4105
R18804 avss.n5993 avss.n5992 3.4105
R18805 avss.n5992 avss.n5991 3.4105
R18806 avss.n5835 avss.n5830 3.4105
R18807 avss.n5800 avss.n5799 3.4105
R18808 avss.n5995 avss.n5994 3.4105
R18809 avss.n5995 avss.n5825 3.4105
R18810 avss.n6004 avss.n6003 3.4105
R18811 avss.n5808 avss.n5801 3.4105
R18812 avss.n5816 avss.n5807 3.4105
R18813 avss.n5807 avss.n5806 3.4105
R18814 avss.n5812 avss.n5809 3.4105
R18815 avss.n5814 avss.n5813 3.4105
R18816 avss.n5820 avss.n5819 3.4105
R18817 avss.n6002 avss.n6001 3.4105
R18818 avss.n6001 avss.n6000 3.4105
R18819 avss.n5997 avss.n5996 3.4105
R18820 avss.n5834 avss.n5833 3.4105
R18821 avss.n5834 avss.n5824 3.4105
R18822 avss.n5988 avss.n5987 3.4105
R18823 avss.n5851 avss.n5850 3.4105
R18824 avss.n5851 avss.n5836 3.4105
R18825 avss.n5978 avss.n5847 3.4105
R18826 avss.n5978 avss.n5977 3.4105
R18827 avss.n5862 avss.n5856 3.4105
R18828 avss.n5860 avss.n5858 3.4105
R18829 avss.n5858 avss.n5857 3.4105
R18830 avss.n5968 avss.n5877 3.4105
R18831 avss.n5960 avss.n5893 3.4105
R18832 avss.n5960 avss.n5881 3.4105
R18833 avss.n5910 avss.n5909 3.4105
R18834 avss.n5914 avss.n5913 3.4105
R18835 avss.n5913 avss.n5905 3.4105
R18836 avss.n5947 avss.n5946 3.4105
R18837 avss.n5942 avss.n5920 3.4105
R18838 avss.n5922 avss.n5920 3.4105
R18839 avss.n5935 avss.n5924 3.4105
R18840 avss.n5924 avss.n5923 3.4105
R18841 avss.n5934 avss.n5933 3.4105
R18842 avss.n5949 avss.n5904 3.4105
R18843 avss.n5949 avss.n5948 3.4105
R18844 avss.n6010 avss.n5798 3.4105
R18845 avss.n6008 avss.n5797 3.4105
R18846 avss.n5823 avss.n5797 3.4105
R18847 avss.n6008 avss.n6007 3.4105
R18848 avss.n5803 avss.n5798 3.4105
R18849 avss.n6011 avss.n6010 3.4105
R18850 avss.n4349 avss.n4343 3.4105
R18851 avss.n6146 avss.n4343 3.4105
R18852 avss.n6140 avss.n6139 3.4105
R18853 avss.n6138 avss.n4353 3.4105
R18854 avss.n6138 avss.n6137 3.4105
R18855 avss.n6131 avss.n6129 3.4105
R18856 avss.n4410 avss.n4409 3.4105
R18857 avss.n4404 avss.n4396 3.4105
R18858 avss.n4408 avss.n4405 3.4105
R18859 avss.n4412 avss.n4403 3.4105
R18860 avss.n4403 avss.n4402 3.4105
R18861 avss.n4416 avss.n4415 3.4105
R18862 avss.n4420 avss.n4419 3.4105
R18863 avss.n4394 avss.n4393 3.4105
R18864 avss.n4393 avss.n4392 3.4105
R18865 avss.n6025 avss.n4390 3.4105
R18866 avss.n6038 avss.n6037 3.4105
R18867 avss.n6018 avss.n6017 3.4105
R18868 avss.n6031 avss.n6030 3.4105
R18869 avss.n6030 avss.n6029 3.4105
R18870 avss.n4387 avss.n4386 3.4105
R18871 avss.n6041 avss.n6040 3.4105
R18872 avss.n6042 avss.n6041 3.4105
R18873 avss.n6027 avss.n6026 3.4105
R18874 avss.n6027 avss.n4385 3.4105
R18875 avss.n6033 avss.n4382 3.4105
R18876 avss.n6035 avss.n6034 3.4105
R18877 avss.n6051 avss.n6050 3.4105
R18878 avss.n6050 avss.n6049 3.4105
R18879 avss.n4383 avss.n4378 3.4105
R18880 avss.n6047 avss.n4384 3.4105
R18881 avss.n6047 avss.n6046 3.4105
R18882 avss.n6057 avss.n4376 3.4105
R18883 avss.n6057 avss.n4371 3.4105
R18884 avss.n6067 avss.n6066 3.4105
R18885 avss.n6056 avss.n6055 3.4105
R18886 avss.n6061 avss.n6060 3.4105
R18887 avss.n6060 avss.n4372 3.4105
R18888 avss.n6069 avss.n6068 3.4105
R18889 avss.n6076 avss.n4370 3.4105
R18890 avss.n6076 avss.n4364 3.4105
R18891 avss.n6085 avss.n4367 3.4105
R18892 avss.n6064 avss.n6063 3.4105
R18893 avss.n6079 avss.n6078 3.4105
R18894 avss.n6078 avss.n6077 3.4105
R18895 avss.n6075 avss.n6074 3.4105
R18896 avss.n6080 avss.n4366 3.4105
R18897 avss.n4366 avss.n4365 3.4105
R18898 avss.n6089 avss.n6088 3.4105
R18899 avss.n6102 avss.n6101 3.4105
R18900 avss.n6082 avss.n6081 3.4105
R18901 avss.n6097 avss.n6096 3.4105
R18902 avss.n6093 avss.n6092 3.4105
R18903 avss.n6105 avss.n6104 3.4105
R18904 avss.n6106 avss.n6105 3.4105
R18905 avss.n4359 avss.n4358 3.4105
R18906 avss.n4358 avss.n4357 3.4105
R18907 avss.n6110 avss.n6109 3.4105
R18908 avss.n6099 avss.n4345 3.4105
R18909 avss.n6144 avss.n4348 3.4105
R18910 avss.n6111 avss.n4348 3.4105
R18911 avss.n6116 avss.n6115 3.4105
R18912 avss.n6144 avss.n4347 3.4105
R18913 avss.n6117 avss.n4347 3.4105
R18914 avss.n6114 avss.n4356 3.4105
R18915 avss.n4356 avss.n4355 3.4105
R18916 avss.n6120 avss.n4342 3.4105
R18917 avss.n6147 avss.n6146 3.4105
R18918 avss.n6121 avss.n4344 3.4105
R18919 avss.n6126 avss.n4352 3.4105
R18920 avss.n6125 avss.n6124 3.4105
R18921 avss.n6125 avss.n4354 3.4105
R18922 avss.n6134 avss.n6130 3.4105
R18923 avss.n6014 avss.n4398 3.4105
R18924 avss.n4398 avss.n4395 3.4105
R18925 avss.n6015 avss.n4395 3.4105
R18926 avss.n6015 avss.n6014 3.4105
R18927 avss.n6019 avss.n4423 3.4105
R18928 avss.n6022 avss.n6021 3.4105
R18929 avss.n5578 avss.n5577 3.4105
R18930 avss.n5584 avss.n5583 3.4105
R18931 avss.n5588 avss.n5587 3.4105
R18932 avss.n5597 avss.n5550 3.4105
R18933 avss.n5592 avss.n5550 3.4105
R18934 avss.n5564 avss.n5563 3.4105
R18935 avss.n5562 avss.n5553 3.4105
R18936 avss.n5599 avss.n5598 3.4105
R18937 avss.n5597 avss.n5547 3.4105
R18938 avss.n5558 avss.n5547 3.4105
R18939 avss.n5602 avss.n5601 3.4105
R18940 avss.n5605 avss.n5604 3.4105
R18941 avss.n5606 avss.n5605 3.4105
R18942 avss.n5609 avss.n5608 3.4105
R18943 avss.n5537 avss.n5536 3.4105
R18944 avss.n5611 avss.n5539 3.4105
R18945 avss.n5534 avss.n5533 3.4105
R18946 avss.n5618 avss.n5617 3.4105
R18947 avss.n5617 avss.n5616 3.4105
R18948 avss.n5526 avss.n5525 3.4105
R18949 avss.n5520 avss.n5519 3.4105
R18950 avss.n5620 avss.n5619 3.4105
R18951 avss.n5621 avss.n5620 3.4105
R18952 avss.n5517 avss.n5516 3.4105
R18953 avss.n5513 avss.n5510 3.4105
R18954 avss.n5513 avss.n5512 3.4105
R18955 avss.n5627 avss.n5626 3.4105
R18956 avss.n5499 avss.n5493 3.4105
R18957 avss.n5491 avss.n5485 3.4105
R18958 avss.n5631 avss.n5486 3.4105
R18959 avss.n5486 avss.n5484 3.4105
R18960 avss.n5488 avss.n5487 3.4105
R18961 avss.n5640 avss.n5639 3.4105
R18962 avss.n5639 avss.n5638 3.4105
R18963 avss.n5482 avss.n5477 3.4105
R18964 avss.n5447 avss.n5446 3.4105
R18965 avss.n5642 avss.n5641 3.4105
R18966 avss.n5642 avss.n5472 3.4105
R18967 avss.n5651 avss.n5650 3.4105
R18968 avss.n5455 avss.n5448 3.4105
R18969 avss.n5463 avss.n5454 3.4105
R18970 avss.n5454 avss.n5453 3.4105
R18971 avss.n5459 avss.n5456 3.4105
R18972 avss.n5461 avss.n5460 3.4105
R18973 avss.n5467 avss.n5466 3.4105
R18974 avss.n5649 avss.n5648 3.4105
R18975 avss.n5648 avss.n5647 3.4105
R18976 avss.n5644 avss.n5643 3.4105
R18977 avss.n5481 avss.n5480 3.4105
R18978 avss.n5481 avss.n5471 3.4105
R18979 avss.n5635 avss.n5634 3.4105
R18980 avss.n5498 avss.n5497 3.4105
R18981 avss.n5498 avss.n5483 3.4105
R18982 avss.n5625 avss.n5494 3.4105
R18983 avss.n5625 avss.n5624 3.4105
R18984 avss.n5509 avss.n5503 3.4105
R18985 avss.n5507 avss.n5505 3.4105
R18986 avss.n5505 avss.n5504 3.4105
R18987 avss.n5615 avss.n5524 3.4105
R18988 avss.n5607 avss.n5540 3.4105
R18989 avss.n5607 avss.n5528 3.4105
R18990 avss.n5557 avss.n5556 3.4105
R18991 avss.n5561 avss.n5560 3.4105
R18992 avss.n5560 avss.n5552 3.4105
R18993 avss.n5594 avss.n5593 3.4105
R18994 avss.n5589 avss.n5567 3.4105
R18995 avss.n5569 avss.n5567 3.4105
R18996 avss.n5582 avss.n5571 3.4105
R18997 avss.n5571 avss.n5570 3.4105
R18998 avss.n5581 avss.n5580 3.4105
R18999 avss.n5596 avss.n5551 3.4105
R19000 avss.n5596 avss.n5595 3.4105
R19001 avss.n5657 avss.n5445 3.4105
R19002 avss.n5655 avss.n5444 3.4105
R19003 avss.n5470 avss.n5444 3.4105
R19004 avss.n5655 avss.n5654 3.4105
R19005 avss.n5450 avss.n5445 3.4105
R19006 avss.n5658 avss.n5657 3.4105
R19007 avss.n4433 avss.n4427 3.4105
R19008 avss.n5793 avss.n4427 3.4105
R19009 avss.n5787 avss.n5786 3.4105
R19010 avss.n5785 avss.n4437 3.4105
R19011 avss.n5785 avss.n5784 3.4105
R19012 avss.n5778 avss.n5776 3.4105
R19013 avss.n4494 avss.n4493 3.4105
R19014 avss.n4488 avss.n4480 3.4105
R19015 avss.n4492 avss.n4489 3.4105
R19016 avss.n4496 avss.n4487 3.4105
R19017 avss.n4487 avss.n4486 3.4105
R19018 avss.n4500 avss.n4499 3.4105
R19019 avss.n4504 avss.n4503 3.4105
R19020 avss.n4478 avss.n4477 3.4105
R19021 avss.n4477 avss.n4476 3.4105
R19022 avss.n5672 avss.n4474 3.4105
R19023 avss.n5685 avss.n5684 3.4105
R19024 avss.n5665 avss.n5664 3.4105
R19025 avss.n5678 avss.n5677 3.4105
R19026 avss.n5677 avss.n5676 3.4105
R19027 avss.n4471 avss.n4470 3.4105
R19028 avss.n5688 avss.n5687 3.4105
R19029 avss.n5689 avss.n5688 3.4105
R19030 avss.n5674 avss.n5673 3.4105
R19031 avss.n5674 avss.n4469 3.4105
R19032 avss.n5680 avss.n4466 3.4105
R19033 avss.n5682 avss.n5681 3.4105
R19034 avss.n5698 avss.n5697 3.4105
R19035 avss.n5697 avss.n5696 3.4105
R19036 avss.n4467 avss.n4462 3.4105
R19037 avss.n5694 avss.n4468 3.4105
R19038 avss.n5694 avss.n5693 3.4105
R19039 avss.n5704 avss.n4460 3.4105
R19040 avss.n5704 avss.n4455 3.4105
R19041 avss.n5714 avss.n5713 3.4105
R19042 avss.n5703 avss.n5702 3.4105
R19043 avss.n5708 avss.n5707 3.4105
R19044 avss.n5707 avss.n4456 3.4105
R19045 avss.n5716 avss.n5715 3.4105
R19046 avss.n5723 avss.n4454 3.4105
R19047 avss.n5723 avss.n4448 3.4105
R19048 avss.n5732 avss.n4451 3.4105
R19049 avss.n5711 avss.n5710 3.4105
R19050 avss.n5726 avss.n5725 3.4105
R19051 avss.n5725 avss.n5724 3.4105
R19052 avss.n5722 avss.n5721 3.4105
R19053 avss.n5727 avss.n4450 3.4105
R19054 avss.n4450 avss.n4449 3.4105
R19055 avss.n5736 avss.n5735 3.4105
R19056 avss.n5749 avss.n5748 3.4105
R19057 avss.n5729 avss.n5728 3.4105
R19058 avss.n5744 avss.n5743 3.4105
R19059 avss.n5740 avss.n5739 3.4105
R19060 avss.n5752 avss.n5751 3.4105
R19061 avss.n5753 avss.n5752 3.4105
R19062 avss.n4443 avss.n4442 3.4105
R19063 avss.n4442 avss.n4441 3.4105
R19064 avss.n5757 avss.n5756 3.4105
R19065 avss.n5746 avss.n4429 3.4105
R19066 avss.n5791 avss.n4432 3.4105
R19067 avss.n5758 avss.n4432 3.4105
R19068 avss.n5763 avss.n5762 3.4105
R19069 avss.n5791 avss.n4431 3.4105
R19070 avss.n5764 avss.n4431 3.4105
R19071 avss.n5761 avss.n4440 3.4105
R19072 avss.n4440 avss.n4439 3.4105
R19073 avss.n5767 avss.n4426 3.4105
R19074 avss.n5794 avss.n5793 3.4105
R19075 avss.n5768 avss.n4428 3.4105
R19076 avss.n5773 avss.n4436 3.4105
R19077 avss.n5772 avss.n5771 3.4105
R19078 avss.n5772 avss.n4438 3.4105
R19079 avss.n5781 avss.n5777 3.4105
R19080 avss.n5661 avss.n4482 3.4105
R19081 avss.n4482 avss.n4479 3.4105
R19082 avss.n5662 avss.n4479 3.4105
R19083 avss.n5662 avss.n5661 3.4105
R19084 avss.n5666 avss.n4507 3.4105
R19085 avss.n5669 avss.n5668 3.4105
R19086 avss.n5237 avss.n5236 3.4105
R19087 avss.n5243 avss.n5242 3.4105
R19088 avss.n5229 avss.n5210 3.4105
R19089 avss.n5222 avss.n5213 3.4105
R19090 avss.n5254 avss.n5253 3.4105
R19091 avss.n5257 avss.n5256 3.4105
R19092 avss.n5260 avss.n5259 3.4105
R19093 avss.n5261 avss.n5260 3.4105
R19094 avss.n5264 avss.n5263 3.4105
R19095 avss.n5191 avss.n5190 3.4105
R19096 avss.n5266 avss.n5193 3.4105
R19097 avss.n5188 avss.n5187 3.4105
R19098 avss.n5273 avss.n5272 3.4105
R19099 avss.n5272 avss.n5271 3.4105
R19100 avss.n5180 avss.n5179 3.4105
R19101 avss.n5174 avss.n5173 3.4105
R19102 avss.n5275 avss.n5274 3.4105
R19103 avss.n5276 avss.n5275 3.4105
R19104 avss.n5171 avss.n5170 3.4105
R19105 avss.n5167 avss.n5164 3.4105
R19106 avss.n5167 avss.n5166 3.4105
R19107 avss.n5282 avss.n5281 3.4105
R19108 avss.n5153 avss.n5147 3.4105
R19109 avss.n5145 avss.n5135 3.4105
R19110 avss.n5286 avss.n5136 3.4105
R19111 avss.n5136 avss.n5134 3.4105
R19112 avss.n5142 avss.n5137 3.4105
R19113 avss.n5139 avss.n5093 3.4105
R19114 avss.n5139 avss.n5132 3.4105
R19115 avss.n5138 avss.n5097 3.4105
R19116 avss.n5301 avss.n5300 3.4105
R19117 avss.n5298 avss.n5297 3.4105
R19118 avss.n5297 avss.n5296 3.4105
R19119 avss.n5091 avss.n5089 3.4105
R19120 avss.n5129 avss.n5091 3.4105
R19121 avss.n5126 avss.n5100 3.4105
R19122 avss.n5116 avss.n5107 3.4105
R19123 avss.n5115 avss.n5105 3.4105
R19124 avss.n5105 avss.n5104 3.4105
R19125 avss.n5111 avss.n5108 3.4105
R19126 avss.n5113 avss.n5112 3.4105
R19127 avss.n5120 avss.n5119 3.4105
R19128 avss.n5128 avss.n5127 3.4105
R19129 avss.n5128 avss.n5099 3.4105
R19130 avss.n5096 avss.n5094 3.4105
R19131 avss.n5294 avss.n5098 3.4105
R19132 avss.n5294 avss.n5293 3.4105
R19133 avss.n5290 avss.n5289 3.4105
R19134 avss.n5152 avss.n5151 3.4105
R19135 avss.n5152 avss.n5133 3.4105
R19136 avss.n5280 avss.n5148 3.4105
R19137 avss.n5280 avss.n5279 3.4105
R19138 avss.n5163 avss.n5157 3.4105
R19139 avss.n5161 avss.n5159 3.4105
R19140 avss.n5159 avss.n5158 3.4105
R19141 avss.n5270 avss.n5178 3.4105
R19142 avss.n5262 avss.n5194 3.4105
R19143 avss.n5262 avss.n5182 3.4105
R19144 avss.n5217 avss.n5216 3.4105
R19145 avss.n5221 avss.n5220 3.4105
R19146 avss.n5220 avss.n5212 3.4105
R19147 avss.n5209 avss.n5208 3.4105
R19148 avss.n5247 avss.n5211 3.4105
R19149 avss.n5247 avss.n5246 3.4105
R19150 avss.n5241 avss.n5228 3.4105
R19151 avss.n5228 avss.n5227 3.4105
R19152 avss.n5240 avss.n5239 3.4105
R19153 avss.n5305 avss.n5090 3.4105
R19154 avss.n5305 avss.n5304 3.4105
R19155 avss.n5250 avss.n5249 3.4105
R19156 avss.n5206 avss.n5200 3.4105
R19157 avss.n5204 avss.n5200 3.4105
R19158 avss.n5224 avss.n5223 3.4105
R19159 avss.n5252 avss.n5201 3.4105
R19160 avss.n5218 avss.n5201 3.4105
R19161 avss.n5204 avss.n5203 3.4105
R19162 avss.n5206 avss.n5203 3.4105
R19163 avss.n4517 avss.n4511 3.4105
R19164 avss.n5440 avss.n4511 3.4105
R19165 avss.n5434 avss.n5433 3.4105
R19166 avss.n5432 avss.n4521 3.4105
R19167 avss.n5432 avss.n5431 3.4105
R19168 avss.n5425 avss.n5423 3.4105
R19169 avss.n4578 avss.n4577 3.4105
R19170 avss.n4572 avss.n4564 3.4105
R19171 avss.n4576 avss.n4573 3.4105
R19172 avss.n4580 avss.n4571 3.4105
R19173 avss.n4571 avss.n4570 3.4105
R19174 avss.n4584 avss.n4583 3.4105
R19175 avss.n4588 avss.n4587 3.4105
R19176 avss.n4562 avss.n4561 3.4105
R19177 avss.n4561 avss.n4560 3.4105
R19178 avss.n5319 avss.n4558 3.4105
R19179 avss.n5332 avss.n5331 3.4105
R19180 avss.n5312 avss.n5311 3.4105
R19181 avss.n5325 avss.n5324 3.4105
R19182 avss.n5324 avss.n5323 3.4105
R19183 avss.n4555 avss.n4554 3.4105
R19184 avss.n5335 avss.n5334 3.4105
R19185 avss.n5336 avss.n5335 3.4105
R19186 avss.n5321 avss.n5320 3.4105
R19187 avss.n5321 avss.n4553 3.4105
R19188 avss.n5327 avss.n4550 3.4105
R19189 avss.n5329 avss.n5328 3.4105
R19190 avss.n5345 avss.n5344 3.4105
R19191 avss.n5344 avss.n5343 3.4105
R19192 avss.n4551 avss.n4546 3.4105
R19193 avss.n5341 avss.n4552 3.4105
R19194 avss.n5341 avss.n5340 3.4105
R19195 avss.n5351 avss.n4544 3.4105
R19196 avss.n5351 avss.n4539 3.4105
R19197 avss.n5361 avss.n5360 3.4105
R19198 avss.n5350 avss.n5349 3.4105
R19199 avss.n5355 avss.n5354 3.4105
R19200 avss.n5354 avss.n4540 3.4105
R19201 avss.n5363 avss.n5362 3.4105
R19202 avss.n5370 avss.n4538 3.4105
R19203 avss.n5370 avss.n4532 3.4105
R19204 avss.n5379 avss.n4535 3.4105
R19205 avss.n5358 avss.n5357 3.4105
R19206 avss.n5373 avss.n5372 3.4105
R19207 avss.n5372 avss.n5371 3.4105
R19208 avss.n5369 avss.n5368 3.4105
R19209 avss.n5374 avss.n4534 3.4105
R19210 avss.n4534 avss.n4533 3.4105
R19211 avss.n5383 avss.n5382 3.4105
R19212 avss.n5396 avss.n5395 3.4105
R19213 avss.n5376 avss.n5375 3.4105
R19214 avss.n5391 avss.n5390 3.4105
R19215 avss.n5387 avss.n5386 3.4105
R19216 avss.n5399 avss.n5398 3.4105
R19217 avss.n5400 avss.n5399 3.4105
R19218 avss.n4527 avss.n4526 3.4105
R19219 avss.n4526 avss.n4525 3.4105
R19220 avss.n5404 avss.n5403 3.4105
R19221 avss.n5393 avss.n4513 3.4105
R19222 avss.n5438 avss.n4516 3.4105
R19223 avss.n5405 avss.n4516 3.4105
R19224 avss.n5410 avss.n5409 3.4105
R19225 avss.n5438 avss.n4515 3.4105
R19226 avss.n5411 avss.n4515 3.4105
R19227 avss.n5408 avss.n4524 3.4105
R19228 avss.n4524 avss.n4523 3.4105
R19229 avss.n5414 avss.n4510 3.4105
R19230 avss.n5441 avss.n5440 3.4105
R19231 avss.n5415 avss.n4512 3.4105
R19232 avss.n5420 avss.n4520 3.4105
R19233 avss.n5419 avss.n5418 3.4105
R19234 avss.n5419 avss.n4522 3.4105
R19235 avss.n5428 avss.n5424 3.4105
R19236 avss.n5308 avss.n4566 3.4105
R19237 avss.n4566 avss.n4563 3.4105
R19238 avss.n5309 avss.n4563 3.4105
R19239 avss.n5309 avss.n5308 3.4105
R19240 avss.n5313 avss.n4591 3.4105
R19241 avss.n5316 avss.n5315 3.4105
R19242 avss.n4883 avss.n4882 3.4105
R19243 avss.n4889 avss.n4888 3.4105
R19244 avss.n4875 avss.n4856 3.4105
R19245 avss.n4868 avss.n4859 3.4105
R19246 avss.n4900 avss.n4899 3.4105
R19247 avss.n4903 avss.n4902 3.4105
R19248 avss.n4906 avss.n4905 3.4105
R19249 avss.n4907 avss.n4906 3.4105
R19250 avss.n4910 avss.n4909 3.4105
R19251 avss.n4837 avss.n4836 3.4105
R19252 avss.n4912 avss.n4839 3.4105
R19253 avss.n4834 avss.n4833 3.4105
R19254 avss.n4919 avss.n4918 3.4105
R19255 avss.n4918 avss.n4917 3.4105
R19256 avss.n4826 avss.n4825 3.4105
R19257 avss.n4820 avss.n4819 3.4105
R19258 avss.n4921 avss.n4920 3.4105
R19259 avss.n4922 avss.n4921 3.4105
R19260 avss.n4817 avss.n4816 3.4105
R19261 avss.n4813 avss.n4810 3.4105
R19262 avss.n4813 avss.n4812 3.4105
R19263 avss.n4928 avss.n4927 3.4105
R19264 avss.n4799 avss.n4793 3.4105
R19265 avss.n4791 avss.n4781 3.4105
R19266 avss.n4932 avss.n4782 3.4105
R19267 avss.n4782 avss.n4780 3.4105
R19268 avss.n4788 avss.n4783 3.4105
R19269 avss.n4785 avss.n4739 3.4105
R19270 avss.n4785 avss.n4778 3.4105
R19271 avss.n4784 avss.n4743 3.4105
R19272 avss.n4947 avss.n4946 3.4105
R19273 avss.n4944 avss.n4943 3.4105
R19274 avss.n4943 avss.n4942 3.4105
R19275 avss.n4737 avss.n4735 3.4105
R19276 avss.n4775 avss.n4737 3.4105
R19277 avss.n4772 avss.n4746 3.4105
R19278 avss.n4762 avss.n4753 3.4105
R19279 avss.n4761 avss.n4751 3.4105
R19280 avss.n4751 avss.n4750 3.4105
R19281 avss.n4757 avss.n4754 3.4105
R19282 avss.n4759 avss.n4758 3.4105
R19283 avss.n4766 avss.n4765 3.4105
R19284 avss.n4774 avss.n4773 3.4105
R19285 avss.n4774 avss.n4745 3.4105
R19286 avss.n4742 avss.n4740 3.4105
R19287 avss.n4940 avss.n4744 3.4105
R19288 avss.n4940 avss.n4939 3.4105
R19289 avss.n4936 avss.n4935 3.4105
R19290 avss.n4798 avss.n4797 3.4105
R19291 avss.n4798 avss.n4779 3.4105
R19292 avss.n4926 avss.n4794 3.4105
R19293 avss.n4926 avss.n4925 3.4105
R19294 avss.n4809 avss.n4803 3.4105
R19295 avss.n4807 avss.n4805 3.4105
R19296 avss.n4805 avss.n4804 3.4105
R19297 avss.n4916 avss.n4824 3.4105
R19298 avss.n4908 avss.n4840 3.4105
R19299 avss.n4908 avss.n4828 3.4105
R19300 avss.n4863 avss.n4862 3.4105
R19301 avss.n4867 avss.n4866 3.4105
R19302 avss.n4866 avss.n4858 3.4105
R19303 avss.n4855 avss.n4854 3.4105
R19304 avss.n4893 avss.n4857 3.4105
R19305 avss.n4893 avss.n4892 3.4105
R19306 avss.n4887 avss.n4874 3.4105
R19307 avss.n4874 avss.n4873 3.4105
R19308 avss.n4886 avss.n4885 3.4105
R19309 avss.n4951 avss.n4736 3.4105
R19310 avss.n4951 avss.n4950 3.4105
R19311 avss.n4896 avss.n4895 3.4105
R19312 avss.n4852 avss.n4846 3.4105
R19313 avss.n4850 avss.n4846 3.4105
R19314 avss.n4870 avss.n4869 3.4105
R19315 avss.n4898 avss.n4847 3.4105
R19316 avss.n4864 avss.n4847 3.4105
R19317 avss.n4850 avss.n4849 3.4105
R19318 avss.n4852 avss.n4849 3.4105
R19319 avss.n4601 avss.n4595 3.4105
R19320 avss.n5086 avss.n4595 3.4105
R19321 avss.n5080 avss.n5079 3.4105
R19322 avss.n5078 avss.n4605 3.4105
R19323 avss.n5078 avss.n5077 3.4105
R19324 avss.n5071 avss.n5069 3.4105
R19325 avss.n4662 avss.n4661 3.4105
R19326 avss.n4656 avss.n4648 3.4105
R19327 avss.n4660 avss.n4657 3.4105
R19328 avss.n4664 avss.n4655 3.4105
R19329 avss.n4655 avss.n4654 3.4105
R19330 avss.n4668 avss.n4667 3.4105
R19331 avss.n4672 avss.n4671 3.4105
R19332 avss.n4646 avss.n4645 3.4105
R19333 avss.n4645 avss.n4644 3.4105
R19334 avss.n4965 avss.n4642 3.4105
R19335 avss.n4978 avss.n4977 3.4105
R19336 avss.n4958 avss.n4957 3.4105
R19337 avss.n4971 avss.n4970 3.4105
R19338 avss.n4970 avss.n4969 3.4105
R19339 avss.n4639 avss.n4638 3.4105
R19340 avss.n4981 avss.n4980 3.4105
R19341 avss.n4982 avss.n4981 3.4105
R19342 avss.n4967 avss.n4966 3.4105
R19343 avss.n4967 avss.n4637 3.4105
R19344 avss.n4973 avss.n4634 3.4105
R19345 avss.n4975 avss.n4974 3.4105
R19346 avss.n4991 avss.n4990 3.4105
R19347 avss.n4990 avss.n4989 3.4105
R19348 avss.n4635 avss.n4630 3.4105
R19349 avss.n4987 avss.n4636 3.4105
R19350 avss.n4987 avss.n4986 3.4105
R19351 avss.n4997 avss.n4628 3.4105
R19352 avss.n4997 avss.n4623 3.4105
R19353 avss.n5007 avss.n5006 3.4105
R19354 avss.n4996 avss.n4995 3.4105
R19355 avss.n5001 avss.n5000 3.4105
R19356 avss.n5000 avss.n4624 3.4105
R19357 avss.n5009 avss.n5008 3.4105
R19358 avss.n5016 avss.n4622 3.4105
R19359 avss.n5016 avss.n4616 3.4105
R19360 avss.n5025 avss.n4619 3.4105
R19361 avss.n5004 avss.n5003 3.4105
R19362 avss.n5019 avss.n5018 3.4105
R19363 avss.n5018 avss.n5017 3.4105
R19364 avss.n5015 avss.n5014 3.4105
R19365 avss.n5020 avss.n4618 3.4105
R19366 avss.n4618 avss.n4617 3.4105
R19367 avss.n5029 avss.n5028 3.4105
R19368 avss.n5042 avss.n5041 3.4105
R19369 avss.n5022 avss.n5021 3.4105
R19370 avss.n5037 avss.n5036 3.4105
R19371 avss.n5033 avss.n5032 3.4105
R19372 avss.n5045 avss.n5044 3.4105
R19373 avss.n5046 avss.n5045 3.4105
R19374 avss.n4611 avss.n4610 3.4105
R19375 avss.n4610 avss.n4609 3.4105
R19376 avss.n5050 avss.n5049 3.4105
R19377 avss.n5039 avss.n4597 3.4105
R19378 avss.n5084 avss.n4600 3.4105
R19379 avss.n5051 avss.n4600 3.4105
R19380 avss.n5056 avss.n5055 3.4105
R19381 avss.n5084 avss.n4599 3.4105
R19382 avss.n5057 avss.n4599 3.4105
R19383 avss.n5054 avss.n4608 3.4105
R19384 avss.n4608 avss.n4607 3.4105
R19385 avss.n5060 avss.n4594 3.4105
R19386 avss.n5087 avss.n5086 3.4105
R19387 avss.n5061 avss.n4596 3.4105
R19388 avss.n5066 avss.n4604 3.4105
R19389 avss.n5065 avss.n5064 3.4105
R19390 avss.n5065 avss.n4606 3.4105
R19391 avss.n5074 avss.n5070 3.4105
R19392 avss.n4954 avss.n4650 3.4105
R19393 avss.n4650 avss.n4647 3.4105
R19394 avss.n4955 avss.n4647 3.4105
R19395 avss.n4955 avss.n4954 3.4105
R19396 avss.n4959 avss.n4675 3.4105
R19397 avss.n4962 avss.n4961 3.4105
R19398 avss.n3344 avss.n3343 3.39706
R19399 avss.n3382 avss.n3277 3.38874
R19400 avss.n3382 avss.n3274 3.38874
R19401 avss.n3014 avss.n2947 3.2005
R19402 avss.n3072 avss.n2931 3.2005
R19403 avss.n3102 avss.n3093 3.2005
R19404 avss.n3663 avss.n2597 3.2005
R19405 avss.n2726 avss.n2660 3.2005
R19406 avss.n2771 avss.n2633 3.2005
R19407 avss.n2876 avss.n2791 3.2005
R19408 avss.n2836 avss.n2827 3.2005
R19409 avss.n3360 avss.n3357 3.16936
R19410 avss.n3383 avss.n3276 3.16936
R19411 avss.n11631 avss 3.09989
R19412 avss.n3355 avss.n3290 3.01226
R19413 avss.n3377 avss.n3277 3.01226
R19414 avss.n3387 avss.n3274 3.01226
R19415 avss.n2976 avss.n2963 3.00679
R19416 avss.n3033 avss.n3020 3.00679
R19417 avss.n2927 avss.n2926 3.00679
R19418 avss.n3625 avss.n2611 3.00679
R19419 avss.n3353 avss.n3285 3.0005
R19420 avss.n3363 avss.n3362 3.0005
R19421 avss.n3392 avss.n3391 3.0005
R19422 avss.n3462 avss.n3461 3.0005
R19423 avss.n3512 avss.n3174 3.0005
R19424 avss.n3348 avss.n3347 3.0005
R19425 avss.n2809 avss.n2794 2.99647
R19426 avss.n2912 avss.n2629 2.99647
R19427 avss.n2657 avss.n2646 2.99647
R19428 avss.n2684 avss.n2673 2.99647
R19429 avss.n3248 avss.t369 2.89714
R19430 avss.n3346 avss.n3290 2.63579
R19431 avss.n3361 avss.n3288 2.63579
R19432 avss.n3013 avss.n2945 2.63064
R19433 avss.n3071 avss.n3070 2.63064
R19434 avss.n3100 avss.n3099 2.63064
R19435 avss.n3662 avss.n2595 2.63064
R19436 avss.n2725 avss.n2658 2.63064
R19437 avss.n2770 avss.n2631 2.63064
R19438 avss.n2874 avss.n2873 2.63064
R19439 avss.n2834 avss.n2833 2.63064
R19440 avss.n3354 avss.n3291 2.25932
R19441 avss.n3369 avss.n3283 2.25932
R19442 avss.n3376 avss.n3279 2.25932
R19443 avss.n3405 avss.n3404 2.25932
R19444 avss.n3420 avss.n3419 2.25932
R19445 avss.n8973 avss 2.19212
R19446 avss avss.n8973 2.16596
R19447 avss.n8645 avss.n8629 2.02873
R19448 avss.n8292 avss.n8276 2.02873
R19449 avss.n7939 avss.n7923 2.02873
R19450 avss.n7586 avss.n7570 2.02873
R19451 avss.n7233 avss.n7217 2.02873
R19452 avss.n6880 avss.n6864 2.02873
R19453 avss.n6527 avss.n6511 2.02873
R19454 avss.n6174 avss.n6158 2.02873
R19455 avss.n5821 avss.n5805 2.02873
R19456 avss.n5468 avss.n5452 2.02873
R19457 avss.n5121 avss.n5103 2.02873
R19458 avss.n4767 avss.n4749 2.02873
R19459 avss.n3745 avss.n3729 2.02855
R19460 avss.n3829 avss.n3813 2.02855
R19461 avss.n3913 avss.n3897 2.02855
R19462 avss.n3997 avss.n3981 2.02855
R19463 avss.n4081 avss.n4065 2.02855
R19464 avss.n4165 avss.n4149 2.02855
R19465 avss.n4249 avss.n4233 2.02855
R19466 avss.n4333 avss.n4317 2.02855
R19467 avss.n4417 avss.n4401 2.02855
R19468 avss.n4501 avss.n4485 2.02855
R19469 avss.n4585 avss.n4569 2.02855
R19470 avss.n4669 avss.n4653 2.02855
R19471 avss.n8751 avss.n8747 2.0141
R19472 avss.n8961 avss.n8960 2.0141
R19473 avss.n8398 avss.n8394 2.0141
R19474 avss.n8608 avss.n8607 2.0141
R19475 avss.n8045 avss.n8041 2.0141
R19476 avss.n8255 avss.n8254 2.0141
R19477 avss.n7692 avss.n7688 2.0141
R19478 avss.n7902 avss.n7901 2.0141
R19479 avss.n7339 avss.n7335 2.0141
R19480 avss.n7549 avss.n7548 2.0141
R19481 avss.n6986 avss.n6982 2.0141
R19482 avss.n7196 avss.n7195 2.0141
R19483 avss.n6633 avss.n6629 2.0141
R19484 avss.n6843 avss.n6842 2.0141
R19485 avss.n6280 avss.n6276 2.0141
R19486 avss.n6490 avss.n6489 2.0141
R19487 avss.n5927 avss.n5923 2.0141
R19488 avss.n6137 avss.n6136 2.0141
R19489 avss.n5574 avss.n5570 2.0141
R19490 avss.n5784 avss.n5783 2.0141
R19491 avss.n5233 avss.n5227 2.0141
R19492 avss.n5431 avss.n5430 2.0141
R19493 avss.n4879 avss.n4873 2.0141
R19494 avss.n5077 avss.n5076 2.0141
R19495 avss.n8770 avss.n8743 1.93672
R19496 avss.n8734 avss.n8732 1.93672
R19497 avss.n8790 avss.n8789 1.93672
R19498 avss.n8792 avss.n8791 1.93672
R19499 avss.n8800 avss.n8680 1.93672
R19500 avss.n8813 avss.n8812 1.93672
R19501 avss.n8822 avss.n8821 1.93672
R19502 avss.n8645 avss.n8644 1.93672
R19503 avss.n8830 avss.n8646 1.93672
R19504 avss.n3745 avss.n3744 1.93672
R19505 avss.n8849 avss.n8848 1.93672
R19506 avss.n8868 avss.n3710 1.93672
R19507 avss.n8894 avss.n8893 1.93672
R19508 avss.n8914 avss.n8913 1.93672
R19509 avss.n8934 avss.n8932 1.93672
R19510 avss.n8944 avss.n8943 1.93672
R19511 avss.n3750 avss.n3746 1.93672
R19512 avss.n8919 avss.n8915 1.93672
R19513 avss.n8417 avss.n8390 1.93672
R19514 avss.n8381 avss.n8379 1.93672
R19515 avss.n8437 avss.n8436 1.93672
R19516 avss.n8439 avss.n8438 1.93672
R19517 avss.n8447 avss.n8327 1.93672
R19518 avss.n8460 avss.n8459 1.93672
R19519 avss.n8469 avss.n8468 1.93672
R19520 avss.n8292 avss.n8291 1.93672
R19521 avss.n8477 avss.n8293 1.93672
R19522 avss.n3829 avss.n3828 1.93672
R19523 avss.n8496 avss.n8495 1.93672
R19524 avss.n8515 avss.n3794 1.93672
R19525 avss.n8541 avss.n8540 1.93672
R19526 avss.n8561 avss.n8560 1.93672
R19527 avss.n8581 avss.n8579 1.93672
R19528 avss.n8591 avss.n8590 1.93672
R19529 avss.n3834 avss.n3830 1.93672
R19530 avss.n8566 avss.n8562 1.93672
R19531 avss.n8064 avss.n8037 1.93672
R19532 avss.n8028 avss.n8026 1.93672
R19533 avss.n8084 avss.n8083 1.93672
R19534 avss.n8086 avss.n8085 1.93672
R19535 avss.n8094 avss.n7974 1.93672
R19536 avss.n8107 avss.n8106 1.93672
R19537 avss.n8116 avss.n8115 1.93672
R19538 avss.n7939 avss.n7938 1.93672
R19539 avss.n8124 avss.n7940 1.93672
R19540 avss.n3913 avss.n3912 1.93672
R19541 avss.n8143 avss.n8142 1.93672
R19542 avss.n8162 avss.n3878 1.93672
R19543 avss.n8188 avss.n8187 1.93672
R19544 avss.n8208 avss.n8207 1.93672
R19545 avss.n8228 avss.n8226 1.93672
R19546 avss.n8238 avss.n8237 1.93672
R19547 avss.n3918 avss.n3914 1.93672
R19548 avss.n8213 avss.n8209 1.93672
R19549 avss.n7711 avss.n7684 1.93672
R19550 avss.n7675 avss.n7673 1.93672
R19551 avss.n7731 avss.n7730 1.93672
R19552 avss.n7733 avss.n7732 1.93672
R19553 avss.n7741 avss.n7621 1.93672
R19554 avss.n7754 avss.n7753 1.93672
R19555 avss.n7763 avss.n7762 1.93672
R19556 avss.n7586 avss.n7585 1.93672
R19557 avss.n7771 avss.n7587 1.93672
R19558 avss.n3997 avss.n3996 1.93672
R19559 avss.n7790 avss.n7789 1.93672
R19560 avss.n7809 avss.n3962 1.93672
R19561 avss.n7835 avss.n7834 1.93672
R19562 avss.n7855 avss.n7854 1.93672
R19563 avss.n7875 avss.n7873 1.93672
R19564 avss.n7885 avss.n7884 1.93672
R19565 avss.n4002 avss.n3998 1.93672
R19566 avss.n7860 avss.n7856 1.93672
R19567 avss.n7358 avss.n7331 1.93672
R19568 avss.n7322 avss.n7320 1.93672
R19569 avss.n7378 avss.n7377 1.93672
R19570 avss.n7380 avss.n7379 1.93672
R19571 avss.n7388 avss.n7268 1.93672
R19572 avss.n7401 avss.n7400 1.93672
R19573 avss.n7410 avss.n7409 1.93672
R19574 avss.n7233 avss.n7232 1.93672
R19575 avss.n7418 avss.n7234 1.93672
R19576 avss.n4081 avss.n4080 1.93672
R19577 avss.n7437 avss.n7436 1.93672
R19578 avss.n7456 avss.n4046 1.93672
R19579 avss.n7482 avss.n7481 1.93672
R19580 avss.n7502 avss.n7501 1.93672
R19581 avss.n7522 avss.n7520 1.93672
R19582 avss.n7532 avss.n7531 1.93672
R19583 avss.n4086 avss.n4082 1.93672
R19584 avss.n7507 avss.n7503 1.93672
R19585 avss.n7005 avss.n6978 1.93672
R19586 avss.n6969 avss.n6967 1.93672
R19587 avss.n7025 avss.n7024 1.93672
R19588 avss.n7027 avss.n7026 1.93672
R19589 avss.n7035 avss.n6915 1.93672
R19590 avss.n7048 avss.n7047 1.93672
R19591 avss.n7057 avss.n7056 1.93672
R19592 avss.n6880 avss.n6879 1.93672
R19593 avss.n7065 avss.n6881 1.93672
R19594 avss.n4165 avss.n4164 1.93672
R19595 avss.n7084 avss.n7083 1.93672
R19596 avss.n7103 avss.n4130 1.93672
R19597 avss.n7129 avss.n7128 1.93672
R19598 avss.n7149 avss.n7148 1.93672
R19599 avss.n7169 avss.n7167 1.93672
R19600 avss.n7179 avss.n7178 1.93672
R19601 avss.n4170 avss.n4166 1.93672
R19602 avss.n7154 avss.n7150 1.93672
R19603 avss.n6652 avss.n6625 1.93672
R19604 avss.n6616 avss.n6614 1.93672
R19605 avss.n6672 avss.n6671 1.93672
R19606 avss.n6674 avss.n6673 1.93672
R19607 avss.n6682 avss.n6562 1.93672
R19608 avss.n6695 avss.n6694 1.93672
R19609 avss.n6704 avss.n6703 1.93672
R19610 avss.n6527 avss.n6526 1.93672
R19611 avss.n6712 avss.n6528 1.93672
R19612 avss.n4249 avss.n4248 1.93672
R19613 avss.n6731 avss.n6730 1.93672
R19614 avss.n6750 avss.n4214 1.93672
R19615 avss.n6776 avss.n6775 1.93672
R19616 avss.n6796 avss.n6795 1.93672
R19617 avss.n6816 avss.n6814 1.93672
R19618 avss.n6826 avss.n6825 1.93672
R19619 avss.n4254 avss.n4250 1.93672
R19620 avss.n6801 avss.n6797 1.93672
R19621 avss.n6299 avss.n6272 1.93672
R19622 avss.n6263 avss.n6261 1.93672
R19623 avss.n6319 avss.n6318 1.93672
R19624 avss.n6321 avss.n6320 1.93672
R19625 avss.n6329 avss.n6209 1.93672
R19626 avss.n6342 avss.n6341 1.93672
R19627 avss.n6351 avss.n6350 1.93672
R19628 avss.n6174 avss.n6173 1.93672
R19629 avss.n6359 avss.n6175 1.93672
R19630 avss.n4333 avss.n4332 1.93672
R19631 avss.n6378 avss.n6377 1.93672
R19632 avss.n6397 avss.n4298 1.93672
R19633 avss.n6423 avss.n6422 1.93672
R19634 avss.n6443 avss.n6442 1.93672
R19635 avss.n6463 avss.n6461 1.93672
R19636 avss.n6473 avss.n6472 1.93672
R19637 avss.n4338 avss.n4334 1.93672
R19638 avss.n6448 avss.n6444 1.93672
R19639 avss.n5946 avss.n5919 1.93672
R19640 avss.n5910 avss.n5908 1.93672
R19641 avss.n5966 avss.n5965 1.93672
R19642 avss.n5968 avss.n5967 1.93672
R19643 avss.n5976 avss.n5856 1.93672
R19644 avss.n5989 avss.n5988 1.93672
R19645 avss.n5998 avss.n5997 1.93672
R19646 avss.n5821 avss.n5820 1.93672
R19647 avss.n6006 avss.n5822 1.93672
R19648 avss.n4417 avss.n4416 1.93672
R19649 avss.n6025 avss.n6024 1.93672
R19650 avss.n6044 avss.n4382 1.93672
R19651 avss.n6070 avss.n6069 1.93672
R19652 avss.n6090 avss.n6089 1.93672
R19653 avss.n6110 avss.n6108 1.93672
R19654 avss.n6120 avss.n6119 1.93672
R19655 avss.n4422 avss.n4418 1.93672
R19656 avss.n6095 avss.n6091 1.93672
R19657 avss.n5593 avss.n5566 1.93672
R19658 avss.n5557 avss.n5555 1.93672
R19659 avss.n5613 avss.n5612 1.93672
R19660 avss.n5615 avss.n5614 1.93672
R19661 avss.n5623 avss.n5503 1.93672
R19662 avss.n5636 avss.n5635 1.93672
R19663 avss.n5645 avss.n5644 1.93672
R19664 avss.n5468 avss.n5467 1.93672
R19665 avss.n5653 avss.n5469 1.93672
R19666 avss.n4501 avss.n4500 1.93672
R19667 avss.n5672 avss.n5671 1.93672
R19668 avss.n5691 avss.n4466 1.93672
R19669 avss.n5717 avss.n5716 1.93672
R19670 avss.n5737 avss.n5736 1.93672
R19671 avss.n5757 avss.n5755 1.93672
R19672 avss.n5767 avss.n5766 1.93672
R19673 avss.n4506 avss.n4502 1.93672
R19674 avss.n5742 avss.n5738 1.93672
R19675 avss.n5226 avss.n5209 1.93672
R19676 avss.n5217 avss.n5215 1.93672
R19677 avss.n5268 avss.n5267 1.93672
R19678 avss.n5270 avss.n5269 1.93672
R19679 avss.n5278 avss.n5157 1.93672
R19680 avss.n5291 avss.n5290 1.93672
R19681 avss.n5131 avss.n5096 1.93672
R19682 avss.n5123 avss.n5122 1.93672
R19683 avss.n5121 avss.n5120 1.93672
R19684 avss.n4585 avss.n4584 1.93672
R19685 avss.n5319 avss.n5318 1.93672
R19686 avss.n5338 avss.n4550 1.93672
R19687 avss.n5364 avss.n5363 1.93672
R19688 avss.n5384 avss.n5383 1.93672
R19689 avss.n5404 avss.n5402 1.93672
R19690 avss.n5414 avss.n5413 1.93672
R19691 avss.n4590 avss.n4586 1.93672
R19692 avss.n5389 avss.n5385 1.93672
R19693 avss.n4872 avss.n4855 1.93672
R19694 avss.n4863 avss.n4861 1.93672
R19695 avss.n4914 avss.n4913 1.93672
R19696 avss.n4916 avss.n4915 1.93672
R19697 avss.n4924 avss.n4803 1.93672
R19698 avss.n4937 avss.n4936 1.93672
R19699 avss.n4777 avss.n4742 1.93672
R19700 avss.n4769 avss.n4768 1.93672
R19701 avss.n4767 avss.n4766 1.93672
R19702 avss.n4669 avss.n4668 1.93672
R19703 avss.n4965 avss.n4964 1.93672
R19704 avss.n4984 avss.n4634 1.93672
R19705 avss.n5010 avss.n5009 1.93672
R19706 avss.n5030 avss.n5029 1.93672
R19707 avss.n5050 avss.n5048 1.93672
R19708 avss.n5060 avss.n5059 1.93672
R19709 avss.n4674 avss.n4670 1.93672
R19710 avss.n5035 avss.n5031 1.93672
R19711 avss.n9109 avss.n9108 1.93672
R19712 avss.n9163 avss.n9162 1.93672
R19713 avss.n9144 avss.n9143 1.93672
R19714 avss.n9129 avss.n9128 1.93672
R19715 avss.n2439 avss.n2438 1.93672
R19716 avss.n2452 avss.n2451 1.93672
R19717 avss.n2471 avss.n2470 1.93672
R19718 avss.n2418 avss.n2417 1.93672
R19719 avss.n2401 avss.n2400 1.93672
R19720 avss.n2565 avss.n2564 1.93672
R19721 avss.n2528 avss.n2527 1.93672
R19722 avss.n2509 avss.n2508 1.93672
R19723 avss.n2496 avss.n2495 1.93672
R19724 avss.n9018 avss.n9017 1.93672
R19725 avss.n9052 avss.n9051 1.93672
R19726 avss.n8997 avss.n8996 1.93672
R19727 avss.n2548 avss.n2547 1.93672
R19728 avss.n9033 avss.n9032 1.93672
R19729 avss.n9330 avss.n9329 1.93672
R19730 avss.n9384 avss.n9383 1.93672
R19731 avss.n9365 avss.n9364 1.93672
R19732 avss.n9350 avss.n9349 1.93672
R19733 avss.n2223 avss.n2222 1.93672
R19734 avss.n2236 avss.n2235 1.93672
R19735 avss.n2255 avss.n2254 1.93672
R19736 avss.n2202 avss.n2201 1.93672
R19737 avss.n2185 avss.n2184 1.93672
R19738 avss.n2349 avss.n2348 1.93672
R19739 avss.n2312 avss.n2311 1.93672
R19740 avss.n2293 avss.n2292 1.93672
R19741 avss.n2280 avss.n2279 1.93672
R19742 avss.n9239 avss.n9238 1.93672
R19743 avss.n9273 avss.n9272 1.93672
R19744 avss.n9218 avss.n9217 1.93672
R19745 avss.n2332 avss.n2331 1.93672
R19746 avss.n9254 avss.n9253 1.93672
R19747 avss.n9551 avss.n9550 1.93672
R19748 avss.n9605 avss.n9604 1.93672
R19749 avss.n9586 avss.n9585 1.93672
R19750 avss.n9571 avss.n9570 1.93672
R19751 avss.n2007 avss.n2006 1.93672
R19752 avss.n2020 avss.n2019 1.93672
R19753 avss.n2039 avss.n2038 1.93672
R19754 avss.n1986 avss.n1985 1.93672
R19755 avss.n1969 avss.n1968 1.93672
R19756 avss.n2133 avss.n2132 1.93672
R19757 avss.n2096 avss.n2095 1.93672
R19758 avss.n2077 avss.n2076 1.93672
R19759 avss.n2064 avss.n2063 1.93672
R19760 avss.n9460 avss.n9459 1.93672
R19761 avss.n9494 avss.n9493 1.93672
R19762 avss.n9439 avss.n9438 1.93672
R19763 avss.n2116 avss.n2115 1.93672
R19764 avss.n9475 avss.n9474 1.93672
R19765 avss.n9772 avss.n9771 1.93672
R19766 avss.n9826 avss.n9825 1.93672
R19767 avss.n9807 avss.n9806 1.93672
R19768 avss.n9792 avss.n9791 1.93672
R19769 avss.n1791 avss.n1790 1.93672
R19770 avss.n1804 avss.n1803 1.93672
R19771 avss.n1823 avss.n1822 1.93672
R19772 avss.n1770 avss.n1769 1.93672
R19773 avss.n1753 avss.n1752 1.93672
R19774 avss.n1917 avss.n1916 1.93672
R19775 avss.n1880 avss.n1879 1.93672
R19776 avss.n1861 avss.n1860 1.93672
R19777 avss.n1848 avss.n1847 1.93672
R19778 avss.n9681 avss.n9680 1.93672
R19779 avss.n9715 avss.n9714 1.93672
R19780 avss.n9660 avss.n9659 1.93672
R19781 avss.n1900 avss.n1899 1.93672
R19782 avss.n9696 avss.n9695 1.93672
R19783 avss.n9993 avss.n9992 1.93672
R19784 avss.n10047 avss.n10046 1.93672
R19785 avss.n10028 avss.n10027 1.93672
R19786 avss.n10013 avss.n10012 1.93672
R19787 avss.n1575 avss.n1574 1.93672
R19788 avss.n1588 avss.n1587 1.93672
R19789 avss.n1607 avss.n1606 1.93672
R19790 avss.n1554 avss.n1553 1.93672
R19791 avss.n1537 avss.n1536 1.93672
R19792 avss.n1701 avss.n1700 1.93672
R19793 avss.n1664 avss.n1663 1.93672
R19794 avss.n1645 avss.n1644 1.93672
R19795 avss.n1632 avss.n1631 1.93672
R19796 avss.n9902 avss.n9901 1.93672
R19797 avss.n9936 avss.n9935 1.93672
R19798 avss.n9881 avss.n9880 1.93672
R19799 avss.n1684 avss.n1683 1.93672
R19800 avss.n9917 avss.n9916 1.93672
R19801 avss.n10214 avss.n10213 1.93672
R19802 avss.n10268 avss.n10267 1.93672
R19803 avss.n10249 avss.n10248 1.93672
R19804 avss.n10234 avss.n10233 1.93672
R19805 avss.n1359 avss.n1358 1.93672
R19806 avss.n1372 avss.n1371 1.93672
R19807 avss.n1391 avss.n1390 1.93672
R19808 avss.n1338 avss.n1337 1.93672
R19809 avss.n1321 avss.n1320 1.93672
R19810 avss.n1485 avss.n1484 1.93672
R19811 avss.n1448 avss.n1447 1.93672
R19812 avss.n1429 avss.n1428 1.93672
R19813 avss.n1416 avss.n1415 1.93672
R19814 avss.n10123 avss.n10122 1.93672
R19815 avss.n10157 avss.n10156 1.93672
R19816 avss.n10102 avss.n10101 1.93672
R19817 avss.n1468 avss.n1467 1.93672
R19818 avss.n10138 avss.n10137 1.93672
R19819 avss.n10435 avss.n10434 1.93672
R19820 avss.n10489 avss.n10488 1.93672
R19821 avss.n10470 avss.n10469 1.93672
R19822 avss.n10455 avss.n10454 1.93672
R19823 avss.n1143 avss.n1142 1.93672
R19824 avss.n1156 avss.n1155 1.93672
R19825 avss.n1175 avss.n1174 1.93672
R19826 avss.n1122 avss.n1121 1.93672
R19827 avss.n1105 avss.n1104 1.93672
R19828 avss.n1269 avss.n1268 1.93672
R19829 avss.n1232 avss.n1231 1.93672
R19830 avss.n1213 avss.n1212 1.93672
R19831 avss.n1200 avss.n1199 1.93672
R19832 avss.n10344 avss.n10343 1.93672
R19833 avss.n10378 avss.n10377 1.93672
R19834 avss.n10323 avss.n10322 1.93672
R19835 avss.n1252 avss.n1251 1.93672
R19836 avss.n10359 avss.n10358 1.93672
R19837 avss.n10656 avss.n10655 1.93672
R19838 avss.n10710 avss.n10709 1.93672
R19839 avss.n10691 avss.n10690 1.93672
R19840 avss.n10676 avss.n10675 1.93672
R19841 avss.n927 avss.n926 1.93672
R19842 avss.n940 avss.n939 1.93672
R19843 avss.n959 avss.n958 1.93672
R19844 avss.n906 avss.n905 1.93672
R19845 avss.n889 avss.n888 1.93672
R19846 avss.n1053 avss.n1052 1.93672
R19847 avss.n1016 avss.n1015 1.93672
R19848 avss.n997 avss.n996 1.93672
R19849 avss.n984 avss.n983 1.93672
R19850 avss.n10565 avss.n10564 1.93672
R19851 avss.n10599 avss.n10598 1.93672
R19852 avss.n10544 avss.n10543 1.93672
R19853 avss.n1036 avss.n1035 1.93672
R19854 avss.n10580 avss.n10579 1.93672
R19855 avss.n10877 avss.n10876 1.93672
R19856 avss.n10931 avss.n10930 1.93672
R19857 avss.n10912 avss.n10911 1.93672
R19858 avss.n10897 avss.n10896 1.93672
R19859 avss.n711 avss.n710 1.93672
R19860 avss.n724 avss.n723 1.93672
R19861 avss.n743 avss.n742 1.93672
R19862 avss.n690 avss.n689 1.93672
R19863 avss.n673 avss.n672 1.93672
R19864 avss.n837 avss.n836 1.93672
R19865 avss.n800 avss.n799 1.93672
R19866 avss.n781 avss.n780 1.93672
R19867 avss.n768 avss.n767 1.93672
R19868 avss.n10786 avss.n10785 1.93672
R19869 avss.n10820 avss.n10819 1.93672
R19870 avss.n10765 avss.n10764 1.93672
R19871 avss.n820 avss.n819 1.93672
R19872 avss.n10801 avss.n10800 1.93672
R19873 avss.n11098 avss.n11097 1.93672
R19874 avss.n11152 avss.n11151 1.93672
R19875 avss.n11133 avss.n11132 1.93672
R19876 avss.n11118 avss.n11117 1.93672
R19877 avss.n495 avss.n494 1.93672
R19878 avss.n508 avss.n507 1.93672
R19879 avss.n527 avss.n526 1.93672
R19880 avss.n474 avss.n473 1.93672
R19881 avss.n457 avss.n456 1.93672
R19882 avss.n621 avss.n620 1.93672
R19883 avss.n584 avss.n583 1.93672
R19884 avss.n565 avss.n564 1.93672
R19885 avss.n552 avss.n551 1.93672
R19886 avss.n11007 avss.n11006 1.93672
R19887 avss.n11041 avss.n11040 1.93672
R19888 avss.n10986 avss.n10985 1.93672
R19889 avss.n604 avss.n603 1.93672
R19890 avss.n11022 avss.n11021 1.93672
R19891 avss.n364 avss.n363 1.93672
R19892 avss.n419 avss.n418 1.93672
R19893 avss.n400 avss.n399 1.93672
R19894 avss.n385 avss.n384 1.93672
R19895 avss.n11324 avss.n11323 1.93672
R19896 avss.n11337 avss.n11336 1.93672
R19897 avss.n11356 avss.n11355 1.93672
R19898 avss.n11375 avss.n11374 1.93672
R19899 avss.n11393 avss.n11392 1.93672
R19900 avss.n296 avss.n295 1.93672
R19901 avss.n259 avss.n258 1.93672
R19902 avss.n240 avss.n239 1.93672
R19903 avss.n227 avss.n226 1.93672
R19904 avss.n11228 avss.n11227 1.93672
R19905 avss.n11262 avss.n11261 1.93672
R19906 avss.n11207 avss.n11206 1.93672
R19907 avss.n279 avss.n278 1.93672
R19908 avss.n11243 avss.n11242 1.93672
R19909 avss.n147 avss.n146 1.93672
R19910 avss.n202 avss.n201 1.93672
R19911 avss.n183 avss.n182 1.93672
R19912 avss.n168 avss.n167 1.93672
R19913 avss.n11545 avss.n11544 1.93672
R19914 avss.n11558 avss.n11557 1.93672
R19915 avss.n11577 avss.n11576 1.93672
R19916 avss.n11596 avss.n11595 1.93672
R19917 avss.n11614 avss.n11613 1.93672
R19918 avss.n79 avss.n78 1.93672
R19919 avss.n42 avss.n41 1.93672
R19920 avss.n23 avss.n22 1.93672
R19921 avss.n10 avss.n9 1.93672
R19922 avss.n11449 avss.n11448 1.93672
R19923 avss.n11483 avss.n11482 1.93672
R19924 avss.n11428 avss.n11427 1.93672
R19925 avss.n62 avss.n61 1.93672
R19926 avss.n11464 avss.n11463 1.93672
R19927 avss.n8789 avss.n8788 1.7055
R19928 avss.n8756 avss.n8750 1.7055
R19929 avss.n8667 avss.n8666 1.7055
R19930 avss.n8807 avss.n8806 1.7055
R19931 avss.n8805 avss.n8669 1.7055
R19932 avss.n8695 avss.n8685 1.7055
R19933 avss.n8712 avss.n8708 1.7055
R19934 avss.n8777 avss.n8720 1.7055
R19935 avss.n8745 avss.n8722 1.7055
R19936 avss.n8752 avss.n8749 1.7055
R19937 avss.n8831 avss.n8830 1.7055
R19938 avss.n8860 avss.n8856 1.7055
R19939 avss.n8877 avss.n8876 1.7055
R19940 avss.n8878 avss.n3703 1.7055
R19941 avss.n8889 avss.n3702 1.7055
R19942 avss.n8908 avss.n8907 1.7055
R19943 avss.n8924 avss.n8922 1.7055
R19944 avss.n8967 avss.n8966 1.7055
R19945 avss.n8965 avss.n3679 1.7055
R19946 avss.n8920 avss.n8919 1.7055
R19947 avss.n8957 avss.n8956 1.7055
R19948 avss.n3751 avss.n3750 1.7055
R19949 avss.n8436 avss.n8435 1.7055
R19950 avss.n8403 avss.n8397 1.7055
R19951 avss.n8314 avss.n8313 1.7055
R19952 avss.n8454 avss.n8453 1.7055
R19953 avss.n8452 avss.n8316 1.7055
R19954 avss.n8342 avss.n8332 1.7055
R19955 avss.n8359 avss.n8355 1.7055
R19956 avss.n8424 avss.n8367 1.7055
R19957 avss.n8392 avss.n8369 1.7055
R19958 avss.n8399 avss.n8396 1.7055
R19959 avss.n8478 avss.n8477 1.7055
R19960 avss.n8507 avss.n8503 1.7055
R19961 avss.n8524 avss.n8523 1.7055
R19962 avss.n8525 avss.n3787 1.7055
R19963 avss.n8536 avss.n3786 1.7055
R19964 avss.n8555 avss.n8554 1.7055
R19965 avss.n8571 avss.n8569 1.7055
R19966 avss.n8614 avss.n8613 1.7055
R19967 avss.n8612 avss.n3763 1.7055
R19968 avss.n8567 avss.n8566 1.7055
R19969 avss.n8604 avss.n8603 1.7055
R19970 avss.n3835 avss.n3834 1.7055
R19971 avss.n8083 avss.n8082 1.7055
R19972 avss.n8050 avss.n8044 1.7055
R19973 avss.n7961 avss.n7960 1.7055
R19974 avss.n8101 avss.n8100 1.7055
R19975 avss.n8099 avss.n7963 1.7055
R19976 avss.n7989 avss.n7979 1.7055
R19977 avss.n8006 avss.n8002 1.7055
R19978 avss.n8071 avss.n8014 1.7055
R19979 avss.n8039 avss.n8016 1.7055
R19980 avss.n8046 avss.n8043 1.7055
R19981 avss.n8125 avss.n8124 1.7055
R19982 avss.n8154 avss.n8150 1.7055
R19983 avss.n8171 avss.n8170 1.7055
R19984 avss.n8172 avss.n3871 1.7055
R19985 avss.n8183 avss.n3870 1.7055
R19986 avss.n8202 avss.n8201 1.7055
R19987 avss.n8218 avss.n8216 1.7055
R19988 avss.n8261 avss.n8260 1.7055
R19989 avss.n8259 avss.n3847 1.7055
R19990 avss.n8214 avss.n8213 1.7055
R19991 avss.n8251 avss.n8250 1.7055
R19992 avss.n3919 avss.n3918 1.7055
R19993 avss.n7730 avss.n7729 1.7055
R19994 avss.n7697 avss.n7691 1.7055
R19995 avss.n7608 avss.n7607 1.7055
R19996 avss.n7748 avss.n7747 1.7055
R19997 avss.n7746 avss.n7610 1.7055
R19998 avss.n7636 avss.n7626 1.7055
R19999 avss.n7653 avss.n7649 1.7055
R20000 avss.n7718 avss.n7661 1.7055
R20001 avss.n7686 avss.n7663 1.7055
R20002 avss.n7693 avss.n7690 1.7055
R20003 avss.n7772 avss.n7771 1.7055
R20004 avss.n7801 avss.n7797 1.7055
R20005 avss.n7818 avss.n7817 1.7055
R20006 avss.n7819 avss.n3955 1.7055
R20007 avss.n7830 avss.n3954 1.7055
R20008 avss.n7849 avss.n7848 1.7055
R20009 avss.n7865 avss.n7863 1.7055
R20010 avss.n7908 avss.n7907 1.7055
R20011 avss.n7906 avss.n3931 1.7055
R20012 avss.n7861 avss.n7860 1.7055
R20013 avss.n7898 avss.n7897 1.7055
R20014 avss.n4003 avss.n4002 1.7055
R20015 avss.n7377 avss.n7376 1.7055
R20016 avss.n7344 avss.n7338 1.7055
R20017 avss.n7255 avss.n7254 1.7055
R20018 avss.n7395 avss.n7394 1.7055
R20019 avss.n7393 avss.n7257 1.7055
R20020 avss.n7283 avss.n7273 1.7055
R20021 avss.n7300 avss.n7296 1.7055
R20022 avss.n7365 avss.n7308 1.7055
R20023 avss.n7333 avss.n7310 1.7055
R20024 avss.n7340 avss.n7337 1.7055
R20025 avss.n7419 avss.n7418 1.7055
R20026 avss.n7448 avss.n7444 1.7055
R20027 avss.n7465 avss.n7464 1.7055
R20028 avss.n7466 avss.n4039 1.7055
R20029 avss.n7477 avss.n4038 1.7055
R20030 avss.n7496 avss.n7495 1.7055
R20031 avss.n7512 avss.n7510 1.7055
R20032 avss.n7555 avss.n7554 1.7055
R20033 avss.n7553 avss.n4015 1.7055
R20034 avss.n7508 avss.n7507 1.7055
R20035 avss.n7545 avss.n7544 1.7055
R20036 avss.n4087 avss.n4086 1.7055
R20037 avss.n7024 avss.n7023 1.7055
R20038 avss.n6991 avss.n6985 1.7055
R20039 avss.n6902 avss.n6901 1.7055
R20040 avss.n7042 avss.n7041 1.7055
R20041 avss.n7040 avss.n6904 1.7055
R20042 avss.n6930 avss.n6920 1.7055
R20043 avss.n6947 avss.n6943 1.7055
R20044 avss.n7012 avss.n6955 1.7055
R20045 avss.n6980 avss.n6957 1.7055
R20046 avss.n6987 avss.n6984 1.7055
R20047 avss.n7066 avss.n7065 1.7055
R20048 avss.n7095 avss.n7091 1.7055
R20049 avss.n7112 avss.n7111 1.7055
R20050 avss.n7113 avss.n4123 1.7055
R20051 avss.n7124 avss.n4122 1.7055
R20052 avss.n7143 avss.n7142 1.7055
R20053 avss.n7159 avss.n7157 1.7055
R20054 avss.n7202 avss.n7201 1.7055
R20055 avss.n7200 avss.n4099 1.7055
R20056 avss.n7155 avss.n7154 1.7055
R20057 avss.n7192 avss.n7191 1.7055
R20058 avss.n4171 avss.n4170 1.7055
R20059 avss.n6671 avss.n6670 1.7055
R20060 avss.n6638 avss.n6632 1.7055
R20061 avss.n6549 avss.n6548 1.7055
R20062 avss.n6689 avss.n6688 1.7055
R20063 avss.n6687 avss.n6551 1.7055
R20064 avss.n6577 avss.n6567 1.7055
R20065 avss.n6594 avss.n6590 1.7055
R20066 avss.n6659 avss.n6602 1.7055
R20067 avss.n6627 avss.n6604 1.7055
R20068 avss.n6634 avss.n6631 1.7055
R20069 avss.n6713 avss.n6712 1.7055
R20070 avss.n6742 avss.n6738 1.7055
R20071 avss.n6759 avss.n6758 1.7055
R20072 avss.n6760 avss.n4207 1.7055
R20073 avss.n6771 avss.n4206 1.7055
R20074 avss.n6790 avss.n6789 1.7055
R20075 avss.n6806 avss.n6804 1.7055
R20076 avss.n6849 avss.n6848 1.7055
R20077 avss.n6847 avss.n4183 1.7055
R20078 avss.n6802 avss.n6801 1.7055
R20079 avss.n6839 avss.n6838 1.7055
R20080 avss.n4255 avss.n4254 1.7055
R20081 avss.n6318 avss.n6317 1.7055
R20082 avss.n6285 avss.n6279 1.7055
R20083 avss.n6196 avss.n6195 1.7055
R20084 avss.n6336 avss.n6335 1.7055
R20085 avss.n6334 avss.n6198 1.7055
R20086 avss.n6224 avss.n6214 1.7055
R20087 avss.n6241 avss.n6237 1.7055
R20088 avss.n6306 avss.n6249 1.7055
R20089 avss.n6274 avss.n6251 1.7055
R20090 avss.n6281 avss.n6278 1.7055
R20091 avss.n6360 avss.n6359 1.7055
R20092 avss.n6389 avss.n6385 1.7055
R20093 avss.n6406 avss.n6405 1.7055
R20094 avss.n6407 avss.n4291 1.7055
R20095 avss.n6418 avss.n4290 1.7055
R20096 avss.n6437 avss.n6436 1.7055
R20097 avss.n6453 avss.n6451 1.7055
R20098 avss.n6496 avss.n6495 1.7055
R20099 avss.n6494 avss.n4267 1.7055
R20100 avss.n6449 avss.n6448 1.7055
R20101 avss.n6486 avss.n6485 1.7055
R20102 avss.n4339 avss.n4338 1.7055
R20103 avss.n5965 avss.n5964 1.7055
R20104 avss.n5932 avss.n5926 1.7055
R20105 avss.n5843 avss.n5842 1.7055
R20106 avss.n5983 avss.n5982 1.7055
R20107 avss.n5981 avss.n5845 1.7055
R20108 avss.n5871 avss.n5861 1.7055
R20109 avss.n5888 avss.n5884 1.7055
R20110 avss.n5953 avss.n5896 1.7055
R20111 avss.n5921 avss.n5898 1.7055
R20112 avss.n5928 avss.n5925 1.7055
R20113 avss.n6007 avss.n6006 1.7055
R20114 avss.n6036 avss.n6032 1.7055
R20115 avss.n6053 avss.n6052 1.7055
R20116 avss.n6054 avss.n4375 1.7055
R20117 avss.n6065 avss.n4374 1.7055
R20118 avss.n6084 avss.n6083 1.7055
R20119 avss.n6100 avss.n6098 1.7055
R20120 avss.n6143 avss.n6142 1.7055
R20121 avss.n6141 avss.n4351 1.7055
R20122 avss.n6096 avss.n6095 1.7055
R20123 avss.n6133 avss.n6132 1.7055
R20124 avss.n4423 avss.n4422 1.7055
R20125 avss.n5612 avss.n5611 1.7055
R20126 avss.n5579 avss.n5573 1.7055
R20127 avss.n5490 avss.n5489 1.7055
R20128 avss.n5630 avss.n5629 1.7055
R20129 avss.n5628 avss.n5492 1.7055
R20130 avss.n5518 avss.n5508 1.7055
R20131 avss.n5535 avss.n5531 1.7055
R20132 avss.n5600 avss.n5543 1.7055
R20133 avss.n5568 avss.n5545 1.7055
R20134 avss.n5575 avss.n5572 1.7055
R20135 avss.n5654 avss.n5653 1.7055
R20136 avss.n5683 avss.n5679 1.7055
R20137 avss.n5700 avss.n5699 1.7055
R20138 avss.n5701 avss.n4459 1.7055
R20139 avss.n5712 avss.n4458 1.7055
R20140 avss.n5731 avss.n5730 1.7055
R20141 avss.n5747 avss.n5745 1.7055
R20142 avss.n5790 avss.n5789 1.7055
R20143 avss.n5788 avss.n4435 1.7055
R20144 avss.n5743 avss.n5742 1.7055
R20145 avss.n5780 avss.n5779 1.7055
R20146 avss.n4507 avss.n4506 1.7055
R20147 avss.n5230 avss.n5199 1.7055
R20148 avss.n5123 avss.n5102 1.7055
R20149 avss.n5267 avss.n5266 1.7055
R20150 avss.n5238 avss.n5232 1.7055
R20151 avss.n5144 avss.n5143 1.7055
R20152 avss.n5285 avss.n5284 1.7055
R20153 avss.n5283 avss.n5146 1.7055
R20154 avss.n5172 avss.n5162 1.7055
R20155 avss.n5189 avss.n5185 1.7055
R20156 avss.n5255 avss.n5197 1.7055
R20157 avss.n5234 avss.n5231 1.7055
R20158 avss.n5330 avss.n5326 1.7055
R20159 avss.n5347 avss.n5346 1.7055
R20160 avss.n5348 avss.n4543 1.7055
R20161 avss.n5359 avss.n4542 1.7055
R20162 avss.n5378 avss.n5377 1.7055
R20163 avss.n5394 avss.n5392 1.7055
R20164 avss.n5437 avss.n5436 1.7055
R20165 avss.n5435 avss.n4519 1.7055
R20166 avss.n5390 avss.n5389 1.7055
R20167 avss.n5427 avss.n5426 1.7055
R20168 avss.n4591 avss.n4590 1.7055
R20169 avss.n4876 avss.n4845 1.7055
R20170 avss.n4769 avss.n4748 1.7055
R20171 avss.n4913 avss.n4912 1.7055
R20172 avss.n4884 avss.n4878 1.7055
R20173 avss.n4790 avss.n4789 1.7055
R20174 avss.n4931 avss.n4930 1.7055
R20175 avss.n4929 avss.n4792 1.7055
R20176 avss.n4818 avss.n4808 1.7055
R20177 avss.n4835 avss.n4831 1.7055
R20178 avss.n4901 avss.n4843 1.7055
R20179 avss.n4880 avss.n4877 1.7055
R20180 avss.n4976 avss.n4972 1.7055
R20181 avss.n4993 avss.n4992 1.7055
R20182 avss.n4994 avss.n4627 1.7055
R20183 avss.n5005 avss.n4626 1.7055
R20184 avss.n5024 avss.n5023 1.7055
R20185 avss.n5040 avss.n5038 1.7055
R20186 avss.n5083 avss.n5082 1.7055
R20187 avss.n5081 avss.n4603 1.7055
R20188 avss.n5036 avss.n5035 1.7055
R20189 avss.n5073 avss.n5072 1.7055
R20190 avss.n4675 avss.n4674 1.7055
R20191 avss.n9096 avss.n9095 1.7055
R20192 avss.n9076 avss.n9075 1.7055
R20193 avss.n9317 avss.n9316 1.7055
R20194 avss.n9297 avss.n9296 1.7055
R20195 avss.n9538 avss.n9537 1.7055
R20196 avss.n9518 avss.n9517 1.7055
R20197 avss.n9759 avss.n9758 1.7055
R20198 avss.n9739 avss.n9738 1.7055
R20199 avss.n9980 avss.n9979 1.7055
R20200 avss.n9960 avss.n9959 1.7055
R20201 avss.n10201 avss.n10200 1.7055
R20202 avss.n10181 avss.n10180 1.7055
R20203 avss.n10422 avss.n10421 1.7055
R20204 avss.n10402 avss.n10401 1.7055
R20205 avss.n10643 avss.n10642 1.7055
R20206 avss.n10623 avss.n10622 1.7055
R20207 avss.n10864 avss.n10863 1.7055
R20208 avss.n10844 avss.n10843 1.7055
R20209 avss.n11085 avss.n11084 1.7055
R20210 avss.n11065 avss.n11064 1.7055
R20211 avss.n336 avss.n335 1.7055
R20212 avss.n11286 avss.n11285 1.7055
R20213 avss.n119 avss.n118 1.7055
R20214 avss.n11507 avss.n11506 1.7055
R20215 avss.n8969 avss.n8968 1.70511
R20216 avss.n8616 avss.n8615 1.70511
R20217 avss.n8263 avss.n8262 1.70511
R20218 avss.n7910 avss.n7909 1.70511
R20219 avss.n7557 avss.n7556 1.70511
R20220 avss.n7204 avss.n7203 1.70511
R20221 avss.n6851 avss.n6850 1.70511
R20222 avss.n6498 avss.n6497 1.70511
R20223 avss.n6145 avss.n6144 1.70511
R20224 avss.n5792 avss.n5791 1.70511
R20225 avss.n5252 avss.n5251 1.70511
R20226 avss.n5439 avss.n5438 1.70511
R20227 avss.n4898 avss.n4897 1.70511
R20228 avss.n5085 avss.n5084 1.70511
R20229 avss.n8772 avss.n8723 1.70483
R20230 avss.n8627 avss.n8620 1.70483
R20231 avss.n3677 avss.n3669 1.70483
R20232 avss.n8419 avss.n8370 1.70483
R20233 avss.n8274 avss.n8267 1.70483
R20234 avss.n3761 avss.n3753 1.70483
R20235 avss.n8066 avss.n8017 1.70483
R20236 avss.n7921 avss.n7914 1.70483
R20237 avss.n3845 avss.n3837 1.70483
R20238 avss.n7713 avss.n7664 1.70483
R20239 avss.n7568 avss.n7561 1.70483
R20240 avss.n3929 avss.n3921 1.70483
R20241 avss.n7360 avss.n7311 1.70483
R20242 avss.n7215 avss.n7208 1.70483
R20243 avss.n4013 avss.n4005 1.70483
R20244 avss.n7007 avss.n6958 1.70483
R20245 avss.n6862 avss.n6855 1.70483
R20246 avss.n4097 avss.n4089 1.70483
R20247 avss.n6654 avss.n6605 1.70483
R20248 avss.n6509 avss.n6502 1.70483
R20249 avss.n4181 avss.n4173 1.70483
R20250 avss.n6301 avss.n6252 1.70483
R20251 avss.n6156 avss.n6149 1.70483
R20252 avss.n4265 avss.n4257 1.70483
R20253 avss.n5948 avss.n5899 1.70483
R20254 avss.n5803 avss.n5796 1.70483
R20255 avss.n4349 avss.n4341 1.70483
R20256 avss.n5595 avss.n5546 1.70483
R20257 avss.n5450 avss.n5443 1.70483
R20258 avss.n4433 avss.n4425 1.70483
R20259 avss.n5304 avss.n5303 1.70483
R20260 avss.n4517 avss.n4509 1.70483
R20261 avss.n4950 avss.n4949 1.70483
R20262 avss.n4601 avss.n4593 1.70483
R20263 avss.n5101 avss.n5089 1.70227
R20264 avss.n4747 avss.n4735 1.70227
R20265 avss.n8844 avss.n8843 1.70192
R20266 avss.n8491 avss.n8490 1.70192
R20267 avss.n8138 avss.n8137 1.70192
R20268 avss.n7785 avss.n7784 1.70192
R20269 avss.n7432 avss.n7431 1.70192
R20270 avss.n7079 avss.n7078 1.70192
R20271 avss.n6726 avss.n6725 1.70192
R20272 avss.n6373 avss.n6372 1.70192
R20273 avss.n6020 avss.n6019 1.70192
R20274 avss.n5667 avss.n5666 1.70192
R20275 avss.n5314 avss.n5313 1.70192
R20276 avss.n4960 avss.n4959 1.70192
R20277 avss.n8774 avss.n8725 1.7005
R20278 avss.n8421 avss.n8372 1.7005
R20279 avss.n8068 avss.n8019 1.7005
R20280 avss.n7715 avss.n7666 1.7005
R20281 avss.n7362 avss.n7313 1.7005
R20282 avss.n7009 avss.n6960 1.7005
R20283 avss.n6656 avss.n6607 1.7005
R20284 avss.n6303 avss.n6254 1.7005
R20285 avss.n5950 avss.n5901 1.7005
R20286 avss.n5597 avss.n5548 1.7005
R20287 avss.n5252 avss.n5205 1.7005
R20288 avss.n4898 avss.n4851 1.7005
R20289 avss.n3511 avss.n3176 1.61892
R20290 avss.n11632 avss.n11631 1.53719
R20291 avss.n8974 avss 1.52724
R20292 avss.n3389 avss.n3270 1.50638
R20293 avss.n3403 avss.n3243 1.50638
R20294 avss.n3411 avss.n3225 1.50638
R20295 avss.n3226 avss.n3222 1.50638
R20296 avss.n3474 avss.n3473 1.50638
R20297 avss.n3194 avss.n3171 1.50638
R20298 avss.n3250 avss.n2619 1.44882
R20299 avss.n3516 avss.n3168 1.18753
R20300 avss.n2980 avss.n2957 1.18311
R20301 avss.n3037 avss.n2941 1.18311
R20302 avss.n3079 avss.n3078 1.18311
R20303 avss.n3629 avss.n2607 1.18311
R20304 avss.n2692 avss.n2670 1.18311
R20305 avss.n2737 avss.n2643 1.18311
R20306 avss.n2777 avss.n2776 1.18311
R20307 avss.n2813 avss.n2812 1.18311
R20308 avss.n9084 avss.n8974 1.15733
R20309 avss.n3014 avss.n3013 1.14023
R20310 avss.n3072 avss.n3071 1.14023
R20311 avss.n3100 avss.n3093 1.14023
R20312 avss.n3663 avss.n3662 1.14023
R20313 avss.n2726 avss.n2725 1.14023
R20314 avss.n2771 avss.n2770 1.14023
R20315 avss.n2874 avss.n2791 1.14023
R20316 avss.n2834 avss.n2827 1.14023
R20317 avss.n8652 avss.n8650 1.13717
R20318 avss.n8774 avss.n8721 1.13717
R20319 avss.n8829 avss.n8628 1.13717
R20320 avss.n8656 avss.n8651 1.13717
R20321 avss.n8673 avss.n8672 1.13717
R20322 avss.n8688 avss.n8679 1.13717
R20323 avss.n8704 avss.n8700 1.13717
R20324 avss.n8787 avss.n8706 1.13717
R20325 avss.n8736 avss.n8731 1.13717
R20326 avss.n8768 avss.n8767 1.13717
R20327 avss.n8635 avss.n8634 1.13717
R20328 avss.n8642 avss.n8641 1.13717
R20329 avss.n8655 avss.n8653 1.13717
R20330 avss.n8810 avss.n8809 1.13717
R20331 avss.n8692 avss.n8691 1.13717
R20332 avss.n8698 avss.n8683 1.13717
R20333 avss.n8709 avss.n8699 1.13717
R20334 avss.n8715 avss.n8707 1.13717
R20335 avss.n8780 avss.n8719 1.13717
R20336 avss.n8968 avss.n3674 1.13717
R20337 avss.n3735 avss.n3734 1.13717
R20338 avss.n3742 avss.n3741 1.13717
R20339 avss.n3749 avss.n3728 1.13717
R20340 avss.n8852 avss.n3719 1.13717
R20341 avss.n8863 avss.n3716 1.13717
R20342 avss.n8840 avss.n3717 1.13717
R20343 avss.n8872 avss.n3709 1.13717
R20344 avss.n3708 avss.n3707 1.13717
R20345 avss.n8883 avss.n8882 1.13717
R20346 avss.n8886 avss.n3701 1.13717
R20347 avss.n8897 avss.n8896 1.13717
R20348 avss.n8911 avss.n8910 1.13717
R20349 avss.n3697 avss.n3696 1.13717
R20350 avss.n8918 avss.n3691 1.13717
R20351 avss.n8927 avss.n3688 1.13717
R20352 avss.n3690 avss.n3689 1.13717
R20353 avss.n8937 avss.n8936 1.13717
R20354 avss.n8947 avss.n8946 1.13717
R20355 avss.n8299 avss.n8297 1.13717
R20356 avss.n8421 avss.n8368 1.13717
R20357 avss.n8476 avss.n8275 1.13717
R20358 avss.n8303 avss.n8298 1.13717
R20359 avss.n8320 avss.n8319 1.13717
R20360 avss.n8335 avss.n8326 1.13717
R20361 avss.n8351 avss.n8347 1.13717
R20362 avss.n8434 avss.n8353 1.13717
R20363 avss.n8383 avss.n8378 1.13717
R20364 avss.n8415 avss.n8414 1.13717
R20365 avss.n8282 avss.n8281 1.13717
R20366 avss.n8289 avss.n8288 1.13717
R20367 avss.n8302 avss.n8300 1.13717
R20368 avss.n8457 avss.n8456 1.13717
R20369 avss.n8339 avss.n8338 1.13717
R20370 avss.n8345 avss.n8330 1.13717
R20371 avss.n8356 avss.n8346 1.13717
R20372 avss.n8362 avss.n8354 1.13717
R20373 avss.n8427 avss.n8366 1.13717
R20374 avss.n8615 avss.n3758 1.13717
R20375 avss.n3819 avss.n3818 1.13717
R20376 avss.n3826 avss.n3825 1.13717
R20377 avss.n3833 avss.n3812 1.13717
R20378 avss.n8499 avss.n3803 1.13717
R20379 avss.n8510 avss.n3800 1.13717
R20380 avss.n8487 avss.n3801 1.13717
R20381 avss.n8519 avss.n3793 1.13717
R20382 avss.n3792 avss.n3791 1.13717
R20383 avss.n8530 avss.n8529 1.13717
R20384 avss.n8533 avss.n3785 1.13717
R20385 avss.n8544 avss.n8543 1.13717
R20386 avss.n8558 avss.n8557 1.13717
R20387 avss.n3781 avss.n3780 1.13717
R20388 avss.n8565 avss.n3775 1.13717
R20389 avss.n8574 avss.n3772 1.13717
R20390 avss.n3774 avss.n3773 1.13717
R20391 avss.n8584 avss.n8583 1.13717
R20392 avss.n8594 avss.n8593 1.13717
R20393 avss.n7946 avss.n7944 1.13717
R20394 avss.n8068 avss.n8015 1.13717
R20395 avss.n8123 avss.n7922 1.13717
R20396 avss.n7950 avss.n7945 1.13717
R20397 avss.n7967 avss.n7966 1.13717
R20398 avss.n7982 avss.n7973 1.13717
R20399 avss.n7998 avss.n7994 1.13717
R20400 avss.n8081 avss.n8000 1.13717
R20401 avss.n8030 avss.n8025 1.13717
R20402 avss.n8062 avss.n8061 1.13717
R20403 avss.n7929 avss.n7928 1.13717
R20404 avss.n7936 avss.n7935 1.13717
R20405 avss.n7949 avss.n7947 1.13717
R20406 avss.n8104 avss.n8103 1.13717
R20407 avss.n7986 avss.n7985 1.13717
R20408 avss.n7992 avss.n7977 1.13717
R20409 avss.n8003 avss.n7993 1.13717
R20410 avss.n8009 avss.n8001 1.13717
R20411 avss.n8074 avss.n8013 1.13717
R20412 avss.n8262 avss.n3842 1.13717
R20413 avss.n3903 avss.n3902 1.13717
R20414 avss.n3910 avss.n3909 1.13717
R20415 avss.n3917 avss.n3896 1.13717
R20416 avss.n8146 avss.n3887 1.13717
R20417 avss.n8157 avss.n3884 1.13717
R20418 avss.n8134 avss.n3885 1.13717
R20419 avss.n8166 avss.n3877 1.13717
R20420 avss.n3876 avss.n3875 1.13717
R20421 avss.n8177 avss.n8176 1.13717
R20422 avss.n8180 avss.n3869 1.13717
R20423 avss.n8191 avss.n8190 1.13717
R20424 avss.n8205 avss.n8204 1.13717
R20425 avss.n3865 avss.n3864 1.13717
R20426 avss.n8212 avss.n3859 1.13717
R20427 avss.n8221 avss.n3856 1.13717
R20428 avss.n3858 avss.n3857 1.13717
R20429 avss.n8231 avss.n8230 1.13717
R20430 avss.n8241 avss.n8240 1.13717
R20431 avss.n7593 avss.n7591 1.13717
R20432 avss.n7715 avss.n7662 1.13717
R20433 avss.n7770 avss.n7569 1.13717
R20434 avss.n7597 avss.n7592 1.13717
R20435 avss.n7614 avss.n7613 1.13717
R20436 avss.n7629 avss.n7620 1.13717
R20437 avss.n7645 avss.n7641 1.13717
R20438 avss.n7728 avss.n7647 1.13717
R20439 avss.n7677 avss.n7672 1.13717
R20440 avss.n7709 avss.n7708 1.13717
R20441 avss.n7576 avss.n7575 1.13717
R20442 avss.n7583 avss.n7582 1.13717
R20443 avss.n7596 avss.n7594 1.13717
R20444 avss.n7751 avss.n7750 1.13717
R20445 avss.n7633 avss.n7632 1.13717
R20446 avss.n7639 avss.n7624 1.13717
R20447 avss.n7650 avss.n7640 1.13717
R20448 avss.n7656 avss.n7648 1.13717
R20449 avss.n7721 avss.n7660 1.13717
R20450 avss.n7909 avss.n3926 1.13717
R20451 avss.n3987 avss.n3986 1.13717
R20452 avss.n3994 avss.n3993 1.13717
R20453 avss.n4001 avss.n3980 1.13717
R20454 avss.n7793 avss.n3971 1.13717
R20455 avss.n7804 avss.n3968 1.13717
R20456 avss.n7781 avss.n3969 1.13717
R20457 avss.n7813 avss.n3961 1.13717
R20458 avss.n3960 avss.n3959 1.13717
R20459 avss.n7824 avss.n7823 1.13717
R20460 avss.n7827 avss.n3953 1.13717
R20461 avss.n7838 avss.n7837 1.13717
R20462 avss.n7852 avss.n7851 1.13717
R20463 avss.n3949 avss.n3948 1.13717
R20464 avss.n7859 avss.n3943 1.13717
R20465 avss.n7868 avss.n3940 1.13717
R20466 avss.n3942 avss.n3941 1.13717
R20467 avss.n7878 avss.n7877 1.13717
R20468 avss.n7888 avss.n7887 1.13717
R20469 avss.n7240 avss.n7238 1.13717
R20470 avss.n7362 avss.n7309 1.13717
R20471 avss.n7417 avss.n7216 1.13717
R20472 avss.n7244 avss.n7239 1.13717
R20473 avss.n7261 avss.n7260 1.13717
R20474 avss.n7276 avss.n7267 1.13717
R20475 avss.n7292 avss.n7288 1.13717
R20476 avss.n7375 avss.n7294 1.13717
R20477 avss.n7324 avss.n7319 1.13717
R20478 avss.n7356 avss.n7355 1.13717
R20479 avss.n7223 avss.n7222 1.13717
R20480 avss.n7230 avss.n7229 1.13717
R20481 avss.n7243 avss.n7241 1.13717
R20482 avss.n7398 avss.n7397 1.13717
R20483 avss.n7280 avss.n7279 1.13717
R20484 avss.n7286 avss.n7271 1.13717
R20485 avss.n7297 avss.n7287 1.13717
R20486 avss.n7303 avss.n7295 1.13717
R20487 avss.n7368 avss.n7307 1.13717
R20488 avss.n7556 avss.n4010 1.13717
R20489 avss.n4071 avss.n4070 1.13717
R20490 avss.n4078 avss.n4077 1.13717
R20491 avss.n4085 avss.n4064 1.13717
R20492 avss.n7440 avss.n4055 1.13717
R20493 avss.n7451 avss.n4052 1.13717
R20494 avss.n7428 avss.n4053 1.13717
R20495 avss.n7460 avss.n4045 1.13717
R20496 avss.n4044 avss.n4043 1.13717
R20497 avss.n7471 avss.n7470 1.13717
R20498 avss.n7474 avss.n4037 1.13717
R20499 avss.n7485 avss.n7484 1.13717
R20500 avss.n7499 avss.n7498 1.13717
R20501 avss.n4033 avss.n4032 1.13717
R20502 avss.n7506 avss.n4027 1.13717
R20503 avss.n7515 avss.n4024 1.13717
R20504 avss.n4026 avss.n4025 1.13717
R20505 avss.n7525 avss.n7524 1.13717
R20506 avss.n7535 avss.n7534 1.13717
R20507 avss.n6887 avss.n6885 1.13717
R20508 avss.n7009 avss.n6956 1.13717
R20509 avss.n7064 avss.n6863 1.13717
R20510 avss.n6891 avss.n6886 1.13717
R20511 avss.n6908 avss.n6907 1.13717
R20512 avss.n6923 avss.n6914 1.13717
R20513 avss.n6939 avss.n6935 1.13717
R20514 avss.n7022 avss.n6941 1.13717
R20515 avss.n6971 avss.n6966 1.13717
R20516 avss.n7003 avss.n7002 1.13717
R20517 avss.n6870 avss.n6869 1.13717
R20518 avss.n6877 avss.n6876 1.13717
R20519 avss.n6890 avss.n6888 1.13717
R20520 avss.n7045 avss.n7044 1.13717
R20521 avss.n6927 avss.n6926 1.13717
R20522 avss.n6933 avss.n6918 1.13717
R20523 avss.n6944 avss.n6934 1.13717
R20524 avss.n6950 avss.n6942 1.13717
R20525 avss.n7015 avss.n6954 1.13717
R20526 avss.n7203 avss.n4094 1.13717
R20527 avss.n4155 avss.n4154 1.13717
R20528 avss.n4162 avss.n4161 1.13717
R20529 avss.n4169 avss.n4148 1.13717
R20530 avss.n7087 avss.n4139 1.13717
R20531 avss.n7098 avss.n4136 1.13717
R20532 avss.n7075 avss.n4137 1.13717
R20533 avss.n7107 avss.n4129 1.13717
R20534 avss.n4128 avss.n4127 1.13717
R20535 avss.n7118 avss.n7117 1.13717
R20536 avss.n7121 avss.n4121 1.13717
R20537 avss.n7132 avss.n7131 1.13717
R20538 avss.n7146 avss.n7145 1.13717
R20539 avss.n4117 avss.n4116 1.13717
R20540 avss.n7153 avss.n4111 1.13717
R20541 avss.n7162 avss.n4108 1.13717
R20542 avss.n4110 avss.n4109 1.13717
R20543 avss.n7172 avss.n7171 1.13717
R20544 avss.n7182 avss.n7181 1.13717
R20545 avss.n6534 avss.n6532 1.13717
R20546 avss.n6656 avss.n6603 1.13717
R20547 avss.n6711 avss.n6510 1.13717
R20548 avss.n6538 avss.n6533 1.13717
R20549 avss.n6555 avss.n6554 1.13717
R20550 avss.n6570 avss.n6561 1.13717
R20551 avss.n6586 avss.n6582 1.13717
R20552 avss.n6669 avss.n6588 1.13717
R20553 avss.n6618 avss.n6613 1.13717
R20554 avss.n6650 avss.n6649 1.13717
R20555 avss.n6517 avss.n6516 1.13717
R20556 avss.n6524 avss.n6523 1.13717
R20557 avss.n6537 avss.n6535 1.13717
R20558 avss.n6692 avss.n6691 1.13717
R20559 avss.n6574 avss.n6573 1.13717
R20560 avss.n6580 avss.n6565 1.13717
R20561 avss.n6591 avss.n6581 1.13717
R20562 avss.n6597 avss.n6589 1.13717
R20563 avss.n6662 avss.n6601 1.13717
R20564 avss.n6850 avss.n4178 1.13717
R20565 avss.n4239 avss.n4238 1.13717
R20566 avss.n4246 avss.n4245 1.13717
R20567 avss.n4253 avss.n4232 1.13717
R20568 avss.n6734 avss.n4223 1.13717
R20569 avss.n6745 avss.n4220 1.13717
R20570 avss.n6722 avss.n4221 1.13717
R20571 avss.n6754 avss.n4213 1.13717
R20572 avss.n4212 avss.n4211 1.13717
R20573 avss.n6765 avss.n6764 1.13717
R20574 avss.n6768 avss.n4205 1.13717
R20575 avss.n6779 avss.n6778 1.13717
R20576 avss.n6793 avss.n6792 1.13717
R20577 avss.n4201 avss.n4200 1.13717
R20578 avss.n6800 avss.n4195 1.13717
R20579 avss.n6809 avss.n4192 1.13717
R20580 avss.n4194 avss.n4193 1.13717
R20581 avss.n6819 avss.n6818 1.13717
R20582 avss.n6829 avss.n6828 1.13717
R20583 avss.n6181 avss.n6179 1.13717
R20584 avss.n6303 avss.n6250 1.13717
R20585 avss.n6358 avss.n6157 1.13717
R20586 avss.n6185 avss.n6180 1.13717
R20587 avss.n6202 avss.n6201 1.13717
R20588 avss.n6217 avss.n6208 1.13717
R20589 avss.n6233 avss.n6229 1.13717
R20590 avss.n6316 avss.n6235 1.13717
R20591 avss.n6265 avss.n6260 1.13717
R20592 avss.n6297 avss.n6296 1.13717
R20593 avss.n6164 avss.n6163 1.13717
R20594 avss.n6171 avss.n6170 1.13717
R20595 avss.n6184 avss.n6182 1.13717
R20596 avss.n6339 avss.n6338 1.13717
R20597 avss.n6221 avss.n6220 1.13717
R20598 avss.n6227 avss.n6212 1.13717
R20599 avss.n6238 avss.n6228 1.13717
R20600 avss.n6244 avss.n6236 1.13717
R20601 avss.n6309 avss.n6248 1.13717
R20602 avss.n6497 avss.n4262 1.13717
R20603 avss.n4323 avss.n4322 1.13717
R20604 avss.n4330 avss.n4329 1.13717
R20605 avss.n4337 avss.n4316 1.13717
R20606 avss.n6381 avss.n4307 1.13717
R20607 avss.n6392 avss.n4304 1.13717
R20608 avss.n6369 avss.n4305 1.13717
R20609 avss.n6401 avss.n4297 1.13717
R20610 avss.n4296 avss.n4295 1.13717
R20611 avss.n6412 avss.n6411 1.13717
R20612 avss.n6415 avss.n4289 1.13717
R20613 avss.n6426 avss.n6425 1.13717
R20614 avss.n6440 avss.n6439 1.13717
R20615 avss.n4285 avss.n4284 1.13717
R20616 avss.n6447 avss.n4279 1.13717
R20617 avss.n6456 avss.n4276 1.13717
R20618 avss.n4278 avss.n4277 1.13717
R20619 avss.n6466 avss.n6465 1.13717
R20620 avss.n6476 avss.n6475 1.13717
R20621 avss.n5828 avss.n5826 1.13717
R20622 avss.n5950 avss.n5897 1.13717
R20623 avss.n6005 avss.n5804 1.13717
R20624 avss.n5832 avss.n5827 1.13717
R20625 avss.n5849 avss.n5848 1.13717
R20626 avss.n5864 avss.n5855 1.13717
R20627 avss.n5880 avss.n5876 1.13717
R20628 avss.n5963 avss.n5882 1.13717
R20629 avss.n5912 avss.n5907 1.13717
R20630 avss.n5944 avss.n5943 1.13717
R20631 avss.n5811 avss.n5810 1.13717
R20632 avss.n5818 avss.n5817 1.13717
R20633 avss.n5831 avss.n5829 1.13717
R20634 avss.n5986 avss.n5985 1.13717
R20635 avss.n5868 avss.n5867 1.13717
R20636 avss.n5874 avss.n5859 1.13717
R20637 avss.n5885 avss.n5875 1.13717
R20638 avss.n5891 avss.n5883 1.13717
R20639 avss.n5956 avss.n5895 1.13717
R20640 avss.n6144 avss.n4346 1.13717
R20641 avss.n4407 avss.n4406 1.13717
R20642 avss.n4414 avss.n4413 1.13717
R20643 avss.n4421 avss.n4400 1.13717
R20644 avss.n6028 avss.n4391 1.13717
R20645 avss.n6039 avss.n4388 1.13717
R20646 avss.n6016 avss.n4389 1.13717
R20647 avss.n6048 avss.n4381 1.13717
R20648 avss.n4380 avss.n4379 1.13717
R20649 avss.n6059 avss.n6058 1.13717
R20650 avss.n6062 avss.n4373 1.13717
R20651 avss.n6073 avss.n6072 1.13717
R20652 avss.n6087 avss.n6086 1.13717
R20653 avss.n4369 avss.n4368 1.13717
R20654 avss.n6094 avss.n4363 1.13717
R20655 avss.n6103 avss.n4360 1.13717
R20656 avss.n4362 avss.n4361 1.13717
R20657 avss.n6113 avss.n6112 1.13717
R20658 avss.n6123 avss.n6122 1.13717
R20659 avss.n5475 avss.n5473 1.13717
R20660 avss.n5597 avss.n5544 1.13717
R20661 avss.n5652 avss.n5451 1.13717
R20662 avss.n5479 avss.n5474 1.13717
R20663 avss.n5496 avss.n5495 1.13717
R20664 avss.n5511 avss.n5502 1.13717
R20665 avss.n5527 avss.n5523 1.13717
R20666 avss.n5610 avss.n5529 1.13717
R20667 avss.n5559 avss.n5554 1.13717
R20668 avss.n5591 avss.n5590 1.13717
R20669 avss.n5458 avss.n5457 1.13717
R20670 avss.n5465 avss.n5464 1.13717
R20671 avss.n5478 avss.n5476 1.13717
R20672 avss.n5633 avss.n5632 1.13717
R20673 avss.n5515 avss.n5514 1.13717
R20674 avss.n5521 avss.n5506 1.13717
R20675 avss.n5532 avss.n5522 1.13717
R20676 avss.n5538 avss.n5530 1.13717
R20677 avss.n5603 avss.n5542 1.13717
R20678 avss.n5791 avss.n4430 1.13717
R20679 avss.n4491 avss.n4490 1.13717
R20680 avss.n4498 avss.n4497 1.13717
R20681 avss.n4505 avss.n4484 1.13717
R20682 avss.n5675 avss.n4475 1.13717
R20683 avss.n5686 avss.n4472 1.13717
R20684 avss.n5663 avss.n4473 1.13717
R20685 avss.n5695 avss.n4465 1.13717
R20686 avss.n4464 avss.n4463 1.13717
R20687 avss.n5706 avss.n5705 1.13717
R20688 avss.n5709 avss.n4457 1.13717
R20689 avss.n5720 avss.n5719 1.13717
R20690 avss.n5734 avss.n5733 1.13717
R20691 avss.n4453 avss.n4452 1.13717
R20692 avss.n5741 avss.n4447 1.13717
R20693 avss.n5750 avss.n4444 1.13717
R20694 avss.n4446 avss.n4445 1.13717
R20695 avss.n5760 avss.n5759 1.13717
R20696 avss.n5770 avss.n5769 1.13717
R20697 avss.n5125 avss.n5124 1.13717
R20698 avss.n5295 avss.n5095 1.13717
R20699 avss.n5150 avss.n5149 1.13717
R20700 avss.n5165 avss.n5156 1.13717
R20701 avss.n5181 avss.n5177 1.13717
R20702 avss.n5265 avss.n5183 1.13717
R20703 avss.n5219 avss.n5214 1.13717
R20704 avss.n5248 avss.n5207 1.13717
R20705 avss.n5110 avss.n5109 1.13717
R20706 avss.n5118 avss.n5117 1.13717
R20707 avss.n5299 avss.n5092 1.13717
R20708 avss.n5141 avss.n5140 1.13717
R20709 avss.n5288 avss.n5287 1.13717
R20710 avss.n5169 avss.n5168 1.13717
R20711 avss.n5175 avss.n5160 1.13717
R20712 avss.n5186 avss.n5176 1.13717
R20713 avss.n5192 avss.n5184 1.13717
R20714 avss.n5258 avss.n5196 1.13717
R20715 avss.n5252 avss.n5198 1.13717
R20716 avss.n5438 avss.n4514 1.13717
R20717 avss.n4575 avss.n4574 1.13717
R20718 avss.n4582 avss.n4581 1.13717
R20719 avss.n4589 avss.n4568 1.13717
R20720 avss.n5322 avss.n4559 1.13717
R20721 avss.n5333 avss.n4556 1.13717
R20722 avss.n5310 avss.n4557 1.13717
R20723 avss.n5342 avss.n4549 1.13717
R20724 avss.n4548 avss.n4547 1.13717
R20725 avss.n5353 avss.n5352 1.13717
R20726 avss.n5356 avss.n4541 1.13717
R20727 avss.n5367 avss.n5366 1.13717
R20728 avss.n5381 avss.n5380 1.13717
R20729 avss.n4537 avss.n4536 1.13717
R20730 avss.n5388 avss.n4531 1.13717
R20731 avss.n5397 avss.n4528 1.13717
R20732 avss.n4530 avss.n4529 1.13717
R20733 avss.n5407 avss.n5406 1.13717
R20734 avss.n5417 avss.n5416 1.13717
R20735 avss.n4771 avss.n4770 1.13717
R20736 avss.n4941 avss.n4741 1.13717
R20737 avss.n4796 avss.n4795 1.13717
R20738 avss.n4811 avss.n4802 1.13717
R20739 avss.n4827 avss.n4823 1.13717
R20740 avss.n4911 avss.n4829 1.13717
R20741 avss.n4865 avss.n4860 1.13717
R20742 avss.n4894 avss.n4853 1.13717
R20743 avss.n4756 avss.n4755 1.13717
R20744 avss.n4764 avss.n4763 1.13717
R20745 avss.n4945 avss.n4738 1.13717
R20746 avss.n4787 avss.n4786 1.13717
R20747 avss.n4934 avss.n4933 1.13717
R20748 avss.n4815 avss.n4814 1.13717
R20749 avss.n4821 avss.n4806 1.13717
R20750 avss.n4832 avss.n4822 1.13717
R20751 avss.n4838 avss.n4830 1.13717
R20752 avss.n4904 avss.n4842 1.13717
R20753 avss.n4898 avss.n4844 1.13717
R20754 avss.n5084 avss.n4598 1.13717
R20755 avss.n4659 avss.n4658 1.13717
R20756 avss.n4666 avss.n4665 1.13717
R20757 avss.n4673 avss.n4652 1.13717
R20758 avss.n4968 avss.n4643 1.13717
R20759 avss.n4979 avss.n4640 1.13717
R20760 avss.n4956 avss.n4641 1.13717
R20761 avss.n4988 avss.n4633 1.13717
R20762 avss.n4632 avss.n4631 1.13717
R20763 avss.n4999 avss.n4998 1.13717
R20764 avss.n5002 avss.n4625 1.13717
R20765 avss.n5013 avss.n5012 1.13717
R20766 avss.n5027 avss.n5026 1.13717
R20767 avss.n4621 avss.n4620 1.13717
R20768 avss.n5034 avss.n4615 1.13717
R20769 avss.n5043 avss.n4612 1.13717
R20770 avss.n4614 avss.n4613 1.13717
R20771 avss.n5053 avss.n5052 1.13717
R20772 avss.n5063 avss.n5062 1.13717
R20773 avss.n2406 avss.n2405 1.13717
R20774 avss.n2477 avss.n2476 1.13717
R20775 avss.n2457 avss.n2456 1.13717
R20776 avss.n2442 avss.n2441 1.13717
R20777 avss.n9132 avss.n9131 1.13717
R20778 avss.n9149 avss.n9148 1.13717
R20779 avss.n9169 avss.n9168 1.13717
R20780 avss.n9114 avss.n9113 1.13717
R20781 avss.n2421 avss.n2420 1.13717
R20782 avss.n2568 avss.n2567 1.13717
R20783 avss.n2553 avss.n2552 1.13717
R20784 avss.n2534 avss.n2533 1.13717
R20785 avss.n2514 avss.n2513 1.13717
R20786 avss.n2499 avss.n2498 1.13717
R20787 avss.n9021 avss.n9020 1.13717
R20788 avss.n9038 avss.n9037 1.13717
R20789 avss.n9058 avss.n9057 1.13717
R20790 avss.n9002 avss.n9001 1.13717
R20791 avss.n2190 avss.n2189 1.13717
R20792 avss.n2261 avss.n2260 1.13717
R20793 avss.n2241 avss.n2240 1.13717
R20794 avss.n2226 avss.n2225 1.13717
R20795 avss.n9353 avss.n9352 1.13717
R20796 avss.n9370 avss.n9369 1.13717
R20797 avss.n9390 avss.n9389 1.13717
R20798 avss.n9335 avss.n9334 1.13717
R20799 avss.n2205 avss.n2204 1.13717
R20800 avss.n2352 avss.n2351 1.13717
R20801 avss.n2337 avss.n2336 1.13717
R20802 avss.n2318 avss.n2317 1.13717
R20803 avss.n2298 avss.n2297 1.13717
R20804 avss.n2283 avss.n2282 1.13717
R20805 avss.n9242 avss.n9241 1.13717
R20806 avss.n9259 avss.n9258 1.13717
R20807 avss.n9279 avss.n9278 1.13717
R20808 avss.n9223 avss.n9222 1.13717
R20809 avss.n1974 avss.n1973 1.13717
R20810 avss.n2045 avss.n2044 1.13717
R20811 avss.n2025 avss.n2024 1.13717
R20812 avss.n2010 avss.n2009 1.13717
R20813 avss.n9574 avss.n9573 1.13717
R20814 avss.n9591 avss.n9590 1.13717
R20815 avss.n9611 avss.n9610 1.13717
R20816 avss.n9556 avss.n9555 1.13717
R20817 avss.n1989 avss.n1988 1.13717
R20818 avss.n2136 avss.n2135 1.13717
R20819 avss.n2121 avss.n2120 1.13717
R20820 avss.n2102 avss.n2101 1.13717
R20821 avss.n2082 avss.n2081 1.13717
R20822 avss.n2067 avss.n2066 1.13717
R20823 avss.n9463 avss.n9462 1.13717
R20824 avss.n9480 avss.n9479 1.13717
R20825 avss.n9500 avss.n9499 1.13717
R20826 avss.n9444 avss.n9443 1.13717
R20827 avss.n1758 avss.n1757 1.13717
R20828 avss.n1829 avss.n1828 1.13717
R20829 avss.n1809 avss.n1808 1.13717
R20830 avss.n1794 avss.n1793 1.13717
R20831 avss.n9795 avss.n9794 1.13717
R20832 avss.n9812 avss.n9811 1.13717
R20833 avss.n9832 avss.n9831 1.13717
R20834 avss.n9777 avss.n9776 1.13717
R20835 avss.n1773 avss.n1772 1.13717
R20836 avss.n1920 avss.n1919 1.13717
R20837 avss.n1905 avss.n1904 1.13717
R20838 avss.n1886 avss.n1885 1.13717
R20839 avss.n1866 avss.n1865 1.13717
R20840 avss.n1851 avss.n1850 1.13717
R20841 avss.n9684 avss.n9683 1.13717
R20842 avss.n9701 avss.n9700 1.13717
R20843 avss.n9721 avss.n9720 1.13717
R20844 avss.n9665 avss.n9664 1.13717
R20845 avss.n1542 avss.n1541 1.13717
R20846 avss.n1613 avss.n1612 1.13717
R20847 avss.n1593 avss.n1592 1.13717
R20848 avss.n1578 avss.n1577 1.13717
R20849 avss.n10016 avss.n10015 1.13717
R20850 avss.n10033 avss.n10032 1.13717
R20851 avss.n10053 avss.n10052 1.13717
R20852 avss.n9998 avss.n9997 1.13717
R20853 avss.n1557 avss.n1556 1.13717
R20854 avss.n1704 avss.n1703 1.13717
R20855 avss.n1689 avss.n1688 1.13717
R20856 avss.n1670 avss.n1669 1.13717
R20857 avss.n1650 avss.n1649 1.13717
R20858 avss.n1635 avss.n1634 1.13717
R20859 avss.n9905 avss.n9904 1.13717
R20860 avss.n9922 avss.n9921 1.13717
R20861 avss.n9942 avss.n9941 1.13717
R20862 avss.n9886 avss.n9885 1.13717
R20863 avss.n1326 avss.n1325 1.13717
R20864 avss.n1397 avss.n1396 1.13717
R20865 avss.n1377 avss.n1376 1.13717
R20866 avss.n1362 avss.n1361 1.13717
R20867 avss.n10237 avss.n10236 1.13717
R20868 avss.n10254 avss.n10253 1.13717
R20869 avss.n10274 avss.n10273 1.13717
R20870 avss.n10219 avss.n10218 1.13717
R20871 avss.n1341 avss.n1340 1.13717
R20872 avss.n1488 avss.n1487 1.13717
R20873 avss.n1473 avss.n1472 1.13717
R20874 avss.n1454 avss.n1453 1.13717
R20875 avss.n1434 avss.n1433 1.13717
R20876 avss.n1419 avss.n1418 1.13717
R20877 avss.n10126 avss.n10125 1.13717
R20878 avss.n10143 avss.n10142 1.13717
R20879 avss.n10163 avss.n10162 1.13717
R20880 avss.n10107 avss.n10106 1.13717
R20881 avss.n1110 avss.n1109 1.13717
R20882 avss.n1181 avss.n1180 1.13717
R20883 avss.n1161 avss.n1160 1.13717
R20884 avss.n1146 avss.n1145 1.13717
R20885 avss.n10458 avss.n10457 1.13717
R20886 avss.n10475 avss.n10474 1.13717
R20887 avss.n10495 avss.n10494 1.13717
R20888 avss.n10440 avss.n10439 1.13717
R20889 avss.n1125 avss.n1124 1.13717
R20890 avss.n1272 avss.n1271 1.13717
R20891 avss.n1257 avss.n1256 1.13717
R20892 avss.n1238 avss.n1237 1.13717
R20893 avss.n1218 avss.n1217 1.13717
R20894 avss.n1203 avss.n1202 1.13717
R20895 avss.n10347 avss.n10346 1.13717
R20896 avss.n10364 avss.n10363 1.13717
R20897 avss.n10384 avss.n10383 1.13717
R20898 avss.n10328 avss.n10327 1.13717
R20899 avss.n894 avss.n893 1.13717
R20900 avss.n965 avss.n964 1.13717
R20901 avss.n945 avss.n944 1.13717
R20902 avss.n930 avss.n929 1.13717
R20903 avss.n10679 avss.n10678 1.13717
R20904 avss.n10696 avss.n10695 1.13717
R20905 avss.n10716 avss.n10715 1.13717
R20906 avss.n10661 avss.n10660 1.13717
R20907 avss.n909 avss.n908 1.13717
R20908 avss.n1056 avss.n1055 1.13717
R20909 avss.n1041 avss.n1040 1.13717
R20910 avss.n1022 avss.n1021 1.13717
R20911 avss.n1002 avss.n1001 1.13717
R20912 avss.n987 avss.n986 1.13717
R20913 avss.n10568 avss.n10567 1.13717
R20914 avss.n10585 avss.n10584 1.13717
R20915 avss.n10605 avss.n10604 1.13717
R20916 avss.n10549 avss.n10548 1.13717
R20917 avss.n678 avss.n677 1.13717
R20918 avss.n749 avss.n748 1.13717
R20919 avss.n729 avss.n728 1.13717
R20920 avss.n714 avss.n713 1.13717
R20921 avss.n10900 avss.n10899 1.13717
R20922 avss.n10917 avss.n10916 1.13717
R20923 avss.n10937 avss.n10936 1.13717
R20924 avss.n10882 avss.n10881 1.13717
R20925 avss.n693 avss.n692 1.13717
R20926 avss.n840 avss.n839 1.13717
R20927 avss.n825 avss.n824 1.13717
R20928 avss.n806 avss.n805 1.13717
R20929 avss.n786 avss.n785 1.13717
R20930 avss.n771 avss.n770 1.13717
R20931 avss.n10789 avss.n10788 1.13717
R20932 avss.n10806 avss.n10805 1.13717
R20933 avss.n10826 avss.n10825 1.13717
R20934 avss.n10770 avss.n10769 1.13717
R20935 avss.n462 avss.n461 1.13717
R20936 avss.n533 avss.n532 1.13717
R20937 avss.n513 avss.n512 1.13717
R20938 avss.n498 avss.n497 1.13717
R20939 avss.n11121 avss.n11120 1.13717
R20940 avss.n11138 avss.n11137 1.13717
R20941 avss.n11158 avss.n11157 1.13717
R20942 avss.n11103 avss.n11102 1.13717
R20943 avss.n477 avss.n476 1.13717
R20944 avss.n624 avss.n623 1.13717
R20945 avss.n609 avss.n608 1.13717
R20946 avss.n590 avss.n589 1.13717
R20947 avss.n570 avss.n569 1.13717
R20948 avss.n555 avss.n554 1.13717
R20949 avss.n11010 avss.n11009 1.13717
R20950 avss.n11027 avss.n11026 1.13717
R20951 avss.n11047 avss.n11046 1.13717
R20952 avss.n10991 avss.n10990 1.13717
R20953 avss.n11380 avss.n11379 1.13717
R20954 avss.n11362 avss.n11361 1.13717
R20955 avss.n11342 avss.n11341 1.13717
R20956 avss.n11327 avss.n11326 1.13717
R20957 avss.n388 avss.n387 1.13717
R20958 avss.n405 avss.n404 1.13717
R20959 avss.n425 avss.n424 1.13717
R20960 avss.n369 avss.n368 1.13717
R20961 avss.n11396 avss.n11395 1.13717
R20962 avss.n299 avss.n298 1.13717
R20963 avss.n284 avss.n283 1.13717
R20964 avss.n265 avss.n264 1.13717
R20965 avss.n245 avss.n244 1.13717
R20966 avss.n230 avss.n229 1.13717
R20967 avss.n11231 avss.n11230 1.13717
R20968 avss.n11248 avss.n11247 1.13717
R20969 avss.n11268 avss.n11267 1.13717
R20970 avss.n11212 avss.n11211 1.13717
R20971 avss.n11601 avss.n11600 1.13717
R20972 avss.n11583 avss.n11582 1.13717
R20973 avss.n11563 avss.n11562 1.13717
R20974 avss.n11548 avss.n11547 1.13717
R20975 avss.n171 avss.n170 1.13717
R20976 avss.n188 avss.n187 1.13717
R20977 avss.n208 avss.n207 1.13717
R20978 avss.n152 avss.n151 1.13717
R20979 avss.n11617 avss.n11616 1.13717
R20980 avss.n82 avss.n81 1.13717
R20981 avss.n67 avss.n66 1.13717
R20982 avss.n48 avss.n47 1.13717
R20983 avss.n28 avss.n27 1.13717
R20984 avss.n13 avss.n12 1.13717
R20985 avss.n11452 avss.n11451 1.13717
R20986 avss.n11469 avss.n11468 1.13717
R20987 avss.n11489 avss.n11488 1.13717
R20988 avss.n11433 avss.n11432 1.13717
R20989 avss.n3457 avss.n3198 1.12991
R20990 avss.n3460 avss.n3458 1.12991
R20991 avss.n8832 avss.n8626 1.12685
R20992 avss.n8479 avss.n8273 1.12685
R20993 avss.n8126 avss.n7920 1.12685
R20994 avss.n7773 avss.n7567 1.12685
R20995 avss.n7420 avss.n7214 1.12685
R20996 avss.n7067 avss.n6861 1.12685
R20997 avss.n6714 avss.n6508 1.12685
R20998 avss.n6361 avss.n6155 1.12685
R20999 avss.n6008 avss.n5802 1.12685
R21000 avss.n5655 avss.n5449 1.12685
R21001 avss.n5106 avss.n5089 1.12685
R21002 avss.n4752 avss.n4735 1.12685
R21003 avss.n8843 avss.n3727 1.12654
R21004 avss.n8490 avss.n3811 1.12654
R21005 avss.n8137 avss.n3895 1.12654
R21006 avss.n7784 avss.n3979 1.12654
R21007 avss.n7431 avss.n4063 1.12654
R21008 avss.n7078 avss.n4147 1.12654
R21009 avss.n6725 avss.n4231 1.12654
R21010 avss.n6372 avss.n4315 1.12654
R21011 avss.n6019 avss.n4399 1.12654
R21012 avss.n5666 avss.n4483 1.12654
R21013 avss.n5302 avss.n5089 1.12654
R21014 avss.n5313 avss.n4567 1.12654
R21015 avss.n4948 avss.n4735 1.12654
R21016 avss.n4959 avss.n4651 1.12654
R21017 avss.n8973 avss.n8972 1.11238
R21018 avss.n3266 avss 0.986602
R21019 avss avss.n3526 0.986602
R21020 avss.n3525 avss 0.986602
R21021 avss.n3267 avss 0.986602
R21022 avss.n2979 avss.n2978 0.974413
R21023 avss.n3036 avss.n3035 0.974413
R21024 avss.n3132 avss.n3131 0.974413
R21025 avss.n3628 avss.n3627 0.974413
R21026 avss.n2691 avss.n2690 0.974413
R21027 avss.n2736 avss.n2735 0.974413
R21028 avss.n2906 avss.n2905 0.974413
R21029 avss.n2866 avss.n2865 0.974413
R21030 avss avss.n11636 0.958395
R21031 avss.n9305 avss.n9195 0.889356
R21032 avss.n8836 avss.n8619 0.889356
R21033 avss.n9526 avss.n9416 0.879776
R21034 avss.n8483 avss.n8266 0.879776
R21035 avss.n7424 avss.n7207 0.870211
R21036 avss.n8130 avss.n7913 0.870211
R21037 avss.n10189 avss.n10079 0.870211
R21038 avss.n9747 avss.n9637 0.870211
R21039 avss.n7777 avss.n7560 0.869861
R21040 avss.n9968 avss.n9858 0.869861
R21041 avss.n7071 avss.n6854 0.860633
R21042 avss.n10410 avss.n10300 0.860633
R21043 avss.n6012 avss.n5795 0.851069
R21044 avss.n6365 avss.n6148 0.851069
R21045 avss.n6718 avss.n6501 0.851069
R21046 avss.n11073 avss.n10963 0.851069
R21047 avss.n10852 avss.n10742 0.851069
R21048 avss.n10631 avss.n10521 0.851069
R21049 avss.n5659 avss.n5442 0.841493
R21050 avss.n11294 avss.n11184 0.841493
R21051 avss.n8833 avss.n8832 0.840061
R21052 avss.n8480 avss.n8479 0.840061
R21053 avss.n8127 avss.n8126 0.840061
R21054 avss.n7774 avss.n7773 0.840061
R21055 avss.n7421 avss.n7420 0.840061
R21056 avss.n7068 avss.n7067 0.840061
R21057 avss.n6715 avss.n6714 0.840061
R21058 avss.n6362 avss.n6361 0.840061
R21059 avss.n6009 avss.n6008 0.840061
R21060 avss.n5656 avss.n5655 0.840061
R21061 avss.n2483 avss.n2482 0.840061
R21062 avss.n2267 avss.n2266 0.840061
R21063 avss.n2051 avss.n2050 0.840061
R21064 avss.n1835 avss.n1834 0.840061
R21065 avss.n1619 avss.n1618 0.840061
R21066 avss.n1403 avss.n1402 0.840061
R21067 avss.n1187 avss.n1186 0.840061
R21068 avss.n971 avss.n970 0.840061
R21069 avss.n755 avss.n754 0.840061
R21070 avss.n539 avss.n538 0.840061
R21071 avss.n8843 avss.n3725 0.839956
R21072 avss.n8490 avss.n3809 0.839956
R21073 avss.n8137 avss.n3893 0.839956
R21074 avss.n7784 avss.n3977 0.839956
R21075 avss.n7431 avss.n4061 0.839956
R21076 avss.n7078 avss.n4145 0.839956
R21077 avss.n6725 avss.n4229 0.839956
R21078 avss.n6372 avss.n4313 0.839956
R21079 avss.n6019 avss.n4397 0.839956
R21080 avss.n5666 avss.n4481 0.839956
R21081 avss.n5313 avss.n4565 0.839956
R21082 avss.n4959 avss.n4649 0.839956
R21083 avss.n5252 avss.n5202 0.836349
R21084 avss.n4898 avss.n4848 0.836349
R21085 avss.n432 avss.n431 0.836349
R21086 avss.n215 avss.n214 0.836349
R21087 avss.n8774 avss.n8726 0.836347
R21088 avss.n8421 avss.n8373 0.836347
R21089 avss.n8068 avss.n8020 0.836347
R21090 avss.n7715 avss.n7667 0.836347
R21091 avss.n7362 avss.n7314 0.836347
R21092 avss.n7009 avss.n6961 0.836347
R21093 avss.n6656 avss.n6608 0.836347
R21094 avss.n6303 avss.n6255 0.836347
R21095 avss.n5950 avss.n5902 0.836347
R21096 avss.n5597 avss.n5549 0.836347
R21097 avss.n9191 avss.n9175 0.836347
R21098 avss.n9412 avss.n9396 0.836347
R21099 avss.n9633 avss.n9617 0.836347
R21100 avss.n9854 avss.n9838 0.836347
R21101 avss.n10075 avss.n10059 0.836347
R21102 avss.n10296 avss.n10280 0.836347
R21103 avss.n10517 avss.n10501 0.836347
R21104 avss.n10738 avss.n10722 0.836347
R21105 avss.n10959 avss.n10943 0.836347
R21106 avss.n11180 avss.n11164 0.836347
R21107 avss.n8968 avss.n3678 0.836346
R21108 avss.n8615 avss.n3762 0.836346
R21109 avss.n8262 avss.n3846 0.836346
R21110 avss.n7909 avss.n3930 0.836346
R21111 avss.n7556 avss.n4014 0.836346
R21112 avss.n7203 avss.n4098 0.836346
R21113 avss.n6850 avss.n4182 0.836346
R21114 avss.n6497 avss.n4266 0.836346
R21115 avss.n6144 avss.n4350 0.836346
R21116 avss.n5791 avss.n4434 0.836346
R21117 avss.n5438 avss.n4518 0.836346
R21118 avss.n5084 avss.n4602 0.836346
R21119 avss.n9081 avss.n9063 0.836346
R21120 avss.n9302 avss.n9284 0.836346
R21121 avss.n9523 avss.n9505 0.836346
R21122 avss.n9744 avss.n9726 0.836346
R21123 avss.n9965 avss.n9947 0.836346
R21124 avss.n10186 avss.n10168 0.836346
R21125 avss.n10407 avss.n10389 0.836346
R21126 avss.n10628 avss.n10610 0.836346
R21127 avss.n10849 avss.n10831 0.836346
R21128 avss.n11070 avss.n11052 0.836346
R21129 avss.n11291 avss.n11273 0.836346
R21130 avss.n11512 avss.n11494 0.836346
R21131 avss.n3009 avss.n2947 0.833377
R21132 avss.n3066 avss.n2931 0.833377
R21133 avss.n3103 avss.n3102 0.833377
R21134 avss.n3658 avss.n2597 0.833377
R21135 avss.n2721 avss.n2660 0.833377
R21136 avss.n2766 avss.n2633 0.833377
R21137 avss.n2877 avss.n2876 0.833377
R21138 avss.n2837 avss.n2836 0.833377
R21139 avss.n11515 avss.n11405 0.831931
R21140 avss.n5306 avss.n5088 0.831931
R21141 avss.n3394 avss.n3196 0.827063
R21142 avss.n3340 avss.n3295 0.753441
R21143 avss.n3346 avss.n3345 0.753441
R21144 avss.n3240 avss.n3239 0.753441
R21145 avss.n3410 avss.n3241 0.753441
R21146 avss.n3435 avss.n3200 0.753441
R21147 avss.n3212 avss.n3201 0.753441
R21148 avss.n3214 avss.n3213 0.753441
R21149 avss.n3519 avss.n3518 0.753441
R21150 avss.n3507 avss.n3172 0.753441
R21151 avss.n8753 avss.n8752 0.738896
R21152 avss.n8400 avss.n8399 0.738896
R21153 avss.n8047 avss.n8046 0.738896
R21154 avss.n7694 avss.n7693 0.738896
R21155 avss.n7341 avss.n7340 0.738896
R21156 avss.n6988 avss.n6987 0.738896
R21157 avss.n6635 avss.n6634 0.738896
R21158 avss.n6282 avss.n6281 0.738896
R21159 avss.n5929 avss.n5928 0.738896
R21160 avss.n5576 avss.n5575 0.738896
R21161 avss.n5235 avss.n5234 0.738896
R21162 avss.n4881 avss.n4880 0.738896
R21163 avss.n9099 avss.n9098 0.738896
R21164 avss.n9320 avss.n9319 0.738896
R21165 avss.n9541 avss.n9540 0.738896
R21166 avss.n9762 avss.n9761 0.738896
R21167 avss.n9983 avss.n9982 0.738896
R21168 avss.n10204 avss.n10203 0.738896
R21169 avss.n10425 avss.n10424 0.738896
R21170 avss.n10646 avss.n10645 0.738896
R21171 avss.n10867 avss.n10866 0.738896
R21172 avss.n11088 avss.n11087 0.738896
R21173 avss.n339 avss.n338 0.738896
R21174 avss.n122 avss.n121 0.738896
R21175 avss.n8959 avss.n3679 0.738877
R21176 avss.n8606 avss.n3763 0.738877
R21177 avss.n8253 avss.n3847 0.738877
R21178 avss.n7900 avss.n3931 0.738877
R21179 avss.n7547 avss.n4015 0.738877
R21180 avss.n7194 avss.n4099 0.738877
R21181 avss.n6841 avss.n4183 0.738877
R21182 avss.n6488 avss.n4267 0.738877
R21183 avss.n6135 avss.n4351 0.738877
R21184 avss.n5782 avss.n4435 0.738877
R21185 avss.n5429 avss.n4519 0.738877
R21186 avss.n5075 avss.n4603 0.738877
R21187 avss.n9079 avss.n9078 0.738877
R21188 avss.n9300 avss.n9299 0.738877
R21189 avss.n9521 avss.n9520 0.738877
R21190 avss.n9742 avss.n9741 0.738877
R21191 avss.n9963 avss.n9962 0.738877
R21192 avss.n10184 avss.n10183 0.738877
R21193 avss.n10405 avss.n10404 0.738877
R21194 avss.n10626 avss.n10625 0.738877
R21195 avss.n10847 avss.n10846 0.738877
R21196 avss.n11068 avss.n11067 0.738877
R21197 avss.n11289 avss.n11288 0.738877
R21198 avss.n11510 avss.n11509 0.738877
R21199 avss avss.n3622 0.704167
R21200 avss avss.n2683 0.704167
R21201 avss avss.n2973 0.703251
R21202 avss avss.n3030 0.703251
R21203 avss.n3137 avss 0.703251
R21204 avss avss.n2808 0.703251
R21205 avss.n2913 avss 0.703251
R21206 avss avss.n2656 0.703251
R21207 avss.n3740 avss.n3739 0.55125
R21208 avss.n3824 avss.n3823 0.55125
R21209 avss.n3908 avss.n3907 0.55125
R21210 avss.n3992 avss.n3991 0.55125
R21211 avss.n4076 avss.n4075 0.55125
R21212 avss.n4160 avss.n4159 0.55125
R21213 avss.n4244 avss.n4243 0.55125
R21214 avss.n4328 avss.n4327 0.55125
R21215 avss.n4412 avss.n4411 0.55125
R21216 avss.n4496 avss.n4495 0.55125
R21217 avss.n4580 avss.n4579 0.55125
R21218 avss.n4664 avss.n4663 0.55125
R21219 avss.n2572 avss.n2571 0.55125
R21220 avss.n2356 avss.n2355 0.55125
R21221 avss.n2140 avss.n2139 0.55125
R21222 avss.n1924 avss.n1923 0.55125
R21223 avss.n1708 avss.n1707 0.55125
R21224 avss.n1492 avss.n1491 0.55125
R21225 avss.n1276 avss.n1275 0.55125
R21226 avss.n1060 avss.n1059 0.55125
R21227 avss.n844 avss.n843 0.55125
R21228 avss.n628 avss.n627 0.55125
R21229 avss.n303 avss.n302 0.55125
R21230 avss.n86 avss.n85 0.55125
R21231 avss.n8640 avss.n8639 0.550534
R21232 avss.n8287 avss.n8286 0.550534
R21233 avss.n7934 avss.n7933 0.550534
R21234 avss.n7581 avss.n7580 0.550534
R21235 avss.n7228 avss.n7227 0.550534
R21236 avss.n6875 avss.n6874 0.550534
R21237 avss.n6522 avss.n6521 0.550534
R21238 avss.n6169 avss.n6168 0.550534
R21239 avss.n5816 avss.n5815 0.550534
R21240 avss.n5463 avss.n5462 0.550534
R21241 avss.n5115 avss.n5114 0.550534
R21242 avss.n4761 avss.n4760 0.550534
R21243 avss.n2425 avss.n2424 0.550534
R21244 avss.n2209 avss.n2208 0.550534
R21245 avss.n1993 avss.n1992 0.550534
R21246 avss.n1777 avss.n1776 0.550534
R21247 avss.n1561 avss.n1560 0.550534
R21248 avss.n1345 avss.n1344 0.550534
R21249 avss.n1129 avss.n1128 0.550534
R21250 avss.n913 avss.n912 0.550534
R21251 avss.n697 avss.n696 0.550534
R21252 avss.n481 avss.n480 0.550534
R21253 avss.n11400 avss.n11399 0.550534
R21254 avss.n11621 avss.n11620 0.550534
R21255 avss.n3010 avss.n3008 0.526527
R21256 avss.n3067 avss.n3065 0.526527
R21257 avss.n3092 avss.n3090 0.526527
R21258 avss.n3659 avss.n3657 0.526527
R21259 avss.n2722 avss.n2720 0.526527
R21260 avss.n2767 avss.n2765 0.526527
R21261 avss.n2790 avss.n2788 0.526527
R21262 avss.n2826 avss.n2824 0.526527
R21263 avss.n3339 avss.n3337 0.440083
R21264 avss.n2961 avss.n2959 0.417891
R21265 avss.n2984 avss.n2957 0.417891
R21266 avss.n3018 avss.n2943 0.417891
R21267 avss.n3041 avss.n2941 0.417891
R21268 avss.n3077 avss.n3076 0.417891
R21269 avss.n3127 avss.n3079 0.417891
R21270 avss.n3095 avss.n2609 0.417891
R21271 avss.n3633 avss.n2607 0.417891
R21272 avss.n2685 avss.n2672 0.417891
R21273 avss.n2696 avss.n2670 0.417891
R21274 avss.n2730 avss.n2645 0.417891
R21275 avss.n2741 avss.n2643 0.417891
R21276 avss.n2908 avss.n2907 0.417891
R21277 avss.n2901 avss.n2777 0.417891
R21278 avss.n2811 avss.n2793 0.417891
R21279 avss.n2861 avss.n2813 0.417891
R21280 avss.n3002 avss.n3001 0.409011
R21281 avss.n3059 avss.n3058 0.409011
R21282 avss.n3112 avss.n3088 0.409011
R21283 avss.n3651 avss.n3650 0.409011
R21284 avss.n2714 avss.n2713 0.409011
R21285 avss.n2759 avss.n2758 0.409011
R21286 avss.n2886 avss.n2786 0.409011
R21287 avss.n2846 avss.n2822 0.409011
R21288 avss.n3509 avss.n3176 0.39052
R21289 avss.n3291 avss.n3287 0.376971
R21290 avss.n3365 avss.n3272 0.3755
R21291 avss.n3348 avss.n3293 0.359875
R21292 avss.n3464 avss.n3175 0.341125
R21293 avss.n8646 avss.n8645 0.329317
R21294 avss.n8791 avss.n8790 0.329317
R21295 avss.n3746 avss.n3745 0.329317
R21296 avss.n8915 avss.n8914 0.329317
R21297 avss.n8293 avss.n8292 0.329317
R21298 avss.n8438 avss.n8437 0.329317
R21299 avss.n3830 avss.n3829 0.329317
R21300 avss.n8562 avss.n8561 0.329317
R21301 avss.n7940 avss.n7939 0.329317
R21302 avss.n8085 avss.n8084 0.329317
R21303 avss.n3914 avss.n3913 0.329317
R21304 avss.n8209 avss.n8208 0.329317
R21305 avss.n7587 avss.n7586 0.329317
R21306 avss.n7732 avss.n7731 0.329317
R21307 avss.n3998 avss.n3997 0.329317
R21308 avss.n7856 avss.n7855 0.329317
R21309 avss.n7234 avss.n7233 0.329317
R21310 avss.n7379 avss.n7378 0.329317
R21311 avss.n4082 avss.n4081 0.329317
R21312 avss.n7503 avss.n7502 0.329317
R21313 avss.n6881 avss.n6880 0.329317
R21314 avss.n7026 avss.n7025 0.329317
R21315 avss.n4166 avss.n4165 0.329317
R21316 avss.n7150 avss.n7149 0.329317
R21317 avss.n6528 avss.n6527 0.329317
R21318 avss.n6673 avss.n6672 0.329317
R21319 avss.n4250 avss.n4249 0.329317
R21320 avss.n6797 avss.n6796 0.329317
R21321 avss.n6175 avss.n6174 0.329317
R21322 avss.n6320 avss.n6319 0.329317
R21323 avss.n4334 avss.n4333 0.329317
R21324 avss.n6444 avss.n6443 0.329317
R21325 avss.n5822 avss.n5821 0.329317
R21326 avss.n5967 avss.n5966 0.329317
R21327 avss.n4418 avss.n4417 0.329317
R21328 avss.n6091 avss.n6090 0.329317
R21329 avss.n5469 avss.n5468 0.329317
R21330 avss.n5614 avss.n5613 0.329317
R21331 avss.n4502 avss.n4501 0.329317
R21332 avss.n5738 avss.n5737 0.329317
R21333 avss.n5122 avss.n5121 0.329317
R21334 avss.n5269 avss.n5268 0.329317
R21335 avss.n4586 avss.n4585 0.329317
R21336 avss.n5385 avss.n5384 0.329317
R21337 avss.n4768 avss.n4767 0.329317
R21338 avss.n4915 avss.n4914 0.329317
R21339 avss.n4670 avss.n4669 0.329317
R21340 avss.n5031 avss.n5030 0.329317
R21341 avss.n8823 avss.n8822 0.306507
R21342 avss.n8814 avss.n8813 0.306507
R21343 avss.n8800 avss.n8799 0.306507
R21344 avss.n8732 avss.n8718 0.306507
R21345 avss.n8743 avss.n8742 0.306507
R21346 avss.n8848 avss.n8847 0.306507
R21347 avss.n8868 avss.n8867 0.306507
R21348 avss.n8895 avss.n8894 0.306507
R21349 avss.n8932 avss.n8931 0.306507
R21350 avss.n8943 avss.n8942 0.306507
R21351 avss.n8470 avss.n8469 0.306507
R21352 avss.n8461 avss.n8460 0.306507
R21353 avss.n8447 avss.n8446 0.306507
R21354 avss.n8379 avss.n8365 0.306507
R21355 avss.n8390 avss.n8389 0.306507
R21356 avss.n8495 avss.n8494 0.306507
R21357 avss.n8515 avss.n8514 0.306507
R21358 avss.n8542 avss.n8541 0.306507
R21359 avss.n8579 avss.n8578 0.306507
R21360 avss.n8590 avss.n8589 0.306507
R21361 avss.n8117 avss.n8116 0.306507
R21362 avss.n8108 avss.n8107 0.306507
R21363 avss.n8094 avss.n8093 0.306507
R21364 avss.n8026 avss.n8012 0.306507
R21365 avss.n8037 avss.n8036 0.306507
R21366 avss.n8142 avss.n8141 0.306507
R21367 avss.n8162 avss.n8161 0.306507
R21368 avss.n8189 avss.n8188 0.306507
R21369 avss.n8226 avss.n8225 0.306507
R21370 avss.n8237 avss.n8236 0.306507
R21371 avss.n7764 avss.n7763 0.306507
R21372 avss.n7755 avss.n7754 0.306507
R21373 avss.n7741 avss.n7740 0.306507
R21374 avss.n7673 avss.n7659 0.306507
R21375 avss.n7684 avss.n7683 0.306507
R21376 avss.n7789 avss.n7788 0.306507
R21377 avss.n7809 avss.n7808 0.306507
R21378 avss.n7836 avss.n7835 0.306507
R21379 avss.n7873 avss.n7872 0.306507
R21380 avss.n7884 avss.n7883 0.306507
R21381 avss.n7411 avss.n7410 0.306507
R21382 avss.n7402 avss.n7401 0.306507
R21383 avss.n7388 avss.n7387 0.306507
R21384 avss.n7320 avss.n7306 0.306507
R21385 avss.n7331 avss.n7330 0.306507
R21386 avss.n7436 avss.n7435 0.306507
R21387 avss.n7456 avss.n7455 0.306507
R21388 avss.n7483 avss.n7482 0.306507
R21389 avss.n7520 avss.n7519 0.306507
R21390 avss.n7531 avss.n7530 0.306507
R21391 avss.n7058 avss.n7057 0.306507
R21392 avss.n7049 avss.n7048 0.306507
R21393 avss.n7035 avss.n7034 0.306507
R21394 avss.n6967 avss.n6953 0.306507
R21395 avss.n6978 avss.n6977 0.306507
R21396 avss.n7083 avss.n7082 0.306507
R21397 avss.n7103 avss.n7102 0.306507
R21398 avss.n7130 avss.n7129 0.306507
R21399 avss.n7167 avss.n7166 0.306507
R21400 avss.n7178 avss.n7177 0.306507
R21401 avss.n6705 avss.n6704 0.306507
R21402 avss.n6696 avss.n6695 0.306507
R21403 avss.n6682 avss.n6681 0.306507
R21404 avss.n6614 avss.n6600 0.306507
R21405 avss.n6625 avss.n6624 0.306507
R21406 avss.n6730 avss.n6729 0.306507
R21407 avss.n6750 avss.n6749 0.306507
R21408 avss.n6777 avss.n6776 0.306507
R21409 avss.n6814 avss.n6813 0.306507
R21410 avss.n6825 avss.n6824 0.306507
R21411 avss.n6352 avss.n6351 0.306507
R21412 avss.n6343 avss.n6342 0.306507
R21413 avss.n6329 avss.n6328 0.306507
R21414 avss.n6261 avss.n6247 0.306507
R21415 avss.n6272 avss.n6271 0.306507
R21416 avss.n6377 avss.n6376 0.306507
R21417 avss.n6397 avss.n6396 0.306507
R21418 avss.n6424 avss.n6423 0.306507
R21419 avss.n6461 avss.n6460 0.306507
R21420 avss.n6472 avss.n6471 0.306507
R21421 avss.n5999 avss.n5998 0.306507
R21422 avss.n5990 avss.n5989 0.306507
R21423 avss.n5976 avss.n5975 0.306507
R21424 avss.n5908 avss.n5894 0.306507
R21425 avss.n5919 avss.n5918 0.306507
R21426 avss.n6024 avss.n6023 0.306507
R21427 avss.n6044 avss.n6043 0.306507
R21428 avss.n6071 avss.n6070 0.306507
R21429 avss.n6108 avss.n6107 0.306507
R21430 avss.n6119 avss.n6118 0.306507
R21431 avss.n5646 avss.n5645 0.306507
R21432 avss.n5637 avss.n5636 0.306507
R21433 avss.n5623 avss.n5622 0.306507
R21434 avss.n5555 avss.n5541 0.306507
R21435 avss.n5566 avss.n5565 0.306507
R21436 avss.n5671 avss.n5670 0.306507
R21437 avss.n5691 avss.n5690 0.306507
R21438 avss.n5718 avss.n5717 0.306507
R21439 avss.n5755 avss.n5754 0.306507
R21440 avss.n5766 avss.n5765 0.306507
R21441 avss.n5131 avss.n5130 0.306507
R21442 avss.n5292 avss.n5291 0.306507
R21443 avss.n5278 avss.n5277 0.306507
R21444 avss.n5215 avss.n5195 0.306507
R21445 avss.n5226 avss.n5225 0.306507
R21446 avss.n5318 avss.n5317 0.306507
R21447 avss.n5338 avss.n5337 0.306507
R21448 avss.n5365 avss.n5364 0.306507
R21449 avss.n5402 avss.n5401 0.306507
R21450 avss.n5413 avss.n5412 0.306507
R21451 avss.n4777 avss.n4776 0.306507
R21452 avss.n4938 avss.n4937 0.306507
R21453 avss.n4924 avss.n4923 0.306507
R21454 avss.n4861 avss.n4841 0.306507
R21455 avss.n4872 avss.n4871 0.306507
R21456 avss.n4964 avss.n4963 0.306507
R21457 avss.n4984 avss.n4983 0.306507
R21458 avss.n5011 avss.n5010 0.306507
R21459 avss.n5048 avss.n5047 0.306507
R21460 avss.n5059 avss.n5058 0.306507
R21461 avss.n8678 avss.n8677 0.283697
R21462 avss.n8869 avss.n3705 0.283697
R21463 avss.n8325 avss.n8324 0.283697
R21464 avss.n8516 avss.n3789 0.283697
R21465 avss.n7972 avss.n7971 0.283697
R21466 avss.n8163 avss.n3873 0.283697
R21467 avss.n7619 avss.n7618 0.283697
R21468 avss.n7810 avss.n3957 0.283697
R21469 avss.n7266 avss.n7265 0.283697
R21470 avss.n7457 avss.n4041 0.283697
R21471 avss.n6913 avss.n6912 0.283697
R21472 avss.n7104 avss.n4125 0.283697
R21473 avss.n6560 avss.n6559 0.283697
R21474 avss.n6751 avss.n4209 0.283697
R21475 avss.n6207 avss.n6206 0.283697
R21476 avss.n6398 avss.n4293 0.283697
R21477 avss.n5854 avss.n5853 0.283697
R21478 avss.n6045 avss.n4377 0.283697
R21479 avss.n5501 avss.n5500 0.283697
R21480 avss.n5692 avss.n4461 0.283697
R21481 avss.n5155 avss.n5154 0.283697
R21482 avss.n5339 avss.n4545 0.283697
R21483 avss.n4801 avss.n4800 0.283697
R21484 avss.n4985 avss.n4629 0.283697
R21485 avss.n8763 avss.n8762 0.266652
R21486 avss.n8952 avss.n8951 0.266652
R21487 avss.n8410 avss.n8409 0.266652
R21488 avss.n8599 avss.n8598 0.266652
R21489 avss.n8057 avss.n8056 0.266652
R21490 avss.n8246 avss.n8245 0.266652
R21491 avss.n7704 avss.n7703 0.266652
R21492 avss.n7893 avss.n7892 0.266652
R21493 avss.n7351 avss.n7350 0.266652
R21494 avss.n7540 avss.n7539 0.266652
R21495 avss.n6998 avss.n6997 0.266652
R21496 avss.n7187 avss.n7186 0.266652
R21497 avss.n6645 avss.n6644 0.266652
R21498 avss.n6834 avss.n6833 0.266652
R21499 avss.n6292 avss.n6291 0.266652
R21500 avss.n6481 avss.n6480 0.266652
R21501 avss.n5939 avss.n5938 0.266652
R21502 avss.n6128 avss.n6127 0.266652
R21503 avss.n5586 avss.n5585 0.266652
R21504 avss.n5775 avss.n5774 0.266652
R21505 avss.n5245 avss.n5244 0.266652
R21506 avss.n5422 avss.n5421 0.266652
R21507 avss.n4891 avss.n4890 0.266652
R21508 avss.n5068 avss.n5067 0.266652
R21509 avss.n9106 avss.n9105 0.266652
R21510 avss.n8994 avss.n8993 0.266652
R21511 avss.n9327 avss.n9326 0.266652
R21512 avss.n9215 avss.n9214 0.266652
R21513 avss.n9548 avss.n9547 0.266652
R21514 avss.n9436 avss.n9435 0.266652
R21515 avss.n9769 avss.n9768 0.266652
R21516 avss.n9657 avss.n9656 0.266652
R21517 avss.n9990 avss.n9989 0.266652
R21518 avss.n9878 avss.n9877 0.266652
R21519 avss.n10211 avss.n10210 0.266652
R21520 avss.n10099 avss.n10098 0.266652
R21521 avss.n10432 avss.n10431 0.266652
R21522 avss.n10320 avss.n10319 0.266652
R21523 avss.n10653 avss.n10652 0.266652
R21524 avss.n10541 avss.n10540 0.266652
R21525 avss.n10874 avss.n10873 0.266652
R21526 avss.n10762 avss.n10761 0.266652
R21527 avss.n11095 avss.n11094 0.266652
R21528 avss.n10983 avss.n10982 0.266652
R21529 avss.n361 avss.n360 0.266652
R21530 avss.n11204 avss.n11203 0.266652
R21531 avss.n144 avss.n143 0.266652
R21532 avss.n11425 avss.n11424 0.266652
R21533 avss.n3017 avss.n2945 0.263514
R21534 avss.n3070 avss.n2929 0.263514
R21535 avss.n3099 avss.n3098 0.263514
R21536 avss.n3666 avss.n2595 0.263514
R21537 avss.n2729 avss.n2658 0.263514
R21538 avss.n2774 avss.n2631 0.263514
R21539 avss.n2873 avss.n2872 0.263514
R21540 avss.n2833 avss.n2832 0.263514
R21541 avss.n2682 avss.n2675 0.260881
R21542 avss.n2655 avss.n2648 0.260881
R21543 avss.n2628 avss.n2625 0.260881
R21544 avss.n2807 avss.n2796 0.260881
R21545 avss.n3138 avss.n2919 0.260872
R21546 avss.n2965 avss.n2964 0.260872
R21547 avss.n3022 avss.n3021 0.260872
R21548 avss.n2613 avss.n2612 0.260872
R21549 avss.n3408 avss.n3407 0.240083
R21550 avss.n3437 avss.n3434 0.240083
R21551 avss.n3469 avss.n3466 0.240083
R21552 avss.t66 avss.n3247 0.233661
R21553 avss.n8773 avss.n3668 0.210867
R21554 avss.n8836 avss.n8835 0.210867
R21555 avss.n8972 avss.n8971 0.210867
R21556 avss.n8839 avss.n8837 0.210867
R21557 avss.n8420 avss.n3752 0.210867
R21558 avss.n8483 avss.n8482 0.210867
R21559 avss.n8619 avss.n8618 0.210867
R21560 avss.n8486 avss.n8484 0.210867
R21561 avss.n8067 avss.n3836 0.210867
R21562 avss.n8130 avss.n8129 0.210867
R21563 avss.n8266 avss.n8265 0.210867
R21564 avss.n8133 avss.n8131 0.210867
R21565 avss.n7714 avss.n3920 0.210867
R21566 avss.n7777 avss.n7776 0.210867
R21567 avss.n7913 avss.n7912 0.210867
R21568 avss.n7780 avss.n7778 0.210867
R21569 avss.n7361 avss.n4004 0.210867
R21570 avss.n7424 avss.n7423 0.210867
R21571 avss.n7560 avss.n7559 0.210867
R21572 avss.n7427 avss.n7425 0.210867
R21573 avss.n7008 avss.n4088 0.210867
R21574 avss.n7071 avss.n7070 0.210867
R21575 avss.n7207 avss.n7206 0.210867
R21576 avss.n7074 avss.n7072 0.210867
R21577 avss.n6655 avss.n4172 0.210867
R21578 avss.n6718 avss.n6717 0.210867
R21579 avss.n6854 avss.n6853 0.210867
R21580 avss.n6721 avss.n6719 0.210867
R21581 avss.n6302 avss.n4256 0.210867
R21582 avss.n6365 avss.n6364 0.210867
R21583 avss.n6501 avss.n6500 0.210867
R21584 avss.n6368 avss.n6366 0.210867
R21585 avss.n5949 avss.n4340 0.210867
R21586 avss.n6012 avss.n6011 0.210867
R21587 avss.n6148 avss.n6147 0.210867
R21588 avss.n6015 avss.n6013 0.210867
R21589 avss.n5596 avss.n4424 0.210867
R21590 avss.n5659 avss.n5658 0.210867
R21591 avss.n5795 avss.n5794 0.210867
R21592 avss.n5662 avss.n5660 0.210867
R21593 avss.n5306 avss.n5305 0.210867
R21594 avss.n5203 avss.n4508 0.210867
R21595 avss.n5442 avss.n5441 0.210867
R21596 avss.n5309 avss.n5307 0.210867
R21597 avss.n4952 avss.n4951 0.210867
R21598 avss.n4849 avss.n4592 0.210867
R21599 avss.n5088 avss.n5087 0.210867
R21600 avss.n4955 avss.n4953 0.210867
R21601 avss.n9193 avss.n9192 0.210867
R21602 avss.n9195 avss.n2485 0.210867
R21603 avss.n9084 avss.n9083 0.210867
R21604 avss.n9194 avss.n2593 0.210867
R21605 avss.n9414 avss.n9413 0.210867
R21606 avss.n9416 avss.n2269 0.210867
R21607 avss.n9305 avss.n9304 0.210867
R21608 avss.n9415 avss.n2377 0.210867
R21609 avss.n9635 avss.n9634 0.210867
R21610 avss.n9637 avss.n2053 0.210867
R21611 avss.n9526 avss.n9525 0.210867
R21612 avss.n9636 avss.n2161 0.210867
R21613 avss.n9856 avss.n9855 0.210867
R21614 avss.n9858 avss.n1837 0.210867
R21615 avss.n9747 avss.n9746 0.210867
R21616 avss.n9857 avss.n1945 0.210867
R21617 avss.n10077 avss.n10076 0.210867
R21618 avss.n10079 avss.n1621 0.210867
R21619 avss.n9968 avss.n9967 0.210867
R21620 avss.n10078 avss.n1729 0.210867
R21621 avss.n10298 avss.n10297 0.210867
R21622 avss.n10300 avss.n1405 0.210867
R21623 avss.n10189 avss.n10188 0.210867
R21624 avss.n10299 avss.n1513 0.210867
R21625 avss.n10519 avss.n10518 0.210867
R21626 avss.n10521 avss.n1189 0.210867
R21627 avss.n10410 avss.n10409 0.210867
R21628 avss.n10520 avss.n1297 0.210867
R21629 avss.n10740 avss.n10739 0.210867
R21630 avss.n10742 avss.n973 0.210867
R21631 avss.n10631 avss.n10630 0.210867
R21632 avss.n10741 avss.n1081 0.210867
R21633 avss.n10961 avss.n10960 0.210867
R21634 avss.n10963 avss.n757 0.210867
R21635 avss.n10852 avss.n10851 0.210867
R21636 avss.n10962 avss.n865 0.210867
R21637 avss.n11182 avss.n11181 0.210867
R21638 avss.n11184 avss.n541 0.210867
R21639 avss.n11073 avss.n11072 0.210867
R21640 avss.n11183 avss.n649 0.210867
R21641 avss.n11405 avss.n11404 0.210867
R21642 avss.n11295 avss.n433 0.210867
R21643 avss.n11294 avss.n11293 0.210867
R21644 avss.n11296 avss.n324 0.210867
R21645 avss.n11626 avss.n11625 0.210867
R21646 avss.n11516 avss.n216 0.210867
R21647 avss.n11515 avss.n11514 0.210867
R21648 avss.n11517 avss.n107 0.210867
R21649 avss.n2981 avss.n2979 0.209196
R21650 avss.n3038 avss.n3036 0.209196
R21651 avss.n3131 avss.n3130 0.209196
R21652 avss.n3630 avss.n3628 0.209196
R21653 avss.n2693 avss.n2691 0.209196
R21654 avss.n2738 avss.n2736 0.209196
R21655 avss.n2905 avss.n2775 0.209196
R21656 avss.n2865 avss.n2864 0.209196
R21657 avss.n2594 avss 0.195812
R21658 avss.n2830 avss 0.195812
R21659 avss.n3368 avss.n3366 0.185917
R21660 avss.n2681 avss.n2621 0.172761
R21661 avss.n2654 avss.n2653 0.172761
R21662 avss.n2916 avss.n2626 0.172761
R21663 avss.n2806 avss.n2805 0.172761
R21664 avss.n3619 avss.n3618 0.172761
R21665 avss.n3027 avss.n3026 0.172761
R21666 avss.n2966 avss.n2620 0.172761
R21667 avss.n3140 avss.n3139 0.172761
R21668 avss.n3249 avss.t187 0.165363
R21669 avss.n3437 avss.n3436 0.146333
R21670 avss.n4694 avss 0.142978
R21671 avss.n3453 avss.n3452 0.142167
R21672 avss avss.n3667 0.140087
R21673 avss.n2829 avss 0.140087
R21674 avss.n3381 avss.n3380 0.133833
R21675 avss.n3531 avss.n3530 0.129298
R21676 avss.n3265 avss.n3264 0.129298
R21677 avss.n4729 avss.n4677 0.120292
R21678 avss.n4724 avss.n4723 0.120292
R21679 avss.n4721 avss.n4681 0.120292
R21680 avss.n4716 avss.n4715 0.120292
R21681 avss.n4713 avss.n4685 0.120292
R21682 avss.n4708 avss.n4707 0.120292
R21683 avss.n4705 avss.n4689 0.120292
R21684 avss.n4700 avss.n4699 0.120292
R21685 avss.n4697 avss.n4693 0.120292
R21686 avss.n2987 avss.n2986 0.120292
R21687 avss.n2988 avss.n2987 0.120292
R21688 avss.n2988 avss.n2954 0.120292
R21689 avss.n2992 avss.n2954 0.120292
R21690 avss.n2994 avss.n2993 0.120292
R21691 avss.n2994 avss.n2951 0.120292
R21692 avss.n2998 avss.n2951 0.120292
R21693 avss.n2999 avss.n2998 0.120292
R21694 avss.n3000 avss.n2949 0.120292
R21695 avss.n3005 avss.n2949 0.120292
R21696 avss.n3006 avss.n3005 0.120292
R21697 avss.n3007 avss.n3006 0.120292
R21698 avss.n3007 avss.n2946 0.120292
R21699 avss.n3015 avss.n2946 0.120292
R21700 avss.n3016 avss.n3015 0.120292
R21701 avss.n3044 avss.n3043 0.120292
R21702 avss.n3045 avss.n3044 0.120292
R21703 avss.n3045 avss.n2938 0.120292
R21704 avss.n3049 avss.n2938 0.120292
R21705 avss.n3051 avss.n3050 0.120292
R21706 avss.n3051 avss.n2935 0.120292
R21707 avss.n3055 avss.n2935 0.120292
R21708 avss.n3056 avss.n3055 0.120292
R21709 avss.n3057 avss.n2933 0.120292
R21710 avss.n3062 avss.n2933 0.120292
R21711 avss.n3063 avss.n3062 0.120292
R21712 avss.n3064 avss.n3063 0.120292
R21713 avss.n3064 avss.n2930 0.120292
R21714 avss.n3073 avss.n2930 0.120292
R21715 avss.n3074 avss.n3073 0.120292
R21716 avss.n3124 avss.n3080 0.120292
R21717 avss.n3124 avss.n3123 0.120292
R21718 avss.n3123 avss.n3122 0.120292
R21719 avss.n3122 avss.n3083 0.120292
R21720 avss.n3117 avss.n3084 0.120292
R21721 avss.n3117 avss.n3116 0.120292
R21722 avss.n3116 avss.n3115 0.120292
R21723 avss.n3115 avss.n3087 0.120292
R21724 avss.n3111 avss.n3110 0.120292
R21725 avss.n3110 avss.n3089 0.120292
R21726 avss.n3106 avss.n3089 0.120292
R21727 avss.n3106 avss.n3105 0.120292
R21728 avss.n3105 avss.n3104 0.120292
R21729 avss.n3104 avss.n3091 0.120292
R21730 avss.n3097 avss.n3091 0.120292
R21731 avss.n3636 avss.n3635 0.120292
R21732 avss.n3637 avss.n3636 0.120292
R21733 avss.n3637 avss.n2604 0.120292
R21734 avss.n3641 avss.n2604 0.120292
R21735 avss.n3643 avss.n3642 0.120292
R21736 avss.n3643 avss.n2601 0.120292
R21737 avss.n3647 avss.n2601 0.120292
R21738 avss.n3648 avss.n3647 0.120292
R21739 avss.n3649 avss.n2599 0.120292
R21740 avss.n3654 avss.n2599 0.120292
R21741 avss.n3655 avss.n3654 0.120292
R21742 avss.n3656 avss.n3655 0.120292
R21743 avss.n3656 avss.n2596 0.120292
R21744 avss.n3664 avss.n2596 0.120292
R21745 avss.n3665 avss.n3664 0.120292
R21746 avss.n2699 avss.n2698 0.120292
R21747 avss.n2700 avss.n2699 0.120292
R21748 avss.n2700 avss.n2667 0.120292
R21749 avss.n2704 avss.n2667 0.120292
R21750 avss.n2706 avss.n2705 0.120292
R21751 avss.n2706 avss.n2664 0.120292
R21752 avss.n2710 avss.n2664 0.120292
R21753 avss.n2711 avss.n2710 0.120292
R21754 avss.n2712 avss.n2662 0.120292
R21755 avss.n2717 avss.n2662 0.120292
R21756 avss.n2718 avss.n2717 0.120292
R21757 avss.n2719 avss.n2718 0.120292
R21758 avss.n2719 avss.n2659 0.120292
R21759 avss.n2727 avss.n2659 0.120292
R21760 avss.n2728 avss.n2727 0.120292
R21761 avss.n2744 avss.n2743 0.120292
R21762 avss.n2745 avss.n2744 0.120292
R21763 avss.n2745 avss.n2640 0.120292
R21764 avss.n2749 avss.n2640 0.120292
R21765 avss.n2751 avss.n2750 0.120292
R21766 avss.n2751 avss.n2637 0.120292
R21767 avss.n2755 avss.n2637 0.120292
R21768 avss.n2756 avss.n2755 0.120292
R21769 avss.n2757 avss.n2635 0.120292
R21770 avss.n2762 avss.n2635 0.120292
R21771 avss.n2763 avss.n2762 0.120292
R21772 avss.n2764 avss.n2763 0.120292
R21773 avss.n2764 avss.n2632 0.120292
R21774 avss.n2772 avss.n2632 0.120292
R21775 avss.n2773 avss.n2772 0.120292
R21776 avss.n2898 avss.n2778 0.120292
R21777 avss.n2898 avss.n2897 0.120292
R21778 avss.n2897 avss.n2896 0.120292
R21779 avss.n2896 avss.n2781 0.120292
R21780 avss.n2891 avss.n2782 0.120292
R21781 avss.n2891 avss.n2890 0.120292
R21782 avss.n2890 avss.n2889 0.120292
R21783 avss.n2889 avss.n2785 0.120292
R21784 avss.n2885 avss.n2884 0.120292
R21785 avss.n2884 avss.n2787 0.120292
R21786 avss.n2880 avss.n2787 0.120292
R21787 avss.n2880 avss.n2879 0.120292
R21788 avss.n2879 avss.n2878 0.120292
R21789 avss.n2878 avss.n2789 0.120292
R21790 avss.n2871 avss.n2789 0.120292
R21791 avss.n2858 avss.n2814 0.120292
R21792 avss.n2858 avss.n2857 0.120292
R21793 avss.n2857 avss.n2856 0.120292
R21794 avss.n2856 avss.n2817 0.120292
R21795 avss.n2851 avss.n2818 0.120292
R21796 avss.n2851 avss.n2850 0.120292
R21797 avss.n2850 avss.n2849 0.120292
R21798 avss.n2849 avss.n2821 0.120292
R21799 avss.n2845 avss.n2844 0.120292
R21800 avss.n2844 avss.n2823 0.120292
R21801 avss.n2840 avss.n2823 0.120292
R21802 avss.n2840 avss.n2839 0.120292
R21803 avss.n2839 avss.n2838 0.120292
R21804 avss.n2838 avss.n2825 0.120292
R21805 avss.n2831 avss.n2825 0.120292
R21806 avss.n3597 avss.n3596 0.120292
R21807 avss.n3596 avss.n3541 0.120292
R21808 avss.n3591 avss.n3542 0.120292
R21809 avss.n3591 avss.n3590 0.120292
R21810 avss.n3589 avss.n3588 0.120292
R21811 avss.n3588 avss.n3545 0.120292
R21812 avss.n3583 avss.n3546 0.120292
R21813 avss.n3583 avss.n3582 0.120292
R21814 avss.n3581 avss.n3580 0.120292
R21815 avss.n3580 avss.n3549 0.120292
R21816 avss.n3575 avss.n3550 0.120292
R21817 avss.n3575 avss.n3574 0.120292
R21818 avss.n3573 avss.n3572 0.120292
R21819 avss.n3572 avss.n3553 0.120292
R21820 avss.n3567 avss.n3554 0.120292
R21821 avss.n3567 avss.n3566 0.120292
R21822 avss.n3565 avss.n3564 0.120292
R21823 avss.n3564 avss.n3557 0.120292
R21824 avss.n2983 avss.n2982 0.116385
R21825 avss.n3040 avss.n3039 0.116385
R21826 avss.n3129 avss.n3128 0.116385
R21827 avss.n3632 avss.n3631 0.116385
R21828 avss.n2695 avss.n2694 0.116385
R21829 avss.n2740 avss.n2739 0.116385
R21830 avss.n2903 avss.n2902 0.116385
R21831 avss.n2863 avss.n2862 0.116385
R21832 avss.n2974 avss 0.114786
R21833 avss.n3031 avss 0.114786
R21834 avss.n3136 avss 0.114786
R21835 avss.n3623 avss 0.114786
R21836 avss.n3378 avss.n3278 0.110917
R21837 avss.n3413 avss.n3412 0.110917
R21838 avss.n4731 avss 0.0994583
R21839 avss avss.n4729 0.0981562
R21840 avss avss.n4724 0.0981562
R21841 avss avss.n4721 0.0981562
R21842 avss avss.n4716 0.0981562
R21843 avss avss.n4713 0.0981562
R21844 avss avss.n4708 0.0981562
R21845 avss avss.n4705 0.0981562
R21846 avss avss.n4700 0.0981562
R21847 avss avss.n4697 0.0981562
R21848 avss.n3467 avss.n3173 0.09425
R21849 avss.n3598 avss 0.0929479
R21850 avss.n3392 avss.n3272 0.0864375
R21851 avss.n2925 avss.n2919 0.0861452
R21852 avss.n2972 avss.n2965 0.0861452
R21853 avss.n3029 avss.n3022 0.0861452
R21854 avss.n3621 avss.n2613 0.0861452
R21855 avss.n3466 avss.n3465 0.0859167
R21856 avss.n2796 avss.n2795 0.0856819
R21857 avss.n2914 avss.n2625 0.0856819
R21858 avss.n2648 avss.n2647 0.0856819
R21859 avss.n2675 avss.n2674 0.0856819
R21860 avss.n3395 avss.n3242 0.0838333
R21861 avss.n8824 avss.n8646 0.082192
R21862 avss.n8822 avss.n8648 0.082192
R21863 avss.n8813 avss.n8660 0.082192
R21864 avss.n8801 avss.n8800 0.082192
R21865 avss.n8791 avss.n8681 0.082192
R21866 avss.n8790 avss.n8705 0.082192
R21867 avss.n8732 avss.n8729 0.082192
R21868 avss.n8746 avss.n8743 0.082192
R21869 avss.n3746 avss.n3720 0.082192
R21870 avss.n8848 avss.n3713 0.082192
R21871 avss.n8870 avss.n8868 0.082192
R21872 avss.n8894 avss.n3699 0.082192
R21873 avss.n8914 avss.n3692 0.082192
R21874 avss.n8915 avss.n3685 0.082192
R21875 avss.n8932 avss.n3683 0.082192
R21876 avss.n8943 avss.n3682 0.082192
R21877 avss.n8471 avss.n8293 0.082192
R21878 avss.n8469 avss.n8295 0.082192
R21879 avss.n8460 avss.n8307 0.082192
R21880 avss.n8448 avss.n8447 0.082192
R21881 avss.n8438 avss.n8328 0.082192
R21882 avss.n8437 avss.n8352 0.082192
R21883 avss.n8379 avss.n8376 0.082192
R21884 avss.n8393 avss.n8390 0.082192
R21885 avss.n3830 avss.n3804 0.082192
R21886 avss.n8495 avss.n3797 0.082192
R21887 avss.n8517 avss.n8515 0.082192
R21888 avss.n8541 avss.n3783 0.082192
R21889 avss.n8561 avss.n3776 0.082192
R21890 avss.n8562 avss.n3769 0.082192
R21891 avss.n8579 avss.n3767 0.082192
R21892 avss.n8590 avss.n3766 0.082192
R21893 avss.n8118 avss.n7940 0.082192
R21894 avss.n8116 avss.n7942 0.082192
R21895 avss.n8107 avss.n7954 0.082192
R21896 avss.n8095 avss.n8094 0.082192
R21897 avss.n8085 avss.n7975 0.082192
R21898 avss.n8084 avss.n7999 0.082192
R21899 avss.n8026 avss.n8023 0.082192
R21900 avss.n8040 avss.n8037 0.082192
R21901 avss.n3914 avss.n3888 0.082192
R21902 avss.n8142 avss.n3881 0.082192
R21903 avss.n8164 avss.n8162 0.082192
R21904 avss.n8188 avss.n3867 0.082192
R21905 avss.n8208 avss.n3860 0.082192
R21906 avss.n8209 avss.n3853 0.082192
R21907 avss.n8226 avss.n3851 0.082192
R21908 avss.n8237 avss.n3850 0.082192
R21909 avss.n7765 avss.n7587 0.082192
R21910 avss.n7763 avss.n7589 0.082192
R21911 avss.n7754 avss.n7601 0.082192
R21912 avss.n7742 avss.n7741 0.082192
R21913 avss.n7732 avss.n7622 0.082192
R21914 avss.n7731 avss.n7646 0.082192
R21915 avss.n7673 avss.n7670 0.082192
R21916 avss.n7687 avss.n7684 0.082192
R21917 avss.n3998 avss.n3972 0.082192
R21918 avss.n7789 avss.n3965 0.082192
R21919 avss.n7811 avss.n7809 0.082192
R21920 avss.n7835 avss.n3951 0.082192
R21921 avss.n7855 avss.n3944 0.082192
R21922 avss.n7856 avss.n3937 0.082192
R21923 avss.n7873 avss.n3935 0.082192
R21924 avss.n7884 avss.n3934 0.082192
R21925 avss.n7412 avss.n7234 0.082192
R21926 avss.n7410 avss.n7236 0.082192
R21927 avss.n7401 avss.n7248 0.082192
R21928 avss.n7389 avss.n7388 0.082192
R21929 avss.n7379 avss.n7269 0.082192
R21930 avss.n7378 avss.n7293 0.082192
R21931 avss.n7320 avss.n7317 0.082192
R21932 avss.n7334 avss.n7331 0.082192
R21933 avss.n4082 avss.n4056 0.082192
R21934 avss.n7436 avss.n4049 0.082192
R21935 avss.n7458 avss.n7456 0.082192
R21936 avss.n7482 avss.n4035 0.082192
R21937 avss.n7502 avss.n4028 0.082192
R21938 avss.n7503 avss.n4021 0.082192
R21939 avss.n7520 avss.n4019 0.082192
R21940 avss.n7531 avss.n4018 0.082192
R21941 avss.n7059 avss.n6881 0.082192
R21942 avss.n7057 avss.n6883 0.082192
R21943 avss.n7048 avss.n6895 0.082192
R21944 avss.n7036 avss.n7035 0.082192
R21945 avss.n7026 avss.n6916 0.082192
R21946 avss.n7025 avss.n6940 0.082192
R21947 avss.n6967 avss.n6964 0.082192
R21948 avss.n6981 avss.n6978 0.082192
R21949 avss.n4166 avss.n4140 0.082192
R21950 avss.n7083 avss.n4133 0.082192
R21951 avss.n7105 avss.n7103 0.082192
R21952 avss.n7129 avss.n4119 0.082192
R21953 avss.n7149 avss.n4112 0.082192
R21954 avss.n7150 avss.n4105 0.082192
R21955 avss.n7167 avss.n4103 0.082192
R21956 avss.n7178 avss.n4102 0.082192
R21957 avss.n6706 avss.n6528 0.082192
R21958 avss.n6704 avss.n6530 0.082192
R21959 avss.n6695 avss.n6542 0.082192
R21960 avss.n6683 avss.n6682 0.082192
R21961 avss.n6673 avss.n6563 0.082192
R21962 avss.n6672 avss.n6587 0.082192
R21963 avss.n6614 avss.n6611 0.082192
R21964 avss.n6628 avss.n6625 0.082192
R21965 avss.n4250 avss.n4224 0.082192
R21966 avss.n6730 avss.n4217 0.082192
R21967 avss.n6752 avss.n6750 0.082192
R21968 avss.n6776 avss.n4203 0.082192
R21969 avss.n6796 avss.n4196 0.082192
R21970 avss.n6797 avss.n4189 0.082192
R21971 avss.n6814 avss.n4187 0.082192
R21972 avss.n6825 avss.n4186 0.082192
R21973 avss.n6353 avss.n6175 0.082192
R21974 avss.n6351 avss.n6177 0.082192
R21975 avss.n6342 avss.n6189 0.082192
R21976 avss.n6330 avss.n6329 0.082192
R21977 avss.n6320 avss.n6210 0.082192
R21978 avss.n6319 avss.n6234 0.082192
R21979 avss.n6261 avss.n6258 0.082192
R21980 avss.n6275 avss.n6272 0.082192
R21981 avss.n4334 avss.n4308 0.082192
R21982 avss.n6377 avss.n4301 0.082192
R21983 avss.n6399 avss.n6397 0.082192
R21984 avss.n6423 avss.n4287 0.082192
R21985 avss.n6443 avss.n4280 0.082192
R21986 avss.n6444 avss.n4273 0.082192
R21987 avss.n6461 avss.n4271 0.082192
R21988 avss.n6472 avss.n4270 0.082192
R21989 avss.n6000 avss.n5822 0.082192
R21990 avss.n5998 avss.n5824 0.082192
R21991 avss.n5989 avss.n5836 0.082192
R21992 avss.n5977 avss.n5976 0.082192
R21993 avss.n5967 avss.n5857 0.082192
R21994 avss.n5966 avss.n5881 0.082192
R21995 avss.n5908 avss.n5905 0.082192
R21996 avss.n5922 avss.n5919 0.082192
R21997 avss.n4418 avss.n4392 0.082192
R21998 avss.n6024 avss.n4385 0.082192
R21999 avss.n6046 avss.n6044 0.082192
R22000 avss.n6070 avss.n4371 0.082192
R22001 avss.n6090 avss.n4364 0.082192
R22002 avss.n6091 avss.n4357 0.082192
R22003 avss.n6108 avss.n4355 0.082192
R22004 avss.n6119 avss.n4354 0.082192
R22005 avss.n5647 avss.n5469 0.082192
R22006 avss.n5645 avss.n5471 0.082192
R22007 avss.n5636 avss.n5483 0.082192
R22008 avss.n5624 avss.n5623 0.082192
R22009 avss.n5614 avss.n5504 0.082192
R22010 avss.n5613 avss.n5528 0.082192
R22011 avss.n5555 avss.n5552 0.082192
R22012 avss.n5569 avss.n5566 0.082192
R22013 avss.n4502 avss.n4476 0.082192
R22014 avss.n5671 avss.n4469 0.082192
R22015 avss.n5693 avss.n5691 0.082192
R22016 avss.n5717 avss.n4455 0.082192
R22017 avss.n5737 avss.n4448 0.082192
R22018 avss.n5738 avss.n4441 0.082192
R22019 avss.n5755 avss.n4439 0.082192
R22020 avss.n5766 avss.n4438 0.082192
R22021 avss.n5122 avss.n5099 0.082192
R22022 avss.n5293 avss.n5131 0.082192
R22023 avss.n5291 avss.n5133 0.082192
R22024 avss.n5279 avss.n5278 0.082192
R22025 avss.n5269 avss.n5158 0.082192
R22026 avss.n5268 avss.n5182 0.082192
R22027 avss.n5215 avss.n5212 0.082192
R22028 avss.n5246 avss.n5226 0.082192
R22029 avss.n4586 avss.n4560 0.082192
R22030 avss.n5318 avss.n4553 0.082192
R22031 avss.n5340 avss.n5338 0.082192
R22032 avss.n5364 avss.n4539 0.082192
R22033 avss.n5384 avss.n4532 0.082192
R22034 avss.n5385 avss.n4525 0.082192
R22035 avss.n5402 avss.n4523 0.082192
R22036 avss.n5413 avss.n4522 0.082192
R22037 avss.n4768 avss.n4745 0.082192
R22038 avss.n4939 avss.n4777 0.082192
R22039 avss.n4937 avss.n4779 0.082192
R22040 avss.n4925 avss.n4924 0.082192
R22041 avss.n4915 avss.n4804 0.082192
R22042 avss.n4914 avss.n4828 0.082192
R22043 avss.n4861 avss.n4858 0.082192
R22044 avss.n4892 avss.n4872 0.082192
R22045 avss.n4670 avss.n4644 0.082192
R22046 avss.n4964 avss.n4637 0.082192
R22047 avss.n4986 avss.n4984 0.082192
R22048 avss.n5010 avss.n4623 0.082192
R22049 avss.n5030 avss.n4616 0.082192
R22050 avss.n5031 avss.n4609 0.082192
R22051 avss.n5048 avss.n4607 0.082192
R22052 avss.n5059 avss.n4606 0.082192
R22053 avss.n2400 avss.n2399 0.082192
R22054 avss.n2470 avss.n2469 0.082192
R22055 avss.n2451 avss.n2450 0.082192
R22056 avss.n2438 avss.n2437 0.082192
R22057 avss.n9128 avss.n9127 0.082192
R22058 avss.n9143 avss.n9142 0.082192
R22059 avss.n9162 avss.n9161 0.082192
R22060 avss.n9108 avss.n9107 0.082192
R22061 avss.n2547 avss.n2546 0.082192
R22062 avss.n2527 avss.n2526 0.082192
R22063 avss.n2508 avss.n2507 0.082192
R22064 avss.n2495 avss.n2494 0.082192
R22065 avss.n9017 avss.n9016 0.082192
R22066 avss.n9032 avss.n9031 0.082192
R22067 avss.n9051 avss.n9050 0.082192
R22068 avss.n8996 avss.n8995 0.082192
R22069 avss.n2184 avss.n2183 0.082192
R22070 avss.n2254 avss.n2253 0.082192
R22071 avss.n2235 avss.n2234 0.082192
R22072 avss.n2222 avss.n2221 0.082192
R22073 avss.n9349 avss.n9348 0.082192
R22074 avss.n9364 avss.n9363 0.082192
R22075 avss.n9383 avss.n9382 0.082192
R22076 avss.n9329 avss.n9328 0.082192
R22077 avss.n2331 avss.n2330 0.082192
R22078 avss.n2311 avss.n2310 0.082192
R22079 avss.n2292 avss.n2291 0.082192
R22080 avss.n2279 avss.n2278 0.082192
R22081 avss.n9238 avss.n9237 0.082192
R22082 avss.n9253 avss.n9252 0.082192
R22083 avss.n9272 avss.n9271 0.082192
R22084 avss.n9217 avss.n9216 0.082192
R22085 avss.n1968 avss.n1967 0.082192
R22086 avss.n2038 avss.n2037 0.082192
R22087 avss.n2019 avss.n2018 0.082192
R22088 avss.n2006 avss.n2005 0.082192
R22089 avss.n9570 avss.n9569 0.082192
R22090 avss.n9585 avss.n9584 0.082192
R22091 avss.n9604 avss.n9603 0.082192
R22092 avss.n9550 avss.n9549 0.082192
R22093 avss.n2115 avss.n2114 0.082192
R22094 avss.n2095 avss.n2094 0.082192
R22095 avss.n2076 avss.n2075 0.082192
R22096 avss.n2063 avss.n2062 0.082192
R22097 avss.n9459 avss.n9458 0.082192
R22098 avss.n9474 avss.n9473 0.082192
R22099 avss.n9493 avss.n9492 0.082192
R22100 avss.n9438 avss.n9437 0.082192
R22101 avss.n1752 avss.n1751 0.082192
R22102 avss.n1822 avss.n1821 0.082192
R22103 avss.n1803 avss.n1802 0.082192
R22104 avss.n1790 avss.n1789 0.082192
R22105 avss.n9791 avss.n9790 0.082192
R22106 avss.n9806 avss.n9805 0.082192
R22107 avss.n9825 avss.n9824 0.082192
R22108 avss.n9771 avss.n9770 0.082192
R22109 avss.n1899 avss.n1898 0.082192
R22110 avss.n1879 avss.n1878 0.082192
R22111 avss.n1860 avss.n1859 0.082192
R22112 avss.n1847 avss.n1846 0.082192
R22113 avss.n9680 avss.n9679 0.082192
R22114 avss.n9695 avss.n9694 0.082192
R22115 avss.n9714 avss.n9713 0.082192
R22116 avss.n9659 avss.n9658 0.082192
R22117 avss.n1536 avss.n1535 0.082192
R22118 avss.n1606 avss.n1605 0.082192
R22119 avss.n1587 avss.n1586 0.082192
R22120 avss.n1574 avss.n1573 0.082192
R22121 avss.n10012 avss.n10011 0.082192
R22122 avss.n10027 avss.n10026 0.082192
R22123 avss.n10046 avss.n10045 0.082192
R22124 avss.n9992 avss.n9991 0.082192
R22125 avss.n1683 avss.n1682 0.082192
R22126 avss.n1663 avss.n1662 0.082192
R22127 avss.n1644 avss.n1643 0.082192
R22128 avss.n1631 avss.n1630 0.082192
R22129 avss.n9901 avss.n9900 0.082192
R22130 avss.n9916 avss.n9915 0.082192
R22131 avss.n9935 avss.n9934 0.082192
R22132 avss.n9880 avss.n9879 0.082192
R22133 avss.n1320 avss.n1319 0.082192
R22134 avss.n1390 avss.n1389 0.082192
R22135 avss.n1371 avss.n1370 0.082192
R22136 avss.n1358 avss.n1357 0.082192
R22137 avss.n10233 avss.n10232 0.082192
R22138 avss.n10248 avss.n10247 0.082192
R22139 avss.n10267 avss.n10266 0.082192
R22140 avss.n10213 avss.n10212 0.082192
R22141 avss.n1467 avss.n1466 0.082192
R22142 avss.n1447 avss.n1446 0.082192
R22143 avss.n1428 avss.n1427 0.082192
R22144 avss.n1415 avss.n1414 0.082192
R22145 avss.n10122 avss.n10121 0.082192
R22146 avss.n10137 avss.n10136 0.082192
R22147 avss.n10156 avss.n10155 0.082192
R22148 avss.n10101 avss.n10100 0.082192
R22149 avss.n1104 avss.n1103 0.082192
R22150 avss.n1174 avss.n1173 0.082192
R22151 avss.n1155 avss.n1154 0.082192
R22152 avss.n1142 avss.n1141 0.082192
R22153 avss.n10454 avss.n10453 0.082192
R22154 avss.n10469 avss.n10468 0.082192
R22155 avss.n10488 avss.n10487 0.082192
R22156 avss.n10434 avss.n10433 0.082192
R22157 avss.n1251 avss.n1250 0.082192
R22158 avss.n1231 avss.n1230 0.082192
R22159 avss.n1212 avss.n1211 0.082192
R22160 avss.n1199 avss.n1198 0.082192
R22161 avss.n10343 avss.n10342 0.082192
R22162 avss.n10358 avss.n10357 0.082192
R22163 avss.n10377 avss.n10376 0.082192
R22164 avss.n10322 avss.n10321 0.082192
R22165 avss.n888 avss.n887 0.082192
R22166 avss.n958 avss.n957 0.082192
R22167 avss.n939 avss.n938 0.082192
R22168 avss.n926 avss.n925 0.082192
R22169 avss.n10675 avss.n10674 0.082192
R22170 avss.n10690 avss.n10689 0.082192
R22171 avss.n10709 avss.n10708 0.082192
R22172 avss.n10655 avss.n10654 0.082192
R22173 avss.n1035 avss.n1034 0.082192
R22174 avss.n1015 avss.n1014 0.082192
R22175 avss.n996 avss.n995 0.082192
R22176 avss.n983 avss.n982 0.082192
R22177 avss.n10564 avss.n10563 0.082192
R22178 avss.n10579 avss.n10578 0.082192
R22179 avss.n10598 avss.n10597 0.082192
R22180 avss.n10543 avss.n10542 0.082192
R22181 avss.n672 avss.n671 0.082192
R22182 avss.n742 avss.n741 0.082192
R22183 avss.n723 avss.n722 0.082192
R22184 avss.n710 avss.n709 0.082192
R22185 avss.n10896 avss.n10895 0.082192
R22186 avss.n10911 avss.n10910 0.082192
R22187 avss.n10930 avss.n10929 0.082192
R22188 avss.n10876 avss.n10875 0.082192
R22189 avss.n819 avss.n818 0.082192
R22190 avss.n799 avss.n798 0.082192
R22191 avss.n780 avss.n779 0.082192
R22192 avss.n767 avss.n766 0.082192
R22193 avss.n10785 avss.n10784 0.082192
R22194 avss.n10800 avss.n10799 0.082192
R22195 avss.n10819 avss.n10818 0.082192
R22196 avss.n10764 avss.n10763 0.082192
R22197 avss.n456 avss.n455 0.082192
R22198 avss.n526 avss.n525 0.082192
R22199 avss.n507 avss.n506 0.082192
R22200 avss.n494 avss.n493 0.082192
R22201 avss.n11117 avss.n11116 0.082192
R22202 avss.n11132 avss.n11131 0.082192
R22203 avss.n11151 avss.n11150 0.082192
R22204 avss.n11097 avss.n11096 0.082192
R22205 avss.n603 avss.n602 0.082192
R22206 avss.n583 avss.n582 0.082192
R22207 avss.n564 avss.n563 0.082192
R22208 avss.n551 avss.n550 0.082192
R22209 avss.n11006 avss.n11005 0.082192
R22210 avss.n11021 avss.n11020 0.082192
R22211 avss.n11040 avss.n11039 0.082192
R22212 avss.n10985 avss.n10984 0.082192
R22213 avss.n11374 avss.n11373 0.082192
R22214 avss.n11355 avss.n11354 0.082192
R22215 avss.n11336 avss.n11335 0.082192
R22216 avss.n11323 avss.n11322 0.082192
R22217 avss.n384 avss.n383 0.082192
R22218 avss.n399 avss.n398 0.082192
R22219 avss.n418 avss.n417 0.082192
R22220 avss.n363 avss.n362 0.082192
R22221 avss.n278 avss.n277 0.082192
R22222 avss.n258 avss.n257 0.082192
R22223 avss.n239 avss.n238 0.082192
R22224 avss.n226 avss.n225 0.082192
R22225 avss.n11227 avss.n11226 0.082192
R22226 avss.n11242 avss.n11241 0.082192
R22227 avss.n11261 avss.n11260 0.082192
R22228 avss.n11206 avss.n11205 0.082192
R22229 avss.n11595 avss.n11594 0.082192
R22230 avss.n11576 avss.n11575 0.082192
R22231 avss.n11557 avss.n11556 0.082192
R22232 avss.n11544 avss.n11543 0.082192
R22233 avss.n167 avss.n166 0.082192
R22234 avss.n182 avss.n181 0.082192
R22235 avss.n201 avss.n200 0.082192
R22236 avss.n146 avss.n145 0.082192
R22237 avss.n61 avss.n60 0.082192
R22238 avss.n41 avss.n40 0.082192
R22239 avss.n22 avss.n21 0.082192
R22240 avss.n9 avss.n8 0.082192
R22241 avss.n11448 avss.n11447 0.082192
R22242 avss.n11463 avss.n11462 0.082192
R22243 avss.n11482 avss.n11481 0.082192
R22244 avss.n11427 avss.n11426 0.082192
R22245 avss.n4734 avss 0.0820789
R22246 avss.n3559 avss 0.0812292
R22247 avss.n3462 avss.n3196 0.078625
R22248 avss avss.n3293 0.0770625
R22249 avss.n3732 avss.n3725 0.072235
R22250 avss.n3816 avss.n3809 0.072235
R22251 avss.n3900 avss.n3893 0.072235
R22252 avss.n3984 avss.n3977 0.072235
R22253 avss.n4068 avss.n4061 0.072235
R22254 avss.n4152 avss.n4145 0.072235
R22255 avss.n4236 avss.n4229 0.072235
R22256 avss.n4320 avss.n4313 0.072235
R22257 avss.n4404 avss.n4397 0.072235
R22258 avss.n4488 avss.n4481 0.072235
R22259 avss.n4572 avss.n4565 0.072235
R22260 avss.n4656 avss.n4649 0.072235
R22261 avss.n2557 avss.n2556 0.072235
R22262 avss.n2341 avss.n2340 0.072235
R22263 avss.n2125 avss.n2124 0.072235
R22264 avss.n1909 avss.n1908 0.072235
R22265 avss.n1693 avss.n1692 0.072235
R22266 avss.n1477 avss.n1476 0.072235
R22267 avss.n1261 avss.n1260 0.072235
R22268 avss.n1045 avss.n1044 0.072235
R22269 avss.n829 avss.n828 0.072235
R22270 avss.n613 avss.n612 0.072235
R22271 avss.n288 avss.n287 0.072235
R22272 avss.n71 avss.n70 0.072235
R22273 avss avss.n3559 0.0721146
R22274 avss.n8833 avss.n8623 0.0715211
R22275 avss.n8480 avss.n8270 0.0715211
R22276 avss.n8127 avss.n7917 0.0715211
R22277 avss.n7774 avss.n7564 0.0715211
R22278 avss.n7421 avss.n7211 0.0715211
R22279 avss.n7068 avss.n6858 0.0715211
R22280 avss.n6715 avss.n6505 0.0715211
R22281 avss.n6362 avss.n6152 0.0715211
R22282 avss.n6009 avss.n5799 0.0715211
R22283 avss.n5656 avss.n5446 0.0715211
R22284 avss.n2482 avss.n2481 0.0715211
R22285 avss.n2266 avss.n2265 0.0715211
R22286 avss.n2050 avss.n2049 0.0715211
R22287 avss.n1834 avss.n1833 0.0715211
R22288 avss.n1618 avss.n1617 0.0715211
R22289 avss.n1402 avss.n1401 0.0715211
R22290 avss.n1186 avss.n1185 0.0715211
R22291 avss.n970 avss.n969 0.0715211
R22292 avss.n754 avss.n753 0.0715211
R22293 avss.n538 avss.n537 0.0715211
R22294 avss.n2963 avss.n2962 0.0713089
R22295 avss.n3020 avss.n3019 0.0713089
R22296 avss.n3075 avss.n2927 0.0713089
R22297 avss.n3096 avss.n2611 0.0713089
R22298 avss.n4694 avss 0.0696335
R22299 avss.n2687 avss.n2686 0.0682083
R22300 avss.n2732 avss.n2731 0.0682083
R22301 avss.n2910 avss.n2909 0.0682083
R22302 avss.n2870 avss.n2869 0.0682083
R22303 avss.n3533 avss.n3532 0.0681222
R22304 avss.n3255 avss.n3250 0.0681222
R22305 avss.n2678 avss.n2677 0.067449
R22306 avss.n2651 avss.n2624 0.067449
R22307 avss.n2800 avss.n2627 0.067449
R22308 avss.n2803 avss.n2616 0.067449
R22309 avss.n3615 avss.n2614 0.067449
R22310 avss.n3023 avss.n2918 0.067449
R22311 avss.n2970 avss.n2969 0.067449
R22312 avss.n2922 avss.n2921 0.067449
R22313 avss.n3337 avss.n3336 0.0671667
R22314 avss.n3380 avss.n3273 0.0671667
R22315 avss.n3454 avss.n3453 0.063
R22316 avss.n8632 avss.n8626 0.0620866
R22317 avss.n8279 avss.n8273 0.0620866
R22318 avss.n7926 avss.n7920 0.0620866
R22319 avss.n7573 avss.n7567 0.0620866
R22320 avss.n7220 avss.n7214 0.0620866
R22321 avss.n6867 avss.n6861 0.0620866
R22322 avss.n6514 avss.n6508 0.0620866
R22323 avss.n6161 avss.n6155 0.0620866
R22324 avss.n5808 avss.n5802 0.0620866
R22325 avss.n5455 avss.n5449 0.0620866
R22326 avss.n5107 avss.n5106 0.0620866
R22327 avss.n4753 avss.n4752 0.0620866
R22328 avss.n2410 avss.n2409 0.0620866
R22329 avss.n2194 avss.n2193 0.0620866
R22330 avss.n1978 avss.n1977 0.0620866
R22331 avss.n1762 avss.n1761 0.0620866
R22332 avss.n1546 avss.n1545 0.0620866
R22333 avss.n1330 avss.n1329 0.0620866
R22334 avss.n1114 avss.n1113 0.0620866
R22335 avss.n898 avss.n897 0.0620866
R22336 avss.n682 avss.n681 0.0620866
R22337 avss.n466 avss.n465 0.0620866
R22338 avss.n11385 avss.n11384 0.0620866
R22339 avss.n11606 avss.n11605 0.0620866
R22340 avss.n2974 avss 0.0612143
R22341 avss.n3031 avss 0.0612143
R22342 avss avss.n3136 0.0612143
R22343 avss.n3623 avss 0.0612143
R22344 avss.n8841 avss.n3727 0.061128
R22345 avss.n8488 avss.n3811 0.061128
R22346 avss.n8135 avss.n3895 0.061128
R22347 avss.n7782 avss.n3979 0.061128
R22348 avss.n7429 avss.n4063 0.061128
R22349 avss.n7076 avss.n4147 0.061128
R22350 avss.n6723 avss.n4231 0.061128
R22351 avss.n6370 avss.n4315 0.061128
R22352 avss.n6017 avss.n4399 0.061128
R22353 avss.n5664 avss.n4483 0.061128
R22354 avss.n5302 avss.n5301 0.061128
R22355 avss.n5311 avss.n4567 0.061128
R22356 avss.n4948 avss.n4947 0.061128
R22357 avss.n4957 avss.n4651 0.061128
R22358 avss.n2539 avss.n2538 0.061128
R22359 avss.n2323 avss.n2322 0.061128
R22360 avss.n2107 avss.n2106 0.061128
R22361 avss.n1891 avss.n1890 0.061128
R22362 avss.n1675 avss.n1674 0.061128
R22363 avss.n1459 avss.n1458 0.061128
R22364 avss.n1243 avss.n1242 0.061128
R22365 avss.n1027 avss.n1026 0.061128
R22366 avss.n811 avss.n810 0.061128
R22367 avss.n595 avss.n594 0.061128
R22368 avss.n11367 avss.n11366 0.061128
R22369 avss.n270 avss.n269 0.061128
R22370 avss.n11588 avss.n11587 0.061128
R22371 avss.n53 avss.n52 0.061128
R22372 avss avss.n4677 0.0603958
R22373 avss.n4723 avss 0.0603958
R22374 avss avss.n4681 0.0603958
R22375 avss.n4715 avss 0.0603958
R22376 avss avss.n4714 0.0603958
R22377 avss avss.n4685 0.0603958
R22378 avss.n4707 avss 0.0603958
R22379 avss avss.n4689 0.0603958
R22380 avss.n4699 avss 0.0603958
R22381 avss avss.n4693 0.0603958
R22382 avss.n2962 avss 0.0603958
R22383 avss.n2986 avss 0.0603958
R22384 avss.n3019 avss 0.0603958
R22385 avss.n3043 avss 0.0603958
R22386 avss.n3075 avss 0.0603958
R22387 avss.n3080 avss 0.0603958
R22388 avss avss.n3096 0.0603958
R22389 avss.n3635 avss 0.0603958
R22390 avss.n2686 avss 0.0603958
R22391 avss.n2698 avss 0.0603958
R22392 avss.n2731 avss 0.0603958
R22393 avss.n2743 avss 0.0603958
R22394 avss.n2909 avss 0.0603958
R22395 avss.n2778 avss 0.0603958
R22396 avss avss.n2870 0.0603958
R22397 avss.n2814 avss 0.0603958
R22398 avss.n3598 avss 0.0603958
R22399 avss.n3550 avss 0.0603958
R22400 avss.n2808 avss.n2795 0.0598606
R22401 avss.n2914 avss.n2913 0.0598606
R22402 avss.n2656 avss.n2647 0.0598606
R22403 avss.n2683 avss.n2674 0.0598606
R22404 avss.n3622 avss.n3621 0.0593974
R22405 avss.n3030 avss.n3029 0.0593974
R22406 avss.n2973 avss.n2972 0.0593974
R22407 avss.n3137 avss.n2925 0.0593974
R22408 avss.n4734 avss.n4733 0.0591735
R22409 avss.n3558 avss 0.0591735
R22410 avss.n4725 avss 0.0590938
R22411 avss.n4717 avss 0.0590938
R22412 avss.n4709 avss 0.0590938
R22413 avss avss.n4706 0.0590938
R22414 avss avss.n4698 0.0590938
R22415 avss.n3542 avss 0.0590938
R22416 avss.n3546 avss 0.0590938
R22417 avss avss.n3581 0.0590938
R22418 avss avss.n3573 0.0590938
R22419 avss avss.n3565 0.0590938
R22420 avss.n11634 avss.n11627 0.0579556
R22421 avss avss.n4722 0.0577917
R22422 avss.n4701 avss 0.0577917
R22423 avss.n3000 avss 0.0577917
R22424 avss.n3057 avss 0.0577917
R22425 avss.n3111 avss 0.0577917
R22426 avss.n3649 avss 0.0577917
R22427 avss.n2712 avss 0.0577917
R22428 avss.n2757 avss 0.0577917
R22429 avss.n2885 avss 0.0577917
R22430 avss.n2845 avss 0.0577917
R22431 avss avss.n3589 0.0577917
R22432 avss.n3554 avss 0.0577917
R22433 avss.n8752 avss.n8722 0.0574697
R22434 avss.n8807 avss.n8669 0.0574697
R22435 avss.n8806 avss.n8805 0.0574697
R22436 avss.n8749 avss.n8745 0.0574697
R22437 avss.n8876 avss.n3703 0.0574697
R22438 avss.n8967 avss.n3679 0.0574697
R22439 avss.n8878 avss.n8877 0.0574697
R22440 avss.n8966 avss.n8965 0.0574697
R22441 avss.n8399 avss.n8369 0.0574697
R22442 avss.n8454 avss.n8316 0.0574697
R22443 avss.n8453 avss.n8452 0.0574697
R22444 avss.n8396 avss.n8392 0.0574697
R22445 avss.n8523 avss.n3787 0.0574697
R22446 avss.n8614 avss.n3763 0.0574697
R22447 avss.n8525 avss.n8524 0.0574697
R22448 avss.n8613 avss.n8612 0.0574697
R22449 avss.n8046 avss.n8016 0.0574697
R22450 avss.n8101 avss.n7963 0.0574697
R22451 avss.n8100 avss.n8099 0.0574697
R22452 avss.n8043 avss.n8039 0.0574697
R22453 avss.n8170 avss.n3871 0.0574697
R22454 avss.n8261 avss.n3847 0.0574697
R22455 avss.n8172 avss.n8171 0.0574697
R22456 avss.n8260 avss.n8259 0.0574697
R22457 avss.n7693 avss.n7663 0.0574697
R22458 avss.n7748 avss.n7610 0.0574697
R22459 avss.n7747 avss.n7746 0.0574697
R22460 avss.n7690 avss.n7686 0.0574697
R22461 avss.n7817 avss.n3955 0.0574697
R22462 avss.n7908 avss.n3931 0.0574697
R22463 avss.n7819 avss.n7818 0.0574697
R22464 avss.n7907 avss.n7906 0.0574697
R22465 avss.n7340 avss.n7310 0.0574697
R22466 avss.n7395 avss.n7257 0.0574697
R22467 avss.n7394 avss.n7393 0.0574697
R22468 avss.n7337 avss.n7333 0.0574697
R22469 avss.n7464 avss.n4039 0.0574697
R22470 avss.n7555 avss.n4015 0.0574697
R22471 avss.n7466 avss.n7465 0.0574697
R22472 avss.n7554 avss.n7553 0.0574697
R22473 avss.n6987 avss.n6957 0.0574697
R22474 avss.n7042 avss.n6904 0.0574697
R22475 avss.n7041 avss.n7040 0.0574697
R22476 avss.n6984 avss.n6980 0.0574697
R22477 avss.n7111 avss.n4123 0.0574697
R22478 avss.n7202 avss.n4099 0.0574697
R22479 avss.n7113 avss.n7112 0.0574697
R22480 avss.n7201 avss.n7200 0.0574697
R22481 avss.n6634 avss.n6604 0.0574697
R22482 avss.n6689 avss.n6551 0.0574697
R22483 avss.n6688 avss.n6687 0.0574697
R22484 avss.n6631 avss.n6627 0.0574697
R22485 avss.n6758 avss.n4207 0.0574697
R22486 avss.n6849 avss.n4183 0.0574697
R22487 avss.n6760 avss.n6759 0.0574697
R22488 avss.n6848 avss.n6847 0.0574697
R22489 avss.n6281 avss.n6251 0.0574697
R22490 avss.n6336 avss.n6198 0.0574697
R22491 avss.n6335 avss.n6334 0.0574697
R22492 avss.n6278 avss.n6274 0.0574697
R22493 avss.n6405 avss.n4291 0.0574697
R22494 avss.n6496 avss.n4267 0.0574697
R22495 avss.n6407 avss.n6406 0.0574697
R22496 avss.n6495 avss.n6494 0.0574697
R22497 avss.n5928 avss.n5898 0.0574697
R22498 avss.n5983 avss.n5845 0.0574697
R22499 avss.n5982 avss.n5981 0.0574697
R22500 avss.n5925 avss.n5921 0.0574697
R22501 avss.n6052 avss.n4375 0.0574697
R22502 avss.n6143 avss.n4351 0.0574697
R22503 avss.n6054 avss.n6053 0.0574697
R22504 avss.n6142 avss.n6141 0.0574697
R22505 avss.n5575 avss.n5545 0.0574697
R22506 avss.n5630 avss.n5492 0.0574697
R22507 avss.n5629 avss.n5628 0.0574697
R22508 avss.n5572 avss.n5568 0.0574697
R22509 avss.n5699 avss.n4459 0.0574697
R22510 avss.n5790 avss.n4435 0.0574697
R22511 avss.n5701 avss.n5700 0.0574697
R22512 avss.n5789 avss.n5788 0.0574697
R22513 avss.n5234 avss.n5199 0.0574697
R22514 avss.n5285 avss.n5146 0.0574697
R22515 avss.n5284 avss.n5283 0.0574697
R22516 avss.n5231 avss.n5230 0.0574697
R22517 avss.n5346 avss.n4543 0.0574697
R22518 avss.n5437 avss.n4519 0.0574697
R22519 avss.n5348 avss.n5347 0.0574697
R22520 avss.n5436 avss.n5435 0.0574697
R22521 avss.n4880 avss.n4845 0.0574697
R22522 avss.n4931 avss.n4792 0.0574697
R22523 avss.n4930 avss.n4929 0.0574697
R22524 avss.n4877 avss.n4876 0.0574697
R22525 avss.n4992 avss.n4627 0.0574697
R22526 avss.n5083 avss.n4603 0.0574697
R22527 avss.n4994 avss.n4993 0.0574697
R22528 avss.n5082 avss.n5081 0.0574697
R22529 avss.n9100 avss.n9099 0.0574697
R22530 avss.n2383 avss.n2382 0.0574697
R22531 avss.n2446 avss.n2445 0.0574697
R22532 avss.n9086 avss.n9085 0.0574697
R22533 avss.n2581 avss.n2580 0.0574697
R22534 avss.n9080 avss.n9079 0.0574697
R22535 avss.n2503 avss.n2502 0.0574697
R22536 avss.n9066 avss.n9065 0.0574697
R22537 avss.n9321 avss.n9320 0.0574697
R22538 avss.n2167 avss.n2166 0.0574697
R22539 avss.n2230 avss.n2229 0.0574697
R22540 avss.n9307 avss.n9306 0.0574697
R22541 avss.n2365 avss.n2364 0.0574697
R22542 avss.n9301 avss.n9300 0.0574697
R22543 avss.n2287 avss.n2286 0.0574697
R22544 avss.n9287 avss.n9286 0.0574697
R22545 avss.n9542 avss.n9541 0.0574697
R22546 avss.n1951 avss.n1950 0.0574697
R22547 avss.n2014 avss.n2013 0.0574697
R22548 avss.n9528 avss.n9527 0.0574697
R22549 avss.n2149 avss.n2148 0.0574697
R22550 avss.n9522 avss.n9521 0.0574697
R22551 avss.n2071 avss.n2070 0.0574697
R22552 avss.n9508 avss.n9507 0.0574697
R22553 avss.n9763 avss.n9762 0.0574697
R22554 avss.n1735 avss.n1734 0.0574697
R22555 avss.n1798 avss.n1797 0.0574697
R22556 avss.n9749 avss.n9748 0.0574697
R22557 avss.n1933 avss.n1932 0.0574697
R22558 avss.n9743 avss.n9742 0.0574697
R22559 avss.n1855 avss.n1854 0.0574697
R22560 avss.n9729 avss.n9728 0.0574697
R22561 avss.n9984 avss.n9983 0.0574697
R22562 avss.n1519 avss.n1518 0.0574697
R22563 avss.n1582 avss.n1581 0.0574697
R22564 avss.n9970 avss.n9969 0.0574697
R22565 avss.n1717 avss.n1716 0.0574697
R22566 avss.n9964 avss.n9963 0.0574697
R22567 avss.n1639 avss.n1638 0.0574697
R22568 avss.n9950 avss.n9949 0.0574697
R22569 avss.n10205 avss.n10204 0.0574697
R22570 avss.n1303 avss.n1302 0.0574697
R22571 avss.n1366 avss.n1365 0.0574697
R22572 avss.n10191 avss.n10190 0.0574697
R22573 avss.n1501 avss.n1500 0.0574697
R22574 avss.n10185 avss.n10184 0.0574697
R22575 avss.n1423 avss.n1422 0.0574697
R22576 avss.n10171 avss.n10170 0.0574697
R22577 avss.n10426 avss.n10425 0.0574697
R22578 avss.n1087 avss.n1086 0.0574697
R22579 avss.n1150 avss.n1149 0.0574697
R22580 avss.n10412 avss.n10411 0.0574697
R22581 avss.n1285 avss.n1284 0.0574697
R22582 avss.n10406 avss.n10405 0.0574697
R22583 avss.n1207 avss.n1206 0.0574697
R22584 avss.n10392 avss.n10391 0.0574697
R22585 avss.n10647 avss.n10646 0.0574697
R22586 avss.n871 avss.n870 0.0574697
R22587 avss.n934 avss.n933 0.0574697
R22588 avss.n10633 avss.n10632 0.0574697
R22589 avss.n1069 avss.n1068 0.0574697
R22590 avss.n10627 avss.n10626 0.0574697
R22591 avss.n991 avss.n990 0.0574697
R22592 avss.n10613 avss.n10612 0.0574697
R22593 avss.n10868 avss.n10867 0.0574697
R22594 avss.n655 avss.n654 0.0574697
R22595 avss.n718 avss.n717 0.0574697
R22596 avss.n10854 avss.n10853 0.0574697
R22597 avss.n853 avss.n852 0.0574697
R22598 avss.n10848 avss.n10847 0.0574697
R22599 avss.n775 avss.n774 0.0574697
R22600 avss.n10834 avss.n10833 0.0574697
R22601 avss.n11089 avss.n11088 0.0574697
R22602 avss.n439 avss.n438 0.0574697
R22603 avss.n502 avss.n501 0.0574697
R22604 avss.n11075 avss.n11074 0.0574697
R22605 avss.n637 avss.n636 0.0574697
R22606 avss.n11069 avss.n11068 0.0574697
R22607 avss.n559 avss.n558 0.0574697
R22608 avss.n11055 avss.n11054 0.0574697
R22609 avss.n340 avss.n339 0.0574697
R22610 avss.n11302 avss.n11301 0.0574697
R22611 avss.n11331 avss.n11330 0.0574697
R22612 avss.n326 avss.n325 0.0574697
R22613 avss.n312 avss.n311 0.0574697
R22614 avss.n11290 avss.n11289 0.0574697
R22615 avss.n234 avss.n233 0.0574697
R22616 avss.n11276 avss.n11275 0.0574697
R22617 avss.n123 avss.n122 0.0574697
R22618 avss.n11523 avss.n11522 0.0574697
R22619 avss.n11552 avss.n11551 0.0574697
R22620 avss.n109 avss.n108 0.0574697
R22621 avss.n95 avss.n94 0.0574697
R22622 avss.n11511 avss.n11510 0.0574697
R22623 avss.n17 avss.n16 0.0574697
R22624 avss.n11497 avss.n11496 0.0574697
R22625 avss.n8667 avss.n8664 0.0567576
R22626 avss.n8666 avss.n8665 0.0567576
R22627 avss.n8862 avss.n8856 0.0567576
R22628 avss.n8861 avss.n8860 0.0567576
R22629 avss.n8314 avss.n8311 0.0567576
R22630 avss.n8313 avss.n8312 0.0567576
R22631 avss.n8509 avss.n8503 0.0567576
R22632 avss.n8508 avss.n8507 0.0567576
R22633 avss.n7961 avss.n7958 0.0567576
R22634 avss.n7960 avss.n7959 0.0567576
R22635 avss.n8156 avss.n8150 0.0567576
R22636 avss.n8155 avss.n8154 0.0567576
R22637 avss.n7608 avss.n7605 0.0567576
R22638 avss.n7607 avss.n7606 0.0567576
R22639 avss.n7803 avss.n7797 0.0567576
R22640 avss.n7802 avss.n7801 0.0567576
R22641 avss.n7255 avss.n7252 0.0567576
R22642 avss.n7254 avss.n7253 0.0567576
R22643 avss.n7450 avss.n7444 0.0567576
R22644 avss.n7449 avss.n7448 0.0567576
R22645 avss.n6902 avss.n6899 0.0567576
R22646 avss.n6901 avss.n6900 0.0567576
R22647 avss.n7097 avss.n7091 0.0567576
R22648 avss.n7096 avss.n7095 0.0567576
R22649 avss.n6549 avss.n6546 0.0567576
R22650 avss.n6548 avss.n6547 0.0567576
R22651 avss.n6744 avss.n6738 0.0567576
R22652 avss.n6743 avss.n6742 0.0567576
R22653 avss.n6196 avss.n6193 0.0567576
R22654 avss.n6195 avss.n6194 0.0567576
R22655 avss.n6391 avss.n6385 0.0567576
R22656 avss.n6390 avss.n6389 0.0567576
R22657 avss.n5843 avss.n5840 0.0567576
R22658 avss.n5842 avss.n5841 0.0567576
R22659 avss.n6038 avss.n6032 0.0567576
R22660 avss.n6037 avss.n6036 0.0567576
R22661 avss.n5490 avss.n5487 0.0567576
R22662 avss.n5489 avss.n5488 0.0567576
R22663 avss.n5685 avss.n5679 0.0567576
R22664 avss.n5684 avss.n5683 0.0567576
R22665 avss.n5144 avss.n5137 0.0567576
R22666 avss.n5143 avss.n5142 0.0567576
R22667 avss.n5332 avss.n5326 0.0567576
R22668 avss.n5331 avss.n5330 0.0567576
R22669 avss.n4790 avss.n4783 0.0567576
R22670 avss.n4789 avss.n4788 0.0567576
R22671 avss.n4978 avss.n4972 0.0567576
R22672 avss.n4977 avss.n4976 0.0567576
R22673 avss.n2388 avss.n2387 0.0567576
R22674 avss.n2463 avss.n2462 0.0567576
R22675 avss.n2586 avss.n2585 0.0567576
R22676 avss.n2520 avss.n2519 0.0567576
R22677 avss.n2172 avss.n2171 0.0567576
R22678 avss.n2247 avss.n2246 0.0567576
R22679 avss.n2370 avss.n2369 0.0567576
R22680 avss.n2304 avss.n2303 0.0567576
R22681 avss.n1956 avss.n1955 0.0567576
R22682 avss.n2031 avss.n2030 0.0567576
R22683 avss.n2154 avss.n2153 0.0567576
R22684 avss.n2088 avss.n2087 0.0567576
R22685 avss.n1740 avss.n1739 0.0567576
R22686 avss.n1815 avss.n1814 0.0567576
R22687 avss.n1938 avss.n1937 0.0567576
R22688 avss.n1872 avss.n1871 0.0567576
R22689 avss.n1524 avss.n1523 0.0567576
R22690 avss.n1599 avss.n1598 0.0567576
R22691 avss.n1722 avss.n1721 0.0567576
R22692 avss.n1656 avss.n1655 0.0567576
R22693 avss.n1308 avss.n1307 0.0567576
R22694 avss.n1383 avss.n1382 0.0567576
R22695 avss.n1506 avss.n1505 0.0567576
R22696 avss.n1440 avss.n1439 0.0567576
R22697 avss.n1092 avss.n1091 0.0567576
R22698 avss.n1167 avss.n1166 0.0567576
R22699 avss.n1290 avss.n1289 0.0567576
R22700 avss.n1224 avss.n1223 0.0567576
R22701 avss.n876 avss.n875 0.0567576
R22702 avss.n951 avss.n950 0.0567576
R22703 avss.n1074 avss.n1073 0.0567576
R22704 avss.n1008 avss.n1007 0.0567576
R22705 avss.n660 avss.n659 0.0567576
R22706 avss.n735 avss.n734 0.0567576
R22707 avss.n858 avss.n857 0.0567576
R22708 avss.n792 avss.n791 0.0567576
R22709 avss.n444 avss.n443 0.0567576
R22710 avss.n519 avss.n518 0.0567576
R22711 avss.n642 avss.n641 0.0567576
R22712 avss.n576 avss.n575 0.0567576
R22713 avss.n11307 avss.n11306 0.0567576
R22714 avss.n11348 avss.n11347 0.0567576
R22715 avss.n317 avss.n316 0.0567576
R22716 avss.n251 avss.n250 0.0567576
R22717 avss.n11528 avss.n11527 0.0567576
R22718 avss.n11569 avss.n11568 0.0567576
R22719 avss.n100 avss.n99 0.0567576
R22720 avss.n34 avss.n33 0.0567576
R22721 avss avss.n4730 0.0564896
R22722 avss avss.n3597 0.0564896
R22723 avss.n3560 avss 0.0564896
R22724 avss.n5208 avss.n5202 0.0555815
R22725 avss.n4854 avss.n4848 0.0555815
R22726 avss.n431 avss.n373 0.0555815
R22727 avss.n214 avss.n156 0.0555815
R22728 avss.n8697 avss.n8685 0.0553333
R22729 avss.n8696 avss.n8695 0.0553333
R22730 avss.n8889 avss.n8888 0.0553333
R22731 avss.n8887 avss.n3702 0.0553333
R22732 avss.n8344 avss.n8332 0.0553333
R22733 avss.n8343 avss.n8342 0.0553333
R22734 avss.n8536 avss.n8535 0.0553333
R22735 avss.n8534 avss.n3786 0.0553333
R22736 avss.n7991 avss.n7979 0.0553333
R22737 avss.n7990 avss.n7989 0.0553333
R22738 avss.n8183 avss.n8182 0.0553333
R22739 avss.n8181 avss.n3870 0.0553333
R22740 avss.n7638 avss.n7626 0.0553333
R22741 avss.n7637 avss.n7636 0.0553333
R22742 avss.n7830 avss.n7829 0.0553333
R22743 avss.n7828 avss.n3954 0.0553333
R22744 avss.n7285 avss.n7273 0.0553333
R22745 avss.n7284 avss.n7283 0.0553333
R22746 avss.n7477 avss.n7476 0.0553333
R22747 avss.n7475 avss.n4038 0.0553333
R22748 avss.n6932 avss.n6920 0.0553333
R22749 avss.n6931 avss.n6930 0.0553333
R22750 avss.n7124 avss.n7123 0.0553333
R22751 avss.n7122 avss.n4122 0.0553333
R22752 avss.n6579 avss.n6567 0.0553333
R22753 avss.n6578 avss.n6577 0.0553333
R22754 avss.n6771 avss.n6770 0.0553333
R22755 avss.n6769 avss.n4206 0.0553333
R22756 avss.n6226 avss.n6214 0.0553333
R22757 avss.n6225 avss.n6224 0.0553333
R22758 avss.n6418 avss.n6417 0.0553333
R22759 avss.n6416 avss.n4290 0.0553333
R22760 avss.n5873 avss.n5861 0.0553333
R22761 avss.n5872 avss.n5871 0.0553333
R22762 avss.n6065 avss.n6064 0.0553333
R22763 avss.n6063 avss.n4374 0.0553333
R22764 avss.n5520 avss.n5508 0.0553333
R22765 avss.n5519 avss.n5518 0.0553333
R22766 avss.n5712 avss.n5711 0.0553333
R22767 avss.n5710 avss.n4458 0.0553333
R22768 avss.n5174 avss.n5162 0.0553333
R22769 avss.n5173 avss.n5172 0.0553333
R22770 avss.n5359 avss.n5358 0.0553333
R22771 avss.n5357 avss.n4542 0.0553333
R22772 avss.n4820 avss.n4808 0.0553333
R22773 avss.n4819 avss.n4818 0.0553333
R22774 avss.n5005 avss.n5004 0.0553333
R22775 avss.n5003 avss.n4626 0.0553333
R22776 avss.n3678 avss.n3670 0.0548345
R22777 avss.n3762 avss.n3754 0.0548345
R22778 avss.n3846 avss.n3838 0.0548345
R22779 avss.n3930 avss.n3922 0.0548345
R22780 avss.n4014 avss.n4006 0.0548345
R22781 avss.n4098 avss.n4090 0.0548345
R22782 avss.n4182 avss.n4174 0.0548345
R22783 avss.n4266 avss.n4258 0.0548345
R22784 avss.n4350 avss.n4342 0.0548345
R22785 avss.n4434 avss.n4426 0.0548345
R22786 avss.n4518 avss.n4510 0.0548345
R22787 avss.n4602 avss.n4594 0.0548345
R22788 avss.n9063 avss.n9006 0.0548345
R22789 avss.n9284 avss.n9227 0.0548345
R22790 avss.n9505 avss.n9448 0.0548345
R22791 avss.n9726 avss.n9669 0.0548345
R22792 avss.n9947 avss.n9890 0.0548345
R22793 avss.n10168 avss.n10111 0.0548345
R22794 avss.n10389 avss.n10332 0.0548345
R22795 avss.n10610 avss.n10553 0.0548345
R22796 avss.n10831 avss.n10774 0.0548345
R22797 avss.n11052 avss.n10995 0.0548345
R22798 avss.n11273 avss.n11216 0.0548345
R22799 avss.n11494 avss.n11437 0.0548345
R22800 avss.n8771 avss.n8726 0.0545704
R22801 avss.n8418 avss.n8373 0.0545704
R22802 avss.n8065 avss.n8020 0.0545704
R22803 avss.n7712 avss.n7667 0.0545704
R22804 avss.n7359 avss.n7314 0.0545704
R22805 avss.n7006 avss.n6961 0.0545704
R22806 avss.n6653 avss.n6608 0.0545704
R22807 avss.n6300 avss.n6255 0.0545704
R22808 avss.n5947 avss.n5902 0.0545704
R22809 avss.n5594 avss.n5549 0.0545704
R22810 avss.n9175 avss.n9117 0.0545704
R22811 avss.n9396 avss.n9338 0.0545704
R22812 avss.n9617 avss.n9559 0.0545704
R22813 avss.n9838 avss.n9780 0.0545704
R22814 avss.n10059 avss.n10001 0.0545704
R22815 avss.n10280 avss.n10222 0.0545704
R22816 avss.n10501 avss.n10443 0.0545704
R22817 avss.n10722 avss.n10664 0.0545704
R22818 avss.n10943 avss.n10885 0.0545704
R22819 avss.n11164 avss.n11106 0.0545704
R22820 avss.n8808 avss.n8807 0.0539091
R22821 avss.n8876 avss.n8875 0.0539091
R22822 avss.n8455 avss.n8454 0.0539091
R22823 avss.n8523 avss.n8522 0.0539091
R22824 avss.n8102 avss.n8101 0.0539091
R22825 avss.n8170 avss.n8169 0.0539091
R22826 avss.n7749 avss.n7748 0.0539091
R22827 avss.n7817 avss.n7816 0.0539091
R22828 avss.n7396 avss.n7395 0.0539091
R22829 avss.n7464 avss.n7463 0.0539091
R22830 avss.n7043 avss.n7042 0.0539091
R22831 avss.n7111 avss.n7110 0.0539091
R22832 avss.n6690 avss.n6689 0.0539091
R22833 avss.n6758 avss.n6757 0.0539091
R22834 avss.n6337 avss.n6336 0.0539091
R22835 avss.n6405 avss.n6404 0.0539091
R22836 avss.n5984 avss.n5983 0.0539091
R22837 avss.n6052 avss.n6051 0.0539091
R22838 avss.n5631 avss.n5630 0.0539091
R22839 avss.n5699 avss.n5698 0.0539091
R22840 avss.n5286 avss.n5285 0.0539091
R22841 avss.n5346 avss.n5345 0.0539091
R22842 avss.n4932 avss.n4931 0.0539091
R22843 avss.n4992 avss.n4991 0.0539091
R22844 avss.n2384 avss.n2383 0.0539091
R22845 avss.n2582 avss.n2581 0.0539091
R22846 avss.n2168 avss.n2167 0.0539091
R22847 avss.n2366 avss.n2365 0.0539091
R22848 avss.n1952 avss.n1951 0.0539091
R22849 avss.n2150 avss.n2149 0.0539091
R22850 avss.n1736 avss.n1735 0.0539091
R22851 avss.n1934 avss.n1933 0.0539091
R22852 avss.n1520 avss.n1519 0.0539091
R22853 avss.n1718 avss.n1717 0.0539091
R22854 avss.n1304 avss.n1303 0.0539091
R22855 avss.n1502 avss.n1501 0.0539091
R22856 avss.n1088 avss.n1087 0.0539091
R22857 avss.n1286 avss.n1285 0.0539091
R22858 avss.n872 avss.n871 0.0539091
R22859 avss.n1070 avss.n1069 0.0539091
R22860 avss.n656 avss.n655 0.0539091
R22861 avss.n854 avss.n853 0.0539091
R22862 avss.n440 avss.n439 0.0539091
R22863 avss.n638 avss.n637 0.0539091
R22864 avss.n11303 avss.n11302 0.0539091
R22865 avss.n313 avss.n312 0.0539091
R22866 avss.n11524 avss.n11523 0.0539091
R22867 avss.n96 avss.n95 0.0539091
R22868 avss.n8728 avss.n8726 0.0532212
R22869 avss.n8375 avss.n8373 0.0532212
R22870 avss.n8022 avss.n8020 0.0532212
R22871 avss.n7669 avss.n7667 0.0532212
R22872 avss.n7316 avss.n7314 0.0532212
R22873 avss.n6963 avss.n6961 0.0532212
R22874 avss.n6610 avss.n6608 0.0532212
R22875 avss.n6257 avss.n6255 0.0532212
R22876 avss.n5904 avss.n5902 0.0532212
R22877 avss.n5551 avss.n5549 0.0532212
R22878 avss.n9175 avss.n9174 0.0532212
R22879 avss.n9396 avss.n9395 0.0532212
R22880 avss.n9617 avss.n9616 0.0532212
R22881 avss.n9838 avss.n9837 0.0532212
R22882 avss.n10059 avss.n10058 0.0532212
R22883 avss.n10280 avss.n10279 0.0532212
R22884 avss.n10501 avss.n10500 0.0532212
R22885 avss.n10722 avss.n10721 0.0532212
R22886 avss.n10943 avss.n10942 0.0532212
R22887 avss.n11164 avss.n11163 0.0532212
R22888 avss.n5204 avss.n5202 0.053194
R22889 avss.n4850 avss.n4848 0.053194
R22890 avss.n431 avss.n430 0.053194
R22891 avss.n214 avss.n213 0.053194
R22892 avss.n3678 avss.n3677 0.0529546
R22893 avss.n3762 avss.n3761 0.0529546
R22894 avss.n3846 avss.n3845 0.0529546
R22895 avss.n3930 avss.n3929 0.0529546
R22896 avss.n4014 avss.n4013 0.0529546
R22897 avss.n4098 avss.n4097 0.0529546
R22898 avss.n4182 avss.n4181 0.0529546
R22899 avss.n4266 avss.n4265 0.0529546
R22900 avss.n4350 avss.n4349 0.0529546
R22901 avss.n4434 avss.n4433 0.0529546
R22902 avss.n4518 avss.n4517 0.0529546
R22903 avss.n4602 avss.n4601 0.0529546
R22904 avss.n9063 avss.n9062 0.0529546
R22905 avss.n9284 avss.n9283 0.0529546
R22906 avss.n9505 avss.n9504 0.0529546
R22907 avss.n9726 avss.n9725 0.0529546
R22908 avss.n9947 avss.n9946 0.0529546
R22909 avss.n10168 avss.n10167 0.0529546
R22910 avss.n10389 avss.n10388 0.0529546
R22911 avss.n10610 avss.n10609 0.0529546
R22912 avss.n10831 avss.n10830 0.0529546
R22913 avss.n11052 avss.n11051 0.0529546
R22914 avss.n11273 avss.n11272 0.0529546
R22915 avss.n11494 avss.n11493 0.0529546
R22916 avss.n8687 avss.n8669 0.0524848
R22917 avss.n8885 avss.n3703 0.0524848
R22918 avss.n8334 avss.n8316 0.0524848
R22919 avss.n8532 avss.n3787 0.0524848
R22920 avss.n7981 avss.n7963 0.0524848
R22921 avss.n8179 avss.n3871 0.0524848
R22922 avss.n7628 avss.n7610 0.0524848
R22923 avss.n7826 avss.n3955 0.0524848
R22924 avss.n7275 avss.n7257 0.0524848
R22925 avss.n7473 avss.n4039 0.0524848
R22926 avss.n6922 avss.n6904 0.0524848
R22927 avss.n7120 avss.n4123 0.0524848
R22928 avss.n6569 avss.n6551 0.0524848
R22929 avss.n6767 avss.n4207 0.0524848
R22930 avss.n6216 avss.n6198 0.0524848
R22931 avss.n6414 avss.n4291 0.0524848
R22932 avss.n5863 avss.n5845 0.0524848
R22933 avss.n6061 avss.n4375 0.0524848
R22934 avss.n5510 avss.n5492 0.0524848
R22935 avss.n5708 avss.n4459 0.0524848
R22936 avss.n5164 avss.n5146 0.0524848
R22937 avss.n5355 avss.n4543 0.0524848
R22938 avss.n4810 avss.n4792 0.0524848
R22939 avss.n5001 avss.n4627 0.0524848
R22940 avss.n2382 avss.n2381 0.0524848
R22941 avss.n2580 avss.n2579 0.0524848
R22942 avss.n2166 avss.n2165 0.0524848
R22943 avss.n2364 avss.n2363 0.0524848
R22944 avss.n1950 avss.n1949 0.0524848
R22945 avss.n2148 avss.n2147 0.0524848
R22946 avss.n1734 avss.n1733 0.0524848
R22947 avss.n1932 avss.n1931 0.0524848
R22948 avss.n1518 avss.n1517 0.0524848
R22949 avss.n1716 avss.n1715 0.0524848
R22950 avss.n1302 avss.n1301 0.0524848
R22951 avss.n1500 avss.n1499 0.0524848
R22952 avss.n1086 avss.n1085 0.0524848
R22953 avss.n1284 avss.n1283 0.0524848
R22954 avss.n870 avss.n869 0.0524848
R22955 avss.n1068 avss.n1067 0.0524848
R22956 avss.n654 avss.n653 0.0524848
R22957 avss.n852 avss.n851 0.0524848
R22958 avss.n438 avss.n437 0.0524848
R22959 avss.n636 avss.n635 0.0524848
R22960 avss.n11301 avss.n11300 0.0524848
R22961 avss.n311 avss.n310 0.0524848
R22962 avss.n11522 avss.n11521 0.0524848
R22963 avss.n94 avss.n93 0.0524848
R22964 avss.n2993 avss 0.0512812
R22965 avss.n3050 avss 0.0512812
R22966 avss.n3084 avss 0.0512812
R22967 avss.n3642 avss 0.0512812
R22968 avss.n2705 avss 0.0512812
R22969 avss.n2750 avss 0.0512812
R22970 avss.n2782 avss 0.0512812
R22971 avss.n2818 avss 0.0512812
R22972 avss.n8779 avss.n8720 0.0510606
R22973 avss.n8926 avss.n8922 0.0510606
R22974 avss.n8426 avss.n8367 0.0510606
R22975 avss.n8573 avss.n8569 0.0510606
R22976 avss.n8073 avss.n8014 0.0510606
R22977 avss.n8220 avss.n8216 0.0510606
R22978 avss.n7720 avss.n7661 0.0510606
R22979 avss.n7867 avss.n7863 0.0510606
R22980 avss.n7367 avss.n7308 0.0510606
R22981 avss.n7514 avss.n7510 0.0510606
R22982 avss.n7014 avss.n6955 0.0510606
R22983 avss.n7161 avss.n7157 0.0510606
R22984 avss.n6661 avss.n6602 0.0510606
R22985 avss.n6808 avss.n6804 0.0510606
R22986 avss.n6308 avss.n6249 0.0510606
R22987 avss.n6455 avss.n6451 0.0510606
R22988 avss.n5955 avss.n5896 0.0510606
R22989 avss.n6102 avss.n6098 0.0510606
R22990 avss.n5602 avss.n5543 0.0510606
R22991 avss.n5749 avss.n5745 0.0510606
R22992 avss.n5257 avss.n5197 0.0510606
R22993 avss.n5396 avss.n5392 0.0510606
R22994 avss.n4903 avss.n4843 0.0510606
R22995 avss.n5042 avss.n5038 0.0510606
R22996 avss.n9189 avss.n9188 0.0510606
R22997 avss.n8988 avss.n8987 0.0510606
R22998 avss.n9410 avss.n9409 0.0510606
R22999 avss.n9209 avss.n9208 0.0510606
R23000 avss.n9631 avss.n9630 0.0510606
R23001 avss.n9430 avss.n9429 0.0510606
R23002 avss.n9852 avss.n9851 0.0510606
R23003 avss.n9651 avss.n9650 0.0510606
R23004 avss.n10073 avss.n10072 0.0510606
R23005 avss.n9872 avss.n9871 0.0510606
R23006 avss.n10294 avss.n10293 0.0510606
R23007 avss.n10093 avss.n10092 0.0510606
R23008 avss.n10515 avss.n10514 0.0510606
R23009 avss.n10314 avss.n10313 0.0510606
R23010 avss.n10736 avss.n10735 0.0510606
R23011 avss.n10535 avss.n10534 0.0510606
R23012 avss.n10957 avss.n10956 0.0510606
R23013 avss.n10756 avss.n10755 0.0510606
R23014 avss.n11178 avss.n11177 0.0510606
R23015 avss.n10977 avss.n10976 0.0510606
R23016 avss.n354 avss.n353 0.0510606
R23017 avss.n11198 avss.n11197 0.0510606
R23018 avss.n137 avss.n136 0.0510606
R23019 avss.n11419 avss.n11418 0.0510606
R23020 avss.n8778 avss.n8777 0.0510606
R23021 avss.n8925 avss.n8924 0.0510606
R23022 avss.n8425 avss.n8424 0.0510606
R23023 avss.n8572 avss.n8571 0.0510606
R23024 avss.n8072 avss.n8071 0.0510606
R23025 avss.n8219 avss.n8218 0.0510606
R23026 avss.n7719 avss.n7718 0.0510606
R23027 avss.n7866 avss.n7865 0.0510606
R23028 avss.n7366 avss.n7365 0.0510606
R23029 avss.n7513 avss.n7512 0.0510606
R23030 avss.n7013 avss.n7012 0.0510606
R23031 avss.n7160 avss.n7159 0.0510606
R23032 avss.n6660 avss.n6659 0.0510606
R23033 avss.n6807 avss.n6806 0.0510606
R23034 avss.n6307 avss.n6306 0.0510606
R23035 avss.n6454 avss.n6453 0.0510606
R23036 avss.n5954 avss.n5953 0.0510606
R23037 avss.n6101 avss.n6100 0.0510606
R23038 avss.n5601 avss.n5600 0.0510606
R23039 avss.n5748 avss.n5747 0.0510606
R23040 avss.n5256 avss.n5255 0.0510606
R23041 avss.n5395 avss.n5394 0.0510606
R23042 avss.n4902 avss.n4901 0.0510606
R23043 avss.n5041 avss.n5040 0.0510606
R23044 avss.n9155 avss.n9154 0.0510606
R23045 avss.n9044 avss.n9043 0.0510606
R23046 avss.n9376 avss.n9375 0.0510606
R23047 avss.n9265 avss.n9264 0.0510606
R23048 avss.n9597 avss.n9596 0.0510606
R23049 avss.n9486 avss.n9485 0.0510606
R23050 avss.n9818 avss.n9817 0.0510606
R23051 avss.n9707 avss.n9706 0.0510606
R23052 avss.n10039 avss.n10038 0.0510606
R23053 avss.n9928 avss.n9927 0.0510606
R23054 avss.n10260 avss.n10259 0.0510606
R23055 avss.n10149 avss.n10148 0.0510606
R23056 avss.n10481 avss.n10480 0.0510606
R23057 avss.n10370 avss.n10369 0.0510606
R23058 avss.n10702 avss.n10701 0.0510606
R23059 avss.n10591 avss.n10590 0.0510606
R23060 avss.n10923 avss.n10922 0.0510606
R23061 avss.n10812 avss.n10811 0.0510606
R23062 avss.n11144 avss.n11143 0.0510606
R23063 avss.n11033 avss.n11032 0.0510606
R23064 avss.n411 avss.n410 0.0510606
R23065 avss.n11254 avss.n11253 0.0510606
R23066 avss.n194 avss.n193 0.0510606
R23067 avss.n11475 avss.n11474 0.0510606
R23068 avss.n2976 avss.n2975 0.0509808
R23069 avss.n3033 avss.n3032 0.0509808
R23070 avss.n3135 avss.n2926 0.0509808
R23071 avss.n3625 avss.n3624 0.0509808
R23072 avss.n8714 avss.n8708 0.0496364
R23073 avss.n8713 avss.n8712 0.0496364
R23074 avss.n8908 avss.n8905 0.0496364
R23075 avss.n8907 avss.n8906 0.0496364
R23076 avss.n8361 avss.n8355 0.0496364
R23077 avss.n8360 avss.n8359 0.0496364
R23078 avss.n8555 avss.n8552 0.0496364
R23079 avss.n8554 avss.n8553 0.0496364
R23080 avss.n8008 avss.n8002 0.0496364
R23081 avss.n8007 avss.n8006 0.0496364
R23082 avss.n8202 avss.n8199 0.0496364
R23083 avss.n8201 avss.n8200 0.0496364
R23084 avss.n7655 avss.n7649 0.0496364
R23085 avss.n7654 avss.n7653 0.0496364
R23086 avss.n7849 avss.n7846 0.0496364
R23087 avss.n7848 avss.n7847 0.0496364
R23088 avss.n7302 avss.n7296 0.0496364
R23089 avss.n7301 avss.n7300 0.0496364
R23090 avss.n7496 avss.n7493 0.0496364
R23091 avss.n7495 avss.n7494 0.0496364
R23092 avss.n6949 avss.n6943 0.0496364
R23093 avss.n6948 avss.n6947 0.0496364
R23094 avss.n7143 avss.n7140 0.0496364
R23095 avss.n7142 avss.n7141 0.0496364
R23096 avss.n6596 avss.n6590 0.0496364
R23097 avss.n6595 avss.n6594 0.0496364
R23098 avss.n6790 avss.n6787 0.0496364
R23099 avss.n6789 avss.n6788 0.0496364
R23100 avss.n6243 avss.n6237 0.0496364
R23101 avss.n6242 avss.n6241 0.0496364
R23102 avss.n6437 avss.n6434 0.0496364
R23103 avss.n6436 avss.n6435 0.0496364
R23104 avss.n5890 avss.n5884 0.0496364
R23105 avss.n5889 avss.n5888 0.0496364
R23106 avss.n6084 avss.n6081 0.0496364
R23107 avss.n6083 avss.n6082 0.0496364
R23108 avss.n5537 avss.n5531 0.0496364
R23109 avss.n5536 avss.n5535 0.0496364
R23110 avss.n5731 avss.n5728 0.0496364
R23111 avss.n5730 avss.n5729 0.0496364
R23112 avss.n5191 avss.n5185 0.0496364
R23113 avss.n5190 avss.n5189 0.0496364
R23114 avss.n5378 avss.n5375 0.0496364
R23115 avss.n5377 avss.n5376 0.0496364
R23116 avss.n4837 avss.n4831 0.0496364
R23117 avss.n4836 avss.n4835 0.0496364
R23118 avss.n5024 avss.n5021 0.0496364
R23119 avss.n5023 avss.n5022 0.0496364
R23120 avss.n9183 avss.n9182 0.0496364
R23121 avss.n9138 avss.n9137 0.0496364
R23122 avss.n8982 avss.n8981 0.0496364
R23123 avss.n9027 avss.n9026 0.0496364
R23124 avss.n9404 avss.n9403 0.0496364
R23125 avss.n9359 avss.n9358 0.0496364
R23126 avss.n9203 avss.n9202 0.0496364
R23127 avss.n9248 avss.n9247 0.0496364
R23128 avss.n9625 avss.n9624 0.0496364
R23129 avss.n9580 avss.n9579 0.0496364
R23130 avss.n9424 avss.n9423 0.0496364
R23131 avss.n9469 avss.n9468 0.0496364
R23132 avss.n9846 avss.n9845 0.0496364
R23133 avss.n9801 avss.n9800 0.0496364
R23134 avss.n9645 avss.n9644 0.0496364
R23135 avss.n9690 avss.n9689 0.0496364
R23136 avss.n10067 avss.n10066 0.0496364
R23137 avss.n10022 avss.n10021 0.0496364
R23138 avss.n9866 avss.n9865 0.0496364
R23139 avss.n9911 avss.n9910 0.0496364
R23140 avss.n10288 avss.n10287 0.0496364
R23141 avss.n10243 avss.n10242 0.0496364
R23142 avss.n10087 avss.n10086 0.0496364
R23143 avss.n10132 avss.n10131 0.0496364
R23144 avss.n10509 avss.n10508 0.0496364
R23145 avss.n10464 avss.n10463 0.0496364
R23146 avss.n10308 avss.n10307 0.0496364
R23147 avss.n10353 avss.n10352 0.0496364
R23148 avss.n10730 avss.n10729 0.0496364
R23149 avss.n10685 avss.n10684 0.0496364
R23150 avss.n10529 avss.n10528 0.0496364
R23151 avss.n10574 avss.n10573 0.0496364
R23152 avss.n10951 avss.n10950 0.0496364
R23153 avss.n10906 avss.n10905 0.0496364
R23154 avss.n10750 avss.n10749 0.0496364
R23155 avss.n10795 avss.n10794 0.0496364
R23156 avss.n11172 avss.n11171 0.0496364
R23157 avss.n11127 avss.n11126 0.0496364
R23158 avss.n10971 avss.n10970 0.0496364
R23159 avss.n11016 avss.n11015 0.0496364
R23160 avss.n348 avss.n347 0.0496364
R23161 avss.n394 avss.n393 0.0496364
R23162 avss.n11192 avss.n11191 0.0496364
R23163 avss.n11237 avss.n11236 0.0496364
R23164 avss.n131 avss.n130 0.0496364
R23165 avss.n177 avss.n176 0.0496364
R23166 avss.n11413 avss.n11412 0.0496364
R23167 avss.n11458 avss.n11457 0.0496364
R23168 avss.n8762 avss.n8747 0.0455026
R23169 avss.n8961 avss.n8952 0.0455026
R23170 avss.n8409 avss.n8394 0.0455026
R23171 avss.n8608 avss.n8599 0.0455026
R23172 avss.n8056 avss.n8041 0.0455026
R23173 avss.n8255 avss.n8246 0.0455026
R23174 avss.n7703 avss.n7688 0.0455026
R23175 avss.n7902 avss.n7893 0.0455026
R23176 avss.n7350 avss.n7335 0.0455026
R23177 avss.n7549 avss.n7540 0.0455026
R23178 avss.n6997 avss.n6982 0.0455026
R23179 avss.n7196 avss.n7187 0.0455026
R23180 avss.n6644 avss.n6629 0.0455026
R23181 avss.n6843 avss.n6834 0.0455026
R23182 avss.n6291 avss.n6276 0.0455026
R23183 avss.n6490 avss.n6481 0.0455026
R23184 avss.n5938 avss.n5923 0.0455026
R23185 avss.n6137 avss.n6128 0.0455026
R23186 avss.n5585 avss.n5570 0.0455026
R23187 avss.n5784 avss.n5775 0.0455026
R23188 avss.n5244 avss.n5227 0.0455026
R23189 avss.n5431 avss.n5422 0.0455026
R23190 avss.n4890 avss.n4873 0.0455026
R23191 avss.n5077 avss.n5068 0.0455026
R23192 avss.n9105 avss.n9104 0.0455026
R23193 avss.n8993 avss.n8992 0.0455026
R23194 avss.n9326 avss.n9325 0.0455026
R23195 avss.n9214 avss.n9213 0.0455026
R23196 avss.n9547 avss.n9546 0.0455026
R23197 avss.n9435 avss.n9434 0.0455026
R23198 avss.n9768 avss.n9767 0.0455026
R23199 avss.n9656 avss.n9655 0.0455026
R23200 avss.n9989 avss.n9988 0.0455026
R23201 avss.n9877 avss.n9876 0.0455026
R23202 avss.n10210 avss.n10209 0.0455026
R23203 avss.n10098 avss.n10097 0.0455026
R23204 avss.n10431 avss.n10430 0.0455026
R23205 avss.n10319 avss.n10318 0.0455026
R23206 avss.n10652 avss.n10651 0.0455026
R23207 avss.n10540 avss.n10539 0.0455026
R23208 avss.n10873 avss.n10872 0.0455026
R23209 avss.n10761 avss.n10760 0.0455026
R23210 avss.n11094 avss.n11093 0.0455026
R23211 avss.n10982 avss.n10981 0.0455026
R23212 avss.n360 avss.n359 0.0455026
R23213 avss.n11203 avss.n11202 0.0455026
R23214 avss.n143 avss.n142 0.0455026
R23215 avss.n11424 avss.n11423 0.0455026
R23216 avss.n8710 avss.n8708 0.0453636
R23217 avss.n8832 avss.n8625 0.0453636
R23218 avss.n8712 avss.n8711 0.0453636
R23219 avss.n8843 avss.n3724 0.0453636
R23220 avss.n8909 avss.n8908 0.0453636
R23221 avss.n8907 avss.n3695 0.0453636
R23222 avss.n8357 avss.n8355 0.0453636
R23223 avss.n8479 avss.n8272 0.0453636
R23224 avss.n8359 avss.n8358 0.0453636
R23225 avss.n8490 avss.n3808 0.0453636
R23226 avss.n8556 avss.n8555 0.0453636
R23227 avss.n8554 avss.n3779 0.0453636
R23228 avss.n8004 avss.n8002 0.0453636
R23229 avss.n8126 avss.n7919 0.0453636
R23230 avss.n8006 avss.n8005 0.0453636
R23231 avss.n8137 avss.n3892 0.0453636
R23232 avss.n8203 avss.n8202 0.0453636
R23233 avss.n8201 avss.n3863 0.0453636
R23234 avss.n7651 avss.n7649 0.0453636
R23235 avss.n7773 avss.n7566 0.0453636
R23236 avss.n7653 avss.n7652 0.0453636
R23237 avss.n7784 avss.n3976 0.0453636
R23238 avss.n7850 avss.n7849 0.0453636
R23239 avss.n7848 avss.n3947 0.0453636
R23240 avss.n7298 avss.n7296 0.0453636
R23241 avss.n7420 avss.n7213 0.0453636
R23242 avss.n7300 avss.n7299 0.0453636
R23243 avss.n7431 avss.n4060 0.0453636
R23244 avss.n7497 avss.n7496 0.0453636
R23245 avss.n7495 avss.n4031 0.0453636
R23246 avss.n6945 avss.n6943 0.0453636
R23247 avss.n7067 avss.n6860 0.0453636
R23248 avss.n6947 avss.n6946 0.0453636
R23249 avss.n7078 avss.n4144 0.0453636
R23250 avss.n7144 avss.n7143 0.0453636
R23251 avss.n7142 avss.n4115 0.0453636
R23252 avss.n6592 avss.n6590 0.0453636
R23253 avss.n6714 avss.n6507 0.0453636
R23254 avss.n6594 avss.n6593 0.0453636
R23255 avss.n6725 avss.n4228 0.0453636
R23256 avss.n6791 avss.n6790 0.0453636
R23257 avss.n6789 avss.n4199 0.0453636
R23258 avss.n6239 avss.n6237 0.0453636
R23259 avss.n6361 avss.n6154 0.0453636
R23260 avss.n6241 avss.n6240 0.0453636
R23261 avss.n6372 avss.n4312 0.0453636
R23262 avss.n6438 avss.n6437 0.0453636
R23263 avss.n6436 avss.n4283 0.0453636
R23264 avss.n5886 avss.n5884 0.0453636
R23265 avss.n6008 avss.n5801 0.0453636
R23266 avss.n5888 avss.n5887 0.0453636
R23267 avss.n6019 avss.n4396 0.0453636
R23268 avss.n6085 avss.n6084 0.0453636
R23269 avss.n6083 avss.n4367 0.0453636
R23270 avss.n5533 avss.n5531 0.0453636
R23271 avss.n5655 avss.n5448 0.0453636
R23272 avss.n5535 avss.n5534 0.0453636
R23273 avss.n5666 avss.n4480 0.0453636
R23274 avss.n5732 avss.n5731 0.0453636
R23275 avss.n5730 avss.n4451 0.0453636
R23276 avss.n5187 avss.n5185 0.0453636
R23277 avss.n5116 avss.n5089 0.0453636
R23278 avss.n5189 avss.n5188 0.0453636
R23279 avss.n5313 avss.n4564 0.0453636
R23280 avss.n5379 avss.n5378 0.0453636
R23281 avss.n5377 avss.n4535 0.0453636
R23282 avss.n4833 avss.n4831 0.0453636
R23283 avss.n4762 avss.n4735 0.0453636
R23284 avss.n4835 avss.n4834 0.0453636
R23285 avss.n4959 avss.n4648 0.0453636
R23286 avss.n5025 avss.n5024 0.0453636
R23287 avss.n5023 avss.n4619 0.0453636
R23288 avss.n9182 avss.n9181 0.0453636
R23289 avss.n2483 avss.n2427 0.0453636
R23290 avss.n9137 avss.n9136 0.0453636
R23291 avss.n2592 avss.n2574 0.0453636
R23292 avss.n8981 avss.n8980 0.0453636
R23293 avss.n9026 avss.n9025 0.0453636
R23294 avss.n9403 avss.n9402 0.0453636
R23295 avss.n2267 avss.n2211 0.0453636
R23296 avss.n9358 avss.n9357 0.0453636
R23297 avss.n2376 avss.n2358 0.0453636
R23298 avss.n9202 avss.n9201 0.0453636
R23299 avss.n9247 avss.n9246 0.0453636
R23300 avss.n9624 avss.n9623 0.0453636
R23301 avss.n2051 avss.n1995 0.0453636
R23302 avss.n9579 avss.n9578 0.0453636
R23303 avss.n2160 avss.n2142 0.0453636
R23304 avss.n9423 avss.n9422 0.0453636
R23305 avss.n9468 avss.n9467 0.0453636
R23306 avss.n9845 avss.n9844 0.0453636
R23307 avss.n1835 avss.n1779 0.0453636
R23308 avss.n9800 avss.n9799 0.0453636
R23309 avss.n1944 avss.n1926 0.0453636
R23310 avss.n9644 avss.n9643 0.0453636
R23311 avss.n9689 avss.n9688 0.0453636
R23312 avss.n10066 avss.n10065 0.0453636
R23313 avss.n1619 avss.n1563 0.0453636
R23314 avss.n10021 avss.n10020 0.0453636
R23315 avss.n1728 avss.n1710 0.0453636
R23316 avss.n9865 avss.n9864 0.0453636
R23317 avss.n9910 avss.n9909 0.0453636
R23318 avss.n10287 avss.n10286 0.0453636
R23319 avss.n1403 avss.n1347 0.0453636
R23320 avss.n10242 avss.n10241 0.0453636
R23321 avss.n1512 avss.n1494 0.0453636
R23322 avss.n10086 avss.n10085 0.0453636
R23323 avss.n10131 avss.n10130 0.0453636
R23324 avss.n10508 avss.n10507 0.0453636
R23325 avss.n1187 avss.n1131 0.0453636
R23326 avss.n10463 avss.n10462 0.0453636
R23327 avss.n1296 avss.n1278 0.0453636
R23328 avss.n10307 avss.n10306 0.0453636
R23329 avss.n10352 avss.n10351 0.0453636
R23330 avss.n10729 avss.n10728 0.0453636
R23331 avss.n971 avss.n915 0.0453636
R23332 avss.n10684 avss.n10683 0.0453636
R23333 avss.n1080 avss.n1062 0.0453636
R23334 avss.n10528 avss.n10527 0.0453636
R23335 avss.n10573 avss.n10572 0.0453636
R23336 avss.n10950 avss.n10949 0.0453636
R23337 avss.n755 avss.n699 0.0453636
R23338 avss.n10905 avss.n10904 0.0453636
R23339 avss.n864 avss.n846 0.0453636
R23340 avss.n10749 avss.n10748 0.0453636
R23341 avss.n10794 avss.n10793 0.0453636
R23342 avss.n11171 avss.n11170 0.0453636
R23343 avss.n539 avss.n483 0.0453636
R23344 avss.n11126 avss.n11125 0.0453636
R23345 avss.n648 avss.n630 0.0453636
R23346 avss.n10970 avss.n10969 0.0453636
R23347 avss.n11015 avss.n11014 0.0453636
R23348 avss.n347 avss.n346 0.0453636
R23349 avss.n11403 avss.n11402 0.0453636
R23350 avss.n393 avss.n392 0.0453636
R23351 avss.n323 avss.n305 0.0453636
R23352 avss.n11191 avss.n11190 0.0453636
R23353 avss.n11236 avss.n11235 0.0453636
R23354 avss.n130 avss.n129 0.0453636
R23355 avss.n11624 avss.n11623 0.0453636
R23356 avss.n176 avss.n175 0.0453636
R23357 avss.n106 avss.n88 0.0453636
R23358 avss.n11412 avss.n11411 0.0453636
R23359 avss.n11457 avss.n11456 0.0453636
R23360 avss avss.n2594 0.0447708
R23361 avss avss.n2830 0.0447708
R23362 avss.n8775 avss.n8720 0.0439394
R23363 avss.n8777 avss.n8776 0.0439394
R23364 avss.n8922 avss.n3673 0.0439394
R23365 avss.n8924 avss.n8923 0.0439394
R23366 avss.n8422 avss.n8367 0.0439394
R23367 avss.n8424 avss.n8423 0.0439394
R23368 avss.n8569 avss.n3757 0.0439394
R23369 avss.n8571 avss.n8570 0.0439394
R23370 avss.n8069 avss.n8014 0.0439394
R23371 avss.n8071 avss.n8070 0.0439394
R23372 avss.n8216 avss.n3841 0.0439394
R23373 avss.n8218 avss.n8217 0.0439394
R23374 avss.n7716 avss.n7661 0.0439394
R23375 avss.n7718 avss.n7717 0.0439394
R23376 avss.n7863 avss.n3925 0.0439394
R23377 avss.n7865 avss.n7864 0.0439394
R23378 avss.n7363 avss.n7308 0.0439394
R23379 avss.n7365 avss.n7364 0.0439394
R23380 avss.n7510 avss.n4009 0.0439394
R23381 avss.n7512 avss.n7511 0.0439394
R23382 avss.n7010 avss.n6955 0.0439394
R23383 avss.n7012 avss.n7011 0.0439394
R23384 avss.n7157 avss.n4093 0.0439394
R23385 avss.n7159 avss.n7158 0.0439394
R23386 avss.n6657 avss.n6602 0.0439394
R23387 avss.n6659 avss.n6658 0.0439394
R23388 avss.n6804 avss.n4177 0.0439394
R23389 avss.n6806 avss.n6805 0.0439394
R23390 avss.n6304 avss.n6249 0.0439394
R23391 avss.n6306 avss.n6305 0.0439394
R23392 avss.n6451 avss.n4261 0.0439394
R23393 avss.n6453 avss.n6452 0.0439394
R23394 avss.n5951 avss.n5896 0.0439394
R23395 avss.n5953 avss.n5952 0.0439394
R23396 avss.n6098 avss.n4345 0.0439394
R23397 avss.n6100 avss.n6099 0.0439394
R23398 avss.n5598 avss.n5543 0.0439394
R23399 avss.n5600 avss.n5599 0.0439394
R23400 avss.n5745 avss.n4429 0.0439394
R23401 avss.n5747 avss.n5746 0.0439394
R23402 avss.n5253 avss.n5197 0.0439394
R23403 avss.n5255 avss.n5254 0.0439394
R23404 avss.n5392 avss.n4513 0.0439394
R23405 avss.n5394 avss.n5393 0.0439394
R23406 avss.n4899 avss.n4843 0.0439394
R23407 avss.n4901 avss.n4900 0.0439394
R23408 avss.n5038 avss.n4597 0.0439394
R23409 avss.n5040 avss.n5039 0.0439394
R23410 avss.n9190 avss.n9189 0.0439394
R23411 avss.n9156 avss.n9155 0.0439394
R23412 avss.n8989 avss.n8988 0.0439394
R23413 avss.n9045 avss.n9044 0.0439394
R23414 avss.n9411 avss.n9410 0.0439394
R23415 avss.n9377 avss.n9376 0.0439394
R23416 avss.n9210 avss.n9209 0.0439394
R23417 avss.n9266 avss.n9265 0.0439394
R23418 avss.n9632 avss.n9631 0.0439394
R23419 avss.n9598 avss.n9597 0.0439394
R23420 avss.n9431 avss.n9430 0.0439394
R23421 avss.n9487 avss.n9486 0.0439394
R23422 avss.n9853 avss.n9852 0.0439394
R23423 avss.n9819 avss.n9818 0.0439394
R23424 avss.n9652 avss.n9651 0.0439394
R23425 avss.n9708 avss.n9707 0.0439394
R23426 avss.n10074 avss.n10073 0.0439394
R23427 avss.n10040 avss.n10039 0.0439394
R23428 avss.n9873 avss.n9872 0.0439394
R23429 avss.n9929 avss.n9928 0.0439394
R23430 avss.n10295 avss.n10294 0.0439394
R23431 avss.n10261 avss.n10260 0.0439394
R23432 avss.n10094 avss.n10093 0.0439394
R23433 avss.n10150 avss.n10149 0.0439394
R23434 avss.n10516 avss.n10515 0.0439394
R23435 avss.n10482 avss.n10481 0.0439394
R23436 avss.n10315 avss.n10314 0.0439394
R23437 avss.n10371 avss.n10370 0.0439394
R23438 avss.n10737 avss.n10736 0.0439394
R23439 avss.n10703 avss.n10702 0.0439394
R23440 avss.n10536 avss.n10535 0.0439394
R23441 avss.n10592 avss.n10591 0.0439394
R23442 avss.n10958 avss.n10957 0.0439394
R23443 avss.n10924 avss.n10923 0.0439394
R23444 avss.n10757 avss.n10756 0.0439394
R23445 avss.n10813 avss.n10812 0.0439394
R23446 avss.n11179 avss.n11178 0.0439394
R23447 avss.n11145 avss.n11144 0.0439394
R23448 avss.n10978 avss.n10977 0.0439394
R23449 avss.n11034 avss.n11033 0.0439394
R23450 avss.n355 avss.n354 0.0439394
R23451 avss.n412 avss.n411 0.0439394
R23452 avss.n11199 avss.n11198 0.0439394
R23453 avss.n11255 avss.n11254 0.0439394
R23454 avss.n138 avss.n137 0.0439394
R23455 avss.n195 avss.n194 0.0439394
R23456 avss.n11420 avss.n11419 0.0439394
R23457 avss.n11476 avss.n11475 0.0439394
R23458 avss.n4953 avss.n4592 0.0425061
R23459 avss.n5307 avss.n4508 0.0425061
R23460 avss.n11517 avss.n11516 0.0425061
R23461 avss.n11296 avss.n11295 0.0425061
R23462 avss.n5660 avss.n4424 0.0421693
R23463 avss.n6013 avss.n4340 0.0421693
R23464 avss.n6366 avss.n4256 0.0421693
R23465 avss.n6719 avss.n4172 0.0421693
R23466 avss.n11183 avss.n11182 0.0421693
R23467 avss.n10962 avss.n10961 0.0421693
R23468 avss.n10741 avss.n10740 0.0421693
R23469 avss.n10520 avss.n10519 0.0421693
R23470 avss.n3347 avss.n3292 0.0421667
R23471 avss.n3353 avss.n3351 0.0421667
R23472 avss.n7072 avss.n4088 0.041838
R23473 avss.n7425 avss.n4004 0.041838
R23474 avss.n7778 avss.n3920 0.041838
R23475 avss.n8131 avss.n3836 0.041838
R23476 avss.n10299 avss.n10298 0.041838
R23477 avss.n10078 avss.n10077 0.041838
R23478 avss.n9857 avss.n9856 0.041838
R23479 avss.n9636 avss.n9635 0.041838
R23480 avss.n8484 avss.n3752 0.0415118
R23481 avss.n8837 avss.n3668 0.0415118
R23482 avss.n9415 avss.n9414 0.0415118
R23483 avss.n9194 avss.n9193 0.0415118
R23484 avss.n8627 avss.n8626 0.0412792
R23485 avss.n8274 avss.n8273 0.0412792
R23486 avss.n7921 avss.n7920 0.0412792
R23487 avss.n7568 avss.n7567 0.0412792
R23488 avss.n7215 avss.n7214 0.0412792
R23489 avss.n6862 avss.n6861 0.0412792
R23490 avss.n6509 avss.n6508 0.0412792
R23491 avss.n6156 avss.n6155 0.0412792
R23492 avss.n5803 avss.n5802 0.0412792
R23493 avss.n5450 avss.n5449 0.0412792
R23494 avss.n5106 avss.n5090 0.0412792
R23495 avss.n4752 avss.n4736 0.0412792
R23496 avss.n2409 avss.n2408 0.0412792
R23497 avss.n2193 avss.n2192 0.0412792
R23498 avss.n1977 avss.n1976 0.0412792
R23499 avss.n1761 avss.n1760 0.0412792
R23500 avss.n1545 avss.n1544 0.0412792
R23501 avss.n1329 avss.n1328 0.0412792
R23502 avss.n1113 avss.n1112 0.0412792
R23503 avss.n897 avss.n896 0.0412792
R23504 avss.n681 avss.n680 0.0412792
R23505 avss.n465 avss.n464 0.0412792
R23506 avss.n11384 avss.n11383 0.0412792
R23507 avss.n11605 avss.n11604 0.0412792
R23508 avss.n3727 avss.n3723 0.0407862
R23509 avss.n3811 avss.n3807 0.0407862
R23510 avss.n3895 avss.n3891 0.0407862
R23511 avss.n3979 avss.n3975 0.0407862
R23512 avss.n4063 avss.n4059 0.0407862
R23513 avss.n4147 avss.n4143 0.0407862
R23514 avss.n4231 avss.n4227 0.0407862
R23515 avss.n4315 avss.n4311 0.0407862
R23516 avss.n4399 avss.n4395 0.0407862
R23517 avss.n4483 avss.n4479 0.0407862
R23518 avss.n5304 avss.n5302 0.0407862
R23519 avss.n4567 avss.n4563 0.0407862
R23520 avss.n4950 avss.n4948 0.0407862
R23521 avss.n4651 avss.n4647 0.0407862
R23522 avss.n2540 avss.n2539 0.0407862
R23523 avss.n2324 avss.n2323 0.0407862
R23524 avss.n2108 avss.n2107 0.0407862
R23525 avss.n1892 avss.n1891 0.0407862
R23526 avss.n1676 avss.n1675 0.0407862
R23527 avss.n1460 avss.n1459 0.0407862
R23528 avss.n1244 avss.n1243 0.0407862
R23529 avss.n1028 avss.n1027 0.0407862
R23530 avss.n812 avss.n811 0.0407862
R23531 avss.n596 avss.n595 0.0407862
R23532 avss.n11368 avss.n11367 0.0407862
R23533 avss.n271 avss.n270 0.0407862
R23534 avss.n11589 avss.n11588 0.0407862
R23535 avss.n54 avss.n53 0.0407862
R23536 avss.n3390 avss.n3273 0.0400833
R23537 avss.n8824 avss.n8823 0.0398017
R23538 avss.n8814 avss.n8648 0.0398017
R23539 avss.n8677 avss.n8660 0.0398017
R23540 avss.n8801 avss.n8678 0.0398017
R23541 avss.n8799 avss.n8681 0.0398017
R23542 avss.n8718 avss.n8705 0.0398017
R23543 avss.n8742 avss.n8729 0.0398017
R23544 avss.n8763 avss.n8746 0.0398017
R23545 avss.n8847 avss.n3720 0.0398017
R23546 avss.n8867 avss.n3713 0.0398017
R23547 avss.n8870 avss.n8869 0.0398017
R23548 avss.n3705 avss.n3699 0.0398017
R23549 avss.n8895 avss.n3692 0.0398017
R23550 avss.n8931 avss.n3685 0.0398017
R23551 avss.n8942 avss.n3683 0.0398017
R23552 avss.n8951 avss.n3682 0.0398017
R23553 avss.n8471 avss.n8470 0.0398017
R23554 avss.n8461 avss.n8295 0.0398017
R23555 avss.n8324 avss.n8307 0.0398017
R23556 avss.n8448 avss.n8325 0.0398017
R23557 avss.n8446 avss.n8328 0.0398017
R23558 avss.n8365 avss.n8352 0.0398017
R23559 avss.n8389 avss.n8376 0.0398017
R23560 avss.n8410 avss.n8393 0.0398017
R23561 avss.n8494 avss.n3804 0.0398017
R23562 avss.n8514 avss.n3797 0.0398017
R23563 avss.n8517 avss.n8516 0.0398017
R23564 avss.n3789 avss.n3783 0.0398017
R23565 avss.n8542 avss.n3776 0.0398017
R23566 avss.n8578 avss.n3769 0.0398017
R23567 avss.n8589 avss.n3767 0.0398017
R23568 avss.n8598 avss.n3766 0.0398017
R23569 avss.n8118 avss.n8117 0.0398017
R23570 avss.n8108 avss.n7942 0.0398017
R23571 avss.n7971 avss.n7954 0.0398017
R23572 avss.n8095 avss.n7972 0.0398017
R23573 avss.n8093 avss.n7975 0.0398017
R23574 avss.n8012 avss.n7999 0.0398017
R23575 avss.n8036 avss.n8023 0.0398017
R23576 avss.n8057 avss.n8040 0.0398017
R23577 avss.n8141 avss.n3888 0.0398017
R23578 avss.n8161 avss.n3881 0.0398017
R23579 avss.n8164 avss.n8163 0.0398017
R23580 avss.n3873 avss.n3867 0.0398017
R23581 avss.n8189 avss.n3860 0.0398017
R23582 avss.n8225 avss.n3853 0.0398017
R23583 avss.n8236 avss.n3851 0.0398017
R23584 avss.n8245 avss.n3850 0.0398017
R23585 avss.n7765 avss.n7764 0.0398017
R23586 avss.n7755 avss.n7589 0.0398017
R23587 avss.n7618 avss.n7601 0.0398017
R23588 avss.n7742 avss.n7619 0.0398017
R23589 avss.n7740 avss.n7622 0.0398017
R23590 avss.n7659 avss.n7646 0.0398017
R23591 avss.n7683 avss.n7670 0.0398017
R23592 avss.n7704 avss.n7687 0.0398017
R23593 avss.n7788 avss.n3972 0.0398017
R23594 avss.n7808 avss.n3965 0.0398017
R23595 avss.n7811 avss.n7810 0.0398017
R23596 avss.n3957 avss.n3951 0.0398017
R23597 avss.n7836 avss.n3944 0.0398017
R23598 avss.n7872 avss.n3937 0.0398017
R23599 avss.n7883 avss.n3935 0.0398017
R23600 avss.n7892 avss.n3934 0.0398017
R23601 avss.n7412 avss.n7411 0.0398017
R23602 avss.n7402 avss.n7236 0.0398017
R23603 avss.n7265 avss.n7248 0.0398017
R23604 avss.n7389 avss.n7266 0.0398017
R23605 avss.n7387 avss.n7269 0.0398017
R23606 avss.n7306 avss.n7293 0.0398017
R23607 avss.n7330 avss.n7317 0.0398017
R23608 avss.n7351 avss.n7334 0.0398017
R23609 avss.n7435 avss.n4056 0.0398017
R23610 avss.n7455 avss.n4049 0.0398017
R23611 avss.n7458 avss.n7457 0.0398017
R23612 avss.n4041 avss.n4035 0.0398017
R23613 avss.n7483 avss.n4028 0.0398017
R23614 avss.n7519 avss.n4021 0.0398017
R23615 avss.n7530 avss.n4019 0.0398017
R23616 avss.n7539 avss.n4018 0.0398017
R23617 avss.n7059 avss.n7058 0.0398017
R23618 avss.n7049 avss.n6883 0.0398017
R23619 avss.n6912 avss.n6895 0.0398017
R23620 avss.n7036 avss.n6913 0.0398017
R23621 avss.n7034 avss.n6916 0.0398017
R23622 avss.n6953 avss.n6940 0.0398017
R23623 avss.n6977 avss.n6964 0.0398017
R23624 avss.n6998 avss.n6981 0.0398017
R23625 avss.n7082 avss.n4140 0.0398017
R23626 avss.n7102 avss.n4133 0.0398017
R23627 avss.n7105 avss.n7104 0.0398017
R23628 avss.n4125 avss.n4119 0.0398017
R23629 avss.n7130 avss.n4112 0.0398017
R23630 avss.n7166 avss.n4105 0.0398017
R23631 avss.n7177 avss.n4103 0.0398017
R23632 avss.n7186 avss.n4102 0.0398017
R23633 avss.n6706 avss.n6705 0.0398017
R23634 avss.n6696 avss.n6530 0.0398017
R23635 avss.n6559 avss.n6542 0.0398017
R23636 avss.n6683 avss.n6560 0.0398017
R23637 avss.n6681 avss.n6563 0.0398017
R23638 avss.n6600 avss.n6587 0.0398017
R23639 avss.n6624 avss.n6611 0.0398017
R23640 avss.n6645 avss.n6628 0.0398017
R23641 avss.n6729 avss.n4224 0.0398017
R23642 avss.n6749 avss.n4217 0.0398017
R23643 avss.n6752 avss.n6751 0.0398017
R23644 avss.n4209 avss.n4203 0.0398017
R23645 avss.n6777 avss.n4196 0.0398017
R23646 avss.n6813 avss.n4189 0.0398017
R23647 avss.n6824 avss.n4187 0.0398017
R23648 avss.n6833 avss.n4186 0.0398017
R23649 avss.n6353 avss.n6352 0.0398017
R23650 avss.n6343 avss.n6177 0.0398017
R23651 avss.n6206 avss.n6189 0.0398017
R23652 avss.n6330 avss.n6207 0.0398017
R23653 avss.n6328 avss.n6210 0.0398017
R23654 avss.n6247 avss.n6234 0.0398017
R23655 avss.n6271 avss.n6258 0.0398017
R23656 avss.n6292 avss.n6275 0.0398017
R23657 avss.n6376 avss.n4308 0.0398017
R23658 avss.n6396 avss.n4301 0.0398017
R23659 avss.n6399 avss.n6398 0.0398017
R23660 avss.n4293 avss.n4287 0.0398017
R23661 avss.n6424 avss.n4280 0.0398017
R23662 avss.n6460 avss.n4273 0.0398017
R23663 avss.n6471 avss.n4271 0.0398017
R23664 avss.n6480 avss.n4270 0.0398017
R23665 avss.n6000 avss.n5999 0.0398017
R23666 avss.n5990 avss.n5824 0.0398017
R23667 avss.n5853 avss.n5836 0.0398017
R23668 avss.n5977 avss.n5854 0.0398017
R23669 avss.n5975 avss.n5857 0.0398017
R23670 avss.n5894 avss.n5881 0.0398017
R23671 avss.n5918 avss.n5905 0.0398017
R23672 avss.n5939 avss.n5922 0.0398017
R23673 avss.n6023 avss.n4392 0.0398017
R23674 avss.n6043 avss.n4385 0.0398017
R23675 avss.n6046 avss.n6045 0.0398017
R23676 avss.n4377 avss.n4371 0.0398017
R23677 avss.n6071 avss.n4364 0.0398017
R23678 avss.n6107 avss.n4357 0.0398017
R23679 avss.n6118 avss.n4355 0.0398017
R23680 avss.n6127 avss.n4354 0.0398017
R23681 avss.n5647 avss.n5646 0.0398017
R23682 avss.n5637 avss.n5471 0.0398017
R23683 avss.n5500 avss.n5483 0.0398017
R23684 avss.n5624 avss.n5501 0.0398017
R23685 avss.n5622 avss.n5504 0.0398017
R23686 avss.n5541 avss.n5528 0.0398017
R23687 avss.n5565 avss.n5552 0.0398017
R23688 avss.n5586 avss.n5569 0.0398017
R23689 avss.n5670 avss.n4476 0.0398017
R23690 avss.n5690 avss.n4469 0.0398017
R23691 avss.n5693 avss.n5692 0.0398017
R23692 avss.n4461 avss.n4455 0.0398017
R23693 avss.n5718 avss.n4448 0.0398017
R23694 avss.n5754 avss.n4441 0.0398017
R23695 avss.n5765 avss.n4439 0.0398017
R23696 avss.n5774 avss.n4438 0.0398017
R23697 avss.n5130 avss.n5099 0.0398017
R23698 avss.n5293 avss.n5292 0.0398017
R23699 avss.n5154 avss.n5133 0.0398017
R23700 avss.n5279 avss.n5155 0.0398017
R23701 avss.n5277 avss.n5158 0.0398017
R23702 avss.n5195 avss.n5182 0.0398017
R23703 avss.n5225 avss.n5212 0.0398017
R23704 avss.n5246 avss.n5245 0.0398017
R23705 avss.n5317 avss.n4560 0.0398017
R23706 avss.n5337 avss.n4553 0.0398017
R23707 avss.n5340 avss.n5339 0.0398017
R23708 avss.n4545 avss.n4539 0.0398017
R23709 avss.n5365 avss.n4532 0.0398017
R23710 avss.n5401 avss.n4525 0.0398017
R23711 avss.n5412 avss.n4523 0.0398017
R23712 avss.n5421 avss.n4522 0.0398017
R23713 avss.n4776 avss.n4745 0.0398017
R23714 avss.n4939 avss.n4938 0.0398017
R23715 avss.n4800 avss.n4779 0.0398017
R23716 avss.n4925 avss.n4801 0.0398017
R23717 avss.n4923 avss.n4804 0.0398017
R23718 avss.n4841 avss.n4828 0.0398017
R23719 avss.n4871 avss.n4858 0.0398017
R23720 avss.n4892 avss.n4891 0.0398017
R23721 avss.n4963 avss.n4644 0.0398017
R23722 avss.n4983 avss.n4637 0.0398017
R23723 avss.n4986 avss.n4985 0.0398017
R23724 avss.n4629 avss.n4623 0.0398017
R23725 avss.n5011 avss.n4616 0.0398017
R23726 avss.n5047 avss.n4609 0.0398017
R23727 avss.n5058 avss.n4607 0.0398017
R23728 avss.n5067 avss.n4606 0.0398017
R23729 avss.n2399 avss.n2398 0.0398017
R23730 avss.n2469 avss.n2468 0.0398017
R23731 avss.n2450 avss.n2449 0.0398017
R23732 avss.n2437 avss.n2436 0.0398017
R23733 avss.n9127 avss.n9126 0.0398017
R23734 avss.n9142 avss.n9141 0.0398017
R23735 avss.n9161 avss.n9160 0.0398017
R23736 avss.n9107 avss.n9106 0.0398017
R23737 avss.n2546 avss.n2545 0.0398017
R23738 avss.n2526 avss.n2525 0.0398017
R23739 avss.n2507 avss.n2506 0.0398017
R23740 avss.n2494 avss.n2493 0.0398017
R23741 avss.n9016 avss.n9015 0.0398017
R23742 avss.n9031 avss.n9030 0.0398017
R23743 avss.n9050 avss.n9049 0.0398017
R23744 avss.n8995 avss.n8994 0.0398017
R23745 avss.n2183 avss.n2182 0.0398017
R23746 avss.n2253 avss.n2252 0.0398017
R23747 avss.n2234 avss.n2233 0.0398017
R23748 avss.n2221 avss.n2220 0.0398017
R23749 avss.n9348 avss.n9347 0.0398017
R23750 avss.n9363 avss.n9362 0.0398017
R23751 avss.n9382 avss.n9381 0.0398017
R23752 avss.n9328 avss.n9327 0.0398017
R23753 avss.n2330 avss.n2329 0.0398017
R23754 avss.n2310 avss.n2309 0.0398017
R23755 avss.n2291 avss.n2290 0.0398017
R23756 avss.n2278 avss.n2277 0.0398017
R23757 avss.n9237 avss.n9236 0.0398017
R23758 avss.n9252 avss.n9251 0.0398017
R23759 avss.n9271 avss.n9270 0.0398017
R23760 avss.n9216 avss.n9215 0.0398017
R23761 avss.n1967 avss.n1966 0.0398017
R23762 avss.n2037 avss.n2036 0.0398017
R23763 avss.n2018 avss.n2017 0.0398017
R23764 avss.n2005 avss.n2004 0.0398017
R23765 avss.n9569 avss.n9568 0.0398017
R23766 avss.n9584 avss.n9583 0.0398017
R23767 avss.n9603 avss.n9602 0.0398017
R23768 avss.n9549 avss.n9548 0.0398017
R23769 avss.n2114 avss.n2113 0.0398017
R23770 avss.n2094 avss.n2093 0.0398017
R23771 avss.n2075 avss.n2074 0.0398017
R23772 avss.n2062 avss.n2061 0.0398017
R23773 avss.n9458 avss.n9457 0.0398017
R23774 avss.n9473 avss.n9472 0.0398017
R23775 avss.n9492 avss.n9491 0.0398017
R23776 avss.n9437 avss.n9436 0.0398017
R23777 avss.n1751 avss.n1750 0.0398017
R23778 avss.n1821 avss.n1820 0.0398017
R23779 avss.n1802 avss.n1801 0.0398017
R23780 avss.n1789 avss.n1788 0.0398017
R23781 avss.n9790 avss.n9789 0.0398017
R23782 avss.n9805 avss.n9804 0.0398017
R23783 avss.n9824 avss.n9823 0.0398017
R23784 avss.n9770 avss.n9769 0.0398017
R23785 avss.n1898 avss.n1897 0.0398017
R23786 avss.n1878 avss.n1877 0.0398017
R23787 avss.n1859 avss.n1858 0.0398017
R23788 avss.n1846 avss.n1845 0.0398017
R23789 avss.n9679 avss.n9678 0.0398017
R23790 avss.n9694 avss.n9693 0.0398017
R23791 avss.n9713 avss.n9712 0.0398017
R23792 avss.n9658 avss.n9657 0.0398017
R23793 avss.n1535 avss.n1534 0.0398017
R23794 avss.n1605 avss.n1604 0.0398017
R23795 avss.n1586 avss.n1585 0.0398017
R23796 avss.n1573 avss.n1572 0.0398017
R23797 avss.n10011 avss.n10010 0.0398017
R23798 avss.n10026 avss.n10025 0.0398017
R23799 avss.n10045 avss.n10044 0.0398017
R23800 avss.n9991 avss.n9990 0.0398017
R23801 avss.n1682 avss.n1681 0.0398017
R23802 avss.n1662 avss.n1661 0.0398017
R23803 avss.n1643 avss.n1642 0.0398017
R23804 avss.n1630 avss.n1629 0.0398017
R23805 avss.n9900 avss.n9899 0.0398017
R23806 avss.n9915 avss.n9914 0.0398017
R23807 avss.n9934 avss.n9933 0.0398017
R23808 avss.n9879 avss.n9878 0.0398017
R23809 avss.n1319 avss.n1318 0.0398017
R23810 avss.n1389 avss.n1388 0.0398017
R23811 avss.n1370 avss.n1369 0.0398017
R23812 avss.n1357 avss.n1356 0.0398017
R23813 avss.n10232 avss.n10231 0.0398017
R23814 avss.n10247 avss.n10246 0.0398017
R23815 avss.n10266 avss.n10265 0.0398017
R23816 avss.n10212 avss.n10211 0.0398017
R23817 avss.n1466 avss.n1465 0.0398017
R23818 avss.n1446 avss.n1445 0.0398017
R23819 avss.n1427 avss.n1426 0.0398017
R23820 avss.n1414 avss.n1413 0.0398017
R23821 avss.n10121 avss.n10120 0.0398017
R23822 avss.n10136 avss.n10135 0.0398017
R23823 avss.n10155 avss.n10154 0.0398017
R23824 avss.n10100 avss.n10099 0.0398017
R23825 avss.n1103 avss.n1102 0.0398017
R23826 avss.n1173 avss.n1172 0.0398017
R23827 avss.n1154 avss.n1153 0.0398017
R23828 avss.n1141 avss.n1140 0.0398017
R23829 avss.n10453 avss.n10452 0.0398017
R23830 avss.n10468 avss.n10467 0.0398017
R23831 avss.n10487 avss.n10486 0.0398017
R23832 avss.n10433 avss.n10432 0.0398017
R23833 avss.n1250 avss.n1249 0.0398017
R23834 avss.n1230 avss.n1229 0.0398017
R23835 avss.n1211 avss.n1210 0.0398017
R23836 avss.n1198 avss.n1197 0.0398017
R23837 avss.n10342 avss.n10341 0.0398017
R23838 avss.n10357 avss.n10356 0.0398017
R23839 avss.n10376 avss.n10375 0.0398017
R23840 avss.n10321 avss.n10320 0.0398017
R23841 avss.n887 avss.n886 0.0398017
R23842 avss.n957 avss.n956 0.0398017
R23843 avss.n938 avss.n937 0.0398017
R23844 avss.n925 avss.n924 0.0398017
R23845 avss.n10674 avss.n10673 0.0398017
R23846 avss.n10689 avss.n10688 0.0398017
R23847 avss.n10708 avss.n10707 0.0398017
R23848 avss.n10654 avss.n10653 0.0398017
R23849 avss.n1034 avss.n1033 0.0398017
R23850 avss.n1014 avss.n1013 0.0398017
R23851 avss.n995 avss.n994 0.0398017
R23852 avss.n982 avss.n981 0.0398017
R23853 avss.n10563 avss.n10562 0.0398017
R23854 avss.n10578 avss.n10577 0.0398017
R23855 avss.n10597 avss.n10596 0.0398017
R23856 avss.n10542 avss.n10541 0.0398017
R23857 avss.n671 avss.n670 0.0398017
R23858 avss.n741 avss.n740 0.0398017
R23859 avss.n722 avss.n721 0.0398017
R23860 avss.n709 avss.n708 0.0398017
R23861 avss.n10895 avss.n10894 0.0398017
R23862 avss.n10910 avss.n10909 0.0398017
R23863 avss.n10929 avss.n10928 0.0398017
R23864 avss.n10875 avss.n10874 0.0398017
R23865 avss.n818 avss.n817 0.0398017
R23866 avss.n798 avss.n797 0.0398017
R23867 avss.n779 avss.n778 0.0398017
R23868 avss.n766 avss.n765 0.0398017
R23869 avss.n10784 avss.n10783 0.0398017
R23870 avss.n10799 avss.n10798 0.0398017
R23871 avss.n10818 avss.n10817 0.0398017
R23872 avss.n10763 avss.n10762 0.0398017
R23873 avss.n455 avss.n454 0.0398017
R23874 avss.n525 avss.n524 0.0398017
R23875 avss.n506 avss.n505 0.0398017
R23876 avss.n493 avss.n492 0.0398017
R23877 avss.n11116 avss.n11115 0.0398017
R23878 avss.n11131 avss.n11130 0.0398017
R23879 avss.n11150 avss.n11149 0.0398017
R23880 avss.n11096 avss.n11095 0.0398017
R23881 avss.n602 avss.n601 0.0398017
R23882 avss.n582 avss.n581 0.0398017
R23883 avss.n563 avss.n562 0.0398017
R23884 avss.n550 avss.n549 0.0398017
R23885 avss.n11005 avss.n11004 0.0398017
R23886 avss.n11020 avss.n11019 0.0398017
R23887 avss.n11039 avss.n11038 0.0398017
R23888 avss.n10984 avss.n10983 0.0398017
R23889 avss.n11373 avss.n11372 0.0398017
R23890 avss.n11354 avss.n11353 0.0398017
R23891 avss.n11335 avss.n11334 0.0398017
R23892 avss.n11322 avss.n11321 0.0398017
R23893 avss.n383 avss.n382 0.0398017
R23894 avss.n398 avss.n397 0.0398017
R23895 avss.n417 avss.n416 0.0398017
R23896 avss.n362 avss.n361 0.0398017
R23897 avss.n277 avss.n276 0.0398017
R23898 avss.n257 avss.n256 0.0398017
R23899 avss.n238 avss.n237 0.0398017
R23900 avss.n225 avss.n224 0.0398017
R23901 avss.n11226 avss.n11225 0.0398017
R23902 avss.n11241 avss.n11240 0.0398017
R23903 avss.n11260 avss.n11259 0.0398017
R23904 avss.n11205 avss.n11204 0.0398017
R23905 avss.n11594 avss.n11593 0.0398017
R23906 avss.n11575 avss.n11574 0.0398017
R23907 avss.n11556 avss.n11555 0.0398017
R23908 avss.n11543 avss.n11542 0.0398017
R23909 avss.n166 avss.n165 0.0398017
R23910 avss.n181 avss.n180 0.0398017
R23911 avss.n200 avss.n199 0.0398017
R23912 avss.n145 avss.n144 0.0398017
R23913 avss.n60 avss.n59 0.0398017
R23914 avss.n40 avss.n39 0.0398017
R23915 avss.n21 avss.n20 0.0398017
R23916 avss.n8 avss.n7 0.0398017
R23917 avss.n11447 avss.n11446 0.0398017
R23918 avss.n11462 avss.n11461 0.0398017
R23919 avss.n11481 avss.n11480 0.0398017
R23920 avss.n11426 avss.n11425 0.0398017
R23921 avss.n8693 avss.n8685 0.0396667
R23922 avss.n8695 avss.n8694 0.0396667
R23923 avss.n8890 avss.n8889 0.0396667
R23924 avss.n8891 avss.n3702 0.0396667
R23925 avss.n8340 avss.n8332 0.0396667
R23926 avss.n8342 avss.n8341 0.0396667
R23927 avss.n8537 avss.n8536 0.0396667
R23928 avss.n8538 avss.n3786 0.0396667
R23929 avss.n7987 avss.n7979 0.0396667
R23930 avss.n7989 avss.n7988 0.0396667
R23931 avss.n8184 avss.n8183 0.0396667
R23932 avss.n8185 avss.n3870 0.0396667
R23933 avss.n7634 avss.n7626 0.0396667
R23934 avss.n7636 avss.n7635 0.0396667
R23935 avss.n7831 avss.n7830 0.0396667
R23936 avss.n7832 avss.n3954 0.0396667
R23937 avss.n7281 avss.n7273 0.0396667
R23938 avss.n7283 avss.n7282 0.0396667
R23939 avss.n7478 avss.n7477 0.0396667
R23940 avss.n7479 avss.n4038 0.0396667
R23941 avss.n6928 avss.n6920 0.0396667
R23942 avss.n6930 avss.n6929 0.0396667
R23943 avss.n7125 avss.n7124 0.0396667
R23944 avss.n7126 avss.n4122 0.0396667
R23945 avss.n6575 avss.n6567 0.0396667
R23946 avss.n6577 avss.n6576 0.0396667
R23947 avss.n6772 avss.n6771 0.0396667
R23948 avss.n6773 avss.n4206 0.0396667
R23949 avss.n6222 avss.n6214 0.0396667
R23950 avss.n6224 avss.n6223 0.0396667
R23951 avss.n6419 avss.n6418 0.0396667
R23952 avss.n6420 avss.n4290 0.0396667
R23953 avss.n5869 avss.n5861 0.0396667
R23954 avss.n5871 avss.n5870 0.0396667
R23955 avss.n6066 avss.n6065 0.0396667
R23956 avss.n6067 avss.n4374 0.0396667
R23957 avss.n5516 avss.n5508 0.0396667
R23958 avss.n5518 avss.n5517 0.0396667
R23959 avss.n5713 avss.n5712 0.0396667
R23960 avss.n5714 avss.n4458 0.0396667
R23961 avss.n5170 avss.n5162 0.0396667
R23962 avss.n5172 avss.n5171 0.0396667
R23963 avss.n5360 avss.n5359 0.0396667
R23964 avss.n5361 avss.n4542 0.0396667
R23965 avss.n4816 avss.n4808 0.0396667
R23966 avss.n4818 avss.n4817 0.0396667
R23967 avss.n5006 avss.n5005 0.0396667
R23968 avss.n5007 avss.n4626 0.0396667
R23969 avss.n2379 avss.n2378 0.0396667
R23970 avss.n2430 avss.n2429 0.0396667
R23971 avss.n2577 avss.n2576 0.0396667
R23972 avss.n2487 avss.n2486 0.0396667
R23973 avss.n2163 avss.n2162 0.0396667
R23974 avss.n2214 avss.n2213 0.0396667
R23975 avss.n2361 avss.n2360 0.0396667
R23976 avss.n2271 avss.n2270 0.0396667
R23977 avss.n1947 avss.n1946 0.0396667
R23978 avss.n1998 avss.n1997 0.0396667
R23979 avss.n2145 avss.n2144 0.0396667
R23980 avss.n2055 avss.n2054 0.0396667
R23981 avss.n1731 avss.n1730 0.0396667
R23982 avss.n1782 avss.n1781 0.0396667
R23983 avss.n1929 avss.n1928 0.0396667
R23984 avss.n1839 avss.n1838 0.0396667
R23985 avss.n1515 avss.n1514 0.0396667
R23986 avss.n1566 avss.n1565 0.0396667
R23987 avss.n1713 avss.n1712 0.0396667
R23988 avss.n1623 avss.n1622 0.0396667
R23989 avss.n1299 avss.n1298 0.0396667
R23990 avss.n1350 avss.n1349 0.0396667
R23991 avss.n1497 avss.n1496 0.0396667
R23992 avss.n1407 avss.n1406 0.0396667
R23993 avss.n1083 avss.n1082 0.0396667
R23994 avss.n1134 avss.n1133 0.0396667
R23995 avss.n1281 avss.n1280 0.0396667
R23996 avss.n1191 avss.n1190 0.0396667
R23997 avss.n867 avss.n866 0.0396667
R23998 avss.n918 avss.n917 0.0396667
R23999 avss.n1065 avss.n1064 0.0396667
R24000 avss.n975 avss.n974 0.0396667
R24001 avss.n651 avss.n650 0.0396667
R24002 avss.n702 avss.n701 0.0396667
R24003 avss.n849 avss.n848 0.0396667
R24004 avss.n759 avss.n758 0.0396667
R24005 avss.n435 avss.n434 0.0396667
R24006 avss.n486 avss.n485 0.0396667
R24007 avss.n633 avss.n632 0.0396667
R24008 avss.n543 avss.n542 0.0396667
R24009 avss.n11298 avss.n11297 0.0396667
R24010 avss.n11315 avss.n11314 0.0396667
R24011 avss.n308 avss.n307 0.0396667
R24012 avss.n218 avss.n217 0.0396667
R24013 avss.n11519 avss.n11518 0.0396667
R24014 avss.n11536 avss.n11535 0.0396667
R24015 avss.n91 avss.n90 0.0396667
R24016 avss.n1 avss.n0 0.0396667
R24017 avss.n8668 avss.n8667 0.0382424
R24018 avss.n8666 avss.n8662 0.0382424
R24019 avss.n8858 avss.n8856 0.0382424
R24020 avss.n8860 avss.n8859 0.0382424
R24021 avss.n8315 avss.n8314 0.0382424
R24022 avss.n8313 avss.n8309 0.0382424
R24023 avss.n8505 avss.n8503 0.0382424
R24024 avss.n8507 avss.n8506 0.0382424
R24025 avss.n7962 avss.n7961 0.0382424
R24026 avss.n7960 avss.n7956 0.0382424
R24027 avss.n8152 avss.n8150 0.0382424
R24028 avss.n8154 avss.n8153 0.0382424
R24029 avss.n7609 avss.n7608 0.0382424
R24030 avss.n7607 avss.n7603 0.0382424
R24031 avss.n7799 avss.n7797 0.0382424
R24032 avss.n7801 avss.n7800 0.0382424
R24033 avss.n7256 avss.n7255 0.0382424
R24034 avss.n7254 avss.n7250 0.0382424
R24035 avss.n7446 avss.n7444 0.0382424
R24036 avss.n7448 avss.n7447 0.0382424
R24037 avss.n6903 avss.n6902 0.0382424
R24038 avss.n6901 avss.n6897 0.0382424
R24039 avss.n7093 avss.n7091 0.0382424
R24040 avss.n7095 avss.n7094 0.0382424
R24041 avss.n6550 avss.n6549 0.0382424
R24042 avss.n6548 avss.n6544 0.0382424
R24043 avss.n6740 avss.n6738 0.0382424
R24044 avss.n6742 avss.n6741 0.0382424
R24045 avss.n6197 avss.n6196 0.0382424
R24046 avss.n6195 avss.n6191 0.0382424
R24047 avss.n6387 avss.n6385 0.0382424
R24048 avss.n6389 avss.n6388 0.0382424
R24049 avss.n5844 avss.n5843 0.0382424
R24050 avss.n5842 avss.n5838 0.0382424
R24051 avss.n6034 avss.n6032 0.0382424
R24052 avss.n6036 avss.n6035 0.0382424
R24053 avss.n5491 avss.n5490 0.0382424
R24054 avss.n5489 avss.n5485 0.0382424
R24055 avss.n5681 avss.n5679 0.0382424
R24056 avss.n5683 avss.n5682 0.0382424
R24057 avss.n5145 avss.n5144 0.0382424
R24058 avss.n5143 avss.n5135 0.0382424
R24059 avss.n5328 avss.n5326 0.0382424
R24060 avss.n5330 avss.n5329 0.0382424
R24061 avss.n4791 avss.n4790 0.0382424
R24062 avss.n4789 avss.n4781 0.0382424
R24063 avss.n4974 avss.n4972 0.0382424
R24064 avss.n4976 avss.n4975 0.0382424
R24065 avss.n2387 avss.n2386 0.0382424
R24066 avss.n2462 avss.n2461 0.0382424
R24067 avss.n2585 avss.n2584 0.0382424
R24068 avss.n2519 avss.n2518 0.0382424
R24069 avss.n2171 avss.n2170 0.0382424
R24070 avss.n2246 avss.n2245 0.0382424
R24071 avss.n2369 avss.n2368 0.0382424
R24072 avss.n2303 avss.n2302 0.0382424
R24073 avss.n1955 avss.n1954 0.0382424
R24074 avss.n2030 avss.n2029 0.0382424
R24075 avss.n2153 avss.n2152 0.0382424
R24076 avss.n2087 avss.n2086 0.0382424
R24077 avss.n1739 avss.n1738 0.0382424
R24078 avss.n1814 avss.n1813 0.0382424
R24079 avss.n1937 avss.n1936 0.0382424
R24080 avss.n1871 avss.n1870 0.0382424
R24081 avss.n1523 avss.n1522 0.0382424
R24082 avss.n1598 avss.n1597 0.0382424
R24083 avss.n1721 avss.n1720 0.0382424
R24084 avss.n1655 avss.n1654 0.0382424
R24085 avss.n1307 avss.n1306 0.0382424
R24086 avss.n1382 avss.n1381 0.0382424
R24087 avss.n1505 avss.n1504 0.0382424
R24088 avss.n1439 avss.n1438 0.0382424
R24089 avss.n1091 avss.n1090 0.0382424
R24090 avss.n1166 avss.n1165 0.0382424
R24091 avss.n1289 avss.n1288 0.0382424
R24092 avss.n1223 avss.n1222 0.0382424
R24093 avss.n875 avss.n874 0.0382424
R24094 avss.n950 avss.n949 0.0382424
R24095 avss.n1073 avss.n1072 0.0382424
R24096 avss.n1007 avss.n1006 0.0382424
R24097 avss.n659 avss.n658 0.0382424
R24098 avss.n734 avss.n733 0.0382424
R24099 avss.n857 avss.n856 0.0382424
R24100 avss.n791 avss.n790 0.0382424
R24101 avss.n443 avss.n442 0.0382424
R24102 avss.n518 avss.n517 0.0382424
R24103 avss.n641 avss.n640 0.0382424
R24104 avss.n575 avss.n574 0.0382424
R24105 avss.n11306 avss.n11305 0.0382424
R24106 avss.n11347 avss.n11346 0.0382424
R24107 avss.n316 avss.n315 0.0382424
R24108 avss.n250 avss.n249 0.0382424
R24109 avss.n11527 avss.n11526 0.0382424
R24110 avss.n11568 avss.n11567 0.0382424
R24111 avss.n99 avss.n98 0.0382424
R24112 avss.n33 avss.n32 0.0382424
R24113 avss.n3510 avss.n3508 0.038
R24114 avss.n3363 avss.n3285 0.0364375
R24115 avss.n4731 avss 0.0356562
R24116 avss.n3607 avss.n3606 0.0352676
R24117 avss.n3537 avss.n3149 0.0352676
R24118 avss.n8806 avss.n8670 0.0339697
R24119 avss.n8765 avss.n8745 0.0339697
R24120 avss.n8877 avss.n3706 0.0339697
R24121 avss.n8966 avss.n3680 0.0339697
R24122 avss.n8453 avss.n8317 0.0339697
R24123 avss.n8412 avss.n8392 0.0339697
R24124 avss.n8524 avss.n3790 0.0339697
R24125 avss.n8613 avss.n3764 0.0339697
R24126 avss.n8100 avss.n7964 0.0339697
R24127 avss.n8059 avss.n8039 0.0339697
R24128 avss.n8171 avss.n3874 0.0339697
R24129 avss.n8260 avss.n3848 0.0339697
R24130 avss.n7747 avss.n7611 0.0339697
R24131 avss.n7706 avss.n7686 0.0339697
R24132 avss.n7818 avss.n3958 0.0339697
R24133 avss.n7907 avss.n3932 0.0339697
R24134 avss.n7394 avss.n7258 0.0339697
R24135 avss.n7353 avss.n7333 0.0339697
R24136 avss.n7465 avss.n4042 0.0339697
R24137 avss.n7554 avss.n4016 0.0339697
R24138 avss.n7041 avss.n6905 0.0339697
R24139 avss.n7000 avss.n6980 0.0339697
R24140 avss.n7112 avss.n4126 0.0339697
R24141 avss.n7201 avss.n4100 0.0339697
R24142 avss.n6688 avss.n6552 0.0339697
R24143 avss.n6647 avss.n6627 0.0339697
R24144 avss.n6759 avss.n4210 0.0339697
R24145 avss.n6848 avss.n4184 0.0339697
R24146 avss.n6335 avss.n6199 0.0339697
R24147 avss.n6294 avss.n6274 0.0339697
R24148 avss.n6406 avss.n4294 0.0339697
R24149 avss.n6495 avss.n4268 0.0339697
R24150 avss.n5982 avss.n5846 0.0339697
R24151 avss.n5941 avss.n5921 0.0339697
R24152 avss.n6053 avss.n4378 0.0339697
R24153 avss.n6142 avss.n4352 0.0339697
R24154 avss.n5629 avss.n5493 0.0339697
R24155 avss.n5588 avss.n5568 0.0339697
R24156 avss.n5700 avss.n4462 0.0339697
R24157 avss.n5789 avss.n4436 0.0339697
R24158 avss.n5284 avss.n5147 0.0339697
R24159 avss.n5230 avss.n5229 0.0339697
R24160 avss.n5347 avss.n4546 0.0339697
R24161 avss.n5436 avss.n4520 0.0339697
R24162 avss.n4930 avss.n4793 0.0339697
R24163 avss.n4876 avss.n4875 0.0339697
R24164 avss.n4993 avss.n4630 0.0339697
R24165 avss.n5082 avss.n4604 0.0339697
R24166 avss.n2447 avss.n2446 0.0339697
R24167 avss.n2504 avss.n2503 0.0339697
R24168 avss.n2231 avss.n2230 0.0339697
R24169 avss.n2288 avss.n2287 0.0339697
R24170 avss.n2015 avss.n2014 0.0339697
R24171 avss.n2072 avss.n2071 0.0339697
R24172 avss.n1799 avss.n1798 0.0339697
R24173 avss.n1856 avss.n1855 0.0339697
R24174 avss.n1583 avss.n1582 0.0339697
R24175 avss.n1640 avss.n1639 0.0339697
R24176 avss.n1367 avss.n1366 0.0339697
R24177 avss.n1424 avss.n1423 0.0339697
R24178 avss.n1151 avss.n1150 0.0339697
R24179 avss.n1208 avss.n1207 0.0339697
R24180 avss.n935 avss.n934 0.0339697
R24181 avss.n992 avss.n991 0.0339697
R24182 avss.n719 avss.n718 0.0339697
R24183 avss.n776 avss.n775 0.0339697
R24184 avss.n503 avss.n502 0.0339697
R24185 avss.n560 avss.n559 0.0339697
R24186 avss.n11332 avss.n11331 0.0339697
R24187 avss.n235 avss.n234 0.0339697
R24188 avss.n11553 avss.n11552 0.0339697
R24189 avss.n18 avss.n17 0.0339697
R24190 avss.n3362 avss.n3286 0.0338333
R24191 avss.n3362 avss.n3284 0.0338333
R24192 avss.n8768 avss.n8744 0.032697
R24193 avss.n8737 avss.n8736 0.032697
R24194 avss.n8789 avss.n8706 0.032697
R24195 avss.n8802 avss.n8679 0.032697
R24196 avss.n8675 avss.n8672 0.032697
R24197 avss.n8658 avss.n8656 0.032697
R24198 avss.n8830 avss.n8829 0.032697
R24199 avss.n3750 avss.n3749 0.032697
R24200 avss.n8852 avss.n8851 0.032697
R24201 avss.n8872 avss.n8871 0.032697
R24202 avss.n8882 avss.n8881 0.032697
R24203 avss.n8919 avss.n8918 0.032697
R24204 avss.n8936 avss.n3684 0.032697
R24205 avss.n8949 avss.n8946 0.032697
R24206 avss.n8415 avss.n8391 0.032697
R24207 avss.n8384 avss.n8383 0.032697
R24208 avss.n8436 avss.n8353 0.032697
R24209 avss.n8449 avss.n8326 0.032697
R24210 avss.n8322 avss.n8319 0.032697
R24211 avss.n8305 avss.n8303 0.032697
R24212 avss.n8477 avss.n8476 0.032697
R24213 avss.n3834 avss.n3833 0.032697
R24214 avss.n8499 avss.n8498 0.032697
R24215 avss.n8519 avss.n8518 0.032697
R24216 avss.n8529 avss.n8528 0.032697
R24217 avss.n8566 avss.n8565 0.032697
R24218 avss.n8583 avss.n3768 0.032697
R24219 avss.n8596 avss.n8593 0.032697
R24220 avss.n8062 avss.n8038 0.032697
R24221 avss.n8031 avss.n8030 0.032697
R24222 avss.n8083 avss.n8000 0.032697
R24223 avss.n8096 avss.n7973 0.032697
R24224 avss.n7969 avss.n7966 0.032697
R24225 avss.n7952 avss.n7950 0.032697
R24226 avss.n8124 avss.n8123 0.032697
R24227 avss.n3918 avss.n3917 0.032697
R24228 avss.n8146 avss.n8145 0.032697
R24229 avss.n8166 avss.n8165 0.032697
R24230 avss.n8176 avss.n8175 0.032697
R24231 avss.n8213 avss.n8212 0.032697
R24232 avss.n8230 avss.n3852 0.032697
R24233 avss.n8243 avss.n8240 0.032697
R24234 avss.n7709 avss.n7685 0.032697
R24235 avss.n7678 avss.n7677 0.032697
R24236 avss.n7730 avss.n7647 0.032697
R24237 avss.n7743 avss.n7620 0.032697
R24238 avss.n7616 avss.n7613 0.032697
R24239 avss.n7599 avss.n7597 0.032697
R24240 avss.n7771 avss.n7770 0.032697
R24241 avss.n4002 avss.n4001 0.032697
R24242 avss.n7793 avss.n7792 0.032697
R24243 avss.n7813 avss.n7812 0.032697
R24244 avss.n7823 avss.n7822 0.032697
R24245 avss.n7860 avss.n7859 0.032697
R24246 avss.n7877 avss.n3936 0.032697
R24247 avss.n7890 avss.n7887 0.032697
R24248 avss.n7356 avss.n7332 0.032697
R24249 avss.n7325 avss.n7324 0.032697
R24250 avss.n7377 avss.n7294 0.032697
R24251 avss.n7390 avss.n7267 0.032697
R24252 avss.n7263 avss.n7260 0.032697
R24253 avss.n7246 avss.n7244 0.032697
R24254 avss.n7418 avss.n7417 0.032697
R24255 avss.n4086 avss.n4085 0.032697
R24256 avss.n7440 avss.n7439 0.032697
R24257 avss.n7460 avss.n7459 0.032697
R24258 avss.n7470 avss.n7469 0.032697
R24259 avss.n7507 avss.n7506 0.032697
R24260 avss.n7524 avss.n4020 0.032697
R24261 avss.n7537 avss.n7534 0.032697
R24262 avss.n7003 avss.n6979 0.032697
R24263 avss.n6972 avss.n6971 0.032697
R24264 avss.n7024 avss.n6941 0.032697
R24265 avss.n7037 avss.n6914 0.032697
R24266 avss.n6910 avss.n6907 0.032697
R24267 avss.n6893 avss.n6891 0.032697
R24268 avss.n7065 avss.n7064 0.032697
R24269 avss.n4170 avss.n4169 0.032697
R24270 avss.n7087 avss.n7086 0.032697
R24271 avss.n7107 avss.n7106 0.032697
R24272 avss.n7117 avss.n7116 0.032697
R24273 avss.n7154 avss.n7153 0.032697
R24274 avss.n7171 avss.n4104 0.032697
R24275 avss.n7184 avss.n7181 0.032697
R24276 avss.n6650 avss.n6626 0.032697
R24277 avss.n6619 avss.n6618 0.032697
R24278 avss.n6671 avss.n6588 0.032697
R24279 avss.n6684 avss.n6561 0.032697
R24280 avss.n6557 avss.n6554 0.032697
R24281 avss.n6540 avss.n6538 0.032697
R24282 avss.n6712 avss.n6711 0.032697
R24283 avss.n4254 avss.n4253 0.032697
R24284 avss.n6734 avss.n6733 0.032697
R24285 avss.n6754 avss.n6753 0.032697
R24286 avss.n6764 avss.n6763 0.032697
R24287 avss.n6801 avss.n6800 0.032697
R24288 avss.n6818 avss.n4188 0.032697
R24289 avss.n6831 avss.n6828 0.032697
R24290 avss.n6297 avss.n6273 0.032697
R24291 avss.n6266 avss.n6265 0.032697
R24292 avss.n6318 avss.n6235 0.032697
R24293 avss.n6331 avss.n6208 0.032697
R24294 avss.n6204 avss.n6201 0.032697
R24295 avss.n6187 avss.n6185 0.032697
R24296 avss.n6359 avss.n6358 0.032697
R24297 avss.n4338 avss.n4337 0.032697
R24298 avss.n6381 avss.n6380 0.032697
R24299 avss.n6401 avss.n6400 0.032697
R24300 avss.n6411 avss.n6410 0.032697
R24301 avss.n6448 avss.n6447 0.032697
R24302 avss.n6465 avss.n4272 0.032697
R24303 avss.n6478 avss.n6475 0.032697
R24304 avss.n5944 avss.n5920 0.032697
R24305 avss.n5913 avss.n5912 0.032697
R24306 avss.n5965 avss.n5882 0.032697
R24307 avss.n5978 avss.n5855 0.032697
R24308 avss.n5851 avss.n5848 0.032697
R24309 avss.n5834 avss.n5832 0.032697
R24310 avss.n6006 avss.n6005 0.032697
R24311 avss.n4422 avss.n4421 0.032697
R24312 avss.n6028 avss.n6027 0.032697
R24313 avss.n6048 avss.n6047 0.032697
R24314 avss.n6058 avss.n6057 0.032697
R24315 avss.n6095 avss.n6094 0.032697
R24316 avss.n6112 avss.n4356 0.032697
R24317 avss.n6125 avss.n6122 0.032697
R24318 avss.n5591 avss.n5567 0.032697
R24319 avss.n5560 avss.n5559 0.032697
R24320 avss.n5612 avss.n5529 0.032697
R24321 avss.n5625 avss.n5502 0.032697
R24322 avss.n5498 avss.n5495 0.032697
R24323 avss.n5481 avss.n5479 0.032697
R24324 avss.n5653 avss.n5652 0.032697
R24325 avss.n4506 avss.n4505 0.032697
R24326 avss.n5675 avss.n5674 0.032697
R24327 avss.n5695 avss.n5694 0.032697
R24328 avss.n5705 avss.n5704 0.032697
R24329 avss.n5742 avss.n5741 0.032697
R24330 avss.n5759 avss.n4440 0.032697
R24331 avss.n5772 avss.n5769 0.032697
R24332 avss.n5248 avss.n5247 0.032697
R24333 avss.n5220 avss.n5219 0.032697
R24334 avss.n5267 avss.n5183 0.032697
R24335 avss.n5280 avss.n5156 0.032697
R24336 avss.n5152 avss.n5149 0.032697
R24337 avss.n5295 avss.n5294 0.032697
R24338 avss.n5124 avss.n5123 0.032697
R24339 avss.n4590 avss.n4589 0.032697
R24340 avss.n5322 avss.n5321 0.032697
R24341 avss.n5342 avss.n5341 0.032697
R24342 avss.n5352 avss.n5351 0.032697
R24343 avss.n5389 avss.n5388 0.032697
R24344 avss.n5406 avss.n4524 0.032697
R24345 avss.n5419 avss.n5416 0.032697
R24346 avss.n4894 avss.n4893 0.032697
R24347 avss.n4866 avss.n4865 0.032697
R24348 avss.n4913 avss.n4829 0.032697
R24349 avss.n4926 avss.n4802 0.032697
R24350 avss.n4798 avss.n4795 0.032697
R24351 avss.n4941 avss.n4940 0.032697
R24352 avss.n4770 avss.n4769 0.032697
R24353 avss.n4674 avss.n4673 0.032697
R24354 avss.n4968 avss.n4967 0.032697
R24355 avss.n4988 avss.n4987 0.032697
R24356 avss.n4998 avss.n4997 0.032697
R24357 avss.n5035 avss.n5034 0.032697
R24358 avss.n5052 avss.n4608 0.032697
R24359 avss.n5065 avss.n5062 0.032697
R24360 avss.n9113 avss.n9112 0.032697
R24361 avss.n9168 avss.n9167 0.032697
R24362 avss.n9148 avss.n9144 0.032697
R24363 avss.n2441 avss.n2435 0.032697
R24364 avss.n2456 avss.n2455 0.032697
R24365 avss.n2476 avss.n2475 0.032697
R24366 avss.n2405 avss.n2401 0.032697
R24367 avss.n2552 avss.n2548 0.032697
R24368 avss.n2533 avss.n2532 0.032697
R24369 avss.n2513 avss.n2512 0.032697
R24370 avss.n2498 avss.n2492 0.032697
R24371 avss.n9037 avss.n9033 0.032697
R24372 avss.n9057 avss.n9056 0.032697
R24373 avss.n9001 avss.n9000 0.032697
R24374 avss.n9334 avss.n9333 0.032697
R24375 avss.n9389 avss.n9388 0.032697
R24376 avss.n9369 avss.n9365 0.032697
R24377 avss.n2225 avss.n2219 0.032697
R24378 avss.n2240 avss.n2239 0.032697
R24379 avss.n2260 avss.n2259 0.032697
R24380 avss.n2189 avss.n2185 0.032697
R24381 avss.n2336 avss.n2332 0.032697
R24382 avss.n2317 avss.n2316 0.032697
R24383 avss.n2297 avss.n2296 0.032697
R24384 avss.n2282 avss.n2276 0.032697
R24385 avss.n9258 avss.n9254 0.032697
R24386 avss.n9278 avss.n9277 0.032697
R24387 avss.n9222 avss.n9221 0.032697
R24388 avss.n9555 avss.n9554 0.032697
R24389 avss.n9610 avss.n9609 0.032697
R24390 avss.n9590 avss.n9586 0.032697
R24391 avss.n2009 avss.n2003 0.032697
R24392 avss.n2024 avss.n2023 0.032697
R24393 avss.n2044 avss.n2043 0.032697
R24394 avss.n1973 avss.n1969 0.032697
R24395 avss.n2120 avss.n2116 0.032697
R24396 avss.n2101 avss.n2100 0.032697
R24397 avss.n2081 avss.n2080 0.032697
R24398 avss.n2066 avss.n2060 0.032697
R24399 avss.n9479 avss.n9475 0.032697
R24400 avss.n9499 avss.n9498 0.032697
R24401 avss.n9443 avss.n9442 0.032697
R24402 avss.n9776 avss.n9775 0.032697
R24403 avss.n9831 avss.n9830 0.032697
R24404 avss.n9811 avss.n9807 0.032697
R24405 avss.n1793 avss.n1787 0.032697
R24406 avss.n1808 avss.n1807 0.032697
R24407 avss.n1828 avss.n1827 0.032697
R24408 avss.n1757 avss.n1753 0.032697
R24409 avss.n1904 avss.n1900 0.032697
R24410 avss.n1885 avss.n1884 0.032697
R24411 avss.n1865 avss.n1864 0.032697
R24412 avss.n1850 avss.n1844 0.032697
R24413 avss.n9700 avss.n9696 0.032697
R24414 avss.n9720 avss.n9719 0.032697
R24415 avss.n9664 avss.n9663 0.032697
R24416 avss.n9997 avss.n9996 0.032697
R24417 avss.n10052 avss.n10051 0.032697
R24418 avss.n10032 avss.n10028 0.032697
R24419 avss.n1577 avss.n1571 0.032697
R24420 avss.n1592 avss.n1591 0.032697
R24421 avss.n1612 avss.n1611 0.032697
R24422 avss.n1541 avss.n1537 0.032697
R24423 avss.n1688 avss.n1684 0.032697
R24424 avss.n1669 avss.n1668 0.032697
R24425 avss.n1649 avss.n1648 0.032697
R24426 avss.n1634 avss.n1628 0.032697
R24427 avss.n9921 avss.n9917 0.032697
R24428 avss.n9941 avss.n9940 0.032697
R24429 avss.n9885 avss.n9884 0.032697
R24430 avss.n10218 avss.n10217 0.032697
R24431 avss.n10273 avss.n10272 0.032697
R24432 avss.n10253 avss.n10249 0.032697
R24433 avss.n1361 avss.n1355 0.032697
R24434 avss.n1376 avss.n1375 0.032697
R24435 avss.n1396 avss.n1395 0.032697
R24436 avss.n1325 avss.n1321 0.032697
R24437 avss.n1472 avss.n1468 0.032697
R24438 avss.n1453 avss.n1452 0.032697
R24439 avss.n1433 avss.n1432 0.032697
R24440 avss.n1418 avss.n1412 0.032697
R24441 avss.n10142 avss.n10138 0.032697
R24442 avss.n10162 avss.n10161 0.032697
R24443 avss.n10106 avss.n10105 0.032697
R24444 avss.n10439 avss.n10438 0.032697
R24445 avss.n10494 avss.n10493 0.032697
R24446 avss.n10474 avss.n10470 0.032697
R24447 avss.n1145 avss.n1139 0.032697
R24448 avss.n1160 avss.n1159 0.032697
R24449 avss.n1180 avss.n1179 0.032697
R24450 avss.n1109 avss.n1105 0.032697
R24451 avss.n1256 avss.n1252 0.032697
R24452 avss.n1237 avss.n1236 0.032697
R24453 avss.n1217 avss.n1216 0.032697
R24454 avss.n1202 avss.n1196 0.032697
R24455 avss.n10363 avss.n10359 0.032697
R24456 avss.n10383 avss.n10382 0.032697
R24457 avss.n10327 avss.n10326 0.032697
R24458 avss.n10660 avss.n10659 0.032697
R24459 avss.n10715 avss.n10714 0.032697
R24460 avss.n10695 avss.n10691 0.032697
R24461 avss.n929 avss.n923 0.032697
R24462 avss.n944 avss.n943 0.032697
R24463 avss.n964 avss.n963 0.032697
R24464 avss.n893 avss.n889 0.032697
R24465 avss.n1040 avss.n1036 0.032697
R24466 avss.n1021 avss.n1020 0.032697
R24467 avss.n1001 avss.n1000 0.032697
R24468 avss.n986 avss.n980 0.032697
R24469 avss.n10584 avss.n10580 0.032697
R24470 avss.n10604 avss.n10603 0.032697
R24471 avss.n10548 avss.n10547 0.032697
R24472 avss.n10881 avss.n10880 0.032697
R24473 avss.n10936 avss.n10935 0.032697
R24474 avss.n10916 avss.n10912 0.032697
R24475 avss.n713 avss.n707 0.032697
R24476 avss.n728 avss.n727 0.032697
R24477 avss.n748 avss.n747 0.032697
R24478 avss.n677 avss.n673 0.032697
R24479 avss.n824 avss.n820 0.032697
R24480 avss.n805 avss.n804 0.032697
R24481 avss.n785 avss.n784 0.032697
R24482 avss.n770 avss.n764 0.032697
R24483 avss.n10805 avss.n10801 0.032697
R24484 avss.n10825 avss.n10824 0.032697
R24485 avss.n10769 avss.n10768 0.032697
R24486 avss.n11102 avss.n11101 0.032697
R24487 avss.n11157 avss.n11156 0.032697
R24488 avss.n11137 avss.n11133 0.032697
R24489 avss.n497 avss.n491 0.032697
R24490 avss.n512 avss.n511 0.032697
R24491 avss.n532 avss.n531 0.032697
R24492 avss.n461 avss.n457 0.032697
R24493 avss.n608 avss.n604 0.032697
R24494 avss.n589 avss.n588 0.032697
R24495 avss.n569 avss.n568 0.032697
R24496 avss.n554 avss.n548 0.032697
R24497 avss.n11026 avss.n11022 0.032697
R24498 avss.n11046 avss.n11045 0.032697
R24499 avss.n10990 avss.n10989 0.032697
R24500 avss.n368 avss.n367 0.032697
R24501 avss.n424 avss.n423 0.032697
R24502 avss.n404 avss.n400 0.032697
R24503 avss.n11326 avss.n11320 0.032697
R24504 avss.n11341 avss.n11340 0.032697
R24505 avss.n11361 avss.n11360 0.032697
R24506 avss.n11379 avss.n11375 0.032697
R24507 avss.n283 avss.n279 0.032697
R24508 avss.n264 avss.n263 0.032697
R24509 avss.n244 avss.n243 0.032697
R24510 avss.n229 avss.n223 0.032697
R24511 avss.n11247 avss.n11243 0.032697
R24512 avss.n11267 avss.n11266 0.032697
R24513 avss.n11211 avss.n11210 0.032697
R24514 avss.n151 avss.n150 0.032697
R24515 avss.n207 avss.n206 0.032697
R24516 avss.n187 avss.n183 0.032697
R24517 avss.n11547 avss.n11541 0.032697
R24518 avss.n11562 avss.n11561 0.032697
R24519 avss.n11582 avss.n11581 0.032697
R24520 avss.n11600 avss.n11596 0.032697
R24521 avss.n66 avss.n62 0.032697
R24522 avss.n47 avss.n46 0.032697
R24523 avss.n27 avss.n26 0.032697
R24524 avss.n12 avss.n6 0.032697
R24525 avss.n11468 avss.n11464 0.032697
R24526 avss.n11488 avss.n11487 0.032697
R24527 avss.n11432 avss.n11431 0.032697
R24528 avss.n8805 avss.n8804 0.0325455
R24529 avss.n8760 avss.n8749 0.0325455
R24530 avss.n8879 avss.n8878 0.0325455
R24531 avss.n8965 avss.n8964 0.0325455
R24532 avss.n8452 avss.n8451 0.0325455
R24533 avss.n8407 avss.n8396 0.0325455
R24534 avss.n8526 avss.n8525 0.0325455
R24535 avss.n8612 avss.n8611 0.0325455
R24536 avss.n8099 avss.n8098 0.0325455
R24537 avss.n8054 avss.n8043 0.0325455
R24538 avss.n8173 avss.n8172 0.0325455
R24539 avss.n8259 avss.n8258 0.0325455
R24540 avss.n7746 avss.n7745 0.0325455
R24541 avss.n7701 avss.n7690 0.0325455
R24542 avss.n7820 avss.n7819 0.0325455
R24543 avss.n7906 avss.n7905 0.0325455
R24544 avss.n7393 avss.n7392 0.0325455
R24545 avss.n7348 avss.n7337 0.0325455
R24546 avss.n7467 avss.n7466 0.0325455
R24547 avss.n7553 avss.n7552 0.0325455
R24548 avss.n7040 avss.n7039 0.0325455
R24549 avss.n6995 avss.n6984 0.0325455
R24550 avss.n7114 avss.n7113 0.0325455
R24551 avss.n7200 avss.n7199 0.0325455
R24552 avss.n6687 avss.n6686 0.0325455
R24553 avss.n6642 avss.n6631 0.0325455
R24554 avss.n6761 avss.n6760 0.0325455
R24555 avss.n6847 avss.n6846 0.0325455
R24556 avss.n6334 avss.n6333 0.0325455
R24557 avss.n6289 avss.n6278 0.0325455
R24558 avss.n6408 avss.n6407 0.0325455
R24559 avss.n6494 avss.n6493 0.0325455
R24560 avss.n5981 avss.n5980 0.0325455
R24561 avss.n5936 avss.n5925 0.0325455
R24562 avss.n6055 avss.n6054 0.0325455
R24563 avss.n6141 avss.n6140 0.0325455
R24564 avss.n5628 avss.n5627 0.0325455
R24565 avss.n5583 avss.n5572 0.0325455
R24566 avss.n5702 avss.n5701 0.0325455
R24567 avss.n5788 avss.n5787 0.0325455
R24568 avss.n5283 avss.n5282 0.0325455
R24569 avss.n5242 avss.n5231 0.0325455
R24570 avss.n5349 avss.n5348 0.0325455
R24571 avss.n5435 avss.n5434 0.0325455
R24572 avss.n4929 avss.n4928 0.0325455
R24573 avss.n4888 avss.n4877 0.0325455
R24574 avss.n4995 avss.n4994 0.0325455
R24575 avss.n5081 avss.n5080 0.0325455
R24576 avss.n2445 avss.n2444 0.0325455
R24577 avss.n9087 avss.n9086 0.0325455
R24578 avss.n2502 avss.n2501 0.0325455
R24579 avss.n9067 avss.n9066 0.0325455
R24580 avss.n2229 avss.n2228 0.0325455
R24581 avss.n9308 avss.n9307 0.0325455
R24582 avss.n2286 avss.n2285 0.0325455
R24583 avss.n9288 avss.n9287 0.0325455
R24584 avss.n2013 avss.n2012 0.0325455
R24585 avss.n9529 avss.n9528 0.0325455
R24586 avss.n2070 avss.n2069 0.0325455
R24587 avss.n9509 avss.n9508 0.0325455
R24588 avss.n1797 avss.n1796 0.0325455
R24589 avss.n9750 avss.n9749 0.0325455
R24590 avss.n1854 avss.n1853 0.0325455
R24591 avss.n9730 avss.n9729 0.0325455
R24592 avss.n1581 avss.n1580 0.0325455
R24593 avss.n9971 avss.n9970 0.0325455
R24594 avss.n1638 avss.n1637 0.0325455
R24595 avss.n9951 avss.n9950 0.0325455
R24596 avss.n1365 avss.n1364 0.0325455
R24597 avss.n10192 avss.n10191 0.0325455
R24598 avss.n1422 avss.n1421 0.0325455
R24599 avss.n10172 avss.n10171 0.0325455
R24600 avss.n1149 avss.n1148 0.0325455
R24601 avss.n10413 avss.n10412 0.0325455
R24602 avss.n1206 avss.n1205 0.0325455
R24603 avss.n10393 avss.n10392 0.0325455
R24604 avss.n933 avss.n932 0.0325455
R24605 avss.n10634 avss.n10633 0.0325455
R24606 avss.n990 avss.n989 0.0325455
R24607 avss.n10614 avss.n10613 0.0325455
R24608 avss.n717 avss.n716 0.0325455
R24609 avss.n10855 avss.n10854 0.0325455
R24610 avss.n774 avss.n773 0.0325455
R24611 avss.n10835 avss.n10834 0.0325455
R24612 avss.n501 avss.n500 0.0325455
R24613 avss.n11076 avss.n11075 0.0325455
R24614 avss.n558 avss.n557 0.0325455
R24615 avss.n11056 avss.n11055 0.0325455
R24616 avss.n11330 avss.n11329 0.0325455
R24617 avss.n327 avss.n326 0.0325455
R24618 avss.n233 avss.n232 0.0325455
R24619 avss.n11277 avss.n11276 0.0325455
R24620 avss.n11551 avss.n11550 0.0325455
R24621 avss.n110 avss.n109 0.0325455
R24622 avss.n16 avss.n15 0.0325455
R24623 avss.n11498 avss.n11497 0.0325455
R24624 avss.n8834 avss.n8833 0.0320239
R24625 avss.n8481 avss.n8480 0.0320239
R24626 avss.n8128 avss.n8127 0.0320239
R24627 avss.n7775 avss.n7774 0.0320239
R24628 avss.n7422 avss.n7421 0.0320239
R24629 avss.n7069 avss.n7068 0.0320239
R24630 avss.n6716 avss.n6715 0.0320239
R24631 avss.n6363 avss.n6362 0.0320239
R24632 avss.n6010 avss.n6009 0.0320239
R24633 avss.n5657 avss.n5656 0.0320239
R24634 avss.n8838 avss.n3725 0.0317611
R24635 avss.n8485 avss.n3809 0.0317611
R24636 avss.n8132 avss.n3893 0.0317611
R24637 avss.n7779 avss.n3977 0.0317611
R24638 avss.n7426 avss.n4061 0.0317611
R24639 avss.n7073 avss.n4145 0.0317611
R24640 avss.n6720 avss.n4229 0.0317611
R24641 avss.n6367 avss.n4313 0.0317611
R24642 avss.n6014 avss.n4397 0.0317611
R24643 avss.n5661 avss.n4481 0.0317611
R24644 avss.n5308 avss.n4565 0.0317611
R24645 avss.n4954 avss.n4649 0.0317611
R24646 avss.n2556 avss.n2555 0.0317611
R24647 avss.n2340 avss.n2339 0.0317611
R24648 avss.n2124 avss.n2123 0.0317611
R24649 avss.n1908 avss.n1907 0.0317611
R24650 avss.n1692 avss.n1691 0.0317611
R24651 avss.n1476 avss.n1475 0.0317611
R24652 avss.n1260 avss.n1259 0.0317611
R24653 avss.n1044 avss.n1043 0.0317611
R24654 avss.n828 avss.n827 0.0317611
R24655 avss.n612 avss.n611 0.0317611
R24656 avss.n287 avss.n286 0.0317611
R24657 avss.n70 avss.n69 0.0317611
R24658 avss.n3349 avss.n3348 0.03175
R24659 avss.n3350 avss.n3285 0.03175
R24660 avss.n3513 avss.n3175 0.03175
R24661 avss.n3512 avss.n3511 0.03175
R24662 avss.n3338 avss.n3294 0.03175
R24663 avss.n3413 avss.n3409 0.03175
R24664 avss.n3452 avss.n3199 0.03175
R24665 avss.n8770 avss.n8769 0.030803
R24666 avss.n8812 avss.n8661 0.030803
R24667 avss.n8873 avss.n3710 0.030803
R24668 avss.n8945 avss.n8944 0.030803
R24669 avss.n8417 avss.n8416 0.030803
R24670 avss.n8459 avss.n8308 0.030803
R24671 avss.n8520 avss.n3794 0.030803
R24672 avss.n8592 avss.n8591 0.030803
R24673 avss.n8064 avss.n8063 0.030803
R24674 avss.n8106 avss.n7955 0.030803
R24675 avss.n8167 avss.n3878 0.030803
R24676 avss.n8239 avss.n8238 0.030803
R24677 avss.n7711 avss.n7710 0.030803
R24678 avss.n7753 avss.n7602 0.030803
R24679 avss.n7814 avss.n3962 0.030803
R24680 avss.n7886 avss.n7885 0.030803
R24681 avss.n7358 avss.n7357 0.030803
R24682 avss.n7400 avss.n7249 0.030803
R24683 avss.n7461 avss.n4046 0.030803
R24684 avss.n7533 avss.n7532 0.030803
R24685 avss.n7005 avss.n7004 0.030803
R24686 avss.n7047 avss.n6896 0.030803
R24687 avss.n7108 avss.n4130 0.030803
R24688 avss.n7180 avss.n7179 0.030803
R24689 avss.n6652 avss.n6651 0.030803
R24690 avss.n6694 avss.n6543 0.030803
R24691 avss.n6755 avss.n4214 0.030803
R24692 avss.n6827 avss.n6826 0.030803
R24693 avss.n6299 avss.n6298 0.030803
R24694 avss.n6341 avss.n6190 0.030803
R24695 avss.n6402 avss.n4298 0.030803
R24696 avss.n6474 avss.n6473 0.030803
R24697 avss.n5946 avss.n5945 0.030803
R24698 avss.n5988 avss.n5837 0.030803
R24699 avss.n6049 avss.n4382 0.030803
R24700 avss.n6121 avss.n6120 0.030803
R24701 avss.n5593 avss.n5592 0.030803
R24702 avss.n5635 avss.n5484 0.030803
R24703 avss.n5696 avss.n4466 0.030803
R24704 avss.n5768 avss.n5767 0.030803
R24705 avss.n5249 avss.n5209 0.030803
R24706 avss.n5290 avss.n5134 0.030803
R24707 avss.n5343 avss.n4550 0.030803
R24708 avss.n5415 avss.n5414 0.030803
R24709 avss.n4895 avss.n4855 0.030803
R24710 avss.n4936 avss.n4780 0.030803
R24711 avss.n4989 avss.n4634 0.030803
R24712 avss.n5061 avss.n5060 0.030803
R24713 avss.n9110 avss.n9109 0.030803
R24714 avss.n2453 avss.n2452 0.030803
R24715 avss.n2510 avss.n2509 0.030803
R24716 avss.n8998 avss.n8997 0.030803
R24717 avss.n9331 avss.n9330 0.030803
R24718 avss.n2237 avss.n2236 0.030803
R24719 avss.n2294 avss.n2293 0.030803
R24720 avss.n9219 avss.n9218 0.030803
R24721 avss.n9552 avss.n9551 0.030803
R24722 avss.n2021 avss.n2020 0.030803
R24723 avss.n2078 avss.n2077 0.030803
R24724 avss.n9440 avss.n9439 0.030803
R24725 avss.n9773 avss.n9772 0.030803
R24726 avss.n1805 avss.n1804 0.030803
R24727 avss.n1862 avss.n1861 0.030803
R24728 avss.n9661 avss.n9660 0.030803
R24729 avss.n9994 avss.n9993 0.030803
R24730 avss.n1589 avss.n1588 0.030803
R24731 avss.n1646 avss.n1645 0.030803
R24732 avss.n9882 avss.n9881 0.030803
R24733 avss.n10215 avss.n10214 0.030803
R24734 avss.n1373 avss.n1372 0.030803
R24735 avss.n1430 avss.n1429 0.030803
R24736 avss.n10103 avss.n10102 0.030803
R24737 avss.n10436 avss.n10435 0.030803
R24738 avss.n1157 avss.n1156 0.030803
R24739 avss.n1214 avss.n1213 0.030803
R24740 avss.n10324 avss.n10323 0.030803
R24741 avss.n10657 avss.n10656 0.030803
R24742 avss.n941 avss.n940 0.030803
R24743 avss.n998 avss.n997 0.030803
R24744 avss.n10545 avss.n10544 0.030803
R24745 avss.n10878 avss.n10877 0.030803
R24746 avss.n725 avss.n724 0.030803
R24747 avss.n782 avss.n781 0.030803
R24748 avss.n10766 avss.n10765 0.030803
R24749 avss.n11099 avss.n11098 0.030803
R24750 avss.n509 avss.n508 0.030803
R24751 avss.n566 avss.n565 0.030803
R24752 avss.n10987 avss.n10986 0.030803
R24753 avss.n365 avss.n364 0.030803
R24754 avss.n11338 avss.n11337 0.030803
R24755 avss.n241 avss.n240 0.030803
R24756 avss.n11208 avss.n11207 0.030803
R24757 avss.n148 avss.n147 0.030803
R24758 avss.n11559 avss.n11558 0.030803
R24759 avss.n24 avss.n23 0.030803
R24760 avss.n11429 avss.n11428 0.030803
R24761 avss.n2977 avss.n2960 0.0304479
R24762 avss.n3034 avss.n2944 0.0304479
R24763 avss.n3134 avss.n3133 0.0304479
R24764 avss.n3626 avss.n2610 0.0304479
R24765 avss.n2689 avss.n2673 0.0304479
R24766 avss.n2734 avss.n2646 0.0304479
R24767 avss.n2630 avss.n2629 0.0304479
R24768 avss.n2867 avss.n2794 0.0304479
R24769 avss.n3456 avss.n3197 0.0296667
R24770 avss.n3461 avss.n3195 0.0296667
R24771 avss.n8785 avss.n8784 0.0289091
R24772 avss.n8828 avss.n8825 0.0289091
R24773 avss.n3748 avss.n3721 0.0289091
R24774 avss.n8917 avss.n3686 0.0289091
R24775 avss.n8432 avss.n8431 0.0289091
R24776 avss.n8475 avss.n8472 0.0289091
R24777 avss.n3832 avss.n3805 0.0289091
R24778 avss.n8564 avss.n3770 0.0289091
R24779 avss.n8079 avss.n8078 0.0289091
R24780 avss.n8122 avss.n8119 0.0289091
R24781 avss.n3916 avss.n3889 0.0289091
R24782 avss.n8211 avss.n3854 0.0289091
R24783 avss.n7726 avss.n7725 0.0289091
R24784 avss.n7769 avss.n7766 0.0289091
R24785 avss.n4000 avss.n3973 0.0289091
R24786 avss.n7858 avss.n3938 0.0289091
R24787 avss.n7373 avss.n7372 0.0289091
R24788 avss.n7416 avss.n7413 0.0289091
R24789 avss.n4084 avss.n4057 0.0289091
R24790 avss.n7505 avss.n4022 0.0289091
R24791 avss.n7020 avss.n7019 0.0289091
R24792 avss.n7063 avss.n7060 0.0289091
R24793 avss.n4168 avss.n4141 0.0289091
R24794 avss.n7152 avss.n4106 0.0289091
R24795 avss.n6667 avss.n6666 0.0289091
R24796 avss.n6710 avss.n6707 0.0289091
R24797 avss.n4252 avss.n4225 0.0289091
R24798 avss.n6799 avss.n4190 0.0289091
R24799 avss.n6314 avss.n6313 0.0289091
R24800 avss.n6357 avss.n6354 0.0289091
R24801 avss.n4336 avss.n4309 0.0289091
R24802 avss.n6446 avss.n4274 0.0289091
R24803 avss.n5961 avss.n5960 0.0289091
R24804 avss.n6004 avss.n6001 0.0289091
R24805 avss.n4420 avss.n4393 0.0289091
R24806 avss.n6093 avss.n4358 0.0289091
R24807 avss.n5608 avss.n5607 0.0289091
R24808 avss.n5651 avss.n5648 0.0289091
R24809 avss.n4504 avss.n4477 0.0289091
R24810 avss.n5740 avss.n4442 0.0289091
R24811 avss.n5263 avss.n5262 0.0289091
R24812 avss.n5128 avss.n5100 0.0289091
R24813 avss.n4588 avss.n4561 0.0289091
R24814 avss.n5387 avss.n4526 0.0289091
R24815 avss.n4909 avss.n4908 0.0289091
R24816 avss.n4774 avss.n4746 0.0289091
R24817 avss.n4672 avss.n4645 0.0289091
R24818 avss.n5033 avss.n4610 0.0289091
R24819 avss.n9147 avss.n9146 0.0289091
R24820 avss.n2404 avss.n2403 0.0289091
R24821 avss.n2551 avss.n2550 0.0289091
R24822 avss.n9036 avss.n9035 0.0289091
R24823 avss.n9368 avss.n9367 0.0289091
R24824 avss.n2188 avss.n2187 0.0289091
R24825 avss.n2335 avss.n2334 0.0289091
R24826 avss.n9257 avss.n9256 0.0289091
R24827 avss.n9589 avss.n9588 0.0289091
R24828 avss.n1972 avss.n1971 0.0289091
R24829 avss.n2119 avss.n2118 0.0289091
R24830 avss.n9478 avss.n9477 0.0289091
R24831 avss.n9810 avss.n9809 0.0289091
R24832 avss.n1756 avss.n1755 0.0289091
R24833 avss.n1903 avss.n1902 0.0289091
R24834 avss.n9699 avss.n9698 0.0289091
R24835 avss.n10031 avss.n10030 0.0289091
R24836 avss.n1540 avss.n1539 0.0289091
R24837 avss.n1687 avss.n1686 0.0289091
R24838 avss.n9920 avss.n9919 0.0289091
R24839 avss.n10252 avss.n10251 0.0289091
R24840 avss.n1324 avss.n1323 0.0289091
R24841 avss.n1471 avss.n1470 0.0289091
R24842 avss.n10141 avss.n10140 0.0289091
R24843 avss.n10473 avss.n10472 0.0289091
R24844 avss.n1108 avss.n1107 0.0289091
R24845 avss.n1255 avss.n1254 0.0289091
R24846 avss.n10362 avss.n10361 0.0289091
R24847 avss.n10694 avss.n10693 0.0289091
R24848 avss.n892 avss.n891 0.0289091
R24849 avss.n1039 avss.n1038 0.0289091
R24850 avss.n10583 avss.n10582 0.0289091
R24851 avss.n10915 avss.n10914 0.0289091
R24852 avss.n676 avss.n675 0.0289091
R24853 avss.n823 avss.n822 0.0289091
R24854 avss.n10804 avss.n10803 0.0289091
R24855 avss.n11136 avss.n11135 0.0289091
R24856 avss.n460 avss.n459 0.0289091
R24857 avss.n607 avss.n606 0.0289091
R24858 avss.n11025 avss.n11024 0.0289091
R24859 avss.n403 avss.n402 0.0289091
R24860 avss.n11378 avss.n11377 0.0289091
R24861 avss.n282 avss.n281 0.0289091
R24862 avss.n11246 avss.n11245 0.0289091
R24863 avss.n186 avss.n185 0.0289091
R24864 avss.n11599 avss.n11598 0.0289091
R24865 avss.n65 avss.n64 0.0289091
R24866 avss.n11467 avss.n11466 0.0289091
R24867 avss.n3667 avss.n2594 0.0286927
R24868 avss.n2830 avss.n2829 0.0286927
R24869 avss.n11633 avss.n11628 0.0278438
R24870 avss.n3560 avss 0.0278438
R24871 avss.n3396 avss.n3395 0.0275833
R24872 avss.n3434 avss.n3224 0.0275833
R24873 avss.n3469 avss.n3468 0.0275833
R24874 avss.n3394 avss.n3393 0.0270625
R24875 avss.n8704 avss.n8703 0.0270152
R24876 avss.n8689 avss.n8680 0.0270152
R24877 avss.n8636 avss.n8635 0.0270152
R24878 avss.n3736 avss.n3735 0.0270152
R24879 avss.n8893 avss.n3700 0.0270152
R24880 avss.n8899 avss.n8896 0.0270152
R24881 avss.n8351 avss.n8350 0.0270152
R24882 avss.n8336 avss.n8327 0.0270152
R24883 avss.n8283 avss.n8282 0.0270152
R24884 avss.n3820 avss.n3819 0.0270152
R24885 avss.n8540 avss.n3784 0.0270152
R24886 avss.n8546 avss.n8543 0.0270152
R24887 avss.n7998 avss.n7997 0.0270152
R24888 avss.n7983 avss.n7974 0.0270152
R24889 avss.n7930 avss.n7929 0.0270152
R24890 avss.n3904 avss.n3903 0.0270152
R24891 avss.n8187 avss.n3868 0.0270152
R24892 avss.n8193 avss.n8190 0.0270152
R24893 avss.n7645 avss.n7644 0.0270152
R24894 avss.n7630 avss.n7621 0.0270152
R24895 avss.n7577 avss.n7576 0.0270152
R24896 avss.n3988 avss.n3987 0.0270152
R24897 avss.n7834 avss.n3952 0.0270152
R24898 avss.n7840 avss.n7837 0.0270152
R24899 avss.n7292 avss.n7291 0.0270152
R24900 avss.n7277 avss.n7268 0.0270152
R24901 avss.n7224 avss.n7223 0.0270152
R24902 avss.n4072 avss.n4071 0.0270152
R24903 avss.n7481 avss.n4036 0.0270152
R24904 avss.n7487 avss.n7484 0.0270152
R24905 avss.n6939 avss.n6938 0.0270152
R24906 avss.n6924 avss.n6915 0.0270152
R24907 avss.n6871 avss.n6870 0.0270152
R24908 avss.n4156 avss.n4155 0.0270152
R24909 avss.n7128 avss.n4120 0.0270152
R24910 avss.n7134 avss.n7131 0.0270152
R24911 avss.n6586 avss.n6585 0.0270152
R24912 avss.n6571 avss.n6562 0.0270152
R24913 avss.n6518 avss.n6517 0.0270152
R24914 avss.n4240 avss.n4239 0.0270152
R24915 avss.n6775 avss.n4204 0.0270152
R24916 avss.n6781 avss.n6778 0.0270152
R24917 avss.n6233 avss.n6232 0.0270152
R24918 avss.n6218 avss.n6209 0.0270152
R24919 avss.n6165 avss.n6164 0.0270152
R24920 avss.n4324 avss.n4323 0.0270152
R24921 avss.n6422 avss.n4288 0.0270152
R24922 avss.n6428 avss.n6425 0.0270152
R24923 avss.n5880 avss.n5879 0.0270152
R24924 avss.n5865 avss.n5856 0.0270152
R24925 avss.n5812 avss.n5811 0.0270152
R24926 avss.n4408 avss.n4407 0.0270152
R24927 avss.n6069 avss.n4372 0.0270152
R24928 avss.n6075 avss.n6072 0.0270152
R24929 avss.n5527 avss.n5526 0.0270152
R24930 avss.n5512 avss.n5503 0.0270152
R24931 avss.n5459 avss.n5458 0.0270152
R24932 avss.n4492 avss.n4491 0.0270152
R24933 avss.n5716 avss.n4456 0.0270152
R24934 avss.n5722 avss.n5719 0.0270152
R24935 avss.n5181 avss.n5180 0.0270152
R24936 avss.n5166 avss.n5157 0.0270152
R24937 avss.n5111 avss.n5110 0.0270152
R24938 avss.n4576 avss.n4575 0.0270152
R24939 avss.n5363 avss.n4540 0.0270152
R24940 avss.n5369 avss.n5366 0.0270152
R24941 avss.n4827 avss.n4826 0.0270152
R24942 avss.n4812 avss.n4803 0.0270152
R24943 avss.n4757 avss.n4756 0.0270152
R24944 avss.n4660 avss.n4659 0.0270152
R24945 avss.n5009 avss.n4624 0.0270152
R24946 avss.n5015 avss.n5012 0.0270152
R24947 avss.n9131 avss.n9125 0.0270152
R24948 avss.n2440 avss.n2439 0.0270152
R24949 avss.n2420 avss.n2416 0.0270152
R24950 avss.n2567 avss.n2563 0.0270152
R24951 avss.n2497 avss.n2496 0.0270152
R24952 avss.n9020 avss.n9014 0.0270152
R24953 avss.n9352 avss.n9346 0.0270152
R24954 avss.n2224 avss.n2223 0.0270152
R24955 avss.n2204 avss.n2200 0.0270152
R24956 avss.n2351 avss.n2347 0.0270152
R24957 avss.n2281 avss.n2280 0.0270152
R24958 avss.n9241 avss.n9235 0.0270152
R24959 avss.n9573 avss.n9567 0.0270152
R24960 avss.n2008 avss.n2007 0.0270152
R24961 avss.n1988 avss.n1984 0.0270152
R24962 avss.n2135 avss.n2131 0.0270152
R24963 avss.n2065 avss.n2064 0.0270152
R24964 avss.n9462 avss.n9456 0.0270152
R24965 avss.n9794 avss.n9788 0.0270152
R24966 avss.n1792 avss.n1791 0.0270152
R24967 avss.n1772 avss.n1768 0.0270152
R24968 avss.n1919 avss.n1915 0.0270152
R24969 avss.n1849 avss.n1848 0.0270152
R24970 avss.n9683 avss.n9677 0.0270152
R24971 avss.n10015 avss.n10009 0.0270152
R24972 avss.n1576 avss.n1575 0.0270152
R24973 avss.n1556 avss.n1552 0.0270152
R24974 avss.n1703 avss.n1699 0.0270152
R24975 avss.n1633 avss.n1632 0.0270152
R24976 avss.n9904 avss.n9898 0.0270152
R24977 avss.n10236 avss.n10230 0.0270152
R24978 avss.n1360 avss.n1359 0.0270152
R24979 avss.n1340 avss.n1336 0.0270152
R24980 avss.n1487 avss.n1483 0.0270152
R24981 avss.n1417 avss.n1416 0.0270152
R24982 avss.n10125 avss.n10119 0.0270152
R24983 avss.n10457 avss.n10451 0.0270152
R24984 avss.n1144 avss.n1143 0.0270152
R24985 avss.n1124 avss.n1120 0.0270152
R24986 avss.n1271 avss.n1267 0.0270152
R24987 avss.n1201 avss.n1200 0.0270152
R24988 avss.n10346 avss.n10340 0.0270152
R24989 avss.n10678 avss.n10672 0.0270152
R24990 avss.n928 avss.n927 0.0270152
R24991 avss.n908 avss.n904 0.0270152
R24992 avss.n1055 avss.n1051 0.0270152
R24993 avss.n985 avss.n984 0.0270152
R24994 avss.n10567 avss.n10561 0.0270152
R24995 avss.n10899 avss.n10893 0.0270152
R24996 avss.n712 avss.n711 0.0270152
R24997 avss.n692 avss.n688 0.0270152
R24998 avss.n839 avss.n835 0.0270152
R24999 avss.n769 avss.n768 0.0270152
R25000 avss.n10788 avss.n10782 0.0270152
R25001 avss.n11120 avss.n11114 0.0270152
R25002 avss.n496 avss.n495 0.0270152
R25003 avss.n476 avss.n472 0.0270152
R25004 avss.n623 avss.n619 0.0270152
R25005 avss.n553 avss.n552 0.0270152
R25006 avss.n11009 avss.n11003 0.0270152
R25007 avss.n387 avss.n381 0.0270152
R25008 avss.n11325 avss.n11324 0.0270152
R25009 avss.n11395 avss.n11391 0.0270152
R25010 avss.n298 avss.n294 0.0270152
R25011 avss.n228 avss.n227 0.0270152
R25012 avss.n11230 avss.n11224 0.0270152
R25013 avss.n170 avss.n164 0.0270152
R25014 avss.n11546 avss.n11545 0.0270152
R25015 avss.n11616 avss.n11612 0.0270152
R25016 avss.n81 avss.n77 0.0270152
R25017 avss.n11 avss.n10 0.0270152
R25018 avss.n11451 avss.n11445 0.0270152
R25019 avss.n8818 avss.n8817 0.0261364
R25020 avss.n8796 avss.n8795 0.0261364
R25021 avss.n8781 avss.n8716 0.0261364
R25022 avss.n8864 avss.n8855 0.0261364
R25023 avss.n8904 avss.n8903 0.0261364
R25024 avss.n8928 avss.n8921 0.0261364
R25025 avss.n8465 avss.n8464 0.0261364
R25026 avss.n8443 avss.n8442 0.0261364
R25027 avss.n8428 avss.n8363 0.0261364
R25028 avss.n8511 avss.n8502 0.0261364
R25029 avss.n8551 avss.n8550 0.0261364
R25030 avss.n8575 avss.n8568 0.0261364
R25031 avss.n8112 avss.n8111 0.0261364
R25032 avss.n8090 avss.n8089 0.0261364
R25033 avss.n8075 avss.n8010 0.0261364
R25034 avss.n8158 avss.n8149 0.0261364
R25035 avss.n8198 avss.n8197 0.0261364
R25036 avss.n8222 avss.n8215 0.0261364
R25037 avss.n7759 avss.n7758 0.0261364
R25038 avss.n7737 avss.n7736 0.0261364
R25039 avss.n7722 avss.n7657 0.0261364
R25040 avss.n7805 avss.n7796 0.0261364
R25041 avss.n7845 avss.n7844 0.0261364
R25042 avss.n7869 avss.n7862 0.0261364
R25043 avss.n7406 avss.n7405 0.0261364
R25044 avss.n7384 avss.n7383 0.0261364
R25045 avss.n7369 avss.n7304 0.0261364
R25046 avss.n7452 avss.n7443 0.0261364
R25047 avss.n7492 avss.n7491 0.0261364
R25048 avss.n7516 avss.n7509 0.0261364
R25049 avss.n7053 avss.n7052 0.0261364
R25050 avss.n7031 avss.n7030 0.0261364
R25051 avss.n7016 avss.n6951 0.0261364
R25052 avss.n7099 avss.n7090 0.0261364
R25053 avss.n7139 avss.n7138 0.0261364
R25054 avss.n7163 avss.n7156 0.0261364
R25055 avss.n6700 avss.n6699 0.0261364
R25056 avss.n6678 avss.n6677 0.0261364
R25057 avss.n6663 avss.n6598 0.0261364
R25058 avss.n6746 avss.n6737 0.0261364
R25059 avss.n6786 avss.n6785 0.0261364
R25060 avss.n6810 avss.n6803 0.0261364
R25061 avss.n6347 avss.n6346 0.0261364
R25062 avss.n6325 avss.n6324 0.0261364
R25063 avss.n6310 avss.n6245 0.0261364
R25064 avss.n6393 avss.n6384 0.0261364
R25065 avss.n6433 avss.n6432 0.0261364
R25066 avss.n6457 avss.n6450 0.0261364
R25067 avss.n5994 avss.n5993 0.0261364
R25068 avss.n5972 avss.n5971 0.0261364
R25069 avss.n5957 avss.n5892 0.0261364
R25070 avss.n6040 avss.n6031 0.0261364
R25071 avss.n6080 avss.n6079 0.0261364
R25072 avss.n6104 avss.n6097 0.0261364
R25073 avss.n5641 avss.n5640 0.0261364
R25074 avss.n5619 avss.n5618 0.0261364
R25075 avss.n5604 avss.n5539 0.0261364
R25076 avss.n5687 avss.n5678 0.0261364
R25077 avss.n5727 avss.n5726 0.0261364
R25078 avss.n5751 avss.n5744 0.0261364
R25079 avss.n5298 avss.n5093 0.0261364
R25080 avss.n5274 avss.n5273 0.0261364
R25081 avss.n5259 avss.n5193 0.0261364
R25082 avss.n5334 avss.n5325 0.0261364
R25083 avss.n5374 avss.n5373 0.0261364
R25084 avss.n5398 avss.n5391 0.0261364
R25085 avss.n4944 avss.n4739 0.0261364
R25086 avss.n4920 avss.n4919 0.0261364
R25087 avss.n4905 avss.n4839 0.0261364
R25088 avss.n4980 avss.n4971 0.0261364
R25089 avss.n5020 avss.n5019 0.0261364
R25090 avss.n5044 avss.n5037 0.0261364
R25091 avss.n2391 avss.n2390 0.0261364
R25092 avss.n9179 avss.n9178 0.0261364
R25093 avss.n9186 avss.n9185 0.0261364
R25094 avss.n2589 avss.n2588 0.0261364
R25095 avss.n8978 avss.n8977 0.0261364
R25096 avss.n8985 avss.n8984 0.0261364
R25097 avss.n2175 avss.n2174 0.0261364
R25098 avss.n9400 avss.n9399 0.0261364
R25099 avss.n9407 avss.n9406 0.0261364
R25100 avss.n2373 avss.n2372 0.0261364
R25101 avss.n9199 avss.n9198 0.0261364
R25102 avss.n9206 avss.n9205 0.0261364
R25103 avss.n1959 avss.n1958 0.0261364
R25104 avss.n9621 avss.n9620 0.0261364
R25105 avss.n9628 avss.n9627 0.0261364
R25106 avss.n2157 avss.n2156 0.0261364
R25107 avss.n9420 avss.n9419 0.0261364
R25108 avss.n9427 avss.n9426 0.0261364
R25109 avss.n1743 avss.n1742 0.0261364
R25110 avss.n9842 avss.n9841 0.0261364
R25111 avss.n9849 avss.n9848 0.0261364
R25112 avss.n1941 avss.n1940 0.0261364
R25113 avss.n9641 avss.n9640 0.0261364
R25114 avss.n9648 avss.n9647 0.0261364
R25115 avss.n1527 avss.n1526 0.0261364
R25116 avss.n10063 avss.n10062 0.0261364
R25117 avss.n10070 avss.n10069 0.0261364
R25118 avss.n1725 avss.n1724 0.0261364
R25119 avss.n9862 avss.n9861 0.0261364
R25120 avss.n9869 avss.n9868 0.0261364
R25121 avss.n1311 avss.n1310 0.0261364
R25122 avss.n10284 avss.n10283 0.0261364
R25123 avss.n10291 avss.n10290 0.0261364
R25124 avss.n1509 avss.n1508 0.0261364
R25125 avss.n10083 avss.n10082 0.0261364
R25126 avss.n10090 avss.n10089 0.0261364
R25127 avss.n1095 avss.n1094 0.0261364
R25128 avss.n10505 avss.n10504 0.0261364
R25129 avss.n10512 avss.n10511 0.0261364
R25130 avss.n1293 avss.n1292 0.0261364
R25131 avss.n10304 avss.n10303 0.0261364
R25132 avss.n10311 avss.n10310 0.0261364
R25133 avss.n879 avss.n878 0.0261364
R25134 avss.n10726 avss.n10725 0.0261364
R25135 avss.n10733 avss.n10732 0.0261364
R25136 avss.n1077 avss.n1076 0.0261364
R25137 avss.n10525 avss.n10524 0.0261364
R25138 avss.n10532 avss.n10531 0.0261364
R25139 avss.n663 avss.n662 0.0261364
R25140 avss.n10947 avss.n10946 0.0261364
R25141 avss.n10954 avss.n10953 0.0261364
R25142 avss.n861 avss.n860 0.0261364
R25143 avss.n10746 avss.n10745 0.0261364
R25144 avss.n10753 avss.n10752 0.0261364
R25145 avss.n447 avss.n446 0.0261364
R25146 avss.n11168 avss.n11167 0.0261364
R25147 avss.n11175 avss.n11174 0.0261364
R25148 avss.n645 avss.n644 0.0261364
R25149 avss.n10967 avss.n10966 0.0261364
R25150 avss.n10974 avss.n10973 0.0261364
R25151 avss.n11310 avss.n11309 0.0261364
R25152 avss.n344 avss.n343 0.0261364
R25153 avss.n351 avss.n350 0.0261364
R25154 avss.n320 avss.n319 0.0261364
R25155 avss.n11188 avss.n11187 0.0261364
R25156 avss.n11195 avss.n11194 0.0261364
R25157 avss.n11531 avss.n11530 0.0261364
R25158 avss.n127 avss.n126 0.0261364
R25159 avss.n134 avss.n133 0.0261364
R25160 avss.n103 avss.n102 0.0261364
R25161 avss.n11409 avss.n11408 0.0261364
R25162 avss.n11416 avss.n11415 0.0261364
R25163 avss.n3364 avss.n3363 0.0255
R25164 avss.n3465 avss.n3195 0.0255
R25165 avss.n3515 avss.n3514 0.0255
R25166 avss.n3367 avss.n3278 0.0234167
R25167 avss.n3407 avss.n3406 0.0234167
R25168 avss.n8757 avss.n8756 0.0232273
R25169 avss.n8956 avss.n8953 0.0232273
R25170 avss.n8404 avss.n8403 0.0232273
R25171 avss.n8603 avss.n8600 0.0232273
R25172 avss.n8051 avss.n8050 0.0232273
R25173 avss.n8250 avss.n8247 0.0232273
R25174 avss.n7698 avss.n7697 0.0232273
R25175 avss.n7897 avss.n7894 0.0232273
R25176 avss.n7345 avss.n7344 0.0232273
R25177 avss.n7544 avss.n7541 0.0232273
R25178 avss.n6992 avss.n6991 0.0232273
R25179 avss.n7191 avss.n7188 0.0232273
R25180 avss.n6639 avss.n6638 0.0232273
R25181 avss.n6838 avss.n6835 0.0232273
R25182 avss.n6286 avss.n6285 0.0232273
R25183 avss.n6485 avss.n6482 0.0232273
R25184 avss.n5933 avss.n5932 0.0232273
R25185 avss.n6132 avss.n6129 0.0232273
R25186 avss.n5580 avss.n5579 0.0232273
R25187 avss.n5779 avss.n5776 0.0232273
R25188 avss.n5239 avss.n5238 0.0232273
R25189 avss.n5426 avss.n5423 0.0232273
R25190 avss.n4885 avss.n4884 0.0232273
R25191 avss.n5072 avss.n5069 0.0232273
R25192 avss.n9095 avss.n9092 0.0232273
R25193 avss.n9075 avss.n9072 0.0232273
R25194 avss.n9316 avss.n9313 0.0232273
R25195 avss.n9296 avss.n9293 0.0232273
R25196 avss.n9537 avss.n9534 0.0232273
R25197 avss.n9517 avss.n9514 0.0232273
R25198 avss.n9758 avss.n9755 0.0232273
R25199 avss.n9738 avss.n9735 0.0232273
R25200 avss.n9979 avss.n9976 0.0232273
R25201 avss.n9959 avss.n9956 0.0232273
R25202 avss.n10200 avss.n10197 0.0232273
R25203 avss.n10180 avss.n10177 0.0232273
R25204 avss.n10421 avss.n10418 0.0232273
R25205 avss.n10401 avss.n10398 0.0232273
R25206 avss.n10642 avss.n10639 0.0232273
R25207 avss.n10622 avss.n10619 0.0232273
R25208 avss.n10863 avss.n10860 0.0232273
R25209 avss.n10843 avss.n10840 0.0232273
R25210 avss.n11084 avss.n11081 0.0232273
R25211 avss.n11064 avss.n11061 0.0232273
R25212 avss.n335 avss.n332 0.0232273
R25213 avss.n11285 avss.n11282 0.0232273
R25214 avss.n118 avss.n115 0.0232273
R25215 avss.n11506 avss.n11503 0.0232273
R25216 avss.n4730 avss 0.0226354
R25217 avss.n4725 avss 0.0226354
R25218 avss.n4722 avss 0.0226354
R25219 avss.n4717 avss 0.0226354
R25220 avss.n4714 avss 0.0226354
R25221 avss.n4709 avss 0.0226354
R25222 avss.n4706 avss 0.0226354
R25223 avss.n4701 avss 0.0226354
R25224 avss.n4698 avss 0.0226354
R25225 avss.n2983 avss 0.0226354
R25226 avss avss.n2992 0.0226354
R25227 avss avss.n2999 0.0226354
R25228 avss.n3016 avss 0.0226354
R25229 avss.n3040 avss 0.0226354
R25230 avss avss.n3049 0.0226354
R25231 avss avss.n3056 0.0226354
R25232 avss avss.n3074 0.0226354
R25233 avss.n3128 avss 0.0226354
R25234 avss avss.n3083 0.0226354
R25235 avss avss.n3087 0.0226354
R25236 avss.n3097 avss 0.0226354
R25237 avss.n3632 avss 0.0226354
R25238 avss avss.n3641 0.0226354
R25239 avss avss.n3648 0.0226354
R25240 avss.n3665 avss 0.0226354
R25241 avss.n2695 avss 0.0226354
R25242 avss avss.n2704 0.0226354
R25243 avss avss.n2711 0.0226354
R25244 avss.n2728 avss 0.0226354
R25245 avss.n2740 avss 0.0226354
R25246 avss avss.n2749 0.0226354
R25247 avss avss.n2756 0.0226354
R25248 avss.n2773 avss 0.0226354
R25249 avss.n2902 avss 0.0226354
R25250 avss avss.n2781 0.0226354
R25251 avss avss.n2785 0.0226354
R25252 avss.n2871 avss 0.0226354
R25253 avss.n2862 avss 0.0226354
R25254 avss avss.n2817 0.0226354
R25255 avss avss.n2821 0.0226354
R25256 avss.n2831 avss 0.0226354
R25257 avss avss.n3541 0.0226354
R25258 avss.n3590 avss 0.0226354
R25259 avss avss.n3545 0.0226354
R25260 avss.n3582 avss 0.0226354
R25261 avss avss.n3549 0.0226354
R25262 avss.n3574 avss 0.0226354
R25263 avss avss.n3553 0.0226354
R25264 avss.n3566 avss 0.0226354
R25265 avss avss.n3557 0.0226354
R25266 avss.n8817 avss.n8653 0.0225758
R25267 avss.n8864 avss.n8863 0.0225758
R25268 avss.n3677 avss.n3675 0.0225758
R25269 avss.n8464 avss.n8300 0.0225758
R25270 avss.n8511 avss.n8510 0.0225758
R25271 avss.n3761 avss.n3759 0.0225758
R25272 avss.n8111 avss.n7947 0.0225758
R25273 avss.n8158 avss.n8157 0.0225758
R25274 avss.n3845 avss.n3843 0.0225758
R25275 avss.n7758 avss.n7594 0.0225758
R25276 avss.n7805 avss.n7804 0.0225758
R25277 avss.n3929 avss.n3927 0.0225758
R25278 avss.n7405 avss.n7241 0.0225758
R25279 avss.n7452 avss.n7451 0.0225758
R25280 avss.n4013 avss.n4011 0.0225758
R25281 avss.n7052 avss.n6888 0.0225758
R25282 avss.n7099 avss.n7098 0.0225758
R25283 avss.n4097 avss.n4095 0.0225758
R25284 avss.n6699 avss.n6535 0.0225758
R25285 avss.n6746 avss.n6745 0.0225758
R25286 avss.n4181 avss.n4179 0.0225758
R25287 avss.n6346 avss.n6182 0.0225758
R25288 avss.n6393 avss.n6392 0.0225758
R25289 avss.n4265 avss.n4263 0.0225758
R25290 avss.n5993 avss.n5829 0.0225758
R25291 avss.n6040 avss.n6039 0.0225758
R25292 avss.n4349 avss.n4347 0.0225758
R25293 avss.n5640 avss.n5476 0.0225758
R25294 avss.n5687 avss.n5686 0.0225758
R25295 avss.n4433 avss.n4431 0.0225758
R25296 avss.n5140 avss.n5093 0.0225758
R25297 avss.n5334 avss.n5333 0.0225758
R25298 avss.n4517 avss.n4515 0.0225758
R25299 avss.n4786 avss.n4739 0.0225758
R25300 avss.n4980 avss.n4979 0.0225758
R25301 avss.n4601 avss.n4599 0.0225758
R25302 avss.n2390 avss.n2389 0.0225758
R25303 avss.n2588 avss.n2587 0.0225758
R25304 avss.n9062 avss.n9061 0.0225758
R25305 avss.n2174 avss.n2173 0.0225758
R25306 avss.n2372 avss.n2371 0.0225758
R25307 avss.n9283 avss.n9282 0.0225758
R25308 avss.n1958 avss.n1957 0.0225758
R25309 avss.n2156 avss.n2155 0.0225758
R25310 avss.n9504 avss.n9503 0.0225758
R25311 avss.n1742 avss.n1741 0.0225758
R25312 avss.n1940 avss.n1939 0.0225758
R25313 avss.n9725 avss.n9724 0.0225758
R25314 avss.n1526 avss.n1525 0.0225758
R25315 avss.n1724 avss.n1723 0.0225758
R25316 avss.n9946 avss.n9945 0.0225758
R25317 avss.n1310 avss.n1309 0.0225758
R25318 avss.n1508 avss.n1507 0.0225758
R25319 avss.n10167 avss.n10166 0.0225758
R25320 avss.n1094 avss.n1093 0.0225758
R25321 avss.n1292 avss.n1291 0.0225758
R25322 avss.n10388 avss.n10387 0.0225758
R25323 avss.n878 avss.n877 0.0225758
R25324 avss.n1076 avss.n1075 0.0225758
R25325 avss.n10609 avss.n10608 0.0225758
R25326 avss.n662 avss.n661 0.0225758
R25327 avss.n860 avss.n859 0.0225758
R25328 avss.n10830 avss.n10829 0.0225758
R25329 avss.n446 avss.n445 0.0225758
R25330 avss.n644 avss.n643 0.0225758
R25331 avss.n11051 avss.n11050 0.0225758
R25332 avss.n11309 avss.n11308 0.0225758
R25333 avss.n319 avss.n318 0.0225758
R25334 avss.n11272 avss.n11271 0.0225758
R25335 avss.n11530 avss.n11529 0.0225758
R25336 avss.n102 avss.n101 0.0225758
R25337 avss.n11493 avss.n11492 0.0225758
R25338 avss.n8816 avss.n8655 0.0225758
R25339 avss.n8865 avss.n3716 0.0225758
R25340 avss.n8463 avss.n8302 0.0225758
R25341 avss.n8512 avss.n3800 0.0225758
R25342 avss.n8110 avss.n7949 0.0225758
R25343 avss.n8159 avss.n3884 0.0225758
R25344 avss.n7757 avss.n7596 0.0225758
R25345 avss.n7806 avss.n3968 0.0225758
R25346 avss.n7404 avss.n7243 0.0225758
R25347 avss.n7453 avss.n4052 0.0225758
R25348 avss.n7051 avss.n6890 0.0225758
R25349 avss.n7100 avss.n4136 0.0225758
R25350 avss.n6698 avss.n6537 0.0225758
R25351 avss.n6747 avss.n4220 0.0225758
R25352 avss.n6345 avss.n6184 0.0225758
R25353 avss.n6394 avss.n4304 0.0225758
R25354 avss.n5992 avss.n5831 0.0225758
R25355 avss.n6041 avss.n4388 0.0225758
R25356 avss.n5639 avss.n5478 0.0225758
R25357 avss.n5688 avss.n4472 0.0225758
R25358 avss.n5141 avss.n5139 0.0225758
R25359 avss.n5335 avss.n4556 0.0225758
R25360 avss.n4787 avss.n4785 0.0225758
R25361 avss.n4981 avss.n4640 0.0225758
R25362 avss.n2465 avss.n2464 0.0225758
R25363 avss.n2522 avss.n2521 0.0225758
R25364 avss.n2249 avss.n2248 0.0225758
R25365 avss.n2306 avss.n2305 0.0225758
R25366 avss.n2033 avss.n2032 0.0225758
R25367 avss.n2090 avss.n2089 0.0225758
R25368 avss.n1817 avss.n1816 0.0225758
R25369 avss.n1874 avss.n1873 0.0225758
R25370 avss.n1601 avss.n1600 0.0225758
R25371 avss.n1658 avss.n1657 0.0225758
R25372 avss.n1385 avss.n1384 0.0225758
R25373 avss.n1442 avss.n1441 0.0225758
R25374 avss.n1169 avss.n1168 0.0225758
R25375 avss.n1226 avss.n1225 0.0225758
R25376 avss.n953 avss.n952 0.0225758
R25377 avss.n1010 avss.n1009 0.0225758
R25378 avss.n737 avss.n736 0.0225758
R25379 avss.n794 avss.n793 0.0225758
R25380 avss.n521 avss.n520 0.0225758
R25381 avss.n578 avss.n577 0.0225758
R25382 avss.n11350 avss.n11349 0.0225758
R25383 avss.n253 avss.n252 0.0225758
R25384 avss.n11571 avss.n11570 0.0225758
R25385 avss.n36 avss.n35 0.0225758
R25386 avss.n11635 avss 0.0225588
R25387 avss.n3463 avss.n3462 0.022375
R25388 avss.n8793 avss.n8704 0.0213333
R25389 avss.n8635 avss.n8630 0.0213333
R25390 avss.n8757 avss.n8748 0.0213333
R25391 avss.n3735 avss.n3730 0.0213333
R25392 avss.n8896 avss.n3693 0.0213333
R25393 avss.n8962 avss.n8953 0.0213333
R25394 avss.n8440 avss.n8351 0.0213333
R25395 avss.n8282 avss.n8277 0.0213333
R25396 avss.n8404 avss.n8395 0.0213333
R25397 avss.n3819 avss.n3814 0.0213333
R25398 avss.n8543 avss.n3777 0.0213333
R25399 avss.n8609 avss.n8600 0.0213333
R25400 avss.n8087 avss.n7998 0.0213333
R25401 avss.n7929 avss.n7924 0.0213333
R25402 avss.n8051 avss.n8042 0.0213333
R25403 avss.n3903 avss.n3898 0.0213333
R25404 avss.n8190 avss.n3861 0.0213333
R25405 avss.n8256 avss.n8247 0.0213333
R25406 avss.n7734 avss.n7645 0.0213333
R25407 avss.n7576 avss.n7571 0.0213333
R25408 avss.n7698 avss.n7689 0.0213333
R25409 avss.n3987 avss.n3982 0.0213333
R25410 avss.n7837 avss.n3945 0.0213333
R25411 avss.n7903 avss.n7894 0.0213333
R25412 avss.n7381 avss.n7292 0.0213333
R25413 avss.n7223 avss.n7218 0.0213333
R25414 avss.n7345 avss.n7336 0.0213333
R25415 avss.n4071 avss.n4066 0.0213333
R25416 avss.n7484 avss.n4029 0.0213333
R25417 avss.n7550 avss.n7541 0.0213333
R25418 avss.n7028 avss.n6939 0.0213333
R25419 avss.n6870 avss.n6865 0.0213333
R25420 avss.n6992 avss.n6983 0.0213333
R25421 avss.n4155 avss.n4150 0.0213333
R25422 avss.n7131 avss.n4113 0.0213333
R25423 avss.n7197 avss.n7188 0.0213333
R25424 avss.n6675 avss.n6586 0.0213333
R25425 avss.n6517 avss.n6512 0.0213333
R25426 avss.n6639 avss.n6630 0.0213333
R25427 avss.n4239 avss.n4234 0.0213333
R25428 avss.n6778 avss.n4197 0.0213333
R25429 avss.n6844 avss.n6835 0.0213333
R25430 avss.n6322 avss.n6233 0.0213333
R25431 avss.n6164 avss.n6159 0.0213333
R25432 avss.n6286 avss.n6277 0.0213333
R25433 avss.n4323 avss.n4318 0.0213333
R25434 avss.n6425 avss.n4281 0.0213333
R25435 avss.n6491 avss.n6482 0.0213333
R25436 avss.n5969 avss.n5880 0.0213333
R25437 avss.n5811 avss.n5806 0.0213333
R25438 avss.n5933 avss.n5924 0.0213333
R25439 avss.n4407 avss.n4402 0.0213333
R25440 avss.n6072 avss.n4365 0.0213333
R25441 avss.n6138 avss.n6129 0.0213333
R25442 avss.n5616 avss.n5527 0.0213333
R25443 avss.n5458 avss.n5453 0.0213333
R25444 avss.n5580 avss.n5571 0.0213333
R25445 avss.n4491 avss.n4486 0.0213333
R25446 avss.n5719 avss.n4449 0.0213333
R25447 avss.n5785 avss.n5776 0.0213333
R25448 avss.n5271 avss.n5181 0.0213333
R25449 avss.n5110 avss.n5104 0.0213333
R25450 avss.n5239 avss.n5228 0.0213333
R25451 avss.n4575 avss.n4570 0.0213333
R25452 avss.n5366 avss.n4533 0.0213333
R25453 avss.n5432 avss.n5423 0.0213333
R25454 avss.n4917 avss.n4827 0.0213333
R25455 avss.n4756 avss.n4750 0.0213333
R25456 avss.n4885 avss.n4874 0.0213333
R25457 avss.n4659 avss.n4654 0.0213333
R25458 avss.n5012 avss.n4617 0.0213333
R25459 avss.n5078 avss.n5069 0.0213333
R25460 avss.n9131 avss.n9130 0.0213333
R25461 avss.n2420 avss.n2419 0.0213333
R25462 avss.n9092 avss.n9091 0.0213333
R25463 avss.n2567 avss.n2566 0.0213333
R25464 avss.n9020 avss.n9019 0.0213333
R25465 avss.n9072 avss.n9071 0.0213333
R25466 avss.n9352 avss.n9351 0.0213333
R25467 avss.n2204 avss.n2203 0.0213333
R25468 avss.n9313 avss.n9312 0.0213333
R25469 avss.n2351 avss.n2350 0.0213333
R25470 avss.n9241 avss.n9240 0.0213333
R25471 avss.n9293 avss.n9292 0.0213333
R25472 avss.n9573 avss.n9572 0.0213333
R25473 avss.n1988 avss.n1987 0.0213333
R25474 avss.n9534 avss.n9533 0.0213333
R25475 avss.n2135 avss.n2134 0.0213333
R25476 avss.n9462 avss.n9461 0.0213333
R25477 avss.n9514 avss.n9513 0.0213333
R25478 avss.n9794 avss.n9793 0.0213333
R25479 avss.n1772 avss.n1771 0.0213333
R25480 avss.n9755 avss.n9754 0.0213333
R25481 avss.n1919 avss.n1918 0.0213333
R25482 avss.n9683 avss.n9682 0.0213333
R25483 avss.n9735 avss.n9734 0.0213333
R25484 avss.n10015 avss.n10014 0.0213333
R25485 avss.n1556 avss.n1555 0.0213333
R25486 avss.n9976 avss.n9975 0.0213333
R25487 avss.n1703 avss.n1702 0.0213333
R25488 avss.n9904 avss.n9903 0.0213333
R25489 avss.n9956 avss.n9955 0.0213333
R25490 avss.n10236 avss.n10235 0.0213333
R25491 avss.n1340 avss.n1339 0.0213333
R25492 avss.n10197 avss.n10196 0.0213333
R25493 avss.n1487 avss.n1486 0.0213333
R25494 avss.n10125 avss.n10124 0.0213333
R25495 avss.n10177 avss.n10176 0.0213333
R25496 avss.n10457 avss.n10456 0.0213333
R25497 avss.n1124 avss.n1123 0.0213333
R25498 avss.n10418 avss.n10417 0.0213333
R25499 avss.n1271 avss.n1270 0.0213333
R25500 avss.n10346 avss.n10345 0.0213333
R25501 avss.n10398 avss.n10397 0.0213333
R25502 avss.n10678 avss.n10677 0.0213333
R25503 avss.n908 avss.n907 0.0213333
R25504 avss.n10639 avss.n10638 0.0213333
R25505 avss.n1055 avss.n1054 0.0213333
R25506 avss.n10567 avss.n10566 0.0213333
R25507 avss.n10619 avss.n10618 0.0213333
R25508 avss.n10899 avss.n10898 0.0213333
R25509 avss.n692 avss.n691 0.0213333
R25510 avss.n10860 avss.n10859 0.0213333
R25511 avss.n839 avss.n838 0.0213333
R25512 avss.n10788 avss.n10787 0.0213333
R25513 avss.n10840 avss.n10839 0.0213333
R25514 avss.n11120 avss.n11119 0.0213333
R25515 avss.n476 avss.n475 0.0213333
R25516 avss.n11081 avss.n11080 0.0213333
R25517 avss.n623 avss.n622 0.0213333
R25518 avss.n11009 avss.n11008 0.0213333
R25519 avss.n11061 avss.n11060 0.0213333
R25520 avss.n387 avss.n386 0.0213333
R25521 avss.n11395 avss.n11394 0.0213333
R25522 avss.n332 avss.n331 0.0213333
R25523 avss.n298 avss.n297 0.0213333
R25524 avss.n11230 avss.n11229 0.0213333
R25525 avss.n11282 avss.n11281 0.0213333
R25526 avss.n170 avss.n169 0.0213333
R25527 avss.n11616 avss.n11615 0.0213333
R25528 avss.n115 avss.n114 0.0213333
R25529 avss.n81 avss.n80 0.0213333
R25530 avss.n11451 avss.n11450 0.0213333
R25531 avss.n11503 avss.n11502 0.0213333
R25532 avss.n3366 avss.n3284 0.0213333
R25533 avss.n8796 avss.n8698 0.0211515
R25534 avss.n8797 avss.n8683 0.0211515
R25535 avss.n8903 avss.n3696 0.0211515
R25536 avss.n8902 avss.n3697 0.0211515
R25537 avss.n8443 avss.n8345 0.0211515
R25538 avss.n8444 avss.n8330 0.0211515
R25539 avss.n8550 avss.n3780 0.0211515
R25540 avss.n8549 avss.n3781 0.0211515
R25541 avss.n8090 avss.n7992 0.0211515
R25542 avss.n8091 avss.n7977 0.0211515
R25543 avss.n8197 avss.n3864 0.0211515
R25544 avss.n8196 avss.n3865 0.0211515
R25545 avss.n7737 avss.n7639 0.0211515
R25546 avss.n7738 avss.n7624 0.0211515
R25547 avss.n7844 avss.n3948 0.0211515
R25548 avss.n7843 avss.n3949 0.0211515
R25549 avss.n7384 avss.n7286 0.0211515
R25550 avss.n7385 avss.n7271 0.0211515
R25551 avss.n7491 avss.n4032 0.0211515
R25552 avss.n7490 avss.n4033 0.0211515
R25553 avss.n7031 avss.n6933 0.0211515
R25554 avss.n7032 avss.n6918 0.0211515
R25555 avss.n7138 avss.n4116 0.0211515
R25556 avss.n7137 avss.n4117 0.0211515
R25557 avss.n6678 avss.n6580 0.0211515
R25558 avss.n6679 avss.n6565 0.0211515
R25559 avss.n6785 avss.n4200 0.0211515
R25560 avss.n6784 avss.n4201 0.0211515
R25561 avss.n6325 avss.n6227 0.0211515
R25562 avss.n6326 avss.n6212 0.0211515
R25563 avss.n6432 avss.n4284 0.0211515
R25564 avss.n6431 avss.n4285 0.0211515
R25565 avss.n5972 avss.n5874 0.0211515
R25566 avss.n5973 avss.n5859 0.0211515
R25567 avss.n6079 avss.n4368 0.0211515
R25568 avss.n6078 avss.n4369 0.0211515
R25569 avss.n5619 avss.n5521 0.0211515
R25570 avss.n5620 avss.n5506 0.0211515
R25571 avss.n5726 avss.n4452 0.0211515
R25572 avss.n5725 avss.n4453 0.0211515
R25573 avss.n5274 avss.n5175 0.0211515
R25574 avss.n5275 avss.n5160 0.0211515
R25575 avss.n5373 avss.n4536 0.0211515
R25576 avss.n5372 avss.n4537 0.0211515
R25577 avss.n4920 avss.n4821 0.0211515
R25578 avss.n4921 avss.n4806 0.0211515
R25579 avss.n5019 avss.n4620 0.0211515
R25580 avss.n5018 avss.n4621 0.0211515
R25581 avss.n9178 avss.n9177 0.0211515
R25582 avss.n9120 avss.n9119 0.0211515
R25583 avss.n8977 avss.n8976 0.0211515
R25584 avss.n9009 avss.n9008 0.0211515
R25585 avss.n9399 avss.n9398 0.0211515
R25586 avss.n9341 avss.n9340 0.0211515
R25587 avss.n9198 avss.n9197 0.0211515
R25588 avss.n9230 avss.n9229 0.0211515
R25589 avss.n9620 avss.n9619 0.0211515
R25590 avss.n9562 avss.n9561 0.0211515
R25591 avss.n9419 avss.n9418 0.0211515
R25592 avss.n9451 avss.n9450 0.0211515
R25593 avss.n9841 avss.n9840 0.0211515
R25594 avss.n9783 avss.n9782 0.0211515
R25595 avss.n9640 avss.n9639 0.0211515
R25596 avss.n9672 avss.n9671 0.0211515
R25597 avss.n10062 avss.n10061 0.0211515
R25598 avss.n10004 avss.n10003 0.0211515
R25599 avss.n9861 avss.n9860 0.0211515
R25600 avss.n9893 avss.n9892 0.0211515
R25601 avss.n10283 avss.n10282 0.0211515
R25602 avss.n10225 avss.n10224 0.0211515
R25603 avss.n10082 avss.n10081 0.0211515
R25604 avss.n10114 avss.n10113 0.0211515
R25605 avss.n10504 avss.n10503 0.0211515
R25606 avss.n10446 avss.n10445 0.0211515
R25607 avss.n10303 avss.n10302 0.0211515
R25608 avss.n10335 avss.n10334 0.0211515
R25609 avss.n10725 avss.n10724 0.0211515
R25610 avss.n10667 avss.n10666 0.0211515
R25611 avss.n10524 avss.n10523 0.0211515
R25612 avss.n10556 avss.n10555 0.0211515
R25613 avss.n10946 avss.n10945 0.0211515
R25614 avss.n10888 avss.n10887 0.0211515
R25615 avss.n10745 avss.n10744 0.0211515
R25616 avss.n10777 avss.n10776 0.0211515
R25617 avss.n11167 avss.n11166 0.0211515
R25618 avss.n11109 avss.n11108 0.0211515
R25619 avss.n10966 avss.n10965 0.0211515
R25620 avss.n10998 avss.n10997 0.0211515
R25621 avss.n343 avss.n342 0.0211515
R25622 avss.n376 avss.n375 0.0211515
R25623 avss.n11187 avss.n11186 0.0211515
R25624 avss.n11219 avss.n11218 0.0211515
R25625 avss.n126 avss.n125 0.0211515
R25626 avss.n159 avss.n158 0.0211515
R25627 avss.n11408 avss.n11407 0.0211515
R25628 avss.n11440 avss.n11439 0.0211515
R25629 avss.n4733 avss 0.0209082
R25630 avss.n3559 avss.n3558 0.0209082
R25631 avss.n8809 avss.n8668 0.0197273
R25632 avss.n8858 avss.n3707 0.0197273
R25633 avss.n8456 avss.n8315 0.0197273
R25634 avss.n8505 avss.n3791 0.0197273
R25635 avss.n8103 avss.n7962 0.0197273
R25636 avss.n8152 avss.n3875 0.0197273
R25637 avss.n7750 avss.n7609 0.0197273
R25638 avss.n7799 avss.n3959 0.0197273
R25639 avss.n7397 avss.n7256 0.0197273
R25640 avss.n7446 avss.n4043 0.0197273
R25641 avss.n7044 avss.n6903 0.0197273
R25642 avss.n7093 avss.n4127 0.0197273
R25643 avss.n6691 avss.n6550 0.0197273
R25644 avss.n6740 avss.n4211 0.0197273
R25645 avss.n6338 avss.n6197 0.0197273
R25646 avss.n6387 avss.n4295 0.0197273
R25647 avss.n5985 avss.n5844 0.0197273
R25648 avss.n6034 avss.n4379 0.0197273
R25649 avss.n5632 avss.n5491 0.0197273
R25650 avss.n5681 avss.n4463 0.0197273
R25651 avss.n5287 avss.n5145 0.0197273
R25652 avss.n5328 avss.n4547 0.0197273
R25653 avss.n4933 avss.n4791 0.0197273
R25654 avss.n4974 avss.n4631 0.0197273
R25655 avss.n2386 avss.n2385 0.0197273
R25656 avss.n2584 avss.n2583 0.0197273
R25657 avss.n2170 avss.n2169 0.0197273
R25658 avss.n2368 avss.n2367 0.0197273
R25659 avss.n1954 avss.n1953 0.0197273
R25660 avss.n2152 avss.n2151 0.0197273
R25661 avss.n1738 avss.n1737 0.0197273
R25662 avss.n1936 avss.n1935 0.0197273
R25663 avss.n1522 avss.n1521 0.0197273
R25664 avss.n1720 avss.n1719 0.0197273
R25665 avss.n1306 avss.n1305 0.0197273
R25666 avss.n1504 avss.n1503 0.0197273
R25667 avss.n1090 avss.n1089 0.0197273
R25668 avss.n1288 avss.n1287 0.0197273
R25669 avss.n874 avss.n873 0.0197273
R25670 avss.n1072 avss.n1071 0.0197273
R25671 avss.n658 avss.n657 0.0197273
R25672 avss.n856 avss.n855 0.0197273
R25673 avss.n442 avss.n441 0.0197273
R25674 avss.n640 avss.n639 0.0197273
R25675 avss.n11305 avss.n11304 0.0197273
R25676 avss.n315 avss.n314 0.0197273
R25677 avss.n11526 avss.n11525 0.0197273
R25678 avss.n98 avss.n97 0.0197273
R25679 avss.n8764 avss.n8744 0.0194394
R25680 avss.n8676 avss.n8675 0.0194394
R25681 avss.n8871 avss.n3711 0.0194394
R25682 avss.n8950 avss.n8949 0.0194394
R25683 avss.n8411 avss.n8391 0.0194394
R25684 avss.n8323 avss.n8322 0.0194394
R25685 avss.n8518 avss.n3795 0.0194394
R25686 avss.n8597 avss.n8596 0.0194394
R25687 avss.n8058 avss.n8038 0.0194394
R25688 avss.n7970 avss.n7969 0.0194394
R25689 avss.n8165 avss.n3879 0.0194394
R25690 avss.n8244 avss.n8243 0.0194394
R25691 avss.n7705 avss.n7685 0.0194394
R25692 avss.n7617 avss.n7616 0.0194394
R25693 avss.n7812 avss.n3963 0.0194394
R25694 avss.n7891 avss.n7890 0.0194394
R25695 avss.n7352 avss.n7332 0.0194394
R25696 avss.n7264 avss.n7263 0.0194394
R25697 avss.n7459 avss.n4047 0.0194394
R25698 avss.n7538 avss.n7537 0.0194394
R25699 avss.n6999 avss.n6979 0.0194394
R25700 avss.n6911 avss.n6910 0.0194394
R25701 avss.n7106 avss.n4131 0.0194394
R25702 avss.n7185 avss.n7184 0.0194394
R25703 avss.n6646 avss.n6626 0.0194394
R25704 avss.n6558 avss.n6557 0.0194394
R25705 avss.n6753 avss.n4215 0.0194394
R25706 avss.n6832 avss.n6831 0.0194394
R25707 avss.n6293 avss.n6273 0.0194394
R25708 avss.n6205 avss.n6204 0.0194394
R25709 avss.n6400 avss.n4299 0.0194394
R25710 avss.n6479 avss.n6478 0.0194394
R25711 avss.n5940 avss.n5920 0.0194394
R25712 avss.n5852 avss.n5851 0.0194394
R25713 avss.n6047 avss.n4383 0.0194394
R25714 avss.n6126 avss.n6125 0.0194394
R25715 avss.n5587 avss.n5567 0.0194394
R25716 avss.n5499 avss.n5498 0.0194394
R25717 avss.n5694 avss.n4467 0.0194394
R25718 avss.n5773 avss.n5772 0.0194394
R25719 avss.n5247 avss.n5210 0.0194394
R25720 avss.n5153 avss.n5152 0.0194394
R25721 avss.n5341 avss.n4551 0.0194394
R25722 avss.n5420 avss.n5419 0.0194394
R25723 avss.n4893 avss.n4856 0.0194394
R25724 avss.n4799 avss.n4798 0.0194394
R25725 avss.n4987 avss.n4635 0.0194394
R25726 avss.n5066 avss.n5065 0.0194394
R25727 avss.n9112 avss.n9111 0.0194394
R25728 avss.n2455 avss.n2454 0.0194394
R25729 avss.n2512 avss.n2511 0.0194394
R25730 avss.n9000 avss.n8999 0.0194394
R25731 avss.n9333 avss.n9332 0.0194394
R25732 avss.n2239 avss.n2238 0.0194394
R25733 avss.n2296 avss.n2295 0.0194394
R25734 avss.n9221 avss.n9220 0.0194394
R25735 avss.n9554 avss.n9553 0.0194394
R25736 avss.n2023 avss.n2022 0.0194394
R25737 avss.n2080 avss.n2079 0.0194394
R25738 avss.n9442 avss.n9441 0.0194394
R25739 avss.n9775 avss.n9774 0.0194394
R25740 avss.n1807 avss.n1806 0.0194394
R25741 avss.n1864 avss.n1863 0.0194394
R25742 avss.n9663 avss.n9662 0.0194394
R25743 avss.n9996 avss.n9995 0.0194394
R25744 avss.n1591 avss.n1590 0.0194394
R25745 avss.n1648 avss.n1647 0.0194394
R25746 avss.n9884 avss.n9883 0.0194394
R25747 avss.n10217 avss.n10216 0.0194394
R25748 avss.n1375 avss.n1374 0.0194394
R25749 avss.n1432 avss.n1431 0.0194394
R25750 avss.n10105 avss.n10104 0.0194394
R25751 avss.n10438 avss.n10437 0.0194394
R25752 avss.n1159 avss.n1158 0.0194394
R25753 avss.n1216 avss.n1215 0.0194394
R25754 avss.n10326 avss.n10325 0.0194394
R25755 avss.n10659 avss.n10658 0.0194394
R25756 avss.n943 avss.n942 0.0194394
R25757 avss.n1000 avss.n999 0.0194394
R25758 avss.n10547 avss.n10546 0.0194394
R25759 avss.n10880 avss.n10879 0.0194394
R25760 avss.n727 avss.n726 0.0194394
R25761 avss.n784 avss.n783 0.0194394
R25762 avss.n10768 avss.n10767 0.0194394
R25763 avss.n11101 avss.n11100 0.0194394
R25764 avss.n511 avss.n510 0.0194394
R25765 avss.n568 avss.n567 0.0194394
R25766 avss.n10989 avss.n10988 0.0194394
R25767 avss.n367 avss.n366 0.0194394
R25768 avss.n11340 avss.n11339 0.0194394
R25769 avss.n243 avss.n242 0.0194394
R25770 avss.n11210 avss.n11209 0.0194394
R25771 avss.n150 avss.n149 0.0194394
R25772 avss.n11561 avss.n11560 0.0194394
R25773 avss.n26 avss.n25 0.0194394
R25774 avss.n11431 avss.n11430 0.0194394
R25775 avss.n3464 avss.n3463 0.01925
R25776 avss.n3381 avss.n3379 0.01925
R25777 avss.n3391 avss.n3271 0.01925
R25778 avss.n3510 avss.n3509 0.01925
R25779 avss.n2977 avss.n2958 0.0187292
R25780 avss.n3034 avss.n2942 0.0187292
R25781 avss.n3133 avss.n2928 0.0187292
R25782 avss.n3626 avss.n2608 0.0187292
R25783 avss.n2689 avss.n2671 0.0187292
R25784 avss.n2734 avss.n2644 0.0187292
R25785 avss.n2904 avss.n2630 0.0187292
R25786 avss.n2867 avss.n2810 0.0187292
R25787 avss.n8693 avss.n8692 0.018303
R25788 avss.n8890 avss.n8886 0.018303
R25789 avss.n8340 avss.n8339 0.018303
R25790 avss.n8537 avss.n8533 0.018303
R25791 avss.n7987 avss.n7986 0.018303
R25792 avss.n8184 avss.n8180 0.018303
R25793 avss.n7634 avss.n7633 0.018303
R25794 avss.n7831 avss.n7827 0.018303
R25795 avss.n7281 avss.n7280 0.018303
R25796 avss.n7478 avss.n7474 0.018303
R25797 avss.n6928 avss.n6927 0.018303
R25798 avss.n7125 avss.n7121 0.018303
R25799 avss.n6575 avss.n6574 0.018303
R25800 avss.n6772 avss.n6768 0.018303
R25801 avss.n6222 avss.n6221 0.018303
R25802 avss.n6419 avss.n6415 0.018303
R25803 avss.n5869 avss.n5868 0.018303
R25804 avss.n6066 avss.n6062 0.018303
R25805 avss.n5516 avss.n5515 0.018303
R25806 avss.n5713 avss.n5709 0.018303
R25807 avss.n5170 avss.n5169 0.018303
R25808 avss.n5360 avss.n5356 0.018303
R25809 avss.n4816 avss.n4815 0.018303
R25810 avss.n5006 avss.n5002 0.018303
R25811 avss.n2380 avss.n2379 0.018303
R25812 avss.n2578 avss.n2577 0.018303
R25813 avss.n2164 avss.n2163 0.018303
R25814 avss.n2362 avss.n2361 0.018303
R25815 avss.n1948 avss.n1947 0.018303
R25816 avss.n2146 avss.n2145 0.018303
R25817 avss.n1732 avss.n1731 0.018303
R25818 avss.n1930 avss.n1929 0.018303
R25819 avss.n1516 avss.n1515 0.018303
R25820 avss.n1714 avss.n1713 0.018303
R25821 avss.n1300 avss.n1299 0.018303
R25822 avss.n1498 avss.n1497 0.018303
R25823 avss.n1084 avss.n1083 0.018303
R25824 avss.n1282 avss.n1281 0.018303
R25825 avss.n868 avss.n867 0.018303
R25826 avss.n1066 avss.n1065 0.018303
R25827 avss.n652 avss.n651 0.018303
R25828 avss.n850 avss.n849 0.018303
R25829 avss.n436 avss.n435 0.018303
R25830 avss.n634 avss.n633 0.018303
R25831 avss.n11299 avss.n11298 0.018303
R25832 avss.n309 avss.n308 0.018303
R25833 avss.n11520 avss.n11519 0.018303
R25834 avss.n92 avss.n91 0.018303
R25835 avss.n2868 avss.n2809 0.0178015
R25836 avss.n2912 avss.n2911 0.0178015
R25837 avss.n2733 avss.n2657 0.0178015
R25838 avss.n2688 avss.n2684 0.0178015
R25839 avss.n8736 avss.n8735 0.0175455
R25840 avss.n8741 avss.n8730 0.0175455
R25841 avss.n8656 avss.n8649 0.0175455
R25842 avss.n8815 avss.n8659 0.0175455
R25843 avss.n8853 avss.n8852 0.0175455
R25844 avss.n8866 avss.n3714 0.0175455
R25845 avss.n8936 avss.n8935 0.0175455
R25846 avss.n8941 avss.n8940 0.0175455
R25847 avss.n8383 avss.n8382 0.0175455
R25848 avss.n8388 avss.n8377 0.0175455
R25849 avss.n8303 avss.n8296 0.0175455
R25850 avss.n8462 avss.n8306 0.0175455
R25851 avss.n8500 avss.n8499 0.0175455
R25852 avss.n8513 avss.n3798 0.0175455
R25853 avss.n8583 avss.n8582 0.0175455
R25854 avss.n8588 avss.n8587 0.0175455
R25855 avss.n8030 avss.n8029 0.0175455
R25856 avss.n8035 avss.n8024 0.0175455
R25857 avss.n7950 avss.n7943 0.0175455
R25858 avss.n8109 avss.n7953 0.0175455
R25859 avss.n8147 avss.n8146 0.0175455
R25860 avss.n8160 avss.n3882 0.0175455
R25861 avss.n8230 avss.n8229 0.0175455
R25862 avss.n8235 avss.n8234 0.0175455
R25863 avss.n7677 avss.n7676 0.0175455
R25864 avss.n7682 avss.n7671 0.0175455
R25865 avss.n7597 avss.n7590 0.0175455
R25866 avss.n7756 avss.n7600 0.0175455
R25867 avss.n7794 avss.n7793 0.0175455
R25868 avss.n7807 avss.n3966 0.0175455
R25869 avss.n7877 avss.n7876 0.0175455
R25870 avss.n7882 avss.n7881 0.0175455
R25871 avss.n7324 avss.n7323 0.0175455
R25872 avss.n7329 avss.n7318 0.0175455
R25873 avss.n7244 avss.n7237 0.0175455
R25874 avss.n7403 avss.n7247 0.0175455
R25875 avss.n7441 avss.n7440 0.0175455
R25876 avss.n7454 avss.n4050 0.0175455
R25877 avss.n7524 avss.n7523 0.0175455
R25878 avss.n7529 avss.n7528 0.0175455
R25879 avss.n6971 avss.n6970 0.0175455
R25880 avss.n6976 avss.n6965 0.0175455
R25881 avss.n6891 avss.n6884 0.0175455
R25882 avss.n7050 avss.n6894 0.0175455
R25883 avss.n7088 avss.n7087 0.0175455
R25884 avss.n7101 avss.n4134 0.0175455
R25885 avss.n7171 avss.n7170 0.0175455
R25886 avss.n7176 avss.n7175 0.0175455
R25887 avss.n6618 avss.n6617 0.0175455
R25888 avss.n6623 avss.n6612 0.0175455
R25889 avss.n6538 avss.n6531 0.0175455
R25890 avss.n6697 avss.n6541 0.0175455
R25891 avss.n6735 avss.n6734 0.0175455
R25892 avss.n6748 avss.n4218 0.0175455
R25893 avss.n6818 avss.n6817 0.0175455
R25894 avss.n6823 avss.n6822 0.0175455
R25895 avss.n6265 avss.n6264 0.0175455
R25896 avss.n6270 avss.n6259 0.0175455
R25897 avss.n6185 avss.n6178 0.0175455
R25898 avss.n6344 avss.n6188 0.0175455
R25899 avss.n6382 avss.n6381 0.0175455
R25900 avss.n6395 avss.n4302 0.0175455
R25901 avss.n6465 avss.n6464 0.0175455
R25902 avss.n6470 avss.n6469 0.0175455
R25903 avss.n5912 avss.n5911 0.0175455
R25904 avss.n5917 avss.n5906 0.0175455
R25905 avss.n5832 avss.n5825 0.0175455
R25906 avss.n5991 avss.n5835 0.0175455
R25907 avss.n6029 avss.n6028 0.0175455
R25908 avss.n6042 avss.n4386 0.0175455
R25909 avss.n6112 avss.n6111 0.0175455
R25910 avss.n6117 avss.n6116 0.0175455
R25911 avss.n5559 avss.n5558 0.0175455
R25912 avss.n5564 avss.n5553 0.0175455
R25913 avss.n5479 avss.n5472 0.0175455
R25914 avss.n5638 avss.n5482 0.0175455
R25915 avss.n5676 avss.n5675 0.0175455
R25916 avss.n5689 avss.n4470 0.0175455
R25917 avss.n5759 avss.n5758 0.0175455
R25918 avss.n5764 avss.n5763 0.0175455
R25919 avss.n5219 avss.n5218 0.0175455
R25920 avss.n5224 avss.n5213 0.0175455
R25921 avss.n5296 avss.n5295 0.0175455
R25922 avss.n5132 avss.n5097 0.0175455
R25923 avss.n5323 avss.n5322 0.0175455
R25924 avss.n5336 avss.n4554 0.0175455
R25925 avss.n5406 avss.n5405 0.0175455
R25926 avss.n5411 avss.n5410 0.0175455
R25927 avss.n4865 avss.n4864 0.0175455
R25928 avss.n4870 avss.n4859 0.0175455
R25929 avss.n4942 avss.n4941 0.0175455
R25930 avss.n4778 avss.n4743 0.0175455
R25931 avss.n4969 avss.n4968 0.0175455
R25932 avss.n4982 avss.n4638 0.0175455
R25933 avss.n5052 avss.n5051 0.0175455
R25934 avss.n5057 avss.n5056 0.0175455
R25935 avss.n9168 avss.n9164 0.0175455
R25936 avss.n9166 avss.n9165 0.0175455
R25937 avss.n2476 avss.n2472 0.0175455
R25938 avss.n2474 avss.n2473 0.0175455
R25939 avss.n2533 avss.n2529 0.0175455
R25940 avss.n2531 avss.n2530 0.0175455
R25941 avss.n9057 avss.n9053 0.0175455
R25942 avss.n9055 avss.n9054 0.0175455
R25943 avss.n9389 avss.n9385 0.0175455
R25944 avss.n9387 avss.n9386 0.0175455
R25945 avss.n2260 avss.n2256 0.0175455
R25946 avss.n2258 avss.n2257 0.0175455
R25947 avss.n2317 avss.n2313 0.0175455
R25948 avss.n2315 avss.n2314 0.0175455
R25949 avss.n9278 avss.n9274 0.0175455
R25950 avss.n9276 avss.n9275 0.0175455
R25951 avss.n9610 avss.n9606 0.0175455
R25952 avss.n9608 avss.n9607 0.0175455
R25953 avss.n2044 avss.n2040 0.0175455
R25954 avss.n2042 avss.n2041 0.0175455
R25955 avss.n2101 avss.n2097 0.0175455
R25956 avss.n2099 avss.n2098 0.0175455
R25957 avss.n9499 avss.n9495 0.0175455
R25958 avss.n9497 avss.n9496 0.0175455
R25959 avss.n9831 avss.n9827 0.0175455
R25960 avss.n9829 avss.n9828 0.0175455
R25961 avss.n1828 avss.n1824 0.0175455
R25962 avss.n1826 avss.n1825 0.0175455
R25963 avss.n1885 avss.n1881 0.0175455
R25964 avss.n1883 avss.n1882 0.0175455
R25965 avss.n9720 avss.n9716 0.0175455
R25966 avss.n9718 avss.n9717 0.0175455
R25967 avss.n10052 avss.n10048 0.0175455
R25968 avss.n10050 avss.n10049 0.0175455
R25969 avss.n1612 avss.n1608 0.0175455
R25970 avss.n1610 avss.n1609 0.0175455
R25971 avss.n1669 avss.n1665 0.0175455
R25972 avss.n1667 avss.n1666 0.0175455
R25973 avss.n9941 avss.n9937 0.0175455
R25974 avss.n9939 avss.n9938 0.0175455
R25975 avss.n10273 avss.n10269 0.0175455
R25976 avss.n10271 avss.n10270 0.0175455
R25977 avss.n1396 avss.n1392 0.0175455
R25978 avss.n1394 avss.n1393 0.0175455
R25979 avss.n1453 avss.n1449 0.0175455
R25980 avss.n1451 avss.n1450 0.0175455
R25981 avss.n10162 avss.n10158 0.0175455
R25982 avss.n10160 avss.n10159 0.0175455
R25983 avss.n10494 avss.n10490 0.0175455
R25984 avss.n10492 avss.n10491 0.0175455
R25985 avss.n1180 avss.n1176 0.0175455
R25986 avss.n1178 avss.n1177 0.0175455
R25987 avss.n1237 avss.n1233 0.0175455
R25988 avss.n1235 avss.n1234 0.0175455
R25989 avss.n10383 avss.n10379 0.0175455
R25990 avss.n10381 avss.n10380 0.0175455
R25991 avss.n10715 avss.n10711 0.0175455
R25992 avss.n10713 avss.n10712 0.0175455
R25993 avss.n964 avss.n960 0.0175455
R25994 avss.n962 avss.n961 0.0175455
R25995 avss.n1021 avss.n1017 0.0175455
R25996 avss.n1019 avss.n1018 0.0175455
R25997 avss.n10604 avss.n10600 0.0175455
R25998 avss.n10602 avss.n10601 0.0175455
R25999 avss.n10936 avss.n10932 0.0175455
R26000 avss.n10934 avss.n10933 0.0175455
R26001 avss.n748 avss.n744 0.0175455
R26002 avss.n746 avss.n745 0.0175455
R26003 avss.n805 avss.n801 0.0175455
R26004 avss.n803 avss.n802 0.0175455
R26005 avss.n10825 avss.n10821 0.0175455
R26006 avss.n10823 avss.n10822 0.0175455
R26007 avss.n11157 avss.n11153 0.0175455
R26008 avss.n11155 avss.n11154 0.0175455
R26009 avss.n532 avss.n528 0.0175455
R26010 avss.n530 avss.n529 0.0175455
R26011 avss.n589 avss.n585 0.0175455
R26012 avss.n587 avss.n586 0.0175455
R26013 avss.n11046 avss.n11042 0.0175455
R26014 avss.n11044 avss.n11043 0.0175455
R26015 avss.n424 avss.n420 0.0175455
R26016 avss.n422 avss.n421 0.0175455
R26017 avss.n11361 avss.n11357 0.0175455
R26018 avss.n11359 avss.n11358 0.0175455
R26019 avss.n264 avss.n260 0.0175455
R26020 avss.n262 avss.n261 0.0175455
R26021 avss.n11267 avss.n11263 0.0175455
R26022 avss.n11265 avss.n11264 0.0175455
R26023 avss.n207 avss.n203 0.0175455
R26024 avss.n205 avss.n204 0.0175455
R26025 avss.n11582 avss.n11578 0.0175455
R26026 avss.n11580 avss.n11579 0.0175455
R26027 avss.n47 avss.n43 0.0175455
R26028 avss.n45 avss.n44 0.0175455
R26029 avss.n11488 avss.n11484 0.0175455
R26030 avss.n11486 avss.n11485 0.0175455
R26031 avss.n3379 avss.n3378 0.0171667
R26032 avss.n3515 avss.n3173 0.0171667
R26033 avss.n8781 avss.n8780 0.0168788
R26034 avss.n8834 avss.n8621 0.0168788
R26035 avss.n8782 avss.n8719 0.0168788
R26036 avss.n8928 avss.n8927 0.0168788
R26037 avss.n8929 avss.n3688 0.0168788
R26038 avss.n8428 avss.n8427 0.0168788
R26039 avss.n8481 avss.n8268 0.0168788
R26040 avss.n8429 avss.n8366 0.0168788
R26041 avss.n8575 avss.n8574 0.0168788
R26042 avss.n8576 avss.n3772 0.0168788
R26043 avss.n8075 avss.n8074 0.0168788
R26044 avss.n8128 avss.n7915 0.0168788
R26045 avss.n8076 avss.n8013 0.0168788
R26046 avss.n8222 avss.n8221 0.0168788
R26047 avss.n8223 avss.n3856 0.0168788
R26048 avss.n7722 avss.n7721 0.0168788
R26049 avss.n7775 avss.n7562 0.0168788
R26050 avss.n7723 avss.n7660 0.0168788
R26051 avss.n7869 avss.n7868 0.0168788
R26052 avss.n7870 avss.n3940 0.0168788
R26053 avss.n7369 avss.n7368 0.0168788
R26054 avss.n7422 avss.n7209 0.0168788
R26055 avss.n7370 avss.n7307 0.0168788
R26056 avss.n7516 avss.n7515 0.0168788
R26057 avss.n7517 avss.n4024 0.0168788
R26058 avss.n7016 avss.n7015 0.0168788
R26059 avss.n7069 avss.n6856 0.0168788
R26060 avss.n7017 avss.n6954 0.0168788
R26061 avss.n7163 avss.n7162 0.0168788
R26062 avss.n7164 avss.n4108 0.0168788
R26063 avss.n6663 avss.n6662 0.0168788
R26064 avss.n6716 avss.n6503 0.0168788
R26065 avss.n6664 avss.n6601 0.0168788
R26066 avss.n6810 avss.n6809 0.0168788
R26067 avss.n6811 avss.n4192 0.0168788
R26068 avss.n6310 avss.n6309 0.0168788
R26069 avss.n6363 avss.n6150 0.0168788
R26070 avss.n6311 avss.n6248 0.0168788
R26071 avss.n6457 avss.n6456 0.0168788
R26072 avss.n6458 avss.n4276 0.0168788
R26073 avss.n5957 avss.n5956 0.0168788
R26074 avss.n6010 avss.n5797 0.0168788
R26075 avss.n5958 avss.n5895 0.0168788
R26076 avss.n6104 avss.n6103 0.0168788
R26077 avss.n6105 avss.n4360 0.0168788
R26078 avss.n5604 avss.n5603 0.0168788
R26079 avss.n5657 avss.n5444 0.0168788
R26080 avss.n5605 avss.n5542 0.0168788
R26081 avss.n5751 avss.n5750 0.0168788
R26082 avss.n5752 avss.n4444 0.0168788
R26083 avss.n5259 avss.n5258 0.0168788
R26084 avss.n5304 avss.n5091 0.0168788
R26085 avss.n5260 avss.n5196 0.0168788
R26086 avss.n5398 avss.n5397 0.0168788
R26087 avss.n5399 avss.n4528 0.0168788
R26088 avss.n4905 avss.n4904 0.0168788
R26089 avss.n4950 avss.n4737 0.0168788
R26090 avss.n4906 avss.n4842 0.0168788
R26091 avss.n5044 avss.n5043 0.0168788
R26092 avss.n5045 avss.n4612 0.0168788
R26093 avss.n9187 avss.n9186 0.0168788
R26094 avss.n2395 avss.n2394 0.0168788
R26095 avss.n9153 avss.n9152 0.0168788
R26096 avss.n8986 avss.n8985 0.0168788
R26097 avss.n9042 avss.n9041 0.0168788
R26098 avss.n9408 avss.n9407 0.0168788
R26099 avss.n2179 avss.n2178 0.0168788
R26100 avss.n9374 avss.n9373 0.0168788
R26101 avss.n9207 avss.n9206 0.0168788
R26102 avss.n9263 avss.n9262 0.0168788
R26103 avss.n9629 avss.n9628 0.0168788
R26104 avss.n1963 avss.n1962 0.0168788
R26105 avss.n9595 avss.n9594 0.0168788
R26106 avss.n9428 avss.n9427 0.0168788
R26107 avss.n9484 avss.n9483 0.0168788
R26108 avss.n9850 avss.n9849 0.0168788
R26109 avss.n1747 avss.n1746 0.0168788
R26110 avss.n9816 avss.n9815 0.0168788
R26111 avss.n9649 avss.n9648 0.0168788
R26112 avss.n9705 avss.n9704 0.0168788
R26113 avss.n10071 avss.n10070 0.0168788
R26114 avss.n1531 avss.n1530 0.0168788
R26115 avss.n10037 avss.n10036 0.0168788
R26116 avss.n9870 avss.n9869 0.0168788
R26117 avss.n9926 avss.n9925 0.0168788
R26118 avss.n10292 avss.n10291 0.0168788
R26119 avss.n1315 avss.n1314 0.0168788
R26120 avss.n10258 avss.n10257 0.0168788
R26121 avss.n10091 avss.n10090 0.0168788
R26122 avss.n10147 avss.n10146 0.0168788
R26123 avss.n10513 avss.n10512 0.0168788
R26124 avss.n1099 avss.n1098 0.0168788
R26125 avss.n10479 avss.n10478 0.0168788
R26126 avss.n10312 avss.n10311 0.0168788
R26127 avss.n10368 avss.n10367 0.0168788
R26128 avss.n10734 avss.n10733 0.0168788
R26129 avss.n883 avss.n882 0.0168788
R26130 avss.n10700 avss.n10699 0.0168788
R26131 avss.n10533 avss.n10532 0.0168788
R26132 avss.n10589 avss.n10588 0.0168788
R26133 avss.n10955 avss.n10954 0.0168788
R26134 avss.n667 avss.n666 0.0168788
R26135 avss.n10921 avss.n10920 0.0168788
R26136 avss.n10754 avss.n10753 0.0168788
R26137 avss.n10810 avss.n10809 0.0168788
R26138 avss.n11176 avss.n11175 0.0168788
R26139 avss.n451 avss.n450 0.0168788
R26140 avss.n11142 avss.n11141 0.0168788
R26141 avss.n10975 avss.n10974 0.0168788
R26142 avss.n11031 avss.n11030 0.0168788
R26143 avss.n352 avss.n351 0.0168788
R26144 avss.n11369 avss.n11368 0.0168788
R26145 avss.n409 avss.n408 0.0168788
R26146 avss.n11196 avss.n11195 0.0168788
R26147 avss.n11252 avss.n11251 0.0168788
R26148 avss.n135 avss.n134 0.0168788
R26149 avss.n11590 avss.n11589 0.0168788
R26150 avss.n192 avss.n191 0.0168788
R26151 avss.n11417 avss.n11416 0.0168788
R26152 avss.n11473 avss.n11472 0.0168788
R26153 avss.n3365 avss.n3364 0.016125
R26154 avss.n8735 avss.n8734 0.0156515
R26155 avss.n8798 avss.n8682 0.0156515
R26156 avss.n8803 avss.n8802 0.0156515
R26157 avss.n8821 avss.n8649 0.0156515
R26158 avss.n8755 avss.n8751 0.0156515
R26159 avss.n8853 avss.n8849 0.0156515
R26160 avss.n8881 avss.n8880 0.0156515
R26161 avss.n8901 avss.n8900 0.0156515
R26162 avss.n8935 avss.n8934 0.0156515
R26163 avss.n8960 avss.n8954 0.0156515
R26164 avss.n8382 avss.n8381 0.0156515
R26165 avss.n8445 avss.n8329 0.0156515
R26166 avss.n8450 avss.n8449 0.0156515
R26167 avss.n8468 avss.n8296 0.0156515
R26168 avss.n8402 avss.n8398 0.0156515
R26169 avss.n8500 avss.n8496 0.0156515
R26170 avss.n8528 avss.n8527 0.0156515
R26171 avss.n8548 avss.n8547 0.0156515
R26172 avss.n8582 avss.n8581 0.0156515
R26173 avss.n8607 avss.n8601 0.0156515
R26174 avss.n8029 avss.n8028 0.0156515
R26175 avss.n8092 avss.n7976 0.0156515
R26176 avss.n8097 avss.n8096 0.0156515
R26177 avss.n8115 avss.n7943 0.0156515
R26178 avss.n8049 avss.n8045 0.0156515
R26179 avss.n8147 avss.n8143 0.0156515
R26180 avss.n8175 avss.n8174 0.0156515
R26181 avss.n8195 avss.n8194 0.0156515
R26182 avss.n8229 avss.n8228 0.0156515
R26183 avss.n8254 avss.n8248 0.0156515
R26184 avss.n7676 avss.n7675 0.0156515
R26185 avss.n7739 avss.n7623 0.0156515
R26186 avss.n7744 avss.n7743 0.0156515
R26187 avss.n7762 avss.n7590 0.0156515
R26188 avss.n7696 avss.n7692 0.0156515
R26189 avss.n7794 avss.n7790 0.0156515
R26190 avss.n7822 avss.n7821 0.0156515
R26191 avss.n7842 avss.n7841 0.0156515
R26192 avss.n7876 avss.n7875 0.0156515
R26193 avss.n7901 avss.n7895 0.0156515
R26194 avss.n7323 avss.n7322 0.0156515
R26195 avss.n7386 avss.n7270 0.0156515
R26196 avss.n7391 avss.n7390 0.0156515
R26197 avss.n7409 avss.n7237 0.0156515
R26198 avss.n7343 avss.n7339 0.0156515
R26199 avss.n7441 avss.n7437 0.0156515
R26200 avss.n7469 avss.n7468 0.0156515
R26201 avss.n7489 avss.n7488 0.0156515
R26202 avss.n7523 avss.n7522 0.0156515
R26203 avss.n7548 avss.n7542 0.0156515
R26204 avss.n6970 avss.n6969 0.0156515
R26205 avss.n7033 avss.n6917 0.0156515
R26206 avss.n7038 avss.n7037 0.0156515
R26207 avss.n7056 avss.n6884 0.0156515
R26208 avss.n6990 avss.n6986 0.0156515
R26209 avss.n7088 avss.n7084 0.0156515
R26210 avss.n7116 avss.n7115 0.0156515
R26211 avss.n7136 avss.n7135 0.0156515
R26212 avss.n7170 avss.n7169 0.0156515
R26213 avss.n7195 avss.n7189 0.0156515
R26214 avss.n6617 avss.n6616 0.0156515
R26215 avss.n6680 avss.n6564 0.0156515
R26216 avss.n6685 avss.n6684 0.0156515
R26217 avss.n6703 avss.n6531 0.0156515
R26218 avss.n6637 avss.n6633 0.0156515
R26219 avss.n6735 avss.n6731 0.0156515
R26220 avss.n6763 avss.n6762 0.0156515
R26221 avss.n6783 avss.n6782 0.0156515
R26222 avss.n6817 avss.n6816 0.0156515
R26223 avss.n6842 avss.n6836 0.0156515
R26224 avss.n6264 avss.n6263 0.0156515
R26225 avss.n6327 avss.n6211 0.0156515
R26226 avss.n6332 avss.n6331 0.0156515
R26227 avss.n6350 avss.n6178 0.0156515
R26228 avss.n6284 avss.n6280 0.0156515
R26229 avss.n6382 avss.n6378 0.0156515
R26230 avss.n6410 avss.n6409 0.0156515
R26231 avss.n6430 avss.n6429 0.0156515
R26232 avss.n6464 avss.n6463 0.0156515
R26233 avss.n6489 avss.n6483 0.0156515
R26234 avss.n5911 avss.n5910 0.0156515
R26235 avss.n5974 avss.n5858 0.0156515
R26236 avss.n5979 avss.n5978 0.0156515
R26237 avss.n5997 avss.n5825 0.0156515
R26238 avss.n5931 avss.n5927 0.0156515
R26239 avss.n6029 avss.n6025 0.0156515
R26240 avss.n6057 avss.n6056 0.0156515
R26241 avss.n6077 avss.n6076 0.0156515
R26242 avss.n6111 avss.n6110 0.0156515
R26243 avss.n6136 avss.n6130 0.0156515
R26244 avss.n5558 avss.n5557 0.0156515
R26245 avss.n5621 avss.n5505 0.0156515
R26246 avss.n5626 avss.n5625 0.0156515
R26247 avss.n5644 avss.n5472 0.0156515
R26248 avss.n5578 avss.n5574 0.0156515
R26249 avss.n5676 avss.n5672 0.0156515
R26250 avss.n5704 avss.n5703 0.0156515
R26251 avss.n5724 avss.n5723 0.0156515
R26252 avss.n5758 avss.n5757 0.0156515
R26253 avss.n5783 avss.n5777 0.0156515
R26254 avss.n5218 avss.n5217 0.0156515
R26255 avss.n5276 avss.n5159 0.0156515
R26256 avss.n5281 avss.n5280 0.0156515
R26257 avss.n5296 avss.n5096 0.0156515
R26258 avss.n5237 avss.n5233 0.0156515
R26259 avss.n5323 avss.n5319 0.0156515
R26260 avss.n5351 avss.n5350 0.0156515
R26261 avss.n5371 avss.n5370 0.0156515
R26262 avss.n5405 avss.n5404 0.0156515
R26263 avss.n5430 avss.n5424 0.0156515
R26264 avss.n4864 avss.n4863 0.0156515
R26265 avss.n4922 avss.n4805 0.0156515
R26266 avss.n4927 avss.n4926 0.0156515
R26267 avss.n4942 avss.n4742 0.0156515
R26268 avss.n4883 avss.n4879 0.0156515
R26269 avss.n4969 avss.n4965 0.0156515
R26270 avss.n4997 avss.n4996 0.0156515
R26271 avss.n5017 avss.n5016 0.0156515
R26272 avss.n5051 avss.n5050 0.0156515
R26273 avss.n5076 avss.n5070 0.0156515
R26274 avss.n9164 avss.n9163 0.0156515
R26275 avss.n9124 avss.n9123 0.0156515
R26276 avss.n2435 avss.n2434 0.0156515
R26277 avss.n2472 avss.n2471 0.0156515
R26278 avss.n9094 avss.n9093 0.0156515
R26279 avss.n2529 avss.n2528 0.0156515
R26280 avss.n2492 avss.n2491 0.0156515
R26281 avss.n9013 avss.n9012 0.0156515
R26282 avss.n9053 avss.n9052 0.0156515
R26283 avss.n9074 avss.n9073 0.0156515
R26284 avss.n9385 avss.n9384 0.0156515
R26285 avss.n9345 avss.n9344 0.0156515
R26286 avss.n2219 avss.n2218 0.0156515
R26287 avss.n2256 avss.n2255 0.0156515
R26288 avss.n9315 avss.n9314 0.0156515
R26289 avss.n2313 avss.n2312 0.0156515
R26290 avss.n2276 avss.n2275 0.0156515
R26291 avss.n9234 avss.n9233 0.0156515
R26292 avss.n9274 avss.n9273 0.0156515
R26293 avss.n9295 avss.n9294 0.0156515
R26294 avss.n9606 avss.n9605 0.0156515
R26295 avss.n9566 avss.n9565 0.0156515
R26296 avss.n2003 avss.n2002 0.0156515
R26297 avss.n2040 avss.n2039 0.0156515
R26298 avss.n9536 avss.n9535 0.0156515
R26299 avss.n2097 avss.n2096 0.0156515
R26300 avss.n2060 avss.n2059 0.0156515
R26301 avss.n9455 avss.n9454 0.0156515
R26302 avss.n9495 avss.n9494 0.0156515
R26303 avss.n9516 avss.n9515 0.0156515
R26304 avss.n9827 avss.n9826 0.0156515
R26305 avss.n9787 avss.n9786 0.0156515
R26306 avss.n1787 avss.n1786 0.0156515
R26307 avss.n1824 avss.n1823 0.0156515
R26308 avss.n9757 avss.n9756 0.0156515
R26309 avss.n1881 avss.n1880 0.0156515
R26310 avss.n1844 avss.n1843 0.0156515
R26311 avss.n9676 avss.n9675 0.0156515
R26312 avss.n9716 avss.n9715 0.0156515
R26313 avss.n9737 avss.n9736 0.0156515
R26314 avss.n10048 avss.n10047 0.0156515
R26315 avss.n10008 avss.n10007 0.0156515
R26316 avss.n1571 avss.n1570 0.0156515
R26317 avss.n1608 avss.n1607 0.0156515
R26318 avss.n9978 avss.n9977 0.0156515
R26319 avss.n1665 avss.n1664 0.0156515
R26320 avss.n1628 avss.n1627 0.0156515
R26321 avss.n9897 avss.n9896 0.0156515
R26322 avss.n9937 avss.n9936 0.0156515
R26323 avss.n9958 avss.n9957 0.0156515
R26324 avss.n10269 avss.n10268 0.0156515
R26325 avss.n10229 avss.n10228 0.0156515
R26326 avss.n1355 avss.n1354 0.0156515
R26327 avss.n1392 avss.n1391 0.0156515
R26328 avss.n10199 avss.n10198 0.0156515
R26329 avss.n1449 avss.n1448 0.0156515
R26330 avss.n1412 avss.n1411 0.0156515
R26331 avss.n10118 avss.n10117 0.0156515
R26332 avss.n10158 avss.n10157 0.0156515
R26333 avss.n10179 avss.n10178 0.0156515
R26334 avss.n10490 avss.n10489 0.0156515
R26335 avss.n10450 avss.n10449 0.0156515
R26336 avss.n1139 avss.n1138 0.0156515
R26337 avss.n1176 avss.n1175 0.0156515
R26338 avss.n10420 avss.n10419 0.0156515
R26339 avss.n1233 avss.n1232 0.0156515
R26340 avss.n1196 avss.n1195 0.0156515
R26341 avss.n10339 avss.n10338 0.0156515
R26342 avss.n10379 avss.n10378 0.0156515
R26343 avss.n10400 avss.n10399 0.0156515
R26344 avss.n10711 avss.n10710 0.0156515
R26345 avss.n10671 avss.n10670 0.0156515
R26346 avss.n923 avss.n922 0.0156515
R26347 avss.n960 avss.n959 0.0156515
R26348 avss.n10641 avss.n10640 0.0156515
R26349 avss.n1017 avss.n1016 0.0156515
R26350 avss.n980 avss.n979 0.0156515
R26351 avss.n10560 avss.n10559 0.0156515
R26352 avss.n10600 avss.n10599 0.0156515
R26353 avss.n10621 avss.n10620 0.0156515
R26354 avss.n10932 avss.n10931 0.0156515
R26355 avss.n10892 avss.n10891 0.0156515
R26356 avss.n707 avss.n706 0.0156515
R26357 avss.n744 avss.n743 0.0156515
R26358 avss.n10862 avss.n10861 0.0156515
R26359 avss.n801 avss.n800 0.0156515
R26360 avss.n764 avss.n763 0.0156515
R26361 avss.n10781 avss.n10780 0.0156515
R26362 avss.n10821 avss.n10820 0.0156515
R26363 avss.n10842 avss.n10841 0.0156515
R26364 avss.n11153 avss.n11152 0.0156515
R26365 avss.n11113 avss.n11112 0.0156515
R26366 avss.n491 avss.n490 0.0156515
R26367 avss.n528 avss.n527 0.0156515
R26368 avss.n11083 avss.n11082 0.0156515
R26369 avss.n585 avss.n584 0.0156515
R26370 avss.n548 avss.n547 0.0156515
R26371 avss.n11002 avss.n11001 0.0156515
R26372 avss.n11042 avss.n11041 0.0156515
R26373 avss.n11063 avss.n11062 0.0156515
R26374 avss.n420 avss.n419 0.0156515
R26375 avss.n380 avss.n379 0.0156515
R26376 avss.n11320 avss.n11319 0.0156515
R26377 avss.n11357 avss.n11356 0.0156515
R26378 avss.n334 avss.n333 0.0156515
R26379 avss.n260 avss.n259 0.0156515
R26380 avss.n223 avss.n222 0.0156515
R26381 avss.n11223 avss.n11222 0.0156515
R26382 avss.n11263 avss.n11262 0.0156515
R26383 avss.n11284 avss.n11283 0.0156515
R26384 avss.n203 avss.n202 0.0156515
R26385 avss.n163 avss.n162 0.0156515
R26386 avss.n11541 avss.n11540 0.0156515
R26387 avss.n11578 avss.n11577 0.0156515
R26388 avss.n117 avss.n116 0.0156515
R26389 avss.n43 avss.n42 0.0156515
R26390 avss.n6 avss.n5 0.0156515
R26391 avss.n11444 avss.n11443 0.0156515
R26392 avss.n11484 avss.n11483 0.0156515
R26393 avss.n11505 avss.n11504 0.0156515
R26394 avss.n8716 avss.n8715 0.0154545
R26395 avss.n8831 avss.n8627 0.0154545
R26396 avss.n8788 avss.n8707 0.0154545
R26397 avss.n8921 avss.n3689 0.0154545
R26398 avss.n8838 avss.n3751 0.0154545
R26399 avss.n8920 avss.n3690 0.0154545
R26400 avss.n8363 avss.n8362 0.0154545
R26401 avss.n8478 avss.n8274 0.0154545
R26402 avss.n8435 avss.n8354 0.0154545
R26403 avss.n8568 avss.n3773 0.0154545
R26404 avss.n8485 avss.n3835 0.0154545
R26405 avss.n8567 avss.n3774 0.0154545
R26406 avss.n8010 avss.n8009 0.0154545
R26407 avss.n8125 avss.n7921 0.0154545
R26408 avss.n8082 avss.n8001 0.0154545
R26409 avss.n8215 avss.n3857 0.0154545
R26410 avss.n8132 avss.n3919 0.0154545
R26411 avss.n8214 avss.n3858 0.0154545
R26412 avss.n7657 avss.n7656 0.0154545
R26413 avss.n7772 avss.n7568 0.0154545
R26414 avss.n7729 avss.n7648 0.0154545
R26415 avss.n7862 avss.n3941 0.0154545
R26416 avss.n7779 avss.n4003 0.0154545
R26417 avss.n7861 avss.n3942 0.0154545
R26418 avss.n7304 avss.n7303 0.0154545
R26419 avss.n7419 avss.n7215 0.0154545
R26420 avss.n7376 avss.n7295 0.0154545
R26421 avss.n7509 avss.n4025 0.0154545
R26422 avss.n7426 avss.n4087 0.0154545
R26423 avss.n7508 avss.n4026 0.0154545
R26424 avss.n6951 avss.n6950 0.0154545
R26425 avss.n7066 avss.n6862 0.0154545
R26426 avss.n7023 avss.n6942 0.0154545
R26427 avss.n7156 avss.n4109 0.0154545
R26428 avss.n7073 avss.n4171 0.0154545
R26429 avss.n7155 avss.n4110 0.0154545
R26430 avss.n6598 avss.n6597 0.0154545
R26431 avss.n6713 avss.n6509 0.0154545
R26432 avss.n6670 avss.n6589 0.0154545
R26433 avss.n6803 avss.n4193 0.0154545
R26434 avss.n6720 avss.n4255 0.0154545
R26435 avss.n6802 avss.n4194 0.0154545
R26436 avss.n6245 avss.n6244 0.0154545
R26437 avss.n6360 avss.n6156 0.0154545
R26438 avss.n6317 avss.n6236 0.0154545
R26439 avss.n6450 avss.n4277 0.0154545
R26440 avss.n6367 avss.n4339 0.0154545
R26441 avss.n6449 avss.n4278 0.0154545
R26442 avss.n5892 avss.n5891 0.0154545
R26443 avss.n6007 avss.n5803 0.0154545
R26444 avss.n5964 avss.n5883 0.0154545
R26445 avss.n6097 avss.n4361 0.0154545
R26446 avss.n6014 avss.n4423 0.0154545
R26447 avss.n6096 avss.n4362 0.0154545
R26448 avss.n5539 avss.n5538 0.0154545
R26449 avss.n5654 avss.n5450 0.0154545
R26450 avss.n5611 avss.n5530 0.0154545
R26451 avss.n5744 avss.n4445 0.0154545
R26452 avss.n5661 avss.n4507 0.0154545
R26453 avss.n5743 avss.n4446 0.0154545
R26454 avss.n5193 avss.n5192 0.0154545
R26455 avss.n5266 avss.n5184 0.0154545
R26456 avss.n5391 avss.n4529 0.0154545
R26457 avss.n5308 avss.n4591 0.0154545
R26458 avss.n5390 avss.n4530 0.0154545
R26459 avss.n4839 avss.n4838 0.0154545
R26460 avss.n4912 avss.n4830 0.0154545
R26461 avss.n5037 avss.n4613 0.0154545
R26462 avss.n4954 avss.n4675 0.0154545
R26463 avss.n5036 avss.n4614 0.0154545
R26464 avss.n9185 avss.n9184 0.0154545
R26465 avss.n2408 avss.n2407 0.0154545
R26466 avss.n9140 avss.n9139 0.0154545
R26467 avss.n8984 avss.n8983 0.0154545
R26468 avss.n2555 avss.n2554 0.0154545
R26469 avss.n9029 avss.n9028 0.0154545
R26470 avss.n9406 avss.n9405 0.0154545
R26471 avss.n2192 avss.n2191 0.0154545
R26472 avss.n9361 avss.n9360 0.0154545
R26473 avss.n9205 avss.n9204 0.0154545
R26474 avss.n2339 avss.n2338 0.0154545
R26475 avss.n9250 avss.n9249 0.0154545
R26476 avss.n9627 avss.n9626 0.0154545
R26477 avss.n1976 avss.n1975 0.0154545
R26478 avss.n9582 avss.n9581 0.0154545
R26479 avss.n9426 avss.n9425 0.0154545
R26480 avss.n2123 avss.n2122 0.0154545
R26481 avss.n9471 avss.n9470 0.0154545
R26482 avss.n9848 avss.n9847 0.0154545
R26483 avss.n1760 avss.n1759 0.0154545
R26484 avss.n9803 avss.n9802 0.0154545
R26485 avss.n9647 avss.n9646 0.0154545
R26486 avss.n1907 avss.n1906 0.0154545
R26487 avss.n9692 avss.n9691 0.0154545
R26488 avss.n10069 avss.n10068 0.0154545
R26489 avss.n1544 avss.n1543 0.0154545
R26490 avss.n10024 avss.n10023 0.0154545
R26491 avss.n9868 avss.n9867 0.0154545
R26492 avss.n1691 avss.n1690 0.0154545
R26493 avss.n9913 avss.n9912 0.0154545
R26494 avss.n10290 avss.n10289 0.0154545
R26495 avss.n1328 avss.n1327 0.0154545
R26496 avss.n10245 avss.n10244 0.0154545
R26497 avss.n10089 avss.n10088 0.0154545
R26498 avss.n1475 avss.n1474 0.0154545
R26499 avss.n10134 avss.n10133 0.0154545
R26500 avss.n10511 avss.n10510 0.0154545
R26501 avss.n1112 avss.n1111 0.0154545
R26502 avss.n10466 avss.n10465 0.0154545
R26503 avss.n10310 avss.n10309 0.0154545
R26504 avss.n1259 avss.n1258 0.0154545
R26505 avss.n10355 avss.n10354 0.0154545
R26506 avss.n10732 avss.n10731 0.0154545
R26507 avss.n896 avss.n895 0.0154545
R26508 avss.n10687 avss.n10686 0.0154545
R26509 avss.n10531 avss.n10530 0.0154545
R26510 avss.n1043 avss.n1042 0.0154545
R26511 avss.n10576 avss.n10575 0.0154545
R26512 avss.n10953 avss.n10952 0.0154545
R26513 avss.n680 avss.n679 0.0154545
R26514 avss.n10908 avss.n10907 0.0154545
R26515 avss.n10752 avss.n10751 0.0154545
R26516 avss.n827 avss.n826 0.0154545
R26517 avss.n10797 avss.n10796 0.0154545
R26518 avss.n11174 avss.n11173 0.0154545
R26519 avss.n464 avss.n463 0.0154545
R26520 avss.n11129 avss.n11128 0.0154545
R26521 avss.n10973 avss.n10972 0.0154545
R26522 avss.n611 avss.n610 0.0154545
R26523 avss.n11018 avss.n11017 0.0154545
R26524 avss.n350 avss.n349 0.0154545
R26525 avss.n396 avss.n395 0.0154545
R26526 avss.n11194 avss.n11193 0.0154545
R26527 avss.n286 avss.n285 0.0154545
R26528 avss.n11239 avss.n11238 0.0154545
R26529 avss.n133 avss.n132 0.0154545
R26530 avss.n179 avss.n178 0.0154545
R26531 avss.n11415 avss.n11414 0.0154545
R26532 avss.n69 avss.n68 0.0154545
R26533 avss.n11460 avss.n11459 0.0154545
R26534 avss.n11635 avss 0.0149231
R26535 avss.n8774 avss.n8722 0.0147424
R26536 avss.n8968 avss.n8967 0.0147424
R26537 avss.n8421 avss.n8369 0.0147424
R26538 avss.n8615 avss.n8614 0.0147424
R26539 avss.n8068 avss.n8016 0.0147424
R26540 avss.n8262 avss.n8261 0.0147424
R26541 avss.n7715 avss.n7663 0.0147424
R26542 avss.n7909 avss.n7908 0.0147424
R26543 avss.n7362 avss.n7310 0.0147424
R26544 avss.n7556 avss.n7555 0.0147424
R26545 avss.n7009 avss.n6957 0.0147424
R26546 avss.n7203 avss.n7202 0.0147424
R26547 avss.n6656 avss.n6604 0.0147424
R26548 avss.n6850 avss.n6849 0.0147424
R26549 avss.n6303 avss.n6251 0.0147424
R26550 avss.n6497 avss.n6496 0.0147424
R26551 avss.n5950 avss.n5898 0.0147424
R26552 avss.n6144 avss.n6143 0.0147424
R26553 avss.n5597 avss.n5545 0.0147424
R26554 avss.n5791 avss.n5790 0.0147424
R26555 avss.n5252 avss.n5199 0.0147424
R26556 avss.n5438 avss.n5437 0.0147424
R26557 avss.n4898 avss.n4845 0.0147424
R26558 avss.n5084 avss.n5083 0.0147424
R26559 avss.n9191 avss.n9100 0.0147424
R26560 avss.n9081 avss.n9080 0.0147424
R26561 avss.n9412 avss.n9321 0.0147424
R26562 avss.n9302 avss.n9301 0.0147424
R26563 avss.n9633 avss.n9542 0.0147424
R26564 avss.n9523 avss.n9522 0.0147424
R26565 avss.n9854 avss.n9763 0.0147424
R26566 avss.n9744 avss.n9743 0.0147424
R26567 avss.n10075 avss.n9984 0.0147424
R26568 avss.n9965 avss.n9964 0.0147424
R26569 avss.n10296 avss.n10205 0.0147424
R26570 avss.n10186 avss.n10185 0.0147424
R26571 avss.n10517 avss.n10426 0.0147424
R26572 avss.n10407 avss.n10406 0.0147424
R26573 avss.n10738 avss.n10647 0.0147424
R26574 avss.n10628 avss.n10627 0.0147424
R26575 avss.n10959 avss.n10868 0.0147424
R26576 avss.n10849 avss.n10848 0.0147424
R26577 avss.n11180 avss.n11089 0.0147424
R26578 avss.n11070 avss.n11069 0.0147424
R26579 avss.n432 avss.n340 0.0147424
R26580 avss.n11291 avss.n11290 0.0147424
R26581 avss.n215 avss.n123 0.0147424
R26582 avss.n11512 avss.n11511 0.0147424
R26583 avss.n3393 avss.n3392 0.0145625
R26584 avss.n2680 avss.n2679 0.0145006
R26585 avss.n2650 avss.n2649 0.0145006
R26586 avss.n2799 avss.n2798 0.0145006
R26587 avss.n2802 avss.n2797 0.0145006
R26588 avss.n3617 avss.n3616 0.0145006
R26589 avss.n3025 avss.n3024 0.0145006
R26590 avss.n2968 avss.n2967 0.0145006
R26591 avss.n2924 avss.n2923 0.0145006
R26592 avss.n8652 avss.n8624 0.0140303
R26593 avss.n8775 avss.n8774 0.0140303
R26594 avss.n8650 avss.n8623 0.0140303
R26595 avss.n8776 avss.n8721 0.0140303
R26596 avss.n8842 avss.n3717 0.0140303
R26597 avss.n8968 avss.n3673 0.0140303
R26598 avss.n8841 avss.n8840 0.0140303
R26599 avss.n8923 avss.n3674 0.0140303
R26600 avss.n8299 avss.n8271 0.0140303
R26601 avss.n8422 avss.n8421 0.0140303
R26602 avss.n8297 avss.n8270 0.0140303
R26603 avss.n8423 avss.n8368 0.0140303
R26604 avss.n8489 avss.n3801 0.0140303
R26605 avss.n8615 avss.n3757 0.0140303
R26606 avss.n8488 avss.n8487 0.0140303
R26607 avss.n8570 avss.n3758 0.0140303
R26608 avss.n7946 avss.n7918 0.0140303
R26609 avss.n8069 avss.n8068 0.0140303
R26610 avss.n7944 avss.n7917 0.0140303
R26611 avss.n8070 avss.n8015 0.0140303
R26612 avss.n8136 avss.n3885 0.0140303
R26613 avss.n8262 avss.n3841 0.0140303
R26614 avss.n8135 avss.n8134 0.0140303
R26615 avss.n8217 avss.n3842 0.0140303
R26616 avss.n7593 avss.n7565 0.0140303
R26617 avss.n7716 avss.n7715 0.0140303
R26618 avss.n7591 avss.n7564 0.0140303
R26619 avss.n7717 avss.n7662 0.0140303
R26620 avss.n7783 avss.n3969 0.0140303
R26621 avss.n7909 avss.n3925 0.0140303
R26622 avss.n7782 avss.n7781 0.0140303
R26623 avss.n7864 avss.n3926 0.0140303
R26624 avss.n7240 avss.n7212 0.0140303
R26625 avss.n7363 avss.n7362 0.0140303
R26626 avss.n7238 avss.n7211 0.0140303
R26627 avss.n7364 avss.n7309 0.0140303
R26628 avss.n7430 avss.n4053 0.0140303
R26629 avss.n7556 avss.n4009 0.0140303
R26630 avss.n7429 avss.n7428 0.0140303
R26631 avss.n7511 avss.n4010 0.0140303
R26632 avss.n6887 avss.n6859 0.0140303
R26633 avss.n7010 avss.n7009 0.0140303
R26634 avss.n6885 avss.n6858 0.0140303
R26635 avss.n7011 avss.n6956 0.0140303
R26636 avss.n7077 avss.n4137 0.0140303
R26637 avss.n7203 avss.n4093 0.0140303
R26638 avss.n7076 avss.n7075 0.0140303
R26639 avss.n7158 avss.n4094 0.0140303
R26640 avss.n6534 avss.n6506 0.0140303
R26641 avss.n6657 avss.n6656 0.0140303
R26642 avss.n6532 avss.n6505 0.0140303
R26643 avss.n6658 avss.n6603 0.0140303
R26644 avss.n6724 avss.n4221 0.0140303
R26645 avss.n6850 avss.n4177 0.0140303
R26646 avss.n6723 avss.n6722 0.0140303
R26647 avss.n6805 avss.n4178 0.0140303
R26648 avss.n6181 avss.n6153 0.0140303
R26649 avss.n6304 avss.n6303 0.0140303
R26650 avss.n6179 avss.n6152 0.0140303
R26651 avss.n6305 avss.n6250 0.0140303
R26652 avss.n6371 avss.n4305 0.0140303
R26653 avss.n6497 avss.n4261 0.0140303
R26654 avss.n6370 avss.n6369 0.0140303
R26655 avss.n6452 avss.n4262 0.0140303
R26656 avss.n5828 avss.n5800 0.0140303
R26657 avss.n5951 avss.n5950 0.0140303
R26658 avss.n5826 avss.n5799 0.0140303
R26659 avss.n5952 avss.n5897 0.0140303
R26660 avss.n6018 avss.n4389 0.0140303
R26661 avss.n6144 avss.n4345 0.0140303
R26662 avss.n6017 avss.n6016 0.0140303
R26663 avss.n6099 avss.n4346 0.0140303
R26664 avss.n5475 avss.n5447 0.0140303
R26665 avss.n5598 avss.n5597 0.0140303
R26666 avss.n5473 avss.n5446 0.0140303
R26667 avss.n5599 avss.n5544 0.0140303
R26668 avss.n5665 avss.n4473 0.0140303
R26669 avss.n5791 avss.n4429 0.0140303
R26670 avss.n5664 avss.n5663 0.0140303
R26671 avss.n5746 avss.n4430 0.0140303
R26672 avss.n5300 avss.n5299 0.0140303
R26673 avss.n5253 avss.n5252 0.0140303
R26674 avss.n5301 avss.n5092 0.0140303
R26675 avss.n5254 avss.n5198 0.0140303
R26676 avss.n5312 avss.n4557 0.0140303
R26677 avss.n5438 avss.n4513 0.0140303
R26678 avss.n5311 avss.n5310 0.0140303
R26679 avss.n5393 avss.n4514 0.0140303
R26680 avss.n4946 avss.n4945 0.0140303
R26681 avss.n4899 avss.n4898 0.0140303
R26682 avss.n4947 avss.n4738 0.0140303
R26683 avss.n4900 avss.n4844 0.0140303
R26684 avss.n4958 avss.n4641 0.0140303
R26685 avss.n5084 avss.n4597 0.0140303
R26686 avss.n4957 avss.n4956 0.0140303
R26687 avss.n5039 avss.n4598 0.0140303
R26688 avss.n2393 avss.n2392 0.0140303
R26689 avss.n9191 avss.n9190 0.0140303
R26690 avss.n2481 avss.n2480 0.0140303
R26691 avss.n9157 avss.n9156 0.0140303
R26692 avss.n2591 avss.n2590 0.0140303
R26693 avss.n9081 avss.n8989 0.0140303
R26694 avss.n2538 avss.n2537 0.0140303
R26695 avss.n9046 avss.n9045 0.0140303
R26696 avss.n2177 avss.n2176 0.0140303
R26697 avss.n9412 avss.n9411 0.0140303
R26698 avss.n2265 avss.n2264 0.0140303
R26699 avss.n9378 avss.n9377 0.0140303
R26700 avss.n2375 avss.n2374 0.0140303
R26701 avss.n9302 avss.n9210 0.0140303
R26702 avss.n2322 avss.n2321 0.0140303
R26703 avss.n9267 avss.n9266 0.0140303
R26704 avss.n1961 avss.n1960 0.0140303
R26705 avss.n9633 avss.n9632 0.0140303
R26706 avss.n2049 avss.n2048 0.0140303
R26707 avss.n9599 avss.n9598 0.0140303
R26708 avss.n2159 avss.n2158 0.0140303
R26709 avss.n9523 avss.n9431 0.0140303
R26710 avss.n2106 avss.n2105 0.0140303
R26711 avss.n9488 avss.n9487 0.0140303
R26712 avss.n1745 avss.n1744 0.0140303
R26713 avss.n9854 avss.n9853 0.0140303
R26714 avss.n1833 avss.n1832 0.0140303
R26715 avss.n9820 avss.n9819 0.0140303
R26716 avss.n1943 avss.n1942 0.0140303
R26717 avss.n9744 avss.n9652 0.0140303
R26718 avss.n1890 avss.n1889 0.0140303
R26719 avss.n9709 avss.n9708 0.0140303
R26720 avss.n1529 avss.n1528 0.0140303
R26721 avss.n10075 avss.n10074 0.0140303
R26722 avss.n1617 avss.n1616 0.0140303
R26723 avss.n10041 avss.n10040 0.0140303
R26724 avss.n1727 avss.n1726 0.0140303
R26725 avss.n9965 avss.n9873 0.0140303
R26726 avss.n1674 avss.n1673 0.0140303
R26727 avss.n9930 avss.n9929 0.0140303
R26728 avss.n1313 avss.n1312 0.0140303
R26729 avss.n10296 avss.n10295 0.0140303
R26730 avss.n1401 avss.n1400 0.0140303
R26731 avss.n10262 avss.n10261 0.0140303
R26732 avss.n1511 avss.n1510 0.0140303
R26733 avss.n10186 avss.n10094 0.0140303
R26734 avss.n1458 avss.n1457 0.0140303
R26735 avss.n10151 avss.n10150 0.0140303
R26736 avss.n1097 avss.n1096 0.0140303
R26737 avss.n10517 avss.n10516 0.0140303
R26738 avss.n1185 avss.n1184 0.0140303
R26739 avss.n10483 avss.n10482 0.0140303
R26740 avss.n1295 avss.n1294 0.0140303
R26741 avss.n10407 avss.n10315 0.0140303
R26742 avss.n1242 avss.n1241 0.0140303
R26743 avss.n10372 avss.n10371 0.0140303
R26744 avss.n881 avss.n880 0.0140303
R26745 avss.n10738 avss.n10737 0.0140303
R26746 avss.n969 avss.n968 0.0140303
R26747 avss.n10704 avss.n10703 0.0140303
R26748 avss.n1079 avss.n1078 0.0140303
R26749 avss.n10628 avss.n10536 0.0140303
R26750 avss.n1026 avss.n1025 0.0140303
R26751 avss.n10593 avss.n10592 0.0140303
R26752 avss.n665 avss.n664 0.0140303
R26753 avss.n10959 avss.n10958 0.0140303
R26754 avss.n753 avss.n752 0.0140303
R26755 avss.n10925 avss.n10924 0.0140303
R26756 avss.n863 avss.n862 0.0140303
R26757 avss.n10849 avss.n10757 0.0140303
R26758 avss.n810 avss.n809 0.0140303
R26759 avss.n10814 avss.n10813 0.0140303
R26760 avss.n449 avss.n448 0.0140303
R26761 avss.n11180 avss.n11179 0.0140303
R26762 avss.n537 avss.n536 0.0140303
R26763 avss.n11146 avss.n11145 0.0140303
R26764 avss.n647 avss.n646 0.0140303
R26765 avss.n11070 avss.n10978 0.0140303
R26766 avss.n594 avss.n593 0.0140303
R26767 avss.n11035 avss.n11034 0.0140303
R26768 avss.n11312 avss.n11311 0.0140303
R26769 avss.n432 avss.n355 0.0140303
R26770 avss.n11366 avss.n11365 0.0140303
R26771 avss.n413 avss.n412 0.0140303
R26772 avss.n322 avss.n321 0.0140303
R26773 avss.n11291 avss.n11199 0.0140303
R26774 avss.n269 avss.n268 0.0140303
R26775 avss.n11256 avss.n11255 0.0140303
R26776 avss.n11533 avss.n11532 0.0140303
R26777 avss.n215 avss.n138 0.0140303
R26778 avss.n11587 avss.n11586 0.0140303
R26779 avss.n196 avss.n195 0.0140303
R26780 avss.n105 avss.n104 0.0140303
R26781 avss.n11512 avss.n11420 0.0140303
R26782 avss.n52 avss.n51 0.0140303
R26783 avss.n11477 avss.n11476 0.0140303
R26784 avss.n8694 avss.n8686 0.0133182
R26785 avss.n8892 avss.n8891 0.0133182
R26786 avss.n8341 avss.n8333 0.0133182
R26787 avss.n8539 avss.n8538 0.0133182
R26788 avss.n7988 avss.n7980 0.0133182
R26789 avss.n8186 avss.n8185 0.0133182
R26790 avss.n7635 avss.n7627 0.0133182
R26791 avss.n7833 avss.n7832 0.0133182
R26792 avss.n7282 avss.n7274 0.0133182
R26793 avss.n7480 avss.n7479 0.0133182
R26794 avss.n6929 avss.n6921 0.0133182
R26795 avss.n7127 avss.n7126 0.0133182
R26796 avss.n6576 avss.n6568 0.0133182
R26797 avss.n6774 avss.n6773 0.0133182
R26798 avss.n6223 avss.n6215 0.0133182
R26799 avss.n6421 avss.n6420 0.0133182
R26800 avss.n5870 avss.n5862 0.0133182
R26801 avss.n6068 avss.n6067 0.0133182
R26802 avss.n5517 avss.n5509 0.0133182
R26803 avss.n5715 avss.n5714 0.0133182
R26804 avss.n5171 avss.n5163 0.0133182
R26805 avss.n5362 avss.n5361 0.0133182
R26806 avss.n4817 avss.n4809 0.0133182
R26807 avss.n5008 avss.n5007 0.0133182
R26808 avss.n2431 avss.n2430 0.0133182
R26809 avss.n2488 avss.n2487 0.0133182
R26810 avss.n2215 avss.n2214 0.0133182
R26811 avss.n2272 avss.n2271 0.0133182
R26812 avss.n1999 avss.n1998 0.0133182
R26813 avss.n2056 avss.n2055 0.0133182
R26814 avss.n1783 avss.n1782 0.0133182
R26815 avss.n1840 avss.n1839 0.0133182
R26816 avss.n1567 avss.n1566 0.0133182
R26817 avss.n1624 avss.n1623 0.0133182
R26818 avss.n1351 avss.n1350 0.0133182
R26819 avss.n1408 avss.n1407 0.0133182
R26820 avss.n1135 avss.n1134 0.0133182
R26821 avss.n1192 avss.n1191 0.0133182
R26822 avss.n919 avss.n918 0.0133182
R26823 avss.n976 avss.n975 0.0133182
R26824 avss.n703 avss.n702 0.0133182
R26825 avss.n760 avss.n759 0.0133182
R26826 avss.n487 avss.n486 0.0133182
R26827 avss.n544 avss.n543 0.0133182
R26828 avss.n11316 avss.n11315 0.0133182
R26829 avss.n219 avss.n218 0.0133182
R26830 avss.n11537 avss.n11536 0.0133182
R26831 avss.n2 avss.n1 0.0133182
R26832 avss.n3353 avss.n3352 0.013
R26833 avss.n3368 avss.n3367 0.013
R26834 avss.n3406 avss.n3242 0.013
R26835 avss.n8710 avss.n8699 0.0126061
R26836 avss.n8641 avss.n8625 0.0126061
R26837 avss.n8642 avss.n8632 0.0126061
R26838 avss.n8831 avss.n8628 0.0126061
R26839 avss.n8657 avss.n8651 0.0126061
R26840 avss.n8674 avss.n8673 0.0126061
R26841 avss.n8688 avss.n8671 0.0126061
R26842 avss.n8711 avss.n8709 0.0126061
R26843 avss.n8788 avss.n8787 0.0126061
R26844 avss.n8738 avss.n8731 0.0126061
R26845 avss.n8767 avss.n8766 0.0126061
R26846 avss.n3741 avss.n3724 0.0126061
R26847 avss.n8910 avss.n8909 0.0126061
R26848 avss.n3742 avss.n3732 0.0126061
R26849 avss.n3751 avss.n3728 0.0126061
R26850 avss.n8850 avss.n3719 0.0126061
R26851 avss.n3712 avss.n3709 0.0126061
R26852 avss.n8883 avss.n3704 0.0126061
R26853 avss.n8911 avss.n3695 0.0126061
R26854 avss.n8920 avss.n3691 0.0126061
R26855 avss.n8938 avss.n8937 0.0126061
R26856 avss.n8948 avss.n8947 0.0126061
R26857 avss.n8357 avss.n8346 0.0126061
R26858 avss.n8288 avss.n8272 0.0126061
R26859 avss.n8289 avss.n8279 0.0126061
R26860 avss.n8478 avss.n8275 0.0126061
R26861 avss.n8304 avss.n8298 0.0126061
R26862 avss.n8321 avss.n8320 0.0126061
R26863 avss.n8335 avss.n8318 0.0126061
R26864 avss.n8358 avss.n8356 0.0126061
R26865 avss.n8435 avss.n8434 0.0126061
R26866 avss.n8385 avss.n8378 0.0126061
R26867 avss.n8414 avss.n8413 0.0126061
R26868 avss.n3825 avss.n3808 0.0126061
R26869 avss.n8557 avss.n8556 0.0126061
R26870 avss.n3826 avss.n3816 0.0126061
R26871 avss.n3835 avss.n3812 0.0126061
R26872 avss.n8497 avss.n3803 0.0126061
R26873 avss.n3796 avss.n3793 0.0126061
R26874 avss.n8530 avss.n3788 0.0126061
R26875 avss.n8558 avss.n3779 0.0126061
R26876 avss.n8567 avss.n3775 0.0126061
R26877 avss.n8585 avss.n8584 0.0126061
R26878 avss.n8595 avss.n8594 0.0126061
R26879 avss.n8004 avss.n7993 0.0126061
R26880 avss.n7935 avss.n7919 0.0126061
R26881 avss.n7936 avss.n7926 0.0126061
R26882 avss.n8125 avss.n7922 0.0126061
R26883 avss.n7951 avss.n7945 0.0126061
R26884 avss.n7968 avss.n7967 0.0126061
R26885 avss.n7982 avss.n7965 0.0126061
R26886 avss.n8005 avss.n8003 0.0126061
R26887 avss.n8082 avss.n8081 0.0126061
R26888 avss.n8032 avss.n8025 0.0126061
R26889 avss.n8061 avss.n8060 0.0126061
R26890 avss.n3909 avss.n3892 0.0126061
R26891 avss.n8204 avss.n8203 0.0126061
R26892 avss.n3910 avss.n3900 0.0126061
R26893 avss.n3919 avss.n3896 0.0126061
R26894 avss.n8144 avss.n3887 0.0126061
R26895 avss.n3880 avss.n3877 0.0126061
R26896 avss.n8177 avss.n3872 0.0126061
R26897 avss.n8205 avss.n3863 0.0126061
R26898 avss.n8214 avss.n3859 0.0126061
R26899 avss.n8232 avss.n8231 0.0126061
R26900 avss.n8242 avss.n8241 0.0126061
R26901 avss.n7651 avss.n7640 0.0126061
R26902 avss.n7582 avss.n7566 0.0126061
R26903 avss.n7583 avss.n7573 0.0126061
R26904 avss.n7772 avss.n7569 0.0126061
R26905 avss.n7598 avss.n7592 0.0126061
R26906 avss.n7615 avss.n7614 0.0126061
R26907 avss.n7629 avss.n7612 0.0126061
R26908 avss.n7652 avss.n7650 0.0126061
R26909 avss.n7729 avss.n7728 0.0126061
R26910 avss.n7679 avss.n7672 0.0126061
R26911 avss.n7708 avss.n7707 0.0126061
R26912 avss.n3993 avss.n3976 0.0126061
R26913 avss.n7851 avss.n7850 0.0126061
R26914 avss.n3994 avss.n3984 0.0126061
R26915 avss.n4003 avss.n3980 0.0126061
R26916 avss.n7791 avss.n3971 0.0126061
R26917 avss.n3964 avss.n3961 0.0126061
R26918 avss.n7824 avss.n3956 0.0126061
R26919 avss.n7852 avss.n3947 0.0126061
R26920 avss.n7861 avss.n3943 0.0126061
R26921 avss.n7879 avss.n7878 0.0126061
R26922 avss.n7889 avss.n7888 0.0126061
R26923 avss.n7298 avss.n7287 0.0126061
R26924 avss.n7229 avss.n7213 0.0126061
R26925 avss.n7230 avss.n7220 0.0126061
R26926 avss.n7419 avss.n7216 0.0126061
R26927 avss.n7245 avss.n7239 0.0126061
R26928 avss.n7262 avss.n7261 0.0126061
R26929 avss.n7276 avss.n7259 0.0126061
R26930 avss.n7299 avss.n7297 0.0126061
R26931 avss.n7376 avss.n7375 0.0126061
R26932 avss.n7326 avss.n7319 0.0126061
R26933 avss.n7355 avss.n7354 0.0126061
R26934 avss.n4077 avss.n4060 0.0126061
R26935 avss.n7498 avss.n7497 0.0126061
R26936 avss.n4078 avss.n4068 0.0126061
R26937 avss.n4087 avss.n4064 0.0126061
R26938 avss.n7438 avss.n4055 0.0126061
R26939 avss.n4048 avss.n4045 0.0126061
R26940 avss.n7471 avss.n4040 0.0126061
R26941 avss.n7499 avss.n4031 0.0126061
R26942 avss.n7508 avss.n4027 0.0126061
R26943 avss.n7526 avss.n7525 0.0126061
R26944 avss.n7536 avss.n7535 0.0126061
R26945 avss.n6945 avss.n6934 0.0126061
R26946 avss.n6876 avss.n6860 0.0126061
R26947 avss.n6877 avss.n6867 0.0126061
R26948 avss.n7066 avss.n6863 0.0126061
R26949 avss.n6892 avss.n6886 0.0126061
R26950 avss.n6909 avss.n6908 0.0126061
R26951 avss.n6923 avss.n6906 0.0126061
R26952 avss.n6946 avss.n6944 0.0126061
R26953 avss.n7023 avss.n7022 0.0126061
R26954 avss.n6973 avss.n6966 0.0126061
R26955 avss.n7002 avss.n7001 0.0126061
R26956 avss.n4161 avss.n4144 0.0126061
R26957 avss.n7145 avss.n7144 0.0126061
R26958 avss.n4162 avss.n4152 0.0126061
R26959 avss.n4171 avss.n4148 0.0126061
R26960 avss.n7085 avss.n4139 0.0126061
R26961 avss.n4132 avss.n4129 0.0126061
R26962 avss.n7118 avss.n4124 0.0126061
R26963 avss.n7146 avss.n4115 0.0126061
R26964 avss.n7155 avss.n4111 0.0126061
R26965 avss.n7173 avss.n7172 0.0126061
R26966 avss.n7183 avss.n7182 0.0126061
R26967 avss.n6592 avss.n6581 0.0126061
R26968 avss.n6523 avss.n6507 0.0126061
R26969 avss.n6524 avss.n6514 0.0126061
R26970 avss.n6713 avss.n6510 0.0126061
R26971 avss.n6539 avss.n6533 0.0126061
R26972 avss.n6556 avss.n6555 0.0126061
R26973 avss.n6570 avss.n6553 0.0126061
R26974 avss.n6593 avss.n6591 0.0126061
R26975 avss.n6670 avss.n6669 0.0126061
R26976 avss.n6620 avss.n6613 0.0126061
R26977 avss.n6649 avss.n6648 0.0126061
R26978 avss.n4245 avss.n4228 0.0126061
R26979 avss.n6792 avss.n6791 0.0126061
R26980 avss.n4246 avss.n4236 0.0126061
R26981 avss.n4255 avss.n4232 0.0126061
R26982 avss.n6732 avss.n4223 0.0126061
R26983 avss.n4216 avss.n4213 0.0126061
R26984 avss.n6765 avss.n4208 0.0126061
R26985 avss.n6793 avss.n4199 0.0126061
R26986 avss.n6802 avss.n4195 0.0126061
R26987 avss.n6820 avss.n6819 0.0126061
R26988 avss.n6830 avss.n6829 0.0126061
R26989 avss.n6239 avss.n6228 0.0126061
R26990 avss.n6170 avss.n6154 0.0126061
R26991 avss.n6171 avss.n6161 0.0126061
R26992 avss.n6360 avss.n6157 0.0126061
R26993 avss.n6186 avss.n6180 0.0126061
R26994 avss.n6203 avss.n6202 0.0126061
R26995 avss.n6217 avss.n6200 0.0126061
R26996 avss.n6240 avss.n6238 0.0126061
R26997 avss.n6317 avss.n6316 0.0126061
R26998 avss.n6267 avss.n6260 0.0126061
R26999 avss.n6296 avss.n6295 0.0126061
R27000 avss.n4329 avss.n4312 0.0126061
R27001 avss.n6439 avss.n6438 0.0126061
R27002 avss.n4330 avss.n4320 0.0126061
R27003 avss.n4339 avss.n4316 0.0126061
R27004 avss.n6379 avss.n4307 0.0126061
R27005 avss.n4300 avss.n4297 0.0126061
R27006 avss.n6412 avss.n4292 0.0126061
R27007 avss.n6440 avss.n4283 0.0126061
R27008 avss.n6449 avss.n4279 0.0126061
R27009 avss.n6467 avss.n6466 0.0126061
R27010 avss.n6477 avss.n6476 0.0126061
R27011 avss.n5886 avss.n5875 0.0126061
R27012 avss.n5817 avss.n5801 0.0126061
R27013 avss.n5818 avss.n5808 0.0126061
R27014 avss.n6007 avss.n5804 0.0126061
R27015 avss.n5833 avss.n5827 0.0126061
R27016 avss.n5850 avss.n5849 0.0126061
R27017 avss.n5864 avss.n5847 0.0126061
R27018 avss.n5887 avss.n5885 0.0126061
R27019 avss.n5964 avss.n5963 0.0126061
R27020 avss.n5914 avss.n5907 0.0126061
R27021 avss.n5943 avss.n5942 0.0126061
R27022 avss.n4413 avss.n4396 0.0126061
R27023 avss.n6086 avss.n6085 0.0126061
R27024 avss.n4414 avss.n4404 0.0126061
R27025 avss.n4423 avss.n4400 0.0126061
R27026 avss.n6026 avss.n4391 0.0126061
R27027 avss.n4384 avss.n4381 0.0126061
R27028 avss.n6059 avss.n4376 0.0126061
R27029 avss.n6087 avss.n4367 0.0126061
R27030 avss.n6096 avss.n4363 0.0126061
R27031 avss.n6114 avss.n6113 0.0126061
R27032 avss.n6124 avss.n6123 0.0126061
R27033 avss.n5533 avss.n5522 0.0126061
R27034 avss.n5464 avss.n5448 0.0126061
R27035 avss.n5465 avss.n5455 0.0126061
R27036 avss.n5654 avss.n5451 0.0126061
R27037 avss.n5480 avss.n5474 0.0126061
R27038 avss.n5497 avss.n5496 0.0126061
R27039 avss.n5511 avss.n5494 0.0126061
R27040 avss.n5534 avss.n5532 0.0126061
R27041 avss.n5611 avss.n5610 0.0126061
R27042 avss.n5561 avss.n5554 0.0126061
R27043 avss.n5590 avss.n5589 0.0126061
R27044 avss.n4497 avss.n4480 0.0126061
R27045 avss.n5733 avss.n5732 0.0126061
R27046 avss.n4498 avss.n4488 0.0126061
R27047 avss.n4507 avss.n4484 0.0126061
R27048 avss.n5673 avss.n4475 0.0126061
R27049 avss.n4468 avss.n4465 0.0126061
R27050 avss.n5706 avss.n4460 0.0126061
R27051 avss.n5734 avss.n4451 0.0126061
R27052 avss.n5743 avss.n4447 0.0126061
R27053 avss.n5761 avss.n5760 0.0126061
R27054 avss.n5771 avss.n5770 0.0126061
R27055 avss.n5187 avss.n5176 0.0126061
R27056 avss.n5117 avss.n5116 0.0126061
R27057 avss.n5118 avss.n5107 0.0126061
R27058 avss.n5125 avss.n5102 0.0126061
R27059 avss.n5098 avss.n5095 0.0126061
R27060 avss.n5151 avss.n5150 0.0126061
R27061 avss.n5165 avss.n5148 0.0126061
R27062 avss.n5188 avss.n5186 0.0126061
R27063 avss.n5266 avss.n5265 0.0126061
R27064 avss.n5221 avss.n5214 0.0126061
R27065 avss.n5211 avss.n5207 0.0126061
R27066 avss.n4581 avss.n4564 0.0126061
R27067 avss.n5380 avss.n5379 0.0126061
R27068 avss.n4582 avss.n4572 0.0126061
R27069 avss.n4591 avss.n4568 0.0126061
R27070 avss.n5320 avss.n4559 0.0126061
R27071 avss.n4552 avss.n4549 0.0126061
R27072 avss.n5353 avss.n4544 0.0126061
R27073 avss.n5381 avss.n4535 0.0126061
R27074 avss.n5390 avss.n4531 0.0126061
R27075 avss.n5408 avss.n5407 0.0126061
R27076 avss.n5418 avss.n5417 0.0126061
R27077 avss.n4833 avss.n4822 0.0126061
R27078 avss.n4763 avss.n4762 0.0126061
R27079 avss.n4764 avss.n4753 0.0126061
R27080 avss.n4771 avss.n4748 0.0126061
R27081 avss.n4744 avss.n4741 0.0126061
R27082 avss.n4797 avss.n4796 0.0126061
R27083 avss.n4811 avss.n4794 0.0126061
R27084 avss.n4834 avss.n4832 0.0126061
R27085 avss.n4912 avss.n4911 0.0126061
R27086 avss.n4867 avss.n4860 0.0126061
R27087 avss.n4857 avss.n4853 0.0126061
R27088 avss.n4665 avss.n4648 0.0126061
R27089 avss.n5026 avss.n5025 0.0126061
R27090 avss.n4666 avss.n4656 0.0126061
R27091 avss.n4675 avss.n4652 0.0126061
R27092 avss.n4966 avss.n4643 0.0126061
R27093 avss.n4636 avss.n4633 0.0126061
R27094 avss.n4999 avss.n4628 0.0126061
R27095 avss.n5027 avss.n4619 0.0126061
R27096 avss.n5036 avss.n4615 0.0126061
R27097 avss.n5054 avss.n5053 0.0126061
R27098 avss.n5064 avss.n5063 0.0126061
R27099 avss.n9181 avss.n9180 0.0126061
R27100 avss.n2427 avss.n2426 0.0126061
R27101 avss.n2411 avss.n2410 0.0126061
R27102 avss.n2407 avss.n2406 0.0126061
R27103 avss.n2477 avss.n2467 0.0126061
R27104 avss.n2457 avss.n2448 0.0126061
R27105 avss.n2443 avss.n2442 0.0126061
R27106 avss.n9136 avss.n9135 0.0126061
R27107 avss.n9149 avss.n9140 0.0126061
R27108 avss.n9170 avss.n9169 0.0126061
R27109 avss.n9114 avss.n9103 0.0126061
R27110 avss.n2574 avss.n2573 0.0126061
R27111 avss.n8980 avss.n8979 0.0126061
R27112 avss.n2558 avss.n2557 0.0126061
R27113 avss.n2554 avss.n2553 0.0126061
R27114 avss.n2534 avss.n2524 0.0126061
R27115 avss.n2514 avss.n2505 0.0126061
R27116 avss.n2500 avss.n2499 0.0126061
R27117 avss.n9025 avss.n9024 0.0126061
R27118 avss.n9038 avss.n9029 0.0126061
R27119 avss.n9059 avss.n9058 0.0126061
R27120 avss.n9002 avss.n8991 0.0126061
R27121 avss.n9402 avss.n9401 0.0126061
R27122 avss.n2211 avss.n2210 0.0126061
R27123 avss.n2195 avss.n2194 0.0126061
R27124 avss.n2191 avss.n2190 0.0126061
R27125 avss.n2261 avss.n2251 0.0126061
R27126 avss.n2241 avss.n2232 0.0126061
R27127 avss.n2227 avss.n2226 0.0126061
R27128 avss.n9357 avss.n9356 0.0126061
R27129 avss.n9370 avss.n9361 0.0126061
R27130 avss.n9391 avss.n9390 0.0126061
R27131 avss.n9335 avss.n9324 0.0126061
R27132 avss.n2358 avss.n2357 0.0126061
R27133 avss.n9201 avss.n9200 0.0126061
R27134 avss.n2342 avss.n2341 0.0126061
R27135 avss.n2338 avss.n2337 0.0126061
R27136 avss.n2318 avss.n2308 0.0126061
R27137 avss.n2298 avss.n2289 0.0126061
R27138 avss.n2284 avss.n2283 0.0126061
R27139 avss.n9246 avss.n9245 0.0126061
R27140 avss.n9259 avss.n9250 0.0126061
R27141 avss.n9280 avss.n9279 0.0126061
R27142 avss.n9223 avss.n9212 0.0126061
R27143 avss.n9623 avss.n9622 0.0126061
R27144 avss.n1995 avss.n1994 0.0126061
R27145 avss.n1979 avss.n1978 0.0126061
R27146 avss.n1975 avss.n1974 0.0126061
R27147 avss.n2045 avss.n2035 0.0126061
R27148 avss.n2025 avss.n2016 0.0126061
R27149 avss.n2011 avss.n2010 0.0126061
R27150 avss.n9578 avss.n9577 0.0126061
R27151 avss.n9591 avss.n9582 0.0126061
R27152 avss.n9612 avss.n9611 0.0126061
R27153 avss.n9556 avss.n9545 0.0126061
R27154 avss.n2142 avss.n2141 0.0126061
R27155 avss.n9422 avss.n9421 0.0126061
R27156 avss.n2126 avss.n2125 0.0126061
R27157 avss.n2122 avss.n2121 0.0126061
R27158 avss.n2102 avss.n2092 0.0126061
R27159 avss.n2082 avss.n2073 0.0126061
R27160 avss.n2068 avss.n2067 0.0126061
R27161 avss.n9467 avss.n9466 0.0126061
R27162 avss.n9480 avss.n9471 0.0126061
R27163 avss.n9501 avss.n9500 0.0126061
R27164 avss.n9444 avss.n9433 0.0126061
R27165 avss.n9844 avss.n9843 0.0126061
R27166 avss.n1779 avss.n1778 0.0126061
R27167 avss.n1763 avss.n1762 0.0126061
R27168 avss.n1759 avss.n1758 0.0126061
R27169 avss.n1829 avss.n1819 0.0126061
R27170 avss.n1809 avss.n1800 0.0126061
R27171 avss.n1795 avss.n1794 0.0126061
R27172 avss.n9799 avss.n9798 0.0126061
R27173 avss.n9812 avss.n9803 0.0126061
R27174 avss.n9833 avss.n9832 0.0126061
R27175 avss.n9777 avss.n9766 0.0126061
R27176 avss.n1926 avss.n1925 0.0126061
R27177 avss.n9643 avss.n9642 0.0126061
R27178 avss.n1910 avss.n1909 0.0126061
R27179 avss.n1906 avss.n1905 0.0126061
R27180 avss.n1886 avss.n1876 0.0126061
R27181 avss.n1866 avss.n1857 0.0126061
R27182 avss.n1852 avss.n1851 0.0126061
R27183 avss.n9688 avss.n9687 0.0126061
R27184 avss.n9701 avss.n9692 0.0126061
R27185 avss.n9722 avss.n9721 0.0126061
R27186 avss.n9665 avss.n9654 0.0126061
R27187 avss.n10065 avss.n10064 0.0126061
R27188 avss.n1563 avss.n1562 0.0126061
R27189 avss.n1547 avss.n1546 0.0126061
R27190 avss.n1543 avss.n1542 0.0126061
R27191 avss.n1613 avss.n1603 0.0126061
R27192 avss.n1593 avss.n1584 0.0126061
R27193 avss.n1579 avss.n1578 0.0126061
R27194 avss.n10020 avss.n10019 0.0126061
R27195 avss.n10033 avss.n10024 0.0126061
R27196 avss.n10054 avss.n10053 0.0126061
R27197 avss.n9998 avss.n9987 0.0126061
R27198 avss.n1710 avss.n1709 0.0126061
R27199 avss.n9864 avss.n9863 0.0126061
R27200 avss.n1694 avss.n1693 0.0126061
R27201 avss.n1690 avss.n1689 0.0126061
R27202 avss.n1670 avss.n1660 0.0126061
R27203 avss.n1650 avss.n1641 0.0126061
R27204 avss.n1636 avss.n1635 0.0126061
R27205 avss.n9909 avss.n9908 0.0126061
R27206 avss.n9922 avss.n9913 0.0126061
R27207 avss.n9943 avss.n9942 0.0126061
R27208 avss.n9886 avss.n9875 0.0126061
R27209 avss.n10286 avss.n10285 0.0126061
R27210 avss.n1347 avss.n1346 0.0126061
R27211 avss.n1331 avss.n1330 0.0126061
R27212 avss.n1327 avss.n1326 0.0126061
R27213 avss.n1397 avss.n1387 0.0126061
R27214 avss.n1377 avss.n1368 0.0126061
R27215 avss.n1363 avss.n1362 0.0126061
R27216 avss.n10241 avss.n10240 0.0126061
R27217 avss.n10254 avss.n10245 0.0126061
R27218 avss.n10275 avss.n10274 0.0126061
R27219 avss.n10219 avss.n10208 0.0126061
R27220 avss.n1494 avss.n1493 0.0126061
R27221 avss.n10085 avss.n10084 0.0126061
R27222 avss.n1478 avss.n1477 0.0126061
R27223 avss.n1474 avss.n1473 0.0126061
R27224 avss.n1454 avss.n1444 0.0126061
R27225 avss.n1434 avss.n1425 0.0126061
R27226 avss.n1420 avss.n1419 0.0126061
R27227 avss.n10130 avss.n10129 0.0126061
R27228 avss.n10143 avss.n10134 0.0126061
R27229 avss.n10164 avss.n10163 0.0126061
R27230 avss.n10107 avss.n10096 0.0126061
R27231 avss.n10507 avss.n10506 0.0126061
R27232 avss.n1131 avss.n1130 0.0126061
R27233 avss.n1115 avss.n1114 0.0126061
R27234 avss.n1111 avss.n1110 0.0126061
R27235 avss.n1181 avss.n1171 0.0126061
R27236 avss.n1161 avss.n1152 0.0126061
R27237 avss.n1147 avss.n1146 0.0126061
R27238 avss.n10462 avss.n10461 0.0126061
R27239 avss.n10475 avss.n10466 0.0126061
R27240 avss.n10496 avss.n10495 0.0126061
R27241 avss.n10440 avss.n10429 0.0126061
R27242 avss.n1278 avss.n1277 0.0126061
R27243 avss.n10306 avss.n10305 0.0126061
R27244 avss.n1262 avss.n1261 0.0126061
R27245 avss.n1258 avss.n1257 0.0126061
R27246 avss.n1238 avss.n1228 0.0126061
R27247 avss.n1218 avss.n1209 0.0126061
R27248 avss.n1204 avss.n1203 0.0126061
R27249 avss.n10351 avss.n10350 0.0126061
R27250 avss.n10364 avss.n10355 0.0126061
R27251 avss.n10385 avss.n10384 0.0126061
R27252 avss.n10328 avss.n10317 0.0126061
R27253 avss.n10728 avss.n10727 0.0126061
R27254 avss.n915 avss.n914 0.0126061
R27255 avss.n899 avss.n898 0.0126061
R27256 avss.n895 avss.n894 0.0126061
R27257 avss.n965 avss.n955 0.0126061
R27258 avss.n945 avss.n936 0.0126061
R27259 avss.n931 avss.n930 0.0126061
R27260 avss.n10683 avss.n10682 0.0126061
R27261 avss.n10696 avss.n10687 0.0126061
R27262 avss.n10717 avss.n10716 0.0126061
R27263 avss.n10661 avss.n10650 0.0126061
R27264 avss.n1062 avss.n1061 0.0126061
R27265 avss.n10527 avss.n10526 0.0126061
R27266 avss.n1046 avss.n1045 0.0126061
R27267 avss.n1042 avss.n1041 0.0126061
R27268 avss.n1022 avss.n1012 0.0126061
R27269 avss.n1002 avss.n993 0.0126061
R27270 avss.n988 avss.n987 0.0126061
R27271 avss.n10572 avss.n10571 0.0126061
R27272 avss.n10585 avss.n10576 0.0126061
R27273 avss.n10606 avss.n10605 0.0126061
R27274 avss.n10549 avss.n10538 0.0126061
R27275 avss.n10949 avss.n10948 0.0126061
R27276 avss.n699 avss.n698 0.0126061
R27277 avss.n683 avss.n682 0.0126061
R27278 avss.n679 avss.n678 0.0126061
R27279 avss.n749 avss.n739 0.0126061
R27280 avss.n729 avss.n720 0.0126061
R27281 avss.n715 avss.n714 0.0126061
R27282 avss.n10904 avss.n10903 0.0126061
R27283 avss.n10917 avss.n10908 0.0126061
R27284 avss.n10938 avss.n10937 0.0126061
R27285 avss.n10882 avss.n10871 0.0126061
R27286 avss.n846 avss.n845 0.0126061
R27287 avss.n10748 avss.n10747 0.0126061
R27288 avss.n830 avss.n829 0.0126061
R27289 avss.n826 avss.n825 0.0126061
R27290 avss.n806 avss.n796 0.0126061
R27291 avss.n786 avss.n777 0.0126061
R27292 avss.n772 avss.n771 0.0126061
R27293 avss.n10793 avss.n10792 0.0126061
R27294 avss.n10806 avss.n10797 0.0126061
R27295 avss.n10827 avss.n10826 0.0126061
R27296 avss.n10770 avss.n10759 0.0126061
R27297 avss.n11170 avss.n11169 0.0126061
R27298 avss.n483 avss.n482 0.0126061
R27299 avss.n467 avss.n466 0.0126061
R27300 avss.n463 avss.n462 0.0126061
R27301 avss.n533 avss.n523 0.0126061
R27302 avss.n513 avss.n504 0.0126061
R27303 avss.n499 avss.n498 0.0126061
R27304 avss.n11125 avss.n11124 0.0126061
R27305 avss.n11138 avss.n11129 0.0126061
R27306 avss.n11159 avss.n11158 0.0126061
R27307 avss.n11103 avss.n11092 0.0126061
R27308 avss.n630 avss.n629 0.0126061
R27309 avss.n10969 avss.n10968 0.0126061
R27310 avss.n614 avss.n613 0.0126061
R27311 avss.n610 avss.n609 0.0126061
R27312 avss.n590 avss.n580 0.0126061
R27313 avss.n570 avss.n561 0.0126061
R27314 avss.n556 avss.n555 0.0126061
R27315 avss.n11014 avss.n11013 0.0126061
R27316 avss.n11027 avss.n11018 0.0126061
R27317 avss.n11048 avss.n11047 0.0126061
R27318 avss.n10991 avss.n10980 0.0126061
R27319 avss.n346 avss.n345 0.0126061
R27320 avss.n11402 avss.n11401 0.0126061
R27321 avss.n11386 avss.n11385 0.0126061
R27322 avss.n11381 avss.n11380 0.0126061
R27323 avss.n11362 avss.n11352 0.0126061
R27324 avss.n11342 avss.n11333 0.0126061
R27325 avss.n11328 avss.n11327 0.0126061
R27326 avss.n392 avss.n391 0.0126061
R27327 avss.n405 avss.n396 0.0126061
R27328 avss.n426 avss.n425 0.0126061
R27329 avss.n369 avss.n358 0.0126061
R27330 avss.n305 avss.n304 0.0126061
R27331 avss.n11190 avss.n11189 0.0126061
R27332 avss.n289 avss.n288 0.0126061
R27333 avss.n285 avss.n284 0.0126061
R27334 avss.n265 avss.n255 0.0126061
R27335 avss.n245 avss.n236 0.0126061
R27336 avss.n231 avss.n230 0.0126061
R27337 avss.n11235 avss.n11234 0.0126061
R27338 avss.n11248 avss.n11239 0.0126061
R27339 avss.n11269 avss.n11268 0.0126061
R27340 avss.n11212 avss.n11201 0.0126061
R27341 avss.n129 avss.n128 0.0126061
R27342 avss.n11623 avss.n11622 0.0126061
R27343 avss.n11607 avss.n11606 0.0126061
R27344 avss.n11602 avss.n11601 0.0126061
R27345 avss.n11583 avss.n11573 0.0126061
R27346 avss.n11563 avss.n11554 0.0126061
R27347 avss.n11549 avss.n11548 0.0126061
R27348 avss.n175 avss.n174 0.0126061
R27349 avss.n188 avss.n179 0.0126061
R27350 avss.n209 avss.n208 0.0126061
R27351 avss.n152 avss.n141 0.0126061
R27352 avss.n88 avss.n87 0.0126061
R27353 avss.n11411 avss.n11410 0.0126061
R27354 avss.n72 avss.n71 0.0126061
R27355 avss.n68 avss.n67 0.0126061
R27356 avss.n48 avss.n38 0.0126061
R27357 avss.n28 avss.n19 0.0126061
R27358 avss.n14 avss.n13 0.0126061
R27359 avss.n11456 avss.n11455 0.0126061
R27360 avss.n11469 avss.n11460 0.0126061
R27361 avss.n11490 avss.n11489 0.0126061
R27362 avss.n11433 avss.n11422 0.0126061
R27363 avss.n8740 avss.n8725 0.0120023
R27364 avss.n8728 avss.n8725 0.0120023
R27365 avss.n8387 avss.n8372 0.0120023
R27366 avss.n8375 avss.n8372 0.0120023
R27367 avss.n8034 avss.n8019 0.0120023
R27368 avss.n8022 avss.n8019 0.0120023
R27369 avss.n7681 avss.n7666 0.0120023
R27370 avss.n7669 avss.n7666 0.0120023
R27371 avss.n7328 avss.n7313 0.0120023
R27372 avss.n7316 avss.n7313 0.0120023
R27373 avss.n6975 avss.n6960 0.0120023
R27374 avss.n6963 avss.n6960 0.0120023
R27375 avss.n6622 avss.n6607 0.0120023
R27376 avss.n6610 avss.n6607 0.0120023
R27377 avss.n6269 avss.n6254 0.0120023
R27378 avss.n6257 avss.n6254 0.0120023
R27379 avss.n5916 avss.n5901 0.0120023
R27380 avss.n5904 avss.n5901 0.0120023
R27381 avss.n5563 avss.n5548 0.0120023
R27382 avss.n5551 avss.n5548 0.0120023
R27383 avss.n5205 avss.n5204 0.0120023
R27384 avss.n5223 avss.n5205 0.0120023
R27385 avss.n4851 avss.n4850 0.0120023
R27386 avss.n4869 avss.n4851 0.0120023
R27387 avss.n9173 avss.n9172 0.0120023
R27388 avss.n9174 avss.n9173 0.0120023
R27389 avss.n9394 avss.n9393 0.0120023
R27390 avss.n9395 avss.n9394 0.0120023
R27391 avss.n9615 avss.n9614 0.0120023
R27392 avss.n9616 avss.n9615 0.0120023
R27393 avss.n9836 avss.n9835 0.0120023
R27394 avss.n9837 avss.n9836 0.0120023
R27395 avss.n10057 avss.n10056 0.0120023
R27396 avss.n10058 avss.n10057 0.0120023
R27397 avss.n10278 avss.n10277 0.0120023
R27398 avss.n10279 avss.n10278 0.0120023
R27399 avss.n10499 avss.n10498 0.0120023
R27400 avss.n10500 avss.n10499 0.0120023
R27401 avss.n10720 avss.n10719 0.0120023
R27402 avss.n10721 avss.n10720 0.0120023
R27403 avss.n10941 avss.n10940 0.0120023
R27404 avss.n10942 avss.n10941 0.0120023
R27405 avss.n11162 avss.n11161 0.0120023
R27406 avss.n11163 avss.n11162 0.0120023
R27407 avss.n430 avss.n429 0.0120023
R27408 avss.n429 avss.n428 0.0120023
R27409 avss.n213 avss.n212 0.0120023
R27410 avss.n212 avss.n211 0.0120023
R27411 avss.n8811 avss.n8662 0.0118939
R27412 avss.n8859 avss.n8857 0.0118939
R27413 avss.n8458 avss.n8309 0.0118939
R27414 avss.n8506 avss.n8504 0.0118939
R27415 avss.n8105 avss.n7956 0.0118939
R27416 avss.n8153 avss.n8151 0.0118939
R27417 avss.n7752 avss.n7603 0.0118939
R27418 avss.n7800 avss.n7798 0.0118939
R27419 avss.n7399 avss.n7250 0.0118939
R27420 avss.n7447 avss.n7445 0.0118939
R27421 avss.n7046 avss.n6897 0.0118939
R27422 avss.n7094 avss.n7092 0.0118939
R27423 avss.n6693 avss.n6544 0.0118939
R27424 avss.n6741 avss.n6739 0.0118939
R27425 avss.n6340 avss.n6191 0.0118939
R27426 avss.n6388 avss.n6386 0.0118939
R27427 avss.n5987 avss.n5838 0.0118939
R27428 avss.n6035 avss.n6033 0.0118939
R27429 avss.n5634 avss.n5485 0.0118939
R27430 avss.n5682 avss.n5680 0.0118939
R27431 avss.n5289 avss.n5135 0.0118939
R27432 avss.n5329 avss.n5327 0.0118939
R27433 avss.n4935 avss.n4781 0.0118939
R27434 avss.n4975 avss.n4973 0.0118939
R27435 avss.n2461 avss.n2460 0.0118939
R27436 avss.n2518 avss.n2517 0.0118939
R27437 avss.n2245 avss.n2244 0.0118939
R27438 avss.n2302 avss.n2301 0.0118939
R27439 avss.n2029 avss.n2028 0.0118939
R27440 avss.n2086 avss.n2085 0.0118939
R27441 avss.n1813 avss.n1812 0.0118939
R27442 avss.n1870 avss.n1869 0.0118939
R27443 avss.n1597 avss.n1596 0.0118939
R27444 avss.n1654 avss.n1653 0.0118939
R27445 avss.n1381 avss.n1380 0.0118939
R27446 avss.n1438 avss.n1437 0.0118939
R27447 avss.n1165 avss.n1164 0.0118939
R27448 avss.n1222 avss.n1221 0.0118939
R27449 avss.n949 avss.n948 0.0118939
R27450 avss.n1006 avss.n1005 0.0118939
R27451 avss.n733 avss.n732 0.0118939
R27452 avss.n790 avss.n789 0.0118939
R27453 avss.n517 avss.n516 0.0118939
R27454 avss.n574 avss.n573 0.0118939
R27455 avss.n11346 avss.n11345 0.0118939
R27456 avss.n249 avss.n248 0.0118939
R27457 avss.n11567 avss.n11566 0.0118939
R27458 avss.n32 avss.n31 0.0118939
R27459 avss.n8793 avss.n8792 0.0118636
R27460 avss.n8644 avss.n8630 0.0118636
R27461 avss.n3744 avss.n3730 0.0118636
R27462 avss.n8913 avss.n3693 0.0118636
R27463 avss.n8440 avss.n8439 0.0118636
R27464 avss.n8291 avss.n8277 0.0118636
R27465 avss.n3828 avss.n3814 0.0118636
R27466 avss.n8560 avss.n3777 0.0118636
R27467 avss.n8087 avss.n8086 0.0118636
R27468 avss.n7938 avss.n7924 0.0118636
R27469 avss.n3912 avss.n3898 0.0118636
R27470 avss.n8207 avss.n3861 0.0118636
R27471 avss.n7734 avss.n7733 0.0118636
R27472 avss.n7585 avss.n7571 0.0118636
R27473 avss.n3996 avss.n3982 0.0118636
R27474 avss.n7854 avss.n3945 0.0118636
R27475 avss.n7381 avss.n7380 0.0118636
R27476 avss.n7232 avss.n7218 0.0118636
R27477 avss.n4080 avss.n4066 0.0118636
R27478 avss.n7501 avss.n4029 0.0118636
R27479 avss.n7028 avss.n7027 0.0118636
R27480 avss.n6879 avss.n6865 0.0118636
R27481 avss.n4164 avss.n4150 0.0118636
R27482 avss.n7148 avss.n4113 0.0118636
R27483 avss.n6675 avss.n6674 0.0118636
R27484 avss.n6526 avss.n6512 0.0118636
R27485 avss.n4248 avss.n4234 0.0118636
R27486 avss.n6795 avss.n4197 0.0118636
R27487 avss.n6322 avss.n6321 0.0118636
R27488 avss.n6173 avss.n6159 0.0118636
R27489 avss.n4332 avss.n4318 0.0118636
R27490 avss.n6442 avss.n4281 0.0118636
R27491 avss.n5969 avss.n5968 0.0118636
R27492 avss.n5820 avss.n5806 0.0118636
R27493 avss.n4416 avss.n4402 0.0118636
R27494 avss.n6089 avss.n4365 0.0118636
R27495 avss.n5616 avss.n5615 0.0118636
R27496 avss.n5467 avss.n5453 0.0118636
R27497 avss.n4500 avss.n4486 0.0118636
R27498 avss.n5736 avss.n4449 0.0118636
R27499 avss.n5271 avss.n5270 0.0118636
R27500 avss.n5120 avss.n5104 0.0118636
R27501 avss.n4584 avss.n4570 0.0118636
R27502 avss.n5383 avss.n4533 0.0118636
R27503 avss.n4917 avss.n4916 0.0118636
R27504 avss.n4766 avss.n4750 0.0118636
R27505 avss.n4668 avss.n4654 0.0118636
R27506 avss.n5029 avss.n4617 0.0118636
R27507 avss.n9130 avss.n9129 0.0118636
R27508 avss.n2419 avss.n2418 0.0118636
R27509 avss.n2566 avss.n2565 0.0118636
R27510 avss.n9019 avss.n9018 0.0118636
R27511 avss.n9351 avss.n9350 0.0118636
R27512 avss.n2203 avss.n2202 0.0118636
R27513 avss.n2350 avss.n2349 0.0118636
R27514 avss.n9240 avss.n9239 0.0118636
R27515 avss.n9572 avss.n9571 0.0118636
R27516 avss.n1987 avss.n1986 0.0118636
R27517 avss.n2134 avss.n2133 0.0118636
R27518 avss.n9461 avss.n9460 0.0118636
R27519 avss.n9793 avss.n9792 0.0118636
R27520 avss.n1771 avss.n1770 0.0118636
R27521 avss.n1918 avss.n1917 0.0118636
R27522 avss.n9682 avss.n9681 0.0118636
R27523 avss.n10014 avss.n10013 0.0118636
R27524 avss.n1555 avss.n1554 0.0118636
R27525 avss.n1702 avss.n1701 0.0118636
R27526 avss.n9903 avss.n9902 0.0118636
R27527 avss.n10235 avss.n10234 0.0118636
R27528 avss.n1339 avss.n1338 0.0118636
R27529 avss.n1486 avss.n1485 0.0118636
R27530 avss.n10124 avss.n10123 0.0118636
R27531 avss.n10456 avss.n10455 0.0118636
R27532 avss.n1123 avss.n1122 0.0118636
R27533 avss.n1270 avss.n1269 0.0118636
R27534 avss.n10345 avss.n10344 0.0118636
R27535 avss.n10677 avss.n10676 0.0118636
R27536 avss.n907 avss.n906 0.0118636
R27537 avss.n1054 avss.n1053 0.0118636
R27538 avss.n10566 avss.n10565 0.0118636
R27539 avss.n10898 avss.n10897 0.0118636
R27540 avss.n691 avss.n690 0.0118636
R27541 avss.n838 avss.n837 0.0118636
R27542 avss.n10787 avss.n10786 0.0118636
R27543 avss.n11119 avss.n11118 0.0118636
R27544 avss.n475 avss.n474 0.0118636
R27545 avss.n622 avss.n621 0.0118636
R27546 avss.n11008 avss.n11007 0.0118636
R27547 avss.n386 avss.n385 0.0118636
R27548 avss.n11394 avss.n11393 0.0118636
R27549 avss.n297 avss.n296 0.0118636
R27550 avss.n11229 avss.n11228 0.0118636
R27551 avss.n169 avss.n168 0.0118636
R27552 avss.n11615 avss.n11614 0.0118636
R27553 avss.n80 avss.n79 0.0118636
R27554 avss.n11450 avss.n11449 0.0118636
R27555 avss.n8795 avss.n8699 0.0111818
R27556 avss.n8641 avss.n8640 0.0111818
R27557 avss.n8827 avss.n8826 0.0111818
R27558 avss.n8786 avss.n8717 0.0111818
R27559 avss.n3741 avss.n3740 0.0111818
R27560 avss.n8910 avss.n8904 0.0111818
R27561 avss.n3747 avss.n3722 0.0111818
R27562 avss.n8916 avss.n3687 0.0111818
R27563 avss.n8442 avss.n8346 0.0111818
R27564 avss.n8288 avss.n8287 0.0111818
R27565 avss.n8474 avss.n8473 0.0111818
R27566 avss.n8433 avss.n8364 0.0111818
R27567 avss.n3825 avss.n3824 0.0111818
R27568 avss.n8557 avss.n8551 0.0111818
R27569 avss.n3831 avss.n3806 0.0111818
R27570 avss.n8563 avss.n3771 0.0111818
R27571 avss.n8089 avss.n7993 0.0111818
R27572 avss.n7935 avss.n7934 0.0111818
R27573 avss.n8121 avss.n8120 0.0111818
R27574 avss.n8080 avss.n8011 0.0111818
R27575 avss.n3909 avss.n3908 0.0111818
R27576 avss.n8204 avss.n8198 0.0111818
R27577 avss.n3915 avss.n3890 0.0111818
R27578 avss.n8210 avss.n3855 0.0111818
R27579 avss.n7736 avss.n7640 0.0111818
R27580 avss.n7582 avss.n7581 0.0111818
R27581 avss.n7768 avss.n7767 0.0111818
R27582 avss.n7727 avss.n7658 0.0111818
R27583 avss.n3993 avss.n3992 0.0111818
R27584 avss.n7851 avss.n7845 0.0111818
R27585 avss.n3999 avss.n3974 0.0111818
R27586 avss.n7857 avss.n3939 0.0111818
R27587 avss.n7383 avss.n7287 0.0111818
R27588 avss.n7229 avss.n7228 0.0111818
R27589 avss.n7415 avss.n7414 0.0111818
R27590 avss.n7374 avss.n7305 0.0111818
R27591 avss.n4077 avss.n4076 0.0111818
R27592 avss.n7498 avss.n7492 0.0111818
R27593 avss.n4083 avss.n4058 0.0111818
R27594 avss.n7504 avss.n4023 0.0111818
R27595 avss.n7030 avss.n6934 0.0111818
R27596 avss.n6876 avss.n6875 0.0111818
R27597 avss.n7062 avss.n7061 0.0111818
R27598 avss.n7021 avss.n6952 0.0111818
R27599 avss.n4161 avss.n4160 0.0111818
R27600 avss.n7145 avss.n7139 0.0111818
R27601 avss.n4167 avss.n4142 0.0111818
R27602 avss.n7151 avss.n4107 0.0111818
R27603 avss.n6677 avss.n6581 0.0111818
R27604 avss.n6523 avss.n6522 0.0111818
R27605 avss.n6709 avss.n6708 0.0111818
R27606 avss.n6668 avss.n6599 0.0111818
R27607 avss.n4245 avss.n4244 0.0111818
R27608 avss.n6792 avss.n6786 0.0111818
R27609 avss.n4251 avss.n4226 0.0111818
R27610 avss.n6798 avss.n4191 0.0111818
R27611 avss.n6324 avss.n6228 0.0111818
R27612 avss.n6170 avss.n6169 0.0111818
R27613 avss.n6356 avss.n6355 0.0111818
R27614 avss.n6315 avss.n6246 0.0111818
R27615 avss.n4329 avss.n4328 0.0111818
R27616 avss.n6439 avss.n6433 0.0111818
R27617 avss.n4335 avss.n4310 0.0111818
R27618 avss.n6445 avss.n4275 0.0111818
R27619 avss.n5971 avss.n5875 0.0111818
R27620 avss.n5817 avss.n5816 0.0111818
R27621 avss.n6003 avss.n6002 0.0111818
R27622 avss.n5962 avss.n5893 0.0111818
R27623 avss.n4413 avss.n4412 0.0111818
R27624 avss.n6086 avss.n6080 0.0111818
R27625 avss.n4419 avss.n4394 0.0111818
R27626 avss.n6092 avss.n4359 0.0111818
R27627 avss.n5618 avss.n5522 0.0111818
R27628 avss.n5464 avss.n5463 0.0111818
R27629 avss.n5650 avss.n5649 0.0111818
R27630 avss.n5609 avss.n5540 0.0111818
R27631 avss.n4497 avss.n4496 0.0111818
R27632 avss.n5733 avss.n5727 0.0111818
R27633 avss.n4503 avss.n4478 0.0111818
R27634 avss.n5739 avss.n4443 0.0111818
R27635 avss.n5273 avss.n5176 0.0111818
R27636 avss.n5117 avss.n5115 0.0111818
R27637 avss.n5127 avss.n5126 0.0111818
R27638 avss.n5264 avss.n5194 0.0111818
R27639 avss.n4581 avss.n4580 0.0111818
R27640 avss.n5380 avss.n5374 0.0111818
R27641 avss.n4587 avss.n4562 0.0111818
R27642 avss.n5386 avss.n4527 0.0111818
R27643 avss.n4919 avss.n4822 0.0111818
R27644 avss.n4763 avss.n4761 0.0111818
R27645 avss.n4773 avss.n4772 0.0111818
R27646 avss.n4910 avss.n4840 0.0111818
R27647 avss.n4665 avss.n4664 0.0111818
R27648 avss.n5026 avss.n5020 0.0111818
R27649 avss.n4671 avss.n4646 0.0111818
R27650 avss.n5032 avss.n4611 0.0111818
R27651 avss.n9180 avss.n9179 0.0111818
R27652 avss.n2426 avss.n2425 0.0111818
R27653 avss.n2397 avss.n2396 0.0111818
R27654 avss.n9151 avss.n9150 0.0111818
R27655 avss.n2573 avss.n2572 0.0111818
R27656 avss.n8979 avss.n8978 0.0111818
R27657 avss.n2544 avss.n2543 0.0111818
R27658 avss.n9040 avss.n9039 0.0111818
R27659 avss.n9401 avss.n9400 0.0111818
R27660 avss.n2210 avss.n2209 0.0111818
R27661 avss.n2181 avss.n2180 0.0111818
R27662 avss.n9372 avss.n9371 0.0111818
R27663 avss.n2357 avss.n2356 0.0111818
R27664 avss.n9200 avss.n9199 0.0111818
R27665 avss.n2328 avss.n2327 0.0111818
R27666 avss.n9261 avss.n9260 0.0111818
R27667 avss.n9622 avss.n9621 0.0111818
R27668 avss.n1994 avss.n1993 0.0111818
R27669 avss.n1965 avss.n1964 0.0111818
R27670 avss.n9593 avss.n9592 0.0111818
R27671 avss.n2141 avss.n2140 0.0111818
R27672 avss.n9421 avss.n9420 0.0111818
R27673 avss.n2112 avss.n2111 0.0111818
R27674 avss.n9482 avss.n9481 0.0111818
R27675 avss.n9843 avss.n9842 0.0111818
R27676 avss.n1778 avss.n1777 0.0111818
R27677 avss.n1749 avss.n1748 0.0111818
R27678 avss.n9814 avss.n9813 0.0111818
R27679 avss.n1925 avss.n1924 0.0111818
R27680 avss.n9642 avss.n9641 0.0111818
R27681 avss.n1896 avss.n1895 0.0111818
R27682 avss.n9703 avss.n9702 0.0111818
R27683 avss.n10064 avss.n10063 0.0111818
R27684 avss.n1562 avss.n1561 0.0111818
R27685 avss.n1533 avss.n1532 0.0111818
R27686 avss.n10035 avss.n10034 0.0111818
R27687 avss.n1709 avss.n1708 0.0111818
R27688 avss.n9863 avss.n9862 0.0111818
R27689 avss.n1680 avss.n1679 0.0111818
R27690 avss.n9924 avss.n9923 0.0111818
R27691 avss.n10285 avss.n10284 0.0111818
R27692 avss.n1346 avss.n1345 0.0111818
R27693 avss.n1317 avss.n1316 0.0111818
R27694 avss.n10256 avss.n10255 0.0111818
R27695 avss.n1493 avss.n1492 0.0111818
R27696 avss.n10084 avss.n10083 0.0111818
R27697 avss.n1464 avss.n1463 0.0111818
R27698 avss.n10145 avss.n10144 0.0111818
R27699 avss.n10506 avss.n10505 0.0111818
R27700 avss.n1130 avss.n1129 0.0111818
R27701 avss.n1101 avss.n1100 0.0111818
R27702 avss.n10477 avss.n10476 0.0111818
R27703 avss.n1277 avss.n1276 0.0111818
R27704 avss.n10305 avss.n10304 0.0111818
R27705 avss.n1248 avss.n1247 0.0111818
R27706 avss.n10366 avss.n10365 0.0111818
R27707 avss.n10727 avss.n10726 0.0111818
R27708 avss.n914 avss.n913 0.0111818
R27709 avss.n885 avss.n884 0.0111818
R27710 avss.n10698 avss.n10697 0.0111818
R27711 avss.n1061 avss.n1060 0.0111818
R27712 avss.n10526 avss.n10525 0.0111818
R27713 avss.n1032 avss.n1031 0.0111818
R27714 avss.n10587 avss.n10586 0.0111818
R27715 avss.n10948 avss.n10947 0.0111818
R27716 avss.n698 avss.n697 0.0111818
R27717 avss.n669 avss.n668 0.0111818
R27718 avss.n10919 avss.n10918 0.0111818
R27719 avss.n845 avss.n844 0.0111818
R27720 avss.n10747 avss.n10746 0.0111818
R27721 avss.n816 avss.n815 0.0111818
R27722 avss.n10808 avss.n10807 0.0111818
R27723 avss.n11169 avss.n11168 0.0111818
R27724 avss.n482 avss.n481 0.0111818
R27725 avss.n453 avss.n452 0.0111818
R27726 avss.n11140 avss.n11139 0.0111818
R27727 avss.n629 avss.n628 0.0111818
R27728 avss.n10968 avss.n10967 0.0111818
R27729 avss.n600 avss.n599 0.0111818
R27730 avss.n11029 avss.n11028 0.0111818
R27731 avss.n345 avss.n344 0.0111818
R27732 avss.n11401 avss.n11400 0.0111818
R27733 avss.n11371 avss.n11370 0.0111818
R27734 avss.n407 avss.n406 0.0111818
R27735 avss.n304 avss.n303 0.0111818
R27736 avss.n11189 avss.n11188 0.0111818
R27737 avss.n275 avss.n274 0.0111818
R27738 avss.n11250 avss.n11249 0.0111818
R27739 avss.n128 avss.n127 0.0111818
R27740 avss.n11622 avss.n11621 0.0111818
R27741 avss.n11592 avss.n11591 0.0111818
R27742 avss.n190 avss.n189 0.0111818
R27743 avss.n87 avss.n86 0.0111818
R27744 avss.n11410 avss.n11409 0.0111818
R27745 avss.n58 avss.n57 0.0111818
R27746 avss.n11471 avss.n11470 0.0111818
R27747 avss.n3351 avss.n3292 0.0109167
R27748 avss.n8634 avss.n8633 0.0104697
R27749 avss.n8702 avss.n8700 0.0104697
R27750 avss.n3734 avss.n3733 0.0104697
R27751 avss.n8898 avss.n8897 0.0104697
R27752 avss.n8281 avss.n8280 0.0104697
R27753 avss.n8349 avss.n8347 0.0104697
R27754 avss.n3818 avss.n3817 0.0104697
R27755 avss.n8545 avss.n8544 0.0104697
R27756 avss.n7928 avss.n7927 0.0104697
R27757 avss.n7996 avss.n7994 0.0104697
R27758 avss.n3902 avss.n3901 0.0104697
R27759 avss.n8192 avss.n8191 0.0104697
R27760 avss.n7575 avss.n7574 0.0104697
R27761 avss.n7643 avss.n7641 0.0104697
R27762 avss.n3986 avss.n3985 0.0104697
R27763 avss.n7839 avss.n7838 0.0104697
R27764 avss.n7222 avss.n7221 0.0104697
R27765 avss.n7290 avss.n7288 0.0104697
R27766 avss.n4070 avss.n4069 0.0104697
R27767 avss.n7486 avss.n7485 0.0104697
R27768 avss.n6869 avss.n6868 0.0104697
R27769 avss.n6937 avss.n6935 0.0104697
R27770 avss.n4154 avss.n4153 0.0104697
R27771 avss.n7133 avss.n7132 0.0104697
R27772 avss.n6516 avss.n6515 0.0104697
R27773 avss.n6584 avss.n6582 0.0104697
R27774 avss.n4238 avss.n4237 0.0104697
R27775 avss.n6780 avss.n6779 0.0104697
R27776 avss.n6163 avss.n6162 0.0104697
R27777 avss.n6231 avss.n6229 0.0104697
R27778 avss.n4322 avss.n4321 0.0104697
R27779 avss.n6427 avss.n6426 0.0104697
R27780 avss.n5810 avss.n5809 0.0104697
R27781 avss.n5878 avss.n5876 0.0104697
R27782 avss.n4406 avss.n4405 0.0104697
R27783 avss.n6074 avss.n6073 0.0104697
R27784 avss.n5457 avss.n5456 0.0104697
R27785 avss.n5525 avss.n5523 0.0104697
R27786 avss.n4490 avss.n4489 0.0104697
R27787 avss.n5721 avss.n5720 0.0104697
R27788 avss.n5109 avss.n5108 0.0104697
R27789 avss.n5179 avss.n5177 0.0104697
R27790 avss.n4574 avss.n4573 0.0104697
R27791 avss.n5368 avss.n5367 0.0104697
R27792 avss.n4755 avss.n4754 0.0104697
R27793 avss.n4825 avss.n4823 0.0104697
R27794 avss.n4658 avss.n4657 0.0104697
R27795 avss.n5014 avss.n5013 0.0104697
R27796 avss.n2422 avss.n2421 0.0104697
R27797 avss.n9132 avss.n9122 0.0104697
R27798 avss.n2569 avss.n2568 0.0104697
R27799 avss.n9021 avss.n9011 0.0104697
R27800 avss.n2206 avss.n2205 0.0104697
R27801 avss.n9353 avss.n9343 0.0104697
R27802 avss.n2353 avss.n2352 0.0104697
R27803 avss.n9242 avss.n9232 0.0104697
R27804 avss.n1990 avss.n1989 0.0104697
R27805 avss.n9574 avss.n9564 0.0104697
R27806 avss.n2137 avss.n2136 0.0104697
R27807 avss.n9463 avss.n9453 0.0104697
R27808 avss.n1774 avss.n1773 0.0104697
R27809 avss.n9795 avss.n9785 0.0104697
R27810 avss.n1921 avss.n1920 0.0104697
R27811 avss.n9684 avss.n9674 0.0104697
R27812 avss.n1558 avss.n1557 0.0104697
R27813 avss.n10016 avss.n10006 0.0104697
R27814 avss.n1705 avss.n1704 0.0104697
R27815 avss.n9905 avss.n9895 0.0104697
R27816 avss.n1342 avss.n1341 0.0104697
R27817 avss.n10237 avss.n10227 0.0104697
R27818 avss.n1489 avss.n1488 0.0104697
R27819 avss.n10126 avss.n10116 0.0104697
R27820 avss.n1126 avss.n1125 0.0104697
R27821 avss.n10458 avss.n10448 0.0104697
R27822 avss.n1273 avss.n1272 0.0104697
R27823 avss.n10347 avss.n10337 0.0104697
R27824 avss.n910 avss.n909 0.0104697
R27825 avss.n10679 avss.n10669 0.0104697
R27826 avss.n1057 avss.n1056 0.0104697
R27827 avss.n10568 avss.n10558 0.0104697
R27828 avss.n694 avss.n693 0.0104697
R27829 avss.n10900 avss.n10890 0.0104697
R27830 avss.n841 avss.n840 0.0104697
R27831 avss.n10789 avss.n10779 0.0104697
R27832 avss.n478 avss.n477 0.0104697
R27833 avss.n11121 avss.n11111 0.0104697
R27834 avss.n625 avss.n624 0.0104697
R27835 avss.n11010 avss.n11000 0.0104697
R27836 avss.n11397 avss.n11396 0.0104697
R27837 avss.n388 avss.n378 0.0104697
R27838 avss.n300 avss.n299 0.0104697
R27839 avss.n11231 avss.n11221 0.0104697
R27840 avss.n11618 avss.n11617 0.0104697
R27841 avss.n171 avss.n161 0.0104697
R27842 avss.n83 avss.n82 0.0104697
R27843 avss.n11452 avss.n11442 0.0104697
R27844 avss.n8974 avss 0.0103377
R27845 avss.n8818 avss.n8652 0.00975758
R27846 avss.n8855 avss.n3717 0.00975758
R27847 avss.n8465 avss.n8299 0.00975758
R27848 avss.n8502 avss.n3801 0.00975758
R27849 avss.n8112 avss.n7946 0.00975758
R27850 avss.n8149 avss.n3885 0.00975758
R27851 avss.n7759 avss.n7593 0.00975758
R27852 avss.n7796 avss.n3969 0.00975758
R27853 avss.n7406 avss.n7240 0.00975758
R27854 avss.n7443 avss.n4053 0.00975758
R27855 avss.n7053 avss.n6887 0.00975758
R27856 avss.n7090 avss.n4137 0.00975758
R27857 avss.n6700 avss.n6534 0.00975758
R27858 avss.n6737 avss.n4221 0.00975758
R27859 avss.n6347 avss.n6181 0.00975758
R27860 avss.n6384 avss.n4305 0.00975758
R27861 avss.n5994 avss.n5828 0.00975758
R27862 avss.n6031 avss.n4389 0.00975758
R27863 avss.n5641 avss.n5475 0.00975758
R27864 avss.n5678 avss.n4473 0.00975758
R27865 avss.n5299 avss.n5298 0.00975758
R27866 avss.n5325 avss.n4557 0.00975758
R27867 avss.n4945 avss.n4944 0.00975758
R27868 avss.n4971 avss.n4641 0.00975758
R27869 avss.n2392 avss.n2391 0.00975758
R27870 avss.n2590 avss.n2589 0.00975758
R27871 avss.n2176 avss.n2175 0.00975758
R27872 avss.n2374 avss.n2373 0.00975758
R27873 avss.n1960 avss.n1959 0.00975758
R27874 avss.n2158 avss.n2157 0.00975758
R27875 avss.n1744 avss.n1743 0.00975758
R27876 avss.n1942 avss.n1941 0.00975758
R27877 avss.n1528 avss.n1527 0.00975758
R27878 avss.n1726 avss.n1725 0.00975758
R27879 avss.n1312 avss.n1311 0.00975758
R27880 avss.n1510 avss.n1509 0.00975758
R27881 avss.n1096 avss.n1095 0.00975758
R27882 avss.n1294 avss.n1293 0.00975758
R27883 avss.n880 avss.n879 0.00975758
R27884 avss.n1078 avss.n1077 0.00975758
R27885 avss.n664 avss.n663 0.00975758
R27886 avss.n862 avss.n861 0.00975758
R27887 avss.n448 avss.n447 0.00975758
R27888 avss.n646 avss.n645 0.00975758
R27889 avss.n11311 avss.n11310 0.00975758
R27890 avss.n321 avss.n320 0.00975758
R27891 avss.n11532 avss.n11531 0.00975758
R27892 avss.n104 avss.n103 0.00975758
R27893 avss.n8845 avss.n8844 0.00916977
R27894 avss.n8844 avss.n3723 0.00916977
R27895 avss.n8492 avss.n8491 0.00916977
R27896 avss.n8491 avss.n3807 0.00916977
R27897 avss.n8139 avss.n8138 0.00916977
R27898 avss.n8138 avss.n3891 0.00916977
R27899 avss.n7786 avss.n7785 0.00916977
R27900 avss.n7785 avss.n3975 0.00916977
R27901 avss.n7433 avss.n7432 0.00916977
R27902 avss.n7432 avss.n4059 0.00916977
R27903 avss.n7080 avss.n7079 0.00916977
R27904 avss.n7079 avss.n4143 0.00916977
R27905 avss.n6727 avss.n6726 0.00916977
R27906 avss.n6726 avss.n4227 0.00916977
R27907 avss.n6374 avss.n6373 0.00916977
R27908 avss.n6373 avss.n4311 0.00916977
R27909 avss.n6021 avss.n6020 0.00916977
R27910 avss.n6020 avss.n4395 0.00916977
R27911 avss.n5668 avss.n5667 0.00916977
R27912 avss.n5667 avss.n4479 0.00916977
R27913 avss.n5315 avss.n5314 0.00916977
R27914 avss.n5314 avss.n4563 0.00916977
R27915 avss.n4961 avss.n4960 0.00916977
R27916 avss.n4960 avss.n4647 0.00916977
R27917 avss.n2542 avss.n2541 0.00916977
R27918 avss.n2541 avss.n2540 0.00916977
R27919 avss.n2326 avss.n2325 0.00916977
R27920 avss.n2325 avss.n2324 0.00916977
R27921 avss.n2110 avss.n2109 0.00916977
R27922 avss.n2109 avss.n2108 0.00916977
R27923 avss.n1894 avss.n1893 0.00916977
R27924 avss.n1893 avss.n1892 0.00916977
R27925 avss.n1678 avss.n1677 0.00916977
R27926 avss.n1677 avss.n1676 0.00916977
R27927 avss.n1462 avss.n1461 0.00916977
R27928 avss.n1461 avss.n1460 0.00916977
R27929 avss.n1246 avss.n1245 0.00916977
R27930 avss.n1245 avss.n1244 0.00916977
R27931 avss.n1030 avss.n1029 0.00916977
R27932 avss.n1029 avss.n1028 0.00916977
R27933 avss.n814 avss.n813 0.00916977
R27934 avss.n813 avss.n812 0.00916977
R27935 avss.n598 avss.n597 0.00916977
R27936 avss.n597 avss.n596 0.00916977
R27937 avss.n273 avss.n272 0.00916977
R27938 avss.n272 avss.n271 0.00916977
R27939 avss.n56 avss.n55 0.00916977
R27940 avss.n55 avss.n54 0.00916977
R27941 avss.n8758 avss.n8750 0.00904545
R27942 avss.n8957 avss.n8955 0.00904545
R27943 avss.n8405 avss.n8397 0.00904545
R27944 avss.n8604 avss.n8602 0.00904545
R27945 avss.n8052 avss.n8044 0.00904545
R27946 avss.n8251 avss.n8249 0.00904545
R27947 avss.n7699 avss.n7691 0.00904545
R27948 avss.n7898 avss.n7896 0.00904545
R27949 avss.n7346 avss.n7338 0.00904545
R27950 avss.n7545 avss.n7543 0.00904545
R27951 avss.n6993 avss.n6985 0.00904545
R27952 avss.n7192 avss.n7190 0.00904545
R27953 avss.n6640 avss.n6632 0.00904545
R27954 avss.n6839 avss.n6837 0.00904545
R27955 avss.n6287 avss.n6279 0.00904545
R27956 avss.n6486 avss.n6484 0.00904545
R27957 avss.n5934 avss.n5926 0.00904545
R27958 avss.n6133 avss.n6131 0.00904545
R27959 avss.n5581 avss.n5573 0.00904545
R27960 avss.n5780 avss.n5778 0.00904545
R27961 avss.n5240 avss.n5232 0.00904545
R27962 avss.n5427 avss.n5425 0.00904545
R27963 avss.n4886 avss.n4878 0.00904545
R27964 avss.n5073 avss.n5071 0.00904545
R27965 avss.n9096 avss.n9089 0.00904545
R27966 avss.n9076 avss.n9069 0.00904545
R27967 avss.n9317 avss.n9310 0.00904545
R27968 avss.n9297 avss.n9290 0.00904545
R27969 avss.n9538 avss.n9531 0.00904545
R27970 avss.n9518 avss.n9511 0.00904545
R27971 avss.n9759 avss.n9752 0.00904545
R27972 avss.n9739 avss.n9732 0.00904545
R27973 avss.n9980 avss.n9973 0.00904545
R27974 avss.n9960 avss.n9953 0.00904545
R27975 avss.n10201 avss.n10194 0.00904545
R27976 avss.n10181 avss.n10174 0.00904545
R27977 avss.n10422 avss.n10415 0.00904545
R27978 avss.n10402 avss.n10395 0.00904545
R27979 avss.n10643 avss.n10636 0.00904545
R27980 avss.n10623 avss.n10616 0.00904545
R27981 avss.n10864 avss.n10857 0.00904545
R27982 avss.n10844 avss.n10837 0.00904545
R27983 avss.n11085 avss.n11078 0.00904545
R27984 avss.n11065 avss.n11058 0.00904545
R27985 avss.n336 avss.n329 0.00904545
R27986 avss.n11286 avss.n11279 0.00904545
R27987 avss.n119 avss.n112 0.00904545
R27988 avss.n11507 avss.n11500 0.00904545
R27989 avss.n3391 avss.n3390 0.00883333
R27990 avss.n3396 avss.n3271 0.00883333
R27991 avss.n3412 avss.n3224 0.00883333
R27992 avss.n3468 avss.n3467 0.00883333
R27993 avss.n5102 avss.n5101 0.00846091
R27994 avss.n5101 avss.n5090 0.00846091
R27995 avss.n4748 avss.n4747 0.00846091
R27996 avss.n4747 avss.n4736 0.00846091
R27997 avss.n11382 avss.n11381 0.00846091
R27998 avss.n11383 avss.n11382 0.00846091
R27999 avss.n11603 avss.n11602 0.00846091
R28000 avss.n11604 avss.n11603 0.00846091
R28001 avss.n8715 avss.n8714 0.00833333
R28002 avss.n8634 avss.n8631 0.00833333
R28003 avss.n8811 avss.n8810 0.00833333
R28004 avss.n8794 avss.n8700 0.00833333
R28005 avss.n8713 avss.n8707 0.00833333
R28006 avss.n8772 avss.n8771 0.00833333
R28007 avss.n8759 avss.n8758 0.00833333
R28008 avss.n8905 avss.n3689 0.00833333
R28009 avss.n3734 avss.n3731 0.00833333
R28010 avss.n8857 avss.n3708 0.00833333
R28011 avss.n8897 avss.n3694 0.00833333
R28012 avss.n8906 avss.n3690 0.00833333
R28013 avss.n8970 avss.n3670 0.00833333
R28014 avss.n8955 avss.n3681 0.00833333
R28015 avss.n8362 avss.n8361 0.00833333
R28016 avss.n8281 avss.n8278 0.00833333
R28017 avss.n8458 avss.n8457 0.00833333
R28018 avss.n8441 avss.n8347 0.00833333
R28019 avss.n8360 avss.n8354 0.00833333
R28020 avss.n8419 avss.n8418 0.00833333
R28021 avss.n8406 avss.n8405 0.00833333
R28022 avss.n8552 avss.n3773 0.00833333
R28023 avss.n3818 avss.n3815 0.00833333
R28024 avss.n8504 avss.n3792 0.00833333
R28025 avss.n8544 avss.n3778 0.00833333
R28026 avss.n8553 avss.n3774 0.00833333
R28027 avss.n8617 avss.n3754 0.00833333
R28028 avss.n8602 avss.n3765 0.00833333
R28029 avss.n8009 avss.n8008 0.00833333
R28030 avss.n7928 avss.n7925 0.00833333
R28031 avss.n8105 avss.n8104 0.00833333
R28032 avss.n8088 avss.n7994 0.00833333
R28033 avss.n8007 avss.n8001 0.00833333
R28034 avss.n8066 avss.n8065 0.00833333
R28035 avss.n8053 avss.n8052 0.00833333
R28036 avss.n8199 avss.n3857 0.00833333
R28037 avss.n3902 avss.n3899 0.00833333
R28038 avss.n8151 avss.n3876 0.00833333
R28039 avss.n8191 avss.n3862 0.00833333
R28040 avss.n8200 avss.n3858 0.00833333
R28041 avss.n8264 avss.n3838 0.00833333
R28042 avss.n8249 avss.n3849 0.00833333
R28043 avss.n7656 avss.n7655 0.00833333
R28044 avss.n7575 avss.n7572 0.00833333
R28045 avss.n7752 avss.n7751 0.00833333
R28046 avss.n7735 avss.n7641 0.00833333
R28047 avss.n7654 avss.n7648 0.00833333
R28048 avss.n7713 avss.n7712 0.00833333
R28049 avss.n7700 avss.n7699 0.00833333
R28050 avss.n7846 avss.n3941 0.00833333
R28051 avss.n3986 avss.n3983 0.00833333
R28052 avss.n7798 avss.n3960 0.00833333
R28053 avss.n7838 avss.n3946 0.00833333
R28054 avss.n7847 avss.n3942 0.00833333
R28055 avss.n7911 avss.n3922 0.00833333
R28056 avss.n7896 avss.n3933 0.00833333
R28057 avss.n7303 avss.n7302 0.00833333
R28058 avss.n7222 avss.n7219 0.00833333
R28059 avss.n7399 avss.n7398 0.00833333
R28060 avss.n7382 avss.n7288 0.00833333
R28061 avss.n7301 avss.n7295 0.00833333
R28062 avss.n7360 avss.n7359 0.00833333
R28063 avss.n7347 avss.n7346 0.00833333
R28064 avss.n7493 avss.n4025 0.00833333
R28065 avss.n4070 avss.n4067 0.00833333
R28066 avss.n7445 avss.n4044 0.00833333
R28067 avss.n7485 avss.n4030 0.00833333
R28068 avss.n7494 avss.n4026 0.00833333
R28069 avss.n7558 avss.n4006 0.00833333
R28070 avss.n7543 avss.n4017 0.00833333
R28071 avss.n6950 avss.n6949 0.00833333
R28072 avss.n6869 avss.n6866 0.00833333
R28073 avss.n7046 avss.n7045 0.00833333
R28074 avss.n7029 avss.n6935 0.00833333
R28075 avss.n6948 avss.n6942 0.00833333
R28076 avss.n7007 avss.n7006 0.00833333
R28077 avss.n6994 avss.n6993 0.00833333
R28078 avss.n7140 avss.n4109 0.00833333
R28079 avss.n4154 avss.n4151 0.00833333
R28080 avss.n7092 avss.n4128 0.00833333
R28081 avss.n7132 avss.n4114 0.00833333
R28082 avss.n7141 avss.n4110 0.00833333
R28083 avss.n7205 avss.n4090 0.00833333
R28084 avss.n7190 avss.n4101 0.00833333
R28085 avss.n6597 avss.n6596 0.00833333
R28086 avss.n6516 avss.n6513 0.00833333
R28087 avss.n6693 avss.n6692 0.00833333
R28088 avss.n6676 avss.n6582 0.00833333
R28089 avss.n6595 avss.n6589 0.00833333
R28090 avss.n6654 avss.n6653 0.00833333
R28091 avss.n6641 avss.n6640 0.00833333
R28092 avss.n6787 avss.n4193 0.00833333
R28093 avss.n4238 avss.n4235 0.00833333
R28094 avss.n6739 avss.n4212 0.00833333
R28095 avss.n6779 avss.n4198 0.00833333
R28096 avss.n6788 avss.n4194 0.00833333
R28097 avss.n6852 avss.n4174 0.00833333
R28098 avss.n6837 avss.n4185 0.00833333
R28099 avss.n6244 avss.n6243 0.00833333
R28100 avss.n6163 avss.n6160 0.00833333
R28101 avss.n6340 avss.n6339 0.00833333
R28102 avss.n6323 avss.n6229 0.00833333
R28103 avss.n6242 avss.n6236 0.00833333
R28104 avss.n6301 avss.n6300 0.00833333
R28105 avss.n6288 avss.n6287 0.00833333
R28106 avss.n6434 avss.n4277 0.00833333
R28107 avss.n4322 avss.n4319 0.00833333
R28108 avss.n6386 avss.n4296 0.00833333
R28109 avss.n6426 avss.n4282 0.00833333
R28110 avss.n6435 avss.n4278 0.00833333
R28111 avss.n6499 avss.n4258 0.00833333
R28112 avss.n6484 avss.n4269 0.00833333
R28113 avss.n5891 avss.n5890 0.00833333
R28114 avss.n5810 avss.n5807 0.00833333
R28115 avss.n5987 avss.n5986 0.00833333
R28116 avss.n5970 avss.n5876 0.00833333
R28117 avss.n5889 avss.n5883 0.00833333
R28118 avss.n5948 avss.n5947 0.00833333
R28119 avss.n5935 avss.n5934 0.00833333
R28120 avss.n6081 avss.n4361 0.00833333
R28121 avss.n4406 avss.n4403 0.00833333
R28122 avss.n6033 avss.n4380 0.00833333
R28123 avss.n6073 avss.n4366 0.00833333
R28124 avss.n6082 avss.n4362 0.00833333
R28125 avss.n6146 avss.n4342 0.00833333
R28126 avss.n6131 avss.n4353 0.00833333
R28127 avss.n5538 avss.n5537 0.00833333
R28128 avss.n5457 avss.n5454 0.00833333
R28129 avss.n5634 avss.n5633 0.00833333
R28130 avss.n5617 avss.n5523 0.00833333
R28131 avss.n5536 avss.n5530 0.00833333
R28132 avss.n5595 avss.n5594 0.00833333
R28133 avss.n5582 avss.n5581 0.00833333
R28134 avss.n5728 avss.n4445 0.00833333
R28135 avss.n4490 avss.n4487 0.00833333
R28136 avss.n5680 avss.n4464 0.00833333
R28137 avss.n5720 avss.n4450 0.00833333
R28138 avss.n5729 avss.n4446 0.00833333
R28139 avss.n5793 avss.n4426 0.00833333
R28140 avss.n5778 avss.n4437 0.00833333
R28141 avss.n5192 avss.n5191 0.00833333
R28142 avss.n5109 avss.n5105 0.00833333
R28143 avss.n5289 avss.n5288 0.00833333
R28144 avss.n5272 avss.n5177 0.00833333
R28145 avss.n5190 avss.n5184 0.00833333
R28146 avss.n5208 avss.n5206 0.00833333
R28147 avss.n5241 avss.n5240 0.00833333
R28148 avss.n5375 avss.n4529 0.00833333
R28149 avss.n4574 avss.n4571 0.00833333
R28150 avss.n5327 avss.n4548 0.00833333
R28151 avss.n5367 avss.n4534 0.00833333
R28152 avss.n5376 avss.n4530 0.00833333
R28153 avss.n5440 avss.n4510 0.00833333
R28154 avss.n5425 avss.n4521 0.00833333
R28155 avss.n4838 avss.n4837 0.00833333
R28156 avss.n4755 avss.n4751 0.00833333
R28157 avss.n4935 avss.n4934 0.00833333
R28158 avss.n4918 avss.n4823 0.00833333
R28159 avss.n4836 avss.n4830 0.00833333
R28160 avss.n4854 avss.n4852 0.00833333
R28161 avss.n4887 avss.n4886 0.00833333
R28162 avss.n5021 avss.n4613 0.00833333
R28163 avss.n4658 avss.n4655 0.00833333
R28164 avss.n4973 avss.n4632 0.00833333
R28165 avss.n5013 avss.n4618 0.00833333
R28166 avss.n5022 avss.n4614 0.00833333
R28167 avss.n5086 avss.n4594 0.00833333
R28168 avss.n5071 avss.n4605 0.00833333
R28169 avss.n9184 avss.n9183 0.00833333
R28170 avss.n2421 avss.n2413 0.00833333
R28171 avss.n2460 avss.n2459 0.00833333
R28172 avss.n9133 avss.n9132 0.00833333
R28173 avss.n9139 avss.n9138 0.00833333
R28174 avss.n9117 avss.n9116 0.00833333
R28175 avss.n9089 avss.n9088 0.00833333
R28176 avss.n8983 avss.n8982 0.00833333
R28177 avss.n2568 avss.n2560 0.00833333
R28178 avss.n2517 avss.n2516 0.00833333
R28179 avss.n9022 avss.n9021 0.00833333
R28180 avss.n9028 avss.n9027 0.00833333
R28181 avss.n9006 avss.n9005 0.00833333
R28182 avss.n9069 avss.n9068 0.00833333
R28183 avss.n9405 avss.n9404 0.00833333
R28184 avss.n2205 avss.n2197 0.00833333
R28185 avss.n2244 avss.n2243 0.00833333
R28186 avss.n9354 avss.n9353 0.00833333
R28187 avss.n9360 avss.n9359 0.00833333
R28188 avss.n9338 avss.n9337 0.00833333
R28189 avss.n9310 avss.n9309 0.00833333
R28190 avss.n9204 avss.n9203 0.00833333
R28191 avss.n2352 avss.n2344 0.00833333
R28192 avss.n2301 avss.n2300 0.00833333
R28193 avss.n9243 avss.n9242 0.00833333
R28194 avss.n9249 avss.n9248 0.00833333
R28195 avss.n9227 avss.n9226 0.00833333
R28196 avss.n9290 avss.n9289 0.00833333
R28197 avss.n9626 avss.n9625 0.00833333
R28198 avss.n1989 avss.n1981 0.00833333
R28199 avss.n2028 avss.n2027 0.00833333
R28200 avss.n9575 avss.n9574 0.00833333
R28201 avss.n9581 avss.n9580 0.00833333
R28202 avss.n9559 avss.n9558 0.00833333
R28203 avss.n9531 avss.n9530 0.00833333
R28204 avss.n9425 avss.n9424 0.00833333
R28205 avss.n2136 avss.n2128 0.00833333
R28206 avss.n2085 avss.n2084 0.00833333
R28207 avss.n9464 avss.n9463 0.00833333
R28208 avss.n9470 avss.n9469 0.00833333
R28209 avss.n9448 avss.n9447 0.00833333
R28210 avss.n9511 avss.n9510 0.00833333
R28211 avss.n9847 avss.n9846 0.00833333
R28212 avss.n1773 avss.n1765 0.00833333
R28213 avss.n1812 avss.n1811 0.00833333
R28214 avss.n9796 avss.n9795 0.00833333
R28215 avss.n9802 avss.n9801 0.00833333
R28216 avss.n9780 avss.n9779 0.00833333
R28217 avss.n9752 avss.n9751 0.00833333
R28218 avss.n9646 avss.n9645 0.00833333
R28219 avss.n1920 avss.n1912 0.00833333
R28220 avss.n1869 avss.n1868 0.00833333
R28221 avss.n9685 avss.n9684 0.00833333
R28222 avss.n9691 avss.n9690 0.00833333
R28223 avss.n9669 avss.n9668 0.00833333
R28224 avss.n9732 avss.n9731 0.00833333
R28225 avss.n10068 avss.n10067 0.00833333
R28226 avss.n1557 avss.n1549 0.00833333
R28227 avss.n1596 avss.n1595 0.00833333
R28228 avss.n10017 avss.n10016 0.00833333
R28229 avss.n10023 avss.n10022 0.00833333
R28230 avss.n10001 avss.n10000 0.00833333
R28231 avss.n9973 avss.n9972 0.00833333
R28232 avss.n9867 avss.n9866 0.00833333
R28233 avss.n1704 avss.n1696 0.00833333
R28234 avss.n1653 avss.n1652 0.00833333
R28235 avss.n9906 avss.n9905 0.00833333
R28236 avss.n9912 avss.n9911 0.00833333
R28237 avss.n9890 avss.n9889 0.00833333
R28238 avss.n9953 avss.n9952 0.00833333
R28239 avss.n10289 avss.n10288 0.00833333
R28240 avss.n1341 avss.n1333 0.00833333
R28241 avss.n1380 avss.n1379 0.00833333
R28242 avss.n10238 avss.n10237 0.00833333
R28243 avss.n10244 avss.n10243 0.00833333
R28244 avss.n10222 avss.n10221 0.00833333
R28245 avss.n10194 avss.n10193 0.00833333
R28246 avss.n10088 avss.n10087 0.00833333
R28247 avss.n1488 avss.n1480 0.00833333
R28248 avss.n1437 avss.n1436 0.00833333
R28249 avss.n10127 avss.n10126 0.00833333
R28250 avss.n10133 avss.n10132 0.00833333
R28251 avss.n10111 avss.n10110 0.00833333
R28252 avss.n10174 avss.n10173 0.00833333
R28253 avss.n10510 avss.n10509 0.00833333
R28254 avss.n1125 avss.n1117 0.00833333
R28255 avss.n1164 avss.n1163 0.00833333
R28256 avss.n10459 avss.n10458 0.00833333
R28257 avss.n10465 avss.n10464 0.00833333
R28258 avss.n10443 avss.n10442 0.00833333
R28259 avss.n10415 avss.n10414 0.00833333
R28260 avss.n10309 avss.n10308 0.00833333
R28261 avss.n1272 avss.n1264 0.00833333
R28262 avss.n1221 avss.n1220 0.00833333
R28263 avss.n10348 avss.n10347 0.00833333
R28264 avss.n10354 avss.n10353 0.00833333
R28265 avss.n10332 avss.n10331 0.00833333
R28266 avss.n10395 avss.n10394 0.00833333
R28267 avss.n10731 avss.n10730 0.00833333
R28268 avss.n909 avss.n901 0.00833333
R28269 avss.n948 avss.n947 0.00833333
R28270 avss.n10680 avss.n10679 0.00833333
R28271 avss.n10686 avss.n10685 0.00833333
R28272 avss.n10664 avss.n10663 0.00833333
R28273 avss.n10636 avss.n10635 0.00833333
R28274 avss.n10530 avss.n10529 0.00833333
R28275 avss.n1056 avss.n1048 0.00833333
R28276 avss.n1005 avss.n1004 0.00833333
R28277 avss.n10569 avss.n10568 0.00833333
R28278 avss.n10575 avss.n10574 0.00833333
R28279 avss.n10553 avss.n10552 0.00833333
R28280 avss.n10616 avss.n10615 0.00833333
R28281 avss.n10952 avss.n10951 0.00833333
R28282 avss.n693 avss.n685 0.00833333
R28283 avss.n732 avss.n731 0.00833333
R28284 avss.n10901 avss.n10900 0.00833333
R28285 avss.n10907 avss.n10906 0.00833333
R28286 avss.n10885 avss.n10884 0.00833333
R28287 avss.n10857 avss.n10856 0.00833333
R28288 avss.n10751 avss.n10750 0.00833333
R28289 avss.n840 avss.n832 0.00833333
R28290 avss.n789 avss.n788 0.00833333
R28291 avss.n10790 avss.n10789 0.00833333
R28292 avss.n10796 avss.n10795 0.00833333
R28293 avss.n10774 avss.n10773 0.00833333
R28294 avss.n10837 avss.n10836 0.00833333
R28295 avss.n11173 avss.n11172 0.00833333
R28296 avss.n477 avss.n469 0.00833333
R28297 avss.n516 avss.n515 0.00833333
R28298 avss.n11122 avss.n11121 0.00833333
R28299 avss.n11128 avss.n11127 0.00833333
R28300 avss.n11106 avss.n11105 0.00833333
R28301 avss.n11078 avss.n11077 0.00833333
R28302 avss.n10972 avss.n10971 0.00833333
R28303 avss.n624 avss.n616 0.00833333
R28304 avss.n573 avss.n572 0.00833333
R28305 avss.n11011 avss.n11010 0.00833333
R28306 avss.n11017 avss.n11016 0.00833333
R28307 avss.n10995 avss.n10994 0.00833333
R28308 avss.n11058 avss.n11057 0.00833333
R28309 avss.n349 avss.n348 0.00833333
R28310 avss.n11396 avss.n11388 0.00833333
R28311 avss.n11345 avss.n11344 0.00833333
R28312 avss.n389 avss.n388 0.00833333
R28313 avss.n395 avss.n394 0.00833333
R28314 avss.n373 avss.n372 0.00833333
R28315 avss.n329 avss.n328 0.00833333
R28316 avss.n11193 avss.n11192 0.00833333
R28317 avss.n299 avss.n291 0.00833333
R28318 avss.n248 avss.n247 0.00833333
R28319 avss.n11232 avss.n11231 0.00833333
R28320 avss.n11238 avss.n11237 0.00833333
R28321 avss.n11216 avss.n11215 0.00833333
R28322 avss.n11279 avss.n11278 0.00833333
R28323 avss.n132 avss.n131 0.00833333
R28324 avss.n11617 avss.n11609 0.00833333
R28325 avss.n11566 avss.n11565 0.00833333
R28326 avss.n172 avss.n171 0.00833333
R28327 avss.n178 avss.n177 0.00833333
R28328 avss.n156 avss.n155 0.00833333
R28329 avss.n112 avss.n111 0.00833333
R28330 avss.n11414 avss.n11413 0.00833333
R28331 avss.n82 avss.n74 0.00833333
R28332 avss.n31 avss.n30 0.00833333
R28333 avss.n11453 avss.n11452 0.00833333
R28334 avss.n11459 avss.n11458 0.00833333
R28335 avss.n11437 avss.n11436 0.00833333
R28336 avss.n11500 avss.n11499 0.00833333
R28337 avss.n3350 avss.n3349 0.0083125
R28338 avss avss.n11634 0.00771154
R28339 avss.n3261 avss 0.00766301
R28340 avss.n3259 avss 0.00766301
R28341 avss.n3527 avss 0.00766301
R28342 avss.n3523 avss 0.00766301
R28343 avss.n8674 avss.n8670 0.00762121
R28344 avss.n8766 avss.n8765 0.00762121
R28345 avss.n3712 avss.n3706 0.00762121
R28346 avss.n8948 avss.n3680 0.00762121
R28347 avss.n8321 avss.n8317 0.00762121
R28348 avss.n8413 avss.n8412 0.00762121
R28349 avss.n3796 avss.n3790 0.00762121
R28350 avss.n8595 avss.n3764 0.00762121
R28351 avss.n7968 avss.n7964 0.00762121
R28352 avss.n8060 avss.n8059 0.00762121
R28353 avss.n3880 avss.n3874 0.00762121
R28354 avss.n8242 avss.n3848 0.00762121
R28355 avss.n7615 avss.n7611 0.00762121
R28356 avss.n7707 avss.n7706 0.00762121
R28357 avss.n3964 avss.n3958 0.00762121
R28358 avss.n7889 avss.n3932 0.00762121
R28359 avss.n7262 avss.n7258 0.00762121
R28360 avss.n7354 avss.n7353 0.00762121
R28361 avss.n4048 avss.n4042 0.00762121
R28362 avss.n7536 avss.n4016 0.00762121
R28363 avss.n6909 avss.n6905 0.00762121
R28364 avss.n7001 avss.n7000 0.00762121
R28365 avss.n4132 avss.n4126 0.00762121
R28366 avss.n7183 avss.n4100 0.00762121
R28367 avss.n6556 avss.n6552 0.00762121
R28368 avss.n6648 avss.n6647 0.00762121
R28369 avss.n4216 avss.n4210 0.00762121
R28370 avss.n6830 avss.n4184 0.00762121
R28371 avss.n6203 avss.n6199 0.00762121
R28372 avss.n6295 avss.n6294 0.00762121
R28373 avss.n4300 avss.n4294 0.00762121
R28374 avss.n6477 avss.n4268 0.00762121
R28375 avss.n5850 avss.n5846 0.00762121
R28376 avss.n5942 avss.n5941 0.00762121
R28377 avss.n4384 avss.n4378 0.00762121
R28378 avss.n6124 avss.n4352 0.00762121
R28379 avss.n5497 avss.n5493 0.00762121
R28380 avss.n5589 avss.n5588 0.00762121
R28381 avss.n4468 avss.n4462 0.00762121
R28382 avss.n5771 avss.n4436 0.00762121
R28383 avss.n5151 avss.n5147 0.00762121
R28384 avss.n5229 avss.n5211 0.00762121
R28385 avss.n4552 avss.n4546 0.00762121
R28386 avss.n5418 avss.n4520 0.00762121
R28387 avss.n4797 avss.n4793 0.00762121
R28388 avss.n4875 avss.n4857 0.00762121
R28389 avss.n4636 avss.n4630 0.00762121
R28390 avss.n5064 avss.n4604 0.00762121
R28391 avss.n2448 avss.n2447 0.00762121
R28392 avss.n9103 avss.n9102 0.00762121
R28393 avss.n2505 avss.n2504 0.00762121
R28394 avss.n8991 avss.n8990 0.00762121
R28395 avss.n2232 avss.n2231 0.00762121
R28396 avss.n9324 avss.n9323 0.00762121
R28397 avss.n2289 avss.n2288 0.00762121
R28398 avss.n9212 avss.n9211 0.00762121
R28399 avss.n2016 avss.n2015 0.00762121
R28400 avss.n9545 avss.n9544 0.00762121
R28401 avss.n2073 avss.n2072 0.00762121
R28402 avss.n9433 avss.n9432 0.00762121
R28403 avss.n1800 avss.n1799 0.00762121
R28404 avss.n9766 avss.n9765 0.00762121
R28405 avss.n1857 avss.n1856 0.00762121
R28406 avss.n9654 avss.n9653 0.00762121
R28407 avss.n1584 avss.n1583 0.00762121
R28408 avss.n9987 avss.n9986 0.00762121
R28409 avss.n1641 avss.n1640 0.00762121
R28410 avss.n9875 avss.n9874 0.00762121
R28411 avss.n1368 avss.n1367 0.00762121
R28412 avss.n10208 avss.n10207 0.00762121
R28413 avss.n1425 avss.n1424 0.00762121
R28414 avss.n10096 avss.n10095 0.00762121
R28415 avss.n1152 avss.n1151 0.00762121
R28416 avss.n10429 avss.n10428 0.00762121
R28417 avss.n1209 avss.n1208 0.00762121
R28418 avss.n10317 avss.n10316 0.00762121
R28419 avss.n936 avss.n935 0.00762121
R28420 avss.n10650 avss.n10649 0.00762121
R28421 avss.n993 avss.n992 0.00762121
R28422 avss.n10538 avss.n10537 0.00762121
R28423 avss.n720 avss.n719 0.00762121
R28424 avss.n10871 avss.n10870 0.00762121
R28425 avss.n777 avss.n776 0.00762121
R28426 avss.n10759 avss.n10758 0.00762121
R28427 avss.n504 avss.n503 0.00762121
R28428 avss.n11092 avss.n11091 0.00762121
R28429 avss.n561 avss.n560 0.00762121
R28430 avss.n10980 avss.n10979 0.00762121
R28431 avss.n11333 avss.n11332 0.00762121
R28432 avss.n358 avss.n357 0.00762121
R28433 avss.n236 avss.n235 0.00762121
R28434 avss.n11201 avss.n11200 0.00762121
R28435 avss.n11554 avss.n11553 0.00762121
R28436 avss.n141 avss.n140 0.00762121
R28437 avss.n19 avss.n18 0.00762121
R28438 avss.n11422 avss.n11421 0.00762121
R28439 avss.n3737 avss.n3729 0.00747678
R28440 avss.n3821 avss.n3813 0.00747678
R28441 avss.n3905 avss.n3897 0.00747678
R28442 avss.n3989 avss.n3981 0.00747678
R28443 avss.n4073 avss.n4065 0.00747678
R28444 avss.n4157 avss.n4149 0.00747678
R28445 avss.n4241 avss.n4233 0.00747678
R28446 avss.n4325 avss.n4317 0.00747678
R28447 avss.n4409 avss.n4401 0.00747678
R28448 avss.n4493 avss.n4485 0.00747678
R28449 avss.n4577 avss.n4569 0.00747678
R28450 avss.n4661 avss.n4653 0.00747678
R28451 avss.n2562 avss.n2561 0.00747678
R28452 avss.n2346 avss.n2345 0.00747678
R28453 avss.n2130 avss.n2129 0.00747678
R28454 avss.n1914 avss.n1913 0.00747678
R28455 avss.n1698 avss.n1697 0.00747678
R28456 avss.n1482 avss.n1481 0.00747678
R28457 avss.n1266 avss.n1265 0.00747678
R28458 avss.n1050 avss.n1049 0.00747678
R28459 avss.n834 avss.n833 0.00747678
R28460 avss.n618 avss.n617 0.00747678
R28461 avss.n293 avss.n292 0.00747678
R28462 avss.n76 avss.n75 0.00747678
R28463 avss.n8637 avss.n8629 0.00747597
R28464 avss.n8284 avss.n8276 0.00747597
R28465 avss.n7931 avss.n7923 0.00747597
R28466 avss.n7578 avss.n7570 0.00747597
R28467 avss.n7225 avss.n7217 0.00747597
R28468 avss.n6872 avss.n6864 0.00747597
R28469 avss.n6519 avss.n6511 0.00747597
R28470 avss.n6166 avss.n6158 0.00747597
R28471 avss.n5813 avss.n5805 0.00747597
R28472 avss.n5460 avss.n5452 0.00747597
R28473 avss.n5112 avss.n5103 0.00747597
R28474 avss.n4758 avss.n4749 0.00747597
R28475 avss.n2415 avss.n2414 0.00747597
R28476 avss.n2199 avss.n2198 0.00747597
R28477 avss.n1983 avss.n1982 0.00747597
R28478 avss.n1767 avss.n1766 0.00747597
R28479 avss.n1551 avss.n1550 0.00747597
R28480 avss.n1335 avss.n1334 0.00747597
R28481 avss.n1119 avss.n1118 0.00747597
R28482 avss.n903 avss.n902 0.00747597
R28483 avss.n687 avss.n686 0.00747597
R28484 avss.n471 avss.n470 0.00747597
R28485 avss.n11390 avss.n11389 0.00747597
R28486 avss.n11611 avss.n11610 0.00747597
R28487 avss.n8780 avss.n8779 0.00690909
R28488 avss.n8643 avss.n8642 0.00690909
R28489 avss.n8819 avss.n8651 0.00690909
R28490 avss.n8816 avss.n8654 0.00690909
R28491 avss.n8709 avss.n8701 0.00690909
R28492 avss.n8778 avss.n8719 0.00690909
R28493 avss.n8731 avss.n8724 0.00690909
R28494 avss.n8740 avss.n8739 0.00690909
R28495 avss.n8927 avss.n8926 0.00690909
R28496 avss.n3743 avss.n3742 0.00690909
R28497 avss.n8854 avss.n3719 0.00690909
R28498 avss.n8865 avss.n3715 0.00690909
R28499 avss.n8912 avss.n8911 0.00690909
R28500 avss.n8925 avss.n3688 0.00690909
R28501 avss.n8937 avss.n3676 0.00690909
R28502 avss.n8939 avss.n3675 0.00690909
R28503 avss.n8427 avss.n8426 0.00690909
R28504 avss.n8290 avss.n8289 0.00690909
R28505 avss.n8466 avss.n8298 0.00690909
R28506 avss.n8463 avss.n8301 0.00690909
R28507 avss.n8356 avss.n8348 0.00690909
R28508 avss.n8425 avss.n8366 0.00690909
R28509 avss.n8378 avss.n8371 0.00690909
R28510 avss.n8387 avss.n8386 0.00690909
R28511 avss.n8574 avss.n8573 0.00690909
R28512 avss.n3827 avss.n3826 0.00690909
R28513 avss.n8501 avss.n3803 0.00690909
R28514 avss.n8512 avss.n3799 0.00690909
R28515 avss.n8559 avss.n8558 0.00690909
R28516 avss.n8572 avss.n3772 0.00690909
R28517 avss.n8584 avss.n3760 0.00690909
R28518 avss.n8586 avss.n3759 0.00690909
R28519 avss.n8074 avss.n8073 0.00690909
R28520 avss.n7937 avss.n7936 0.00690909
R28521 avss.n8113 avss.n7945 0.00690909
R28522 avss.n8110 avss.n7948 0.00690909
R28523 avss.n8003 avss.n7995 0.00690909
R28524 avss.n8072 avss.n8013 0.00690909
R28525 avss.n8025 avss.n8018 0.00690909
R28526 avss.n8034 avss.n8033 0.00690909
R28527 avss.n8221 avss.n8220 0.00690909
R28528 avss.n3911 avss.n3910 0.00690909
R28529 avss.n8148 avss.n3887 0.00690909
R28530 avss.n8159 avss.n3883 0.00690909
R28531 avss.n8206 avss.n8205 0.00690909
R28532 avss.n8219 avss.n3856 0.00690909
R28533 avss.n8231 avss.n3844 0.00690909
R28534 avss.n8233 avss.n3843 0.00690909
R28535 avss.n7721 avss.n7720 0.00690909
R28536 avss.n7584 avss.n7583 0.00690909
R28537 avss.n7760 avss.n7592 0.00690909
R28538 avss.n7757 avss.n7595 0.00690909
R28539 avss.n7650 avss.n7642 0.00690909
R28540 avss.n7719 avss.n7660 0.00690909
R28541 avss.n7672 avss.n7665 0.00690909
R28542 avss.n7681 avss.n7680 0.00690909
R28543 avss.n7868 avss.n7867 0.00690909
R28544 avss.n3995 avss.n3994 0.00690909
R28545 avss.n7795 avss.n3971 0.00690909
R28546 avss.n7806 avss.n3967 0.00690909
R28547 avss.n7853 avss.n7852 0.00690909
R28548 avss.n7866 avss.n3940 0.00690909
R28549 avss.n7878 avss.n3928 0.00690909
R28550 avss.n7880 avss.n3927 0.00690909
R28551 avss.n7368 avss.n7367 0.00690909
R28552 avss.n7231 avss.n7230 0.00690909
R28553 avss.n7407 avss.n7239 0.00690909
R28554 avss.n7404 avss.n7242 0.00690909
R28555 avss.n7297 avss.n7289 0.00690909
R28556 avss.n7366 avss.n7307 0.00690909
R28557 avss.n7319 avss.n7312 0.00690909
R28558 avss.n7328 avss.n7327 0.00690909
R28559 avss.n7515 avss.n7514 0.00690909
R28560 avss.n4079 avss.n4078 0.00690909
R28561 avss.n7442 avss.n4055 0.00690909
R28562 avss.n7453 avss.n4051 0.00690909
R28563 avss.n7500 avss.n7499 0.00690909
R28564 avss.n7513 avss.n4024 0.00690909
R28565 avss.n7525 avss.n4012 0.00690909
R28566 avss.n7527 avss.n4011 0.00690909
R28567 avss.n7015 avss.n7014 0.00690909
R28568 avss.n6878 avss.n6877 0.00690909
R28569 avss.n7054 avss.n6886 0.00690909
R28570 avss.n7051 avss.n6889 0.00690909
R28571 avss.n6944 avss.n6936 0.00690909
R28572 avss.n7013 avss.n6954 0.00690909
R28573 avss.n6966 avss.n6959 0.00690909
R28574 avss.n6975 avss.n6974 0.00690909
R28575 avss.n7162 avss.n7161 0.00690909
R28576 avss.n4163 avss.n4162 0.00690909
R28577 avss.n7089 avss.n4139 0.00690909
R28578 avss.n7100 avss.n4135 0.00690909
R28579 avss.n7147 avss.n7146 0.00690909
R28580 avss.n7160 avss.n4108 0.00690909
R28581 avss.n7172 avss.n4096 0.00690909
R28582 avss.n7174 avss.n4095 0.00690909
R28583 avss.n6662 avss.n6661 0.00690909
R28584 avss.n6525 avss.n6524 0.00690909
R28585 avss.n6701 avss.n6533 0.00690909
R28586 avss.n6698 avss.n6536 0.00690909
R28587 avss.n6591 avss.n6583 0.00690909
R28588 avss.n6660 avss.n6601 0.00690909
R28589 avss.n6613 avss.n6606 0.00690909
R28590 avss.n6622 avss.n6621 0.00690909
R28591 avss.n6809 avss.n6808 0.00690909
R28592 avss.n4247 avss.n4246 0.00690909
R28593 avss.n6736 avss.n4223 0.00690909
R28594 avss.n6747 avss.n4219 0.00690909
R28595 avss.n6794 avss.n6793 0.00690909
R28596 avss.n6807 avss.n4192 0.00690909
R28597 avss.n6819 avss.n4180 0.00690909
R28598 avss.n6821 avss.n4179 0.00690909
R28599 avss.n6309 avss.n6308 0.00690909
R28600 avss.n6172 avss.n6171 0.00690909
R28601 avss.n6348 avss.n6180 0.00690909
R28602 avss.n6345 avss.n6183 0.00690909
R28603 avss.n6238 avss.n6230 0.00690909
R28604 avss.n6307 avss.n6248 0.00690909
R28605 avss.n6260 avss.n6253 0.00690909
R28606 avss.n6269 avss.n6268 0.00690909
R28607 avss.n6456 avss.n6455 0.00690909
R28608 avss.n4331 avss.n4330 0.00690909
R28609 avss.n6383 avss.n4307 0.00690909
R28610 avss.n6394 avss.n4303 0.00690909
R28611 avss.n6441 avss.n6440 0.00690909
R28612 avss.n6454 avss.n4276 0.00690909
R28613 avss.n6466 avss.n4264 0.00690909
R28614 avss.n6468 avss.n4263 0.00690909
R28615 avss.n5956 avss.n5955 0.00690909
R28616 avss.n5819 avss.n5818 0.00690909
R28617 avss.n5995 avss.n5827 0.00690909
R28618 avss.n5992 avss.n5830 0.00690909
R28619 avss.n5885 avss.n5877 0.00690909
R28620 avss.n5954 avss.n5895 0.00690909
R28621 avss.n5907 avss.n5900 0.00690909
R28622 avss.n5916 avss.n5915 0.00690909
R28623 avss.n6103 avss.n6102 0.00690909
R28624 avss.n4415 avss.n4414 0.00690909
R28625 avss.n6030 avss.n4391 0.00690909
R28626 avss.n6041 avss.n4387 0.00690909
R28627 avss.n6088 avss.n6087 0.00690909
R28628 avss.n6101 avss.n4360 0.00690909
R28629 avss.n6113 avss.n4348 0.00690909
R28630 avss.n6115 avss.n4347 0.00690909
R28631 avss.n5603 avss.n5602 0.00690909
R28632 avss.n5466 avss.n5465 0.00690909
R28633 avss.n5642 avss.n5474 0.00690909
R28634 avss.n5639 avss.n5477 0.00690909
R28635 avss.n5532 avss.n5524 0.00690909
R28636 avss.n5601 avss.n5542 0.00690909
R28637 avss.n5554 avss.n5547 0.00690909
R28638 avss.n5563 avss.n5562 0.00690909
R28639 avss.n5750 avss.n5749 0.00690909
R28640 avss.n4499 avss.n4498 0.00690909
R28641 avss.n5677 avss.n4475 0.00690909
R28642 avss.n5688 avss.n4471 0.00690909
R28643 avss.n5735 avss.n5734 0.00690909
R28644 avss.n5748 avss.n4444 0.00690909
R28645 avss.n5760 avss.n4432 0.00690909
R28646 avss.n5762 avss.n4431 0.00690909
R28647 avss.n5258 avss.n5257 0.00690909
R28648 avss.n5119 avss.n5118 0.00690909
R28649 avss.n5297 avss.n5095 0.00690909
R28650 avss.n5139 avss.n5138 0.00690909
R28651 avss.n5186 avss.n5178 0.00690909
R28652 avss.n5256 avss.n5196 0.00690909
R28653 avss.n5214 avss.n5201 0.00690909
R28654 avss.n5223 avss.n5222 0.00690909
R28655 avss.n5397 avss.n5396 0.00690909
R28656 avss.n4583 avss.n4582 0.00690909
R28657 avss.n5324 avss.n4559 0.00690909
R28658 avss.n5335 avss.n4555 0.00690909
R28659 avss.n5382 avss.n5381 0.00690909
R28660 avss.n5395 avss.n4528 0.00690909
R28661 avss.n5407 avss.n4516 0.00690909
R28662 avss.n5409 avss.n4515 0.00690909
R28663 avss.n4904 avss.n4903 0.00690909
R28664 avss.n4765 avss.n4764 0.00690909
R28665 avss.n4943 avss.n4741 0.00690909
R28666 avss.n4785 avss.n4784 0.00690909
R28667 avss.n4832 avss.n4824 0.00690909
R28668 avss.n4902 avss.n4842 0.00690909
R28669 avss.n4860 avss.n4847 0.00690909
R28670 avss.n4869 avss.n4868 0.00690909
R28671 avss.n5043 avss.n5042 0.00690909
R28672 avss.n4667 avss.n4666 0.00690909
R28673 avss.n4970 avss.n4643 0.00690909
R28674 avss.n4981 avss.n4639 0.00690909
R28675 avss.n5028 avss.n5027 0.00690909
R28676 avss.n5041 avss.n4612 0.00690909
R28677 avss.n5053 avss.n4600 0.00690909
R28678 avss.n5055 avss.n4599 0.00690909
R28679 avss.n9188 avss.n9187 0.00690909
R28680 avss.n2412 avss.n2411 0.00690909
R28681 avss.n2478 avss.n2477 0.00690909
R28682 avss.n2466 avss.n2465 0.00690909
R28683 avss.n9135 avss.n9134 0.00690909
R28684 avss.n9154 avss.n9153 0.00690909
R28685 avss.n9169 avss.n9159 0.00690909
R28686 avss.n9172 avss.n9171 0.00690909
R28687 avss.n8987 avss.n8986 0.00690909
R28688 avss.n2559 avss.n2558 0.00690909
R28689 avss.n2535 avss.n2534 0.00690909
R28690 avss.n2523 avss.n2522 0.00690909
R28691 avss.n9024 avss.n9023 0.00690909
R28692 avss.n9043 avss.n9042 0.00690909
R28693 avss.n9058 avss.n9048 0.00690909
R28694 avss.n9061 avss.n9060 0.00690909
R28695 avss.n9409 avss.n9408 0.00690909
R28696 avss.n2196 avss.n2195 0.00690909
R28697 avss.n2262 avss.n2261 0.00690909
R28698 avss.n2250 avss.n2249 0.00690909
R28699 avss.n9356 avss.n9355 0.00690909
R28700 avss.n9375 avss.n9374 0.00690909
R28701 avss.n9390 avss.n9380 0.00690909
R28702 avss.n9393 avss.n9392 0.00690909
R28703 avss.n9208 avss.n9207 0.00690909
R28704 avss.n2343 avss.n2342 0.00690909
R28705 avss.n2319 avss.n2318 0.00690909
R28706 avss.n2307 avss.n2306 0.00690909
R28707 avss.n9245 avss.n9244 0.00690909
R28708 avss.n9264 avss.n9263 0.00690909
R28709 avss.n9279 avss.n9269 0.00690909
R28710 avss.n9282 avss.n9281 0.00690909
R28711 avss.n9630 avss.n9629 0.00690909
R28712 avss.n1980 avss.n1979 0.00690909
R28713 avss.n2046 avss.n2045 0.00690909
R28714 avss.n2034 avss.n2033 0.00690909
R28715 avss.n9577 avss.n9576 0.00690909
R28716 avss.n9596 avss.n9595 0.00690909
R28717 avss.n9611 avss.n9601 0.00690909
R28718 avss.n9614 avss.n9613 0.00690909
R28719 avss.n9429 avss.n9428 0.00690909
R28720 avss.n2127 avss.n2126 0.00690909
R28721 avss.n2103 avss.n2102 0.00690909
R28722 avss.n2091 avss.n2090 0.00690909
R28723 avss.n9466 avss.n9465 0.00690909
R28724 avss.n9485 avss.n9484 0.00690909
R28725 avss.n9500 avss.n9490 0.00690909
R28726 avss.n9503 avss.n9502 0.00690909
R28727 avss.n9851 avss.n9850 0.00690909
R28728 avss.n1764 avss.n1763 0.00690909
R28729 avss.n1830 avss.n1829 0.00690909
R28730 avss.n1818 avss.n1817 0.00690909
R28731 avss.n9798 avss.n9797 0.00690909
R28732 avss.n9817 avss.n9816 0.00690909
R28733 avss.n9832 avss.n9822 0.00690909
R28734 avss.n9835 avss.n9834 0.00690909
R28735 avss.n9650 avss.n9649 0.00690909
R28736 avss.n1911 avss.n1910 0.00690909
R28737 avss.n1887 avss.n1886 0.00690909
R28738 avss.n1875 avss.n1874 0.00690909
R28739 avss.n9687 avss.n9686 0.00690909
R28740 avss.n9706 avss.n9705 0.00690909
R28741 avss.n9721 avss.n9711 0.00690909
R28742 avss.n9724 avss.n9723 0.00690909
R28743 avss.n10072 avss.n10071 0.00690909
R28744 avss.n1548 avss.n1547 0.00690909
R28745 avss.n1614 avss.n1613 0.00690909
R28746 avss.n1602 avss.n1601 0.00690909
R28747 avss.n10019 avss.n10018 0.00690909
R28748 avss.n10038 avss.n10037 0.00690909
R28749 avss.n10053 avss.n10043 0.00690909
R28750 avss.n10056 avss.n10055 0.00690909
R28751 avss.n9871 avss.n9870 0.00690909
R28752 avss.n1695 avss.n1694 0.00690909
R28753 avss.n1671 avss.n1670 0.00690909
R28754 avss.n1659 avss.n1658 0.00690909
R28755 avss.n9908 avss.n9907 0.00690909
R28756 avss.n9927 avss.n9926 0.00690909
R28757 avss.n9942 avss.n9932 0.00690909
R28758 avss.n9945 avss.n9944 0.00690909
R28759 avss.n10293 avss.n10292 0.00690909
R28760 avss.n1332 avss.n1331 0.00690909
R28761 avss.n1398 avss.n1397 0.00690909
R28762 avss.n1386 avss.n1385 0.00690909
R28763 avss.n10240 avss.n10239 0.00690909
R28764 avss.n10259 avss.n10258 0.00690909
R28765 avss.n10274 avss.n10264 0.00690909
R28766 avss.n10277 avss.n10276 0.00690909
R28767 avss.n10092 avss.n10091 0.00690909
R28768 avss.n1479 avss.n1478 0.00690909
R28769 avss.n1455 avss.n1454 0.00690909
R28770 avss.n1443 avss.n1442 0.00690909
R28771 avss.n10129 avss.n10128 0.00690909
R28772 avss.n10148 avss.n10147 0.00690909
R28773 avss.n10163 avss.n10153 0.00690909
R28774 avss.n10166 avss.n10165 0.00690909
R28775 avss.n10514 avss.n10513 0.00690909
R28776 avss.n1116 avss.n1115 0.00690909
R28777 avss.n1182 avss.n1181 0.00690909
R28778 avss.n1170 avss.n1169 0.00690909
R28779 avss.n10461 avss.n10460 0.00690909
R28780 avss.n10480 avss.n10479 0.00690909
R28781 avss.n10495 avss.n10485 0.00690909
R28782 avss.n10498 avss.n10497 0.00690909
R28783 avss.n10313 avss.n10312 0.00690909
R28784 avss.n1263 avss.n1262 0.00690909
R28785 avss.n1239 avss.n1238 0.00690909
R28786 avss.n1227 avss.n1226 0.00690909
R28787 avss.n10350 avss.n10349 0.00690909
R28788 avss.n10369 avss.n10368 0.00690909
R28789 avss.n10384 avss.n10374 0.00690909
R28790 avss.n10387 avss.n10386 0.00690909
R28791 avss.n10735 avss.n10734 0.00690909
R28792 avss.n900 avss.n899 0.00690909
R28793 avss.n966 avss.n965 0.00690909
R28794 avss.n954 avss.n953 0.00690909
R28795 avss.n10682 avss.n10681 0.00690909
R28796 avss.n10701 avss.n10700 0.00690909
R28797 avss.n10716 avss.n10706 0.00690909
R28798 avss.n10719 avss.n10718 0.00690909
R28799 avss.n10534 avss.n10533 0.00690909
R28800 avss.n1047 avss.n1046 0.00690909
R28801 avss.n1023 avss.n1022 0.00690909
R28802 avss.n1011 avss.n1010 0.00690909
R28803 avss.n10571 avss.n10570 0.00690909
R28804 avss.n10590 avss.n10589 0.00690909
R28805 avss.n10605 avss.n10595 0.00690909
R28806 avss.n10608 avss.n10607 0.00690909
R28807 avss.n10956 avss.n10955 0.00690909
R28808 avss.n684 avss.n683 0.00690909
R28809 avss.n750 avss.n749 0.00690909
R28810 avss.n738 avss.n737 0.00690909
R28811 avss.n10903 avss.n10902 0.00690909
R28812 avss.n10922 avss.n10921 0.00690909
R28813 avss.n10937 avss.n10927 0.00690909
R28814 avss.n10940 avss.n10939 0.00690909
R28815 avss.n10755 avss.n10754 0.00690909
R28816 avss.n831 avss.n830 0.00690909
R28817 avss.n807 avss.n806 0.00690909
R28818 avss.n795 avss.n794 0.00690909
R28819 avss.n10792 avss.n10791 0.00690909
R28820 avss.n10811 avss.n10810 0.00690909
R28821 avss.n10826 avss.n10816 0.00690909
R28822 avss.n10829 avss.n10828 0.00690909
R28823 avss.n11177 avss.n11176 0.00690909
R28824 avss.n468 avss.n467 0.00690909
R28825 avss.n534 avss.n533 0.00690909
R28826 avss.n522 avss.n521 0.00690909
R28827 avss.n11124 avss.n11123 0.00690909
R28828 avss.n11143 avss.n11142 0.00690909
R28829 avss.n11158 avss.n11148 0.00690909
R28830 avss.n11161 avss.n11160 0.00690909
R28831 avss.n10976 avss.n10975 0.00690909
R28832 avss.n615 avss.n614 0.00690909
R28833 avss.n591 avss.n590 0.00690909
R28834 avss.n579 avss.n578 0.00690909
R28835 avss.n11013 avss.n11012 0.00690909
R28836 avss.n11032 avss.n11031 0.00690909
R28837 avss.n11047 avss.n11037 0.00690909
R28838 avss.n11050 avss.n11049 0.00690909
R28839 avss.n353 avss.n352 0.00690909
R28840 avss.n11387 avss.n11386 0.00690909
R28841 avss.n11363 avss.n11362 0.00690909
R28842 avss.n11351 avss.n11350 0.00690909
R28843 avss.n391 avss.n390 0.00690909
R28844 avss.n410 avss.n409 0.00690909
R28845 avss.n425 avss.n415 0.00690909
R28846 avss.n428 avss.n427 0.00690909
R28847 avss.n11197 avss.n11196 0.00690909
R28848 avss.n290 avss.n289 0.00690909
R28849 avss.n266 avss.n265 0.00690909
R28850 avss.n254 avss.n253 0.00690909
R28851 avss.n11234 avss.n11233 0.00690909
R28852 avss.n11253 avss.n11252 0.00690909
R28853 avss.n11268 avss.n11258 0.00690909
R28854 avss.n11271 avss.n11270 0.00690909
R28855 avss.n136 avss.n135 0.00690909
R28856 avss.n11608 avss.n11607 0.00690909
R28857 avss.n11584 avss.n11583 0.00690909
R28858 avss.n11572 avss.n11571 0.00690909
R28859 avss.n174 avss.n173 0.00690909
R28860 avss.n193 avss.n192 0.00690909
R28861 avss.n208 avss.n198 0.00690909
R28862 avss.n211 avss.n210 0.00690909
R28863 avss.n11418 avss.n11417 0.00690909
R28864 avss.n73 avss.n72 0.00690909
R28865 avss.n49 avss.n48 0.00690909
R28866 avss.n37 avss.n36 0.00690909
R28867 avss.n11455 avss.n11454 0.00690909
R28868 avss.n11474 avss.n11473 0.00690909
R28869 avss.n11489 avss.n11479 0.00690909
R28870 avss.n11492 avss.n11491 0.00690909
R28871 avss.n3461 avss.n3197 0.00675
R28872 avss.n3514 avss.n3174 0.00675
R28873 avss.n8639 avss.n8638 0.00619697
R28874 avss.n8820 avss.n8819 0.00619697
R28875 avss.n8804 avss.n8671 0.00619697
R28876 avss.n8797 avss.n8684 0.00619697
R28877 avss.n8733 avss.n8724 0.00619697
R28878 avss.n3739 avss.n3738 0.00619697
R28879 avss.n8854 avss.n3718 0.00619697
R28880 avss.n8879 avss.n3704 0.00619697
R28881 avss.n8902 avss.n3698 0.00619697
R28882 avss.n8933 avss.n3676 0.00619697
R28883 avss.n8286 avss.n8285 0.00619697
R28884 avss.n8467 avss.n8466 0.00619697
R28885 avss.n8451 avss.n8318 0.00619697
R28886 avss.n8444 avss.n8331 0.00619697
R28887 avss.n8380 avss.n8371 0.00619697
R28888 avss.n3823 avss.n3822 0.00619697
R28889 avss.n8501 avss.n3802 0.00619697
R28890 avss.n8526 avss.n3788 0.00619697
R28891 avss.n8549 avss.n3782 0.00619697
R28892 avss.n8580 avss.n3760 0.00619697
R28893 avss.n7933 avss.n7932 0.00619697
R28894 avss.n8114 avss.n8113 0.00619697
R28895 avss.n8098 avss.n7965 0.00619697
R28896 avss.n8091 avss.n7978 0.00619697
R28897 avss.n8027 avss.n8018 0.00619697
R28898 avss.n3907 avss.n3906 0.00619697
R28899 avss.n8148 avss.n3886 0.00619697
R28900 avss.n8173 avss.n3872 0.00619697
R28901 avss.n8196 avss.n3866 0.00619697
R28902 avss.n8227 avss.n3844 0.00619697
R28903 avss.n7580 avss.n7579 0.00619697
R28904 avss.n7761 avss.n7760 0.00619697
R28905 avss.n7745 avss.n7612 0.00619697
R28906 avss.n7738 avss.n7625 0.00619697
R28907 avss.n7674 avss.n7665 0.00619697
R28908 avss.n3991 avss.n3990 0.00619697
R28909 avss.n7795 avss.n3970 0.00619697
R28910 avss.n7820 avss.n3956 0.00619697
R28911 avss.n7843 avss.n3950 0.00619697
R28912 avss.n7874 avss.n3928 0.00619697
R28913 avss.n7227 avss.n7226 0.00619697
R28914 avss.n7408 avss.n7407 0.00619697
R28915 avss.n7392 avss.n7259 0.00619697
R28916 avss.n7385 avss.n7272 0.00619697
R28917 avss.n7321 avss.n7312 0.00619697
R28918 avss.n4075 avss.n4074 0.00619697
R28919 avss.n7442 avss.n4054 0.00619697
R28920 avss.n7467 avss.n4040 0.00619697
R28921 avss.n7490 avss.n4034 0.00619697
R28922 avss.n7521 avss.n4012 0.00619697
R28923 avss.n6874 avss.n6873 0.00619697
R28924 avss.n7055 avss.n7054 0.00619697
R28925 avss.n7039 avss.n6906 0.00619697
R28926 avss.n7032 avss.n6919 0.00619697
R28927 avss.n6968 avss.n6959 0.00619697
R28928 avss.n4159 avss.n4158 0.00619697
R28929 avss.n7089 avss.n4138 0.00619697
R28930 avss.n7114 avss.n4124 0.00619697
R28931 avss.n7137 avss.n4118 0.00619697
R28932 avss.n7168 avss.n4096 0.00619697
R28933 avss.n6521 avss.n6520 0.00619697
R28934 avss.n6702 avss.n6701 0.00619697
R28935 avss.n6686 avss.n6553 0.00619697
R28936 avss.n6679 avss.n6566 0.00619697
R28937 avss.n6615 avss.n6606 0.00619697
R28938 avss.n4243 avss.n4242 0.00619697
R28939 avss.n6736 avss.n4222 0.00619697
R28940 avss.n6761 avss.n4208 0.00619697
R28941 avss.n6784 avss.n4202 0.00619697
R28942 avss.n6815 avss.n4180 0.00619697
R28943 avss.n6168 avss.n6167 0.00619697
R28944 avss.n6349 avss.n6348 0.00619697
R28945 avss.n6333 avss.n6200 0.00619697
R28946 avss.n6326 avss.n6213 0.00619697
R28947 avss.n6262 avss.n6253 0.00619697
R28948 avss.n4327 avss.n4326 0.00619697
R28949 avss.n6383 avss.n4306 0.00619697
R28950 avss.n6408 avss.n4292 0.00619697
R28951 avss.n6431 avss.n4286 0.00619697
R28952 avss.n6462 avss.n4264 0.00619697
R28953 avss.n5815 avss.n5814 0.00619697
R28954 avss.n5996 avss.n5995 0.00619697
R28955 avss.n5980 avss.n5847 0.00619697
R28956 avss.n5973 avss.n5860 0.00619697
R28957 avss.n5909 avss.n5900 0.00619697
R28958 avss.n4411 avss.n4410 0.00619697
R28959 avss.n6030 avss.n4390 0.00619697
R28960 avss.n6055 avss.n4376 0.00619697
R28961 avss.n6078 avss.n4370 0.00619697
R28962 avss.n6109 avss.n4348 0.00619697
R28963 avss.n5462 avss.n5461 0.00619697
R28964 avss.n5643 avss.n5642 0.00619697
R28965 avss.n5627 avss.n5494 0.00619697
R28966 avss.n5620 avss.n5507 0.00619697
R28967 avss.n5556 avss.n5547 0.00619697
R28968 avss.n4495 avss.n4494 0.00619697
R28969 avss.n5677 avss.n4474 0.00619697
R28970 avss.n5702 avss.n4460 0.00619697
R28971 avss.n5725 avss.n4454 0.00619697
R28972 avss.n5756 avss.n4432 0.00619697
R28973 avss.n5114 avss.n5113 0.00619697
R28974 avss.n5297 avss.n5094 0.00619697
R28975 avss.n5282 avss.n5148 0.00619697
R28976 avss.n5275 avss.n5161 0.00619697
R28977 avss.n5216 avss.n5201 0.00619697
R28978 avss.n4579 avss.n4578 0.00619697
R28979 avss.n5324 avss.n4558 0.00619697
R28980 avss.n5349 avss.n4544 0.00619697
R28981 avss.n5372 avss.n4538 0.00619697
R28982 avss.n5403 avss.n4516 0.00619697
R28983 avss.n4760 avss.n4759 0.00619697
R28984 avss.n4943 avss.n4740 0.00619697
R28985 avss.n4928 avss.n4794 0.00619697
R28986 avss.n4921 avss.n4807 0.00619697
R28987 avss.n4862 avss.n4847 0.00619697
R28988 avss.n4663 avss.n4662 0.00619697
R28989 avss.n4970 avss.n4642 0.00619697
R28990 avss.n4995 avss.n4628 0.00619697
R28991 avss.n5018 avss.n4622 0.00619697
R28992 avss.n5049 avss.n4600 0.00619697
R28993 avss.n2424 avss.n2423 0.00619697
R28994 avss.n2479 avss.n2478 0.00619697
R28995 avss.n2444 avss.n2443 0.00619697
R28996 avss.n9121 avss.n9120 0.00619697
R28997 avss.n9159 avss.n9158 0.00619697
R28998 avss.n2571 avss.n2570 0.00619697
R28999 avss.n2536 avss.n2535 0.00619697
R29000 avss.n2501 avss.n2500 0.00619697
R29001 avss.n9010 avss.n9009 0.00619697
R29002 avss.n9048 avss.n9047 0.00619697
R29003 avss.n2208 avss.n2207 0.00619697
R29004 avss.n2263 avss.n2262 0.00619697
R29005 avss.n2228 avss.n2227 0.00619697
R29006 avss.n9342 avss.n9341 0.00619697
R29007 avss.n9380 avss.n9379 0.00619697
R29008 avss.n2355 avss.n2354 0.00619697
R29009 avss.n2320 avss.n2319 0.00619697
R29010 avss.n2285 avss.n2284 0.00619697
R29011 avss.n9231 avss.n9230 0.00619697
R29012 avss.n9269 avss.n9268 0.00619697
R29013 avss.n1992 avss.n1991 0.00619697
R29014 avss.n2047 avss.n2046 0.00619697
R29015 avss.n2012 avss.n2011 0.00619697
R29016 avss.n9563 avss.n9562 0.00619697
R29017 avss.n9601 avss.n9600 0.00619697
R29018 avss.n2139 avss.n2138 0.00619697
R29019 avss.n2104 avss.n2103 0.00619697
R29020 avss.n2069 avss.n2068 0.00619697
R29021 avss.n9452 avss.n9451 0.00619697
R29022 avss.n9490 avss.n9489 0.00619697
R29023 avss.n1776 avss.n1775 0.00619697
R29024 avss.n1831 avss.n1830 0.00619697
R29025 avss.n1796 avss.n1795 0.00619697
R29026 avss.n9784 avss.n9783 0.00619697
R29027 avss.n9822 avss.n9821 0.00619697
R29028 avss.n1923 avss.n1922 0.00619697
R29029 avss.n1888 avss.n1887 0.00619697
R29030 avss.n1853 avss.n1852 0.00619697
R29031 avss.n9673 avss.n9672 0.00619697
R29032 avss.n9711 avss.n9710 0.00619697
R29033 avss.n1560 avss.n1559 0.00619697
R29034 avss.n1615 avss.n1614 0.00619697
R29035 avss.n1580 avss.n1579 0.00619697
R29036 avss.n10005 avss.n10004 0.00619697
R29037 avss.n10043 avss.n10042 0.00619697
R29038 avss.n1707 avss.n1706 0.00619697
R29039 avss.n1672 avss.n1671 0.00619697
R29040 avss.n1637 avss.n1636 0.00619697
R29041 avss.n9894 avss.n9893 0.00619697
R29042 avss.n9932 avss.n9931 0.00619697
R29043 avss.n1344 avss.n1343 0.00619697
R29044 avss.n1399 avss.n1398 0.00619697
R29045 avss.n1364 avss.n1363 0.00619697
R29046 avss.n10226 avss.n10225 0.00619697
R29047 avss.n10264 avss.n10263 0.00619697
R29048 avss.n1491 avss.n1490 0.00619697
R29049 avss.n1456 avss.n1455 0.00619697
R29050 avss.n1421 avss.n1420 0.00619697
R29051 avss.n10115 avss.n10114 0.00619697
R29052 avss.n10153 avss.n10152 0.00619697
R29053 avss.n1128 avss.n1127 0.00619697
R29054 avss.n1183 avss.n1182 0.00619697
R29055 avss.n1148 avss.n1147 0.00619697
R29056 avss.n10447 avss.n10446 0.00619697
R29057 avss.n10485 avss.n10484 0.00619697
R29058 avss.n1275 avss.n1274 0.00619697
R29059 avss.n1240 avss.n1239 0.00619697
R29060 avss.n1205 avss.n1204 0.00619697
R29061 avss.n10336 avss.n10335 0.00619697
R29062 avss.n10374 avss.n10373 0.00619697
R29063 avss.n912 avss.n911 0.00619697
R29064 avss.n967 avss.n966 0.00619697
R29065 avss.n932 avss.n931 0.00619697
R29066 avss.n10668 avss.n10667 0.00619697
R29067 avss.n10706 avss.n10705 0.00619697
R29068 avss.n1059 avss.n1058 0.00619697
R29069 avss.n1024 avss.n1023 0.00619697
R29070 avss.n989 avss.n988 0.00619697
R29071 avss.n10557 avss.n10556 0.00619697
R29072 avss.n10595 avss.n10594 0.00619697
R29073 avss.n696 avss.n695 0.00619697
R29074 avss.n751 avss.n750 0.00619697
R29075 avss.n716 avss.n715 0.00619697
R29076 avss.n10889 avss.n10888 0.00619697
R29077 avss.n10927 avss.n10926 0.00619697
R29078 avss.n843 avss.n842 0.00619697
R29079 avss.n808 avss.n807 0.00619697
R29080 avss.n773 avss.n772 0.00619697
R29081 avss.n10778 avss.n10777 0.00619697
R29082 avss.n10816 avss.n10815 0.00619697
R29083 avss.n480 avss.n479 0.00619697
R29084 avss.n535 avss.n534 0.00619697
R29085 avss.n500 avss.n499 0.00619697
R29086 avss.n11110 avss.n11109 0.00619697
R29087 avss.n11148 avss.n11147 0.00619697
R29088 avss.n627 avss.n626 0.00619697
R29089 avss.n592 avss.n591 0.00619697
R29090 avss.n557 avss.n556 0.00619697
R29091 avss.n10999 avss.n10998 0.00619697
R29092 avss.n11037 avss.n11036 0.00619697
R29093 avss.n11399 avss.n11398 0.00619697
R29094 avss.n11364 avss.n11363 0.00619697
R29095 avss.n11329 avss.n11328 0.00619697
R29096 avss.n377 avss.n376 0.00619697
R29097 avss.n415 avss.n414 0.00619697
R29098 avss.n302 avss.n301 0.00619697
R29099 avss.n267 avss.n266 0.00619697
R29100 avss.n232 avss.n231 0.00619697
R29101 avss.n11220 avss.n11219 0.00619697
R29102 avss.n11258 avss.n11257 0.00619697
R29103 avss.n11620 avss.n11619 0.00619697
R29104 avss.n11585 avss.n11584 0.00619697
R29105 avss.n11550 avss.n11549 0.00619697
R29106 avss.n160 avss.n159 0.00619697
R29107 avss.n198 avss.n197 0.00619697
R29108 avss.n85 avss.n84 0.00619697
R29109 avss.n50 avss.n49 0.00619697
R29110 avss.n15 avss.n14 0.00619697
R29111 avss.n11441 avss.n11440 0.00619697
R29112 avss.n11479 avss.n11478 0.00619697
R29113 avss.n8703 avss.n8682 0.00618182
R29114 avss.n8689 avss.n8679 0.00618182
R29115 avss.n8637 avss.n8636 0.00618182
R29116 avss.n8756 avss.n8755 0.00618182
R29117 avss.n3737 avss.n3736 0.00618182
R29118 avss.n8882 avss.n3700 0.00618182
R29119 avss.n8900 avss.n8899 0.00618182
R29120 avss.n8956 avss.n8954 0.00618182
R29121 avss.n8350 avss.n8329 0.00618182
R29122 avss.n8336 avss.n8326 0.00618182
R29123 avss.n8284 avss.n8283 0.00618182
R29124 avss.n8403 avss.n8402 0.00618182
R29125 avss.n3821 avss.n3820 0.00618182
R29126 avss.n8529 avss.n3784 0.00618182
R29127 avss.n8547 avss.n8546 0.00618182
R29128 avss.n8603 avss.n8601 0.00618182
R29129 avss.n7997 avss.n7976 0.00618182
R29130 avss.n7983 avss.n7973 0.00618182
R29131 avss.n7931 avss.n7930 0.00618182
R29132 avss.n8050 avss.n8049 0.00618182
R29133 avss.n3905 avss.n3904 0.00618182
R29134 avss.n8176 avss.n3868 0.00618182
R29135 avss.n8194 avss.n8193 0.00618182
R29136 avss.n8250 avss.n8248 0.00618182
R29137 avss.n7644 avss.n7623 0.00618182
R29138 avss.n7630 avss.n7620 0.00618182
R29139 avss.n7578 avss.n7577 0.00618182
R29140 avss.n7697 avss.n7696 0.00618182
R29141 avss.n3989 avss.n3988 0.00618182
R29142 avss.n7823 avss.n3952 0.00618182
R29143 avss.n7841 avss.n7840 0.00618182
R29144 avss.n7897 avss.n7895 0.00618182
R29145 avss.n7291 avss.n7270 0.00618182
R29146 avss.n7277 avss.n7267 0.00618182
R29147 avss.n7225 avss.n7224 0.00618182
R29148 avss.n7344 avss.n7343 0.00618182
R29149 avss.n4073 avss.n4072 0.00618182
R29150 avss.n7470 avss.n4036 0.00618182
R29151 avss.n7488 avss.n7487 0.00618182
R29152 avss.n7544 avss.n7542 0.00618182
R29153 avss.n6938 avss.n6917 0.00618182
R29154 avss.n6924 avss.n6914 0.00618182
R29155 avss.n6872 avss.n6871 0.00618182
R29156 avss.n6991 avss.n6990 0.00618182
R29157 avss.n4157 avss.n4156 0.00618182
R29158 avss.n7117 avss.n4120 0.00618182
R29159 avss.n7135 avss.n7134 0.00618182
R29160 avss.n7191 avss.n7189 0.00618182
R29161 avss.n6585 avss.n6564 0.00618182
R29162 avss.n6571 avss.n6561 0.00618182
R29163 avss.n6519 avss.n6518 0.00618182
R29164 avss.n6638 avss.n6637 0.00618182
R29165 avss.n4241 avss.n4240 0.00618182
R29166 avss.n6764 avss.n4204 0.00618182
R29167 avss.n6782 avss.n6781 0.00618182
R29168 avss.n6838 avss.n6836 0.00618182
R29169 avss.n6232 avss.n6211 0.00618182
R29170 avss.n6218 avss.n6208 0.00618182
R29171 avss.n6166 avss.n6165 0.00618182
R29172 avss.n6285 avss.n6284 0.00618182
R29173 avss.n4325 avss.n4324 0.00618182
R29174 avss.n6411 avss.n4288 0.00618182
R29175 avss.n6429 avss.n6428 0.00618182
R29176 avss.n6485 avss.n6483 0.00618182
R29177 avss.n5879 avss.n5858 0.00618182
R29178 avss.n5865 avss.n5855 0.00618182
R29179 avss.n5813 avss.n5812 0.00618182
R29180 avss.n5932 avss.n5931 0.00618182
R29181 avss.n4409 avss.n4408 0.00618182
R29182 avss.n6058 avss.n4372 0.00618182
R29183 avss.n6076 avss.n6075 0.00618182
R29184 avss.n6132 avss.n6130 0.00618182
R29185 avss.n5526 avss.n5505 0.00618182
R29186 avss.n5512 avss.n5502 0.00618182
R29187 avss.n5460 avss.n5459 0.00618182
R29188 avss.n5579 avss.n5578 0.00618182
R29189 avss.n4493 avss.n4492 0.00618182
R29190 avss.n5705 avss.n4456 0.00618182
R29191 avss.n5723 avss.n5722 0.00618182
R29192 avss.n5779 avss.n5777 0.00618182
R29193 avss.n5180 avss.n5159 0.00618182
R29194 avss.n5166 avss.n5156 0.00618182
R29195 avss.n5112 avss.n5111 0.00618182
R29196 avss.n5238 avss.n5237 0.00618182
R29197 avss.n4577 avss.n4576 0.00618182
R29198 avss.n5352 avss.n4540 0.00618182
R29199 avss.n5370 avss.n5369 0.00618182
R29200 avss.n5426 avss.n5424 0.00618182
R29201 avss.n4826 avss.n4805 0.00618182
R29202 avss.n4812 avss.n4802 0.00618182
R29203 avss.n4758 avss.n4757 0.00618182
R29204 avss.n4884 avss.n4883 0.00618182
R29205 avss.n4661 avss.n4660 0.00618182
R29206 avss.n4998 avss.n4624 0.00618182
R29207 avss.n5016 avss.n5015 0.00618182
R29208 avss.n5072 avss.n5070 0.00618182
R29209 avss.n9125 avss.n9124 0.00618182
R29210 avss.n2441 avss.n2440 0.00618182
R29211 avss.n2416 avss.n2415 0.00618182
R29212 avss.n9095 avss.n9094 0.00618182
R29213 avss.n2563 avss.n2562 0.00618182
R29214 avss.n2498 avss.n2497 0.00618182
R29215 avss.n9014 avss.n9013 0.00618182
R29216 avss.n9075 avss.n9074 0.00618182
R29217 avss.n9346 avss.n9345 0.00618182
R29218 avss.n2225 avss.n2224 0.00618182
R29219 avss.n2200 avss.n2199 0.00618182
R29220 avss.n9316 avss.n9315 0.00618182
R29221 avss.n2347 avss.n2346 0.00618182
R29222 avss.n2282 avss.n2281 0.00618182
R29223 avss.n9235 avss.n9234 0.00618182
R29224 avss.n9296 avss.n9295 0.00618182
R29225 avss.n9567 avss.n9566 0.00618182
R29226 avss.n2009 avss.n2008 0.00618182
R29227 avss.n1984 avss.n1983 0.00618182
R29228 avss.n9537 avss.n9536 0.00618182
R29229 avss.n2131 avss.n2130 0.00618182
R29230 avss.n2066 avss.n2065 0.00618182
R29231 avss.n9456 avss.n9455 0.00618182
R29232 avss.n9517 avss.n9516 0.00618182
R29233 avss.n9788 avss.n9787 0.00618182
R29234 avss.n1793 avss.n1792 0.00618182
R29235 avss.n1768 avss.n1767 0.00618182
R29236 avss.n9758 avss.n9757 0.00618182
R29237 avss.n1915 avss.n1914 0.00618182
R29238 avss.n1850 avss.n1849 0.00618182
R29239 avss.n9677 avss.n9676 0.00618182
R29240 avss.n9738 avss.n9737 0.00618182
R29241 avss.n10009 avss.n10008 0.00618182
R29242 avss.n1577 avss.n1576 0.00618182
R29243 avss.n1552 avss.n1551 0.00618182
R29244 avss.n9979 avss.n9978 0.00618182
R29245 avss.n1699 avss.n1698 0.00618182
R29246 avss.n1634 avss.n1633 0.00618182
R29247 avss.n9898 avss.n9897 0.00618182
R29248 avss.n9959 avss.n9958 0.00618182
R29249 avss.n10230 avss.n10229 0.00618182
R29250 avss.n1361 avss.n1360 0.00618182
R29251 avss.n1336 avss.n1335 0.00618182
R29252 avss.n10200 avss.n10199 0.00618182
R29253 avss.n1483 avss.n1482 0.00618182
R29254 avss.n1418 avss.n1417 0.00618182
R29255 avss.n10119 avss.n10118 0.00618182
R29256 avss.n10180 avss.n10179 0.00618182
R29257 avss.n10451 avss.n10450 0.00618182
R29258 avss.n1145 avss.n1144 0.00618182
R29259 avss.n1120 avss.n1119 0.00618182
R29260 avss.n10421 avss.n10420 0.00618182
R29261 avss.n1267 avss.n1266 0.00618182
R29262 avss.n1202 avss.n1201 0.00618182
R29263 avss.n10340 avss.n10339 0.00618182
R29264 avss.n10401 avss.n10400 0.00618182
R29265 avss.n10672 avss.n10671 0.00618182
R29266 avss.n929 avss.n928 0.00618182
R29267 avss.n904 avss.n903 0.00618182
R29268 avss.n10642 avss.n10641 0.00618182
R29269 avss.n1051 avss.n1050 0.00618182
R29270 avss.n986 avss.n985 0.00618182
R29271 avss.n10561 avss.n10560 0.00618182
R29272 avss.n10622 avss.n10621 0.00618182
R29273 avss.n10893 avss.n10892 0.00618182
R29274 avss.n713 avss.n712 0.00618182
R29275 avss.n688 avss.n687 0.00618182
R29276 avss.n10863 avss.n10862 0.00618182
R29277 avss.n835 avss.n834 0.00618182
R29278 avss.n770 avss.n769 0.00618182
R29279 avss.n10782 avss.n10781 0.00618182
R29280 avss.n10843 avss.n10842 0.00618182
R29281 avss.n11114 avss.n11113 0.00618182
R29282 avss.n497 avss.n496 0.00618182
R29283 avss.n472 avss.n471 0.00618182
R29284 avss.n11084 avss.n11083 0.00618182
R29285 avss.n619 avss.n618 0.00618182
R29286 avss.n554 avss.n553 0.00618182
R29287 avss.n11003 avss.n11002 0.00618182
R29288 avss.n11064 avss.n11063 0.00618182
R29289 avss.n381 avss.n380 0.00618182
R29290 avss.n11326 avss.n11325 0.00618182
R29291 avss.n11391 avss.n11390 0.00618182
R29292 avss.n335 avss.n334 0.00618182
R29293 avss.n294 avss.n293 0.00618182
R29294 avss.n229 avss.n228 0.00618182
R29295 avss.n11224 avss.n11223 0.00618182
R29296 avss.n11285 avss.n11284 0.00618182
R29297 avss.n164 avss.n163 0.00618182
R29298 avss.n11547 avss.n11546 0.00618182
R29299 avss.n11612 avss.n11611 0.00618182
R29300 avss.n118 avss.n117 0.00618182
R29301 avss.n77 avss.n76 0.00618182
R29302 avss.n12 avss.n11 0.00618182
R29303 avss.n11445 avss.n11444 0.00618182
R29304 avss.n11506 avss.n11505 0.00618182
R29305 avss.n8754 avss.n8753 0.0060117
R29306 avss.n8401 avss.n8400 0.0060117
R29307 avss.n8048 avss.n8047 0.0060117
R29308 avss.n7695 avss.n7694 0.0060117
R29309 avss.n7342 avss.n7341 0.0060117
R29310 avss.n6989 avss.n6988 0.0060117
R29311 avss.n6636 avss.n6635 0.0060117
R29312 avss.n6283 avss.n6282 0.0060117
R29313 avss.n5930 avss.n5929 0.0060117
R29314 avss.n5577 avss.n5576 0.0060117
R29315 avss.n5236 avss.n5235 0.0060117
R29316 avss.n4882 avss.n4881 0.0060117
R29317 avss.n9098 avss.n9097 0.0060117
R29318 avss.n9319 avss.n9318 0.0060117
R29319 avss.n9540 avss.n9539 0.0060117
R29320 avss.n9761 avss.n9760 0.0060117
R29321 avss.n9982 avss.n9981 0.0060117
R29322 avss.n10203 avss.n10202 0.0060117
R29323 avss.n10424 avss.n10423 0.0060117
R29324 avss.n10645 avss.n10644 0.0060117
R29325 avss.n10866 avss.n10865 0.0060117
R29326 avss.n11087 avss.n11086 0.0060117
R29327 avss.n338 avss.n337 0.0060117
R29328 avss.n121 avss.n120 0.0060117
R29329 avss.n8959 avss.n8958 0.00551524
R29330 avss.n8606 avss.n8605 0.00551524
R29331 avss.n8253 avss.n8252 0.00551524
R29332 avss.n7900 avss.n7899 0.00551524
R29333 avss.n7547 avss.n7546 0.00551524
R29334 avss.n7194 avss.n7193 0.00551524
R29335 avss.n6841 avss.n6840 0.00551524
R29336 avss.n6488 avss.n6487 0.00551524
R29337 avss.n6135 avss.n6134 0.00551524
R29338 avss.n5782 avss.n5781 0.00551524
R29339 avss.n5429 avss.n5428 0.00551524
R29340 avss.n5075 avss.n5074 0.00551524
R29341 avss.n9078 avss.n9077 0.00551524
R29342 avss.n9299 avss.n9298 0.00551524
R29343 avss.n9520 avss.n9519 0.00551524
R29344 avss.n9741 avss.n9740 0.00551524
R29345 avss.n9962 avss.n9961 0.00551524
R29346 avss.n10183 avss.n10182 0.00551524
R29347 avss.n10404 avss.n10403 0.00551524
R29348 avss.n10625 avss.n10624 0.00551524
R29349 avss.n10846 avss.n10845 0.00551524
R29350 avss.n11067 avss.n11066 0.00551524
R29351 avss.n11288 avss.n11287 0.00551524
R29352 avss.n11509 avss.n11508 0.00551524
R29353 avss.n8692 avss.n8687 0.00548485
R29354 avss.n8691 avss.n8690 0.00548485
R29355 avss.n8691 avss.n8686 0.00548485
R29356 avss.n8886 avss.n8885 0.00548485
R29357 avss.n8884 avss.n3701 0.00548485
R29358 avss.n8892 avss.n3701 0.00548485
R29359 avss.n8339 avss.n8334 0.00548485
R29360 avss.n8338 avss.n8337 0.00548485
R29361 avss.n8338 avss.n8333 0.00548485
R29362 avss.n8533 avss.n8532 0.00548485
R29363 avss.n8531 avss.n3785 0.00548485
R29364 avss.n8539 avss.n3785 0.00548485
R29365 avss.n7986 avss.n7981 0.00548485
R29366 avss.n7985 avss.n7984 0.00548485
R29367 avss.n7985 avss.n7980 0.00548485
R29368 avss.n8180 avss.n8179 0.00548485
R29369 avss.n8178 avss.n3869 0.00548485
R29370 avss.n8186 avss.n3869 0.00548485
R29371 avss.n7633 avss.n7628 0.00548485
R29372 avss.n7632 avss.n7631 0.00548485
R29373 avss.n7632 avss.n7627 0.00548485
R29374 avss.n7827 avss.n7826 0.00548485
R29375 avss.n7825 avss.n3953 0.00548485
R29376 avss.n7833 avss.n3953 0.00548485
R29377 avss.n7280 avss.n7275 0.00548485
R29378 avss.n7279 avss.n7278 0.00548485
R29379 avss.n7279 avss.n7274 0.00548485
R29380 avss.n7474 avss.n7473 0.00548485
R29381 avss.n7472 avss.n4037 0.00548485
R29382 avss.n7480 avss.n4037 0.00548485
R29383 avss.n6927 avss.n6922 0.00548485
R29384 avss.n6926 avss.n6925 0.00548485
R29385 avss.n6926 avss.n6921 0.00548485
R29386 avss.n7121 avss.n7120 0.00548485
R29387 avss.n7119 avss.n4121 0.00548485
R29388 avss.n7127 avss.n4121 0.00548485
R29389 avss.n6574 avss.n6569 0.00548485
R29390 avss.n6573 avss.n6572 0.00548485
R29391 avss.n6573 avss.n6568 0.00548485
R29392 avss.n6768 avss.n6767 0.00548485
R29393 avss.n6766 avss.n4205 0.00548485
R29394 avss.n6774 avss.n4205 0.00548485
R29395 avss.n6221 avss.n6216 0.00548485
R29396 avss.n6220 avss.n6219 0.00548485
R29397 avss.n6220 avss.n6215 0.00548485
R29398 avss.n6415 avss.n6414 0.00548485
R29399 avss.n6413 avss.n4289 0.00548485
R29400 avss.n6421 avss.n4289 0.00548485
R29401 avss.n5868 avss.n5863 0.00548485
R29402 avss.n5867 avss.n5866 0.00548485
R29403 avss.n5867 avss.n5862 0.00548485
R29404 avss.n6062 avss.n6061 0.00548485
R29405 avss.n6060 avss.n4373 0.00548485
R29406 avss.n6068 avss.n4373 0.00548485
R29407 avss.n5515 avss.n5510 0.00548485
R29408 avss.n5514 avss.n5513 0.00548485
R29409 avss.n5514 avss.n5509 0.00548485
R29410 avss.n5709 avss.n5708 0.00548485
R29411 avss.n5707 avss.n4457 0.00548485
R29412 avss.n5715 avss.n4457 0.00548485
R29413 avss.n5169 avss.n5164 0.00548485
R29414 avss.n5168 avss.n5167 0.00548485
R29415 avss.n5168 avss.n5163 0.00548485
R29416 avss.n5356 avss.n5355 0.00548485
R29417 avss.n5354 avss.n4541 0.00548485
R29418 avss.n5362 avss.n4541 0.00548485
R29419 avss.n4815 avss.n4810 0.00548485
R29420 avss.n4814 avss.n4813 0.00548485
R29421 avss.n4814 avss.n4809 0.00548485
R29422 avss.n5002 avss.n5001 0.00548485
R29423 avss.n5000 avss.n4625 0.00548485
R29424 avss.n5008 avss.n4625 0.00548485
R29425 avss.n2381 avss.n2380 0.00548485
R29426 avss.n2433 avss.n2432 0.00548485
R29427 avss.n2432 avss.n2431 0.00548485
R29428 avss.n2579 avss.n2578 0.00548485
R29429 avss.n2490 avss.n2489 0.00548485
R29430 avss.n2489 avss.n2488 0.00548485
R29431 avss.n2165 avss.n2164 0.00548485
R29432 avss.n2217 avss.n2216 0.00548485
R29433 avss.n2216 avss.n2215 0.00548485
R29434 avss.n2363 avss.n2362 0.00548485
R29435 avss.n2274 avss.n2273 0.00548485
R29436 avss.n2273 avss.n2272 0.00548485
R29437 avss.n1949 avss.n1948 0.00548485
R29438 avss.n2001 avss.n2000 0.00548485
R29439 avss.n2000 avss.n1999 0.00548485
R29440 avss.n2147 avss.n2146 0.00548485
R29441 avss.n2058 avss.n2057 0.00548485
R29442 avss.n2057 avss.n2056 0.00548485
R29443 avss.n1733 avss.n1732 0.00548485
R29444 avss.n1785 avss.n1784 0.00548485
R29445 avss.n1784 avss.n1783 0.00548485
R29446 avss.n1931 avss.n1930 0.00548485
R29447 avss.n1842 avss.n1841 0.00548485
R29448 avss.n1841 avss.n1840 0.00548485
R29449 avss.n1517 avss.n1516 0.00548485
R29450 avss.n1569 avss.n1568 0.00548485
R29451 avss.n1568 avss.n1567 0.00548485
R29452 avss.n1715 avss.n1714 0.00548485
R29453 avss.n1626 avss.n1625 0.00548485
R29454 avss.n1625 avss.n1624 0.00548485
R29455 avss.n1301 avss.n1300 0.00548485
R29456 avss.n1353 avss.n1352 0.00548485
R29457 avss.n1352 avss.n1351 0.00548485
R29458 avss.n1499 avss.n1498 0.00548485
R29459 avss.n1410 avss.n1409 0.00548485
R29460 avss.n1409 avss.n1408 0.00548485
R29461 avss.n1085 avss.n1084 0.00548485
R29462 avss.n1137 avss.n1136 0.00548485
R29463 avss.n1136 avss.n1135 0.00548485
R29464 avss.n1283 avss.n1282 0.00548485
R29465 avss.n1194 avss.n1193 0.00548485
R29466 avss.n1193 avss.n1192 0.00548485
R29467 avss.n869 avss.n868 0.00548485
R29468 avss.n921 avss.n920 0.00548485
R29469 avss.n920 avss.n919 0.00548485
R29470 avss.n1067 avss.n1066 0.00548485
R29471 avss.n978 avss.n977 0.00548485
R29472 avss.n977 avss.n976 0.00548485
R29473 avss.n653 avss.n652 0.00548485
R29474 avss.n705 avss.n704 0.00548485
R29475 avss.n704 avss.n703 0.00548485
R29476 avss.n851 avss.n850 0.00548485
R29477 avss.n762 avss.n761 0.00548485
R29478 avss.n761 avss.n760 0.00548485
R29479 avss.n437 avss.n436 0.00548485
R29480 avss.n489 avss.n488 0.00548485
R29481 avss.n488 avss.n487 0.00548485
R29482 avss.n635 avss.n634 0.00548485
R29483 avss.n546 avss.n545 0.00548485
R29484 avss.n545 avss.n544 0.00548485
R29485 avss.n11300 avss.n11299 0.00548485
R29486 avss.n11318 avss.n11317 0.00548485
R29487 avss.n11317 avss.n11316 0.00548485
R29488 avss.n310 avss.n309 0.00548485
R29489 avss.n221 avss.n220 0.00548485
R29490 avss.n220 avss.n219 0.00548485
R29491 avss.n11521 avss.n11520 0.00548485
R29492 avss.n11539 avss.n11538 0.00548485
R29493 avss.n11538 avss.n11537 0.00548485
R29494 avss.n93 avss.n92 0.00548485
R29495 avss.n4 avss.n3 0.00548485
R29496 avss.n3 avss.n2 0.00548485
R29497 avss.n8774 avss.n8773 0.0052
R29498 avss.n8832 avss.n8622 0.0052
R29499 avss.n8968 avss.n3671 0.0052
R29500 avss.n8843 avss.n8839 0.0052
R29501 avss.n8843 avss.n3726 0.0052
R29502 avss.n8421 avss.n8420 0.0052
R29503 avss.n8479 avss.n8269 0.0052
R29504 avss.n8615 avss.n3755 0.0052
R29505 avss.n8490 avss.n8486 0.0052
R29506 avss.n8490 avss.n3810 0.0052
R29507 avss.n8068 avss.n8067 0.0052
R29508 avss.n8126 avss.n7916 0.0052
R29509 avss.n8262 avss.n3839 0.0052
R29510 avss.n8137 avss.n8133 0.0052
R29511 avss.n8137 avss.n3894 0.0052
R29512 avss.n7715 avss.n7714 0.0052
R29513 avss.n7773 avss.n7563 0.0052
R29514 avss.n7909 avss.n3923 0.0052
R29515 avss.n7784 avss.n7780 0.0052
R29516 avss.n7784 avss.n3978 0.0052
R29517 avss.n7362 avss.n7361 0.0052
R29518 avss.n7420 avss.n7210 0.0052
R29519 avss.n7556 avss.n4007 0.0052
R29520 avss.n7431 avss.n7427 0.0052
R29521 avss.n7431 avss.n4062 0.0052
R29522 avss.n7009 avss.n7008 0.0052
R29523 avss.n7067 avss.n6857 0.0052
R29524 avss.n7203 avss.n4091 0.0052
R29525 avss.n7078 avss.n7074 0.0052
R29526 avss.n7078 avss.n4146 0.0052
R29527 avss.n6656 avss.n6655 0.0052
R29528 avss.n6714 avss.n6504 0.0052
R29529 avss.n6850 avss.n4175 0.0052
R29530 avss.n6725 avss.n6721 0.0052
R29531 avss.n6725 avss.n4230 0.0052
R29532 avss.n6303 avss.n6302 0.0052
R29533 avss.n6361 avss.n6151 0.0052
R29534 avss.n6497 avss.n4259 0.0052
R29535 avss.n6372 avss.n6368 0.0052
R29536 avss.n6372 avss.n4314 0.0052
R29537 avss.n5950 avss.n5949 0.0052
R29538 avss.n6008 avss.n5798 0.0052
R29539 avss.n6144 avss.n4343 0.0052
R29540 avss.n6019 avss.n6015 0.0052
R29541 avss.n6019 avss.n4398 0.0052
R29542 avss.n5597 avss.n5596 0.0052
R29543 avss.n5655 avss.n5445 0.0052
R29544 avss.n5791 avss.n4427 0.0052
R29545 avss.n5666 avss.n5662 0.0052
R29546 avss.n5666 avss.n4482 0.0052
R29547 avss.n5305 avss.n5089 0.0052
R29548 avss.n5252 avss.n5200 0.0052
R29549 avss.n5252 avss.n5203 0.0052
R29550 avss.n5438 avss.n4511 0.0052
R29551 avss.n5313 avss.n5309 0.0052
R29552 avss.n5313 avss.n4566 0.0052
R29553 avss.n4951 avss.n4735 0.0052
R29554 avss.n4898 avss.n4846 0.0052
R29555 avss.n4898 avss.n4849 0.0052
R29556 avss.n5084 avss.n4595 0.0052
R29557 avss.n4959 avss.n4955 0.0052
R29558 avss.n4959 avss.n4650 0.0052
R29559 avss.n9192 avss.n9191 0.0052
R29560 avss.n2483 avss.n2428 0.0052
R29561 avss.n9081 avss.n9064 0.0052
R29562 avss.n2593 avss.n2592 0.0052
R29563 avss.n2592 avss.n2575 0.0052
R29564 avss.n9413 avss.n9412 0.0052
R29565 avss.n2267 avss.n2212 0.0052
R29566 avss.n9302 avss.n9285 0.0052
R29567 avss.n2377 avss.n2376 0.0052
R29568 avss.n2376 avss.n2359 0.0052
R29569 avss.n9634 avss.n9633 0.0052
R29570 avss.n2051 avss.n1996 0.0052
R29571 avss.n9523 avss.n9506 0.0052
R29572 avss.n2161 avss.n2160 0.0052
R29573 avss.n2160 avss.n2143 0.0052
R29574 avss.n9855 avss.n9854 0.0052
R29575 avss.n1835 avss.n1780 0.0052
R29576 avss.n9744 avss.n9727 0.0052
R29577 avss.n1945 avss.n1944 0.0052
R29578 avss.n1944 avss.n1927 0.0052
R29579 avss.n10076 avss.n10075 0.0052
R29580 avss.n1619 avss.n1564 0.0052
R29581 avss.n9965 avss.n9948 0.0052
R29582 avss.n1729 avss.n1728 0.0052
R29583 avss.n1728 avss.n1711 0.0052
R29584 avss.n10297 avss.n10296 0.0052
R29585 avss.n1403 avss.n1348 0.0052
R29586 avss.n10186 avss.n10169 0.0052
R29587 avss.n1513 avss.n1512 0.0052
R29588 avss.n1512 avss.n1495 0.0052
R29589 avss.n10518 avss.n10517 0.0052
R29590 avss.n1187 avss.n1132 0.0052
R29591 avss.n10407 avss.n10390 0.0052
R29592 avss.n1297 avss.n1296 0.0052
R29593 avss.n1296 avss.n1279 0.0052
R29594 avss.n10739 avss.n10738 0.0052
R29595 avss.n971 avss.n916 0.0052
R29596 avss.n10628 avss.n10611 0.0052
R29597 avss.n1081 avss.n1080 0.0052
R29598 avss.n1080 avss.n1063 0.0052
R29599 avss.n10960 avss.n10959 0.0052
R29600 avss.n755 avss.n700 0.0052
R29601 avss.n10849 avss.n10832 0.0052
R29602 avss.n865 avss.n864 0.0052
R29603 avss.n864 avss.n847 0.0052
R29604 avss.n11181 avss.n11180 0.0052
R29605 avss.n539 avss.n484 0.0052
R29606 avss.n11070 avss.n11053 0.0052
R29607 avss.n649 avss.n648 0.0052
R29608 avss.n648 avss.n631 0.0052
R29609 avss.n11404 avss.n11403 0.0052
R29610 avss.n432 avss.n356 0.0052
R29611 avss.n433 avss.n432 0.0052
R29612 avss.n11291 avss.n11274 0.0052
R29613 avss.n324 avss.n323 0.0052
R29614 avss.n323 avss.n306 0.0052
R29615 avss.n11625 avss.n11624 0.0052
R29616 avss.n215 avss.n139 0.0052
R29617 avss.n216 avss.n215 0.0052
R29618 avss.n11512 avss.n11495 0.0052
R29619 avss.n107 avss.n106 0.0052
R29620 avss.n106 avss.n89 0.0052
R29621 avss.n3513 avss.n3512 0.0051875
R29622 avss.n8794 avss.n8701 0.00477273
R29623 avss.n8912 avss.n3694 0.00477273
R29624 avss.n8441 avss.n8348 0.00477273
R29625 avss.n8559 avss.n3778 0.00477273
R29626 avss.n8088 avss.n7995 0.00477273
R29627 avss.n8206 avss.n3862 0.00477273
R29628 avss.n7735 avss.n7642 0.00477273
R29629 avss.n7853 avss.n3946 0.00477273
R29630 avss.n7382 avss.n7289 0.00477273
R29631 avss.n7500 avss.n4030 0.00477273
R29632 avss.n7029 avss.n6936 0.00477273
R29633 avss.n7147 avss.n4114 0.00477273
R29634 avss.n6676 avss.n6583 0.00477273
R29635 avss.n6794 avss.n4198 0.00477273
R29636 avss.n6323 avss.n6230 0.00477273
R29637 avss.n6441 avss.n4282 0.00477273
R29638 avss.n5970 avss.n5877 0.00477273
R29639 avss.n6088 avss.n4366 0.00477273
R29640 avss.n5617 avss.n5524 0.00477273
R29641 avss.n5735 avss.n4450 0.00477273
R29642 avss.n5272 avss.n5178 0.00477273
R29643 avss.n5382 avss.n4534 0.00477273
R29644 avss.n4918 avss.n4824 0.00477273
R29645 avss.n5028 avss.n4618 0.00477273
R29646 avss.n9134 avss.n9133 0.00477273
R29647 avss.n9023 avss.n9022 0.00477273
R29648 avss.n9355 avss.n9354 0.00477273
R29649 avss.n9244 avss.n9243 0.00477273
R29650 avss.n9576 avss.n9575 0.00477273
R29651 avss.n9465 avss.n9464 0.00477273
R29652 avss.n9797 avss.n9796 0.00477273
R29653 avss.n9686 avss.n9685 0.00477273
R29654 avss.n10018 avss.n10017 0.00477273
R29655 avss.n9907 avss.n9906 0.00477273
R29656 avss.n10239 avss.n10238 0.00477273
R29657 avss.n10128 avss.n10127 0.00477273
R29658 avss.n10460 avss.n10459 0.00477273
R29659 avss.n10349 avss.n10348 0.00477273
R29660 avss.n10681 avss.n10680 0.00477273
R29661 avss.n10570 avss.n10569 0.00477273
R29662 avss.n10902 avss.n10901 0.00477273
R29663 avss.n10791 avss.n10790 0.00477273
R29664 avss.n11123 avss.n11122 0.00477273
R29665 avss.n11012 avss.n11011 0.00477273
R29666 avss.n390 avss.n389 0.00477273
R29667 avss.n11233 avss.n11232 0.00477273
R29668 avss.n173 avss.n172 0.00477273
R29669 avss.n11454 avss.n11453 0.00477273
R29670 avss.n8643 avss.n8631 0.00477273
R29671 avss.n3743 avss.n3731 0.00477273
R29672 avss.n8290 avss.n8278 0.00477273
R29673 avss.n3827 avss.n3815 0.00477273
R29674 avss.n7937 avss.n7925 0.00477273
R29675 avss.n3911 avss.n3899 0.00477273
R29676 avss.n7584 avss.n7572 0.00477273
R29677 avss.n3995 avss.n3983 0.00477273
R29678 avss.n7231 avss.n7219 0.00477273
R29679 avss.n4079 avss.n4067 0.00477273
R29680 avss.n6878 avss.n6866 0.00477273
R29681 avss.n4163 avss.n4151 0.00477273
R29682 avss.n6525 avss.n6513 0.00477273
R29683 avss.n4247 avss.n4235 0.00477273
R29684 avss.n6172 avss.n6160 0.00477273
R29685 avss.n4331 avss.n4319 0.00477273
R29686 avss.n5819 avss.n5807 0.00477273
R29687 avss.n4415 avss.n4403 0.00477273
R29688 avss.n5466 avss.n5454 0.00477273
R29689 avss.n4499 avss.n4487 0.00477273
R29690 avss.n5119 avss.n5105 0.00477273
R29691 avss.n4583 avss.n4571 0.00477273
R29692 avss.n4765 avss.n4751 0.00477273
R29693 avss.n4667 avss.n4655 0.00477273
R29694 avss.n2413 avss.n2412 0.00477273
R29695 avss.n2560 avss.n2559 0.00477273
R29696 avss.n2197 avss.n2196 0.00477273
R29697 avss.n2344 avss.n2343 0.00477273
R29698 avss.n1981 avss.n1980 0.00477273
R29699 avss.n2128 avss.n2127 0.00477273
R29700 avss.n1765 avss.n1764 0.00477273
R29701 avss.n1912 avss.n1911 0.00477273
R29702 avss.n1549 avss.n1548 0.00477273
R29703 avss.n1696 avss.n1695 0.00477273
R29704 avss.n1333 avss.n1332 0.00477273
R29705 avss.n1480 avss.n1479 0.00477273
R29706 avss.n1117 avss.n1116 0.00477273
R29707 avss.n1264 avss.n1263 0.00477273
R29708 avss.n901 avss.n900 0.00477273
R29709 avss.n1048 avss.n1047 0.00477273
R29710 avss.n685 avss.n684 0.00477273
R29711 avss.n832 avss.n831 0.00477273
R29712 avss.n469 avss.n468 0.00477273
R29713 avss.n616 avss.n615 0.00477273
R29714 avss.n11388 avss.n11387 0.00477273
R29715 avss.n291 avss.n290 0.00477273
R29716 avss.n11609 avss.n11608 0.00477273
R29717 avss.n74 avss.n73 0.00477273
R29718 avss.n3339 avss.n3338 0.00466667
R29719 avss.n3347 avss.n3294 0.00466667
R29720 avss.n3409 avss.n3408 0.00466667
R29721 avss.n3436 avss.n3199 0.00466667
R29722 avss.n3455 avss.n3454 0.00466667
R29723 avss.n3508 avss.n3174 0.00466667
R29724 avss.n2982 avss.n2958 0.00440625
R29725 avss.n3039 avss.n2942 0.00440625
R29726 avss.n3129 avss.n2928 0.00440625
R29727 avss.n3631 avss.n2608 0.00440625
R29728 avss.n2687 avss.n2673 0.00440625
R29729 avss.n2694 avss.n2671 0.00440625
R29730 avss.n2732 avss.n2646 0.00440625
R29731 avss.n2739 avss.n2644 0.00440625
R29732 avss.n2910 avss.n2629 0.00440625
R29733 avss.n2904 avss.n2903 0.00440625
R29734 avss.n2869 avss.n2794 0.00440625
R29735 avss.n2863 avss.n2810 0.00440625
R29736 avss.n8785 avss.n8706 0.00428788
R29737 avss.n8784 avss.n8783 0.00428788
R29738 avss.n8829 avss.n8828 0.00428788
R29739 avss.n8825 avss.n8647 0.00428788
R29740 avss.n8761 avss.n8748 0.00428788
R29741 avss.n3749 avss.n3748 0.00428788
R29742 avss.n8846 avss.n3721 0.00428788
R29743 avss.n8918 avss.n8917 0.00428788
R29744 avss.n8930 avss.n3686 0.00428788
R29745 avss.n8963 avss.n8962 0.00428788
R29746 avss.n8432 avss.n8353 0.00428788
R29747 avss.n8431 avss.n8430 0.00428788
R29748 avss.n8476 avss.n8475 0.00428788
R29749 avss.n8472 avss.n8294 0.00428788
R29750 avss.n8408 avss.n8395 0.00428788
R29751 avss.n3833 avss.n3832 0.00428788
R29752 avss.n8493 avss.n3805 0.00428788
R29753 avss.n8565 avss.n8564 0.00428788
R29754 avss.n8577 avss.n3770 0.00428788
R29755 avss.n8610 avss.n8609 0.00428788
R29756 avss.n8079 avss.n8000 0.00428788
R29757 avss.n8078 avss.n8077 0.00428788
R29758 avss.n8123 avss.n8122 0.00428788
R29759 avss.n8119 avss.n7941 0.00428788
R29760 avss.n8055 avss.n8042 0.00428788
R29761 avss.n3917 avss.n3916 0.00428788
R29762 avss.n8140 avss.n3889 0.00428788
R29763 avss.n8212 avss.n8211 0.00428788
R29764 avss.n8224 avss.n3854 0.00428788
R29765 avss.n8257 avss.n8256 0.00428788
R29766 avss.n7726 avss.n7647 0.00428788
R29767 avss.n7725 avss.n7724 0.00428788
R29768 avss.n7770 avss.n7769 0.00428788
R29769 avss.n7766 avss.n7588 0.00428788
R29770 avss.n7702 avss.n7689 0.00428788
R29771 avss.n4001 avss.n4000 0.00428788
R29772 avss.n7787 avss.n3973 0.00428788
R29773 avss.n7859 avss.n7858 0.00428788
R29774 avss.n7871 avss.n3938 0.00428788
R29775 avss.n7904 avss.n7903 0.00428788
R29776 avss.n7373 avss.n7294 0.00428788
R29777 avss.n7372 avss.n7371 0.00428788
R29778 avss.n7417 avss.n7416 0.00428788
R29779 avss.n7413 avss.n7235 0.00428788
R29780 avss.n7349 avss.n7336 0.00428788
R29781 avss.n4085 avss.n4084 0.00428788
R29782 avss.n7434 avss.n4057 0.00428788
R29783 avss.n7506 avss.n7505 0.00428788
R29784 avss.n7518 avss.n4022 0.00428788
R29785 avss.n7551 avss.n7550 0.00428788
R29786 avss.n7020 avss.n6941 0.00428788
R29787 avss.n7019 avss.n7018 0.00428788
R29788 avss.n7064 avss.n7063 0.00428788
R29789 avss.n7060 avss.n6882 0.00428788
R29790 avss.n6996 avss.n6983 0.00428788
R29791 avss.n4169 avss.n4168 0.00428788
R29792 avss.n7081 avss.n4141 0.00428788
R29793 avss.n7153 avss.n7152 0.00428788
R29794 avss.n7165 avss.n4106 0.00428788
R29795 avss.n7198 avss.n7197 0.00428788
R29796 avss.n6667 avss.n6588 0.00428788
R29797 avss.n6666 avss.n6665 0.00428788
R29798 avss.n6711 avss.n6710 0.00428788
R29799 avss.n6707 avss.n6529 0.00428788
R29800 avss.n6643 avss.n6630 0.00428788
R29801 avss.n4253 avss.n4252 0.00428788
R29802 avss.n6728 avss.n4225 0.00428788
R29803 avss.n6800 avss.n6799 0.00428788
R29804 avss.n6812 avss.n4190 0.00428788
R29805 avss.n6845 avss.n6844 0.00428788
R29806 avss.n6314 avss.n6235 0.00428788
R29807 avss.n6313 avss.n6312 0.00428788
R29808 avss.n6358 avss.n6357 0.00428788
R29809 avss.n6354 avss.n6176 0.00428788
R29810 avss.n6290 avss.n6277 0.00428788
R29811 avss.n4337 avss.n4336 0.00428788
R29812 avss.n6375 avss.n4309 0.00428788
R29813 avss.n6447 avss.n6446 0.00428788
R29814 avss.n6459 avss.n4274 0.00428788
R29815 avss.n6492 avss.n6491 0.00428788
R29816 avss.n5961 avss.n5882 0.00428788
R29817 avss.n5960 avss.n5959 0.00428788
R29818 avss.n6005 avss.n6004 0.00428788
R29819 avss.n6001 avss.n5823 0.00428788
R29820 avss.n5937 avss.n5924 0.00428788
R29821 avss.n4421 avss.n4420 0.00428788
R29822 avss.n6022 avss.n4393 0.00428788
R29823 avss.n6094 avss.n6093 0.00428788
R29824 avss.n6106 avss.n4358 0.00428788
R29825 avss.n6139 avss.n6138 0.00428788
R29826 avss.n5608 avss.n5529 0.00428788
R29827 avss.n5607 avss.n5606 0.00428788
R29828 avss.n5652 avss.n5651 0.00428788
R29829 avss.n5648 avss.n5470 0.00428788
R29830 avss.n5584 avss.n5571 0.00428788
R29831 avss.n4505 avss.n4504 0.00428788
R29832 avss.n5669 avss.n4477 0.00428788
R29833 avss.n5741 avss.n5740 0.00428788
R29834 avss.n5753 avss.n4442 0.00428788
R29835 avss.n5786 avss.n5785 0.00428788
R29836 avss.n5263 avss.n5183 0.00428788
R29837 avss.n5262 avss.n5261 0.00428788
R29838 avss.n5124 avss.n5100 0.00428788
R29839 avss.n5129 avss.n5128 0.00428788
R29840 avss.n5243 avss.n5228 0.00428788
R29841 avss.n4589 avss.n4588 0.00428788
R29842 avss.n5316 avss.n4561 0.00428788
R29843 avss.n5388 avss.n5387 0.00428788
R29844 avss.n5400 avss.n4526 0.00428788
R29845 avss.n5433 avss.n5432 0.00428788
R29846 avss.n4909 avss.n4829 0.00428788
R29847 avss.n4908 avss.n4907 0.00428788
R29848 avss.n4770 avss.n4746 0.00428788
R29849 avss.n4775 avss.n4774 0.00428788
R29850 avss.n4889 avss.n4874 0.00428788
R29851 avss.n4673 avss.n4672 0.00428788
R29852 avss.n4962 avss.n4645 0.00428788
R29853 avss.n5034 avss.n5033 0.00428788
R29854 avss.n5046 avss.n4610 0.00428788
R29855 avss.n5079 avss.n5078 0.00428788
R29856 avss.n9148 avss.n9147 0.00428788
R29857 avss.n9146 avss.n9145 0.00428788
R29858 avss.n2405 avss.n2404 0.00428788
R29859 avss.n2403 avss.n2402 0.00428788
R29860 avss.n9091 avss.n9090 0.00428788
R29861 avss.n2552 avss.n2551 0.00428788
R29862 avss.n2550 avss.n2549 0.00428788
R29863 avss.n9037 avss.n9036 0.00428788
R29864 avss.n9035 avss.n9034 0.00428788
R29865 avss.n9071 avss.n9070 0.00428788
R29866 avss.n9369 avss.n9368 0.00428788
R29867 avss.n9367 avss.n9366 0.00428788
R29868 avss.n2189 avss.n2188 0.00428788
R29869 avss.n2187 avss.n2186 0.00428788
R29870 avss.n9312 avss.n9311 0.00428788
R29871 avss.n2336 avss.n2335 0.00428788
R29872 avss.n2334 avss.n2333 0.00428788
R29873 avss.n9258 avss.n9257 0.00428788
R29874 avss.n9256 avss.n9255 0.00428788
R29875 avss.n9292 avss.n9291 0.00428788
R29876 avss.n9590 avss.n9589 0.00428788
R29877 avss.n9588 avss.n9587 0.00428788
R29878 avss.n1973 avss.n1972 0.00428788
R29879 avss.n1971 avss.n1970 0.00428788
R29880 avss.n9533 avss.n9532 0.00428788
R29881 avss.n2120 avss.n2119 0.00428788
R29882 avss.n2118 avss.n2117 0.00428788
R29883 avss.n9479 avss.n9478 0.00428788
R29884 avss.n9477 avss.n9476 0.00428788
R29885 avss.n9513 avss.n9512 0.00428788
R29886 avss.n9811 avss.n9810 0.00428788
R29887 avss.n9809 avss.n9808 0.00428788
R29888 avss.n1757 avss.n1756 0.00428788
R29889 avss.n1755 avss.n1754 0.00428788
R29890 avss.n9754 avss.n9753 0.00428788
R29891 avss.n1904 avss.n1903 0.00428788
R29892 avss.n1902 avss.n1901 0.00428788
R29893 avss.n9700 avss.n9699 0.00428788
R29894 avss.n9698 avss.n9697 0.00428788
R29895 avss.n9734 avss.n9733 0.00428788
R29896 avss.n10032 avss.n10031 0.00428788
R29897 avss.n10030 avss.n10029 0.00428788
R29898 avss.n1541 avss.n1540 0.00428788
R29899 avss.n1539 avss.n1538 0.00428788
R29900 avss.n9975 avss.n9974 0.00428788
R29901 avss.n1688 avss.n1687 0.00428788
R29902 avss.n1686 avss.n1685 0.00428788
R29903 avss.n9921 avss.n9920 0.00428788
R29904 avss.n9919 avss.n9918 0.00428788
R29905 avss.n9955 avss.n9954 0.00428788
R29906 avss.n10253 avss.n10252 0.00428788
R29907 avss.n10251 avss.n10250 0.00428788
R29908 avss.n1325 avss.n1324 0.00428788
R29909 avss.n1323 avss.n1322 0.00428788
R29910 avss.n10196 avss.n10195 0.00428788
R29911 avss.n1472 avss.n1471 0.00428788
R29912 avss.n1470 avss.n1469 0.00428788
R29913 avss.n10142 avss.n10141 0.00428788
R29914 avss.n10140 avss.n10139 0.00428788
R29915 avss.n10176 avss.n10175 0.00428788
R29916 avss.n10474 avss.n10473 0.00428788
R29917 avss.n10472 avss.n10471 0.00428788
R29918 avss.n1109 avss.n1108 0.00428788
R29919 avss.n1107 avss.n1106 0.00428788
R29920 avss.n10417 avss.n10416 0.00428788
R29921 avss.n1256 avss.n1255 0.00428788
R29922 avss.n1254 avss.n1253 0.00428788
R29923 avss.n10363 avss.n10362 0.00428788
R29924 avss.n10361 avss.n10360 0.00428788
R29925 avss.n10397 avss.n10396 0.00428788
R29926 avss.n10695 avss.n10694 0.00428788
R29927 avss.n10693 avss.n10692 0.00428788
R29928 avss.n893 avss.n892 0.00428788
R29929 avss.n891 avss.n890 0.00428788
R29930 avss.n10638 avss.n10637 0.00428788
R29931 avss.n1040 avss.n1039 0.00428788
R29932 avss.n1038 avss.n1037 0.00428788
R29933 avss.n10584 avss.n10583 0.00428788
R29934 avss.n10582 avss.n10581 0.00428788
R29935 avss.n10618 avss.n10617 0.00428788
R29936 avss.n10916 avss.n10915 0.00428788
R29937 avss.n10914 avss.n10913 0.00428788
R29938 avss.n677 avss.n676 0.00428788
R29939 avss.n675 avss.n674 0.00428788
R29940 avss.n10859 avss.n10858 0.00428788
R29941 avss.n824 avss.n823 0.00428788
R29942 avss.n822 avss.n821 0.00428788
R29943 avss.n10805 avss.n10804 0.00428788
R29944 avss.n10803 avss.n10802 0.00428788
R29945 avss.n10839 avss.n10838 0.00428788
R29946 avss.n11137 avss.n11136 0.00428788
R29947 avss.n11135 avss.n11134 0.00428788
R29948 avss.n461 avss.n460 0.00428788
R29949 avss.n459 avss.n458 0.00428788
R29950 avss.n11080 avss.n11079 0.00428788
R29951 avss.n608 avss.n607 0.00428788
R29952 avss.n606 avss.n605 0.00428788
R29953 avss.n11026 avss.n11025 0.00428788
R29954 avss.n11024 avss.n11023 0.00428788
R29955 avss.n11060 avss.n11059 0.00428788
R29956 avss.n404 avss.n403 0.00428788
R29957 avss.n402 avss.n401 0.00428788
R29958 avss.n11379 avss.n11378 0.00428788
R29959 avss.n11377 avss.n11376 0.00428788
R29960 avss.n331 avss.n330 0.00428788
R29961 avss.n283 avss.n282 0.00428788
R29962 avss.n281 avss.n280 0.00428788
R29963 avss.n11247 avss.n11246 0.00428788
R29964 avss.n11245 avss.n11244 0.00428788
R29965 avss.n11281 avss.n11280 0.00428788
R29966 avss.n187 avss.n186 0.00428788
R29967 avss.n185 avss.n184 0.00428788
R29968 avss.n11600 avss.n11599 0.00428788
R29969 avss.n11598 avss.n11597 0.00428788
R29970 avss.n114 avss.n113 0.00428788
R29971 avss.n66 avss.n65 0.00428788
R29972 avss.n64 avss.n63 0.00428788
R29973 avss.n11468 avss.n11467 0.00428788
R29974 avss.n11466 avss.n11465 0.00428788
R29975 avss.n11502 avss.n11501 0.00428788
R29976 avss.n8809 avss.n8808 0.00406061
R29977 avss.n8820 avss.n8650 0.00406061
R29978 avss.n8810 avss.n8663 0.00406061
R29979 avss.n8733 avss.n8721 0.00406061
R29980 avss.n8772 avss.n8727 0.00406061
R29981 avss.n8875 avss.n3707 0.00406061
R29982 avss.n8840 avss.n3718 0.00406061
R29983 avss.n8874 avss.n3708 0.00406061
R29984 avss.n8933 avss.n3674 0.00406061
R29985 avss.n8456 avss.n8455 0.00406061
R29986 avss.n8467 avss.n8297 0.00406061
R29987 avss.n8457 avss.n8310 0.00406061
R29988 avss.n8380 avss.n8368 0.00406061
R29989 avss.n8419 avss.n8374 0.00406061
R29990 avss.n8522 avss.n3791 0.00406061
R29991 avss.n8487 avss.n3802 0.00406061
R29992 avss.n8521 avss.n3792 0.00406061
R29993 avss.n8580 avss.n3758 0.00406061
R29994 avss.n8103 avss.n8102 0.00406061
R29995 avss.n8114 avss.n7944 0.00406061
R29996 avss.n8104 avss.n7957 0.00406061
R29997 avss.n8027 avss.n8015 0.00406061
R29998 avss.n8066 avss.n8021 0.00406061
R29999 avss.n8169 avss.n3875 0.00406061
R30000 avss.n8134 avss.n3886 0.00406061
R30001 avss.n8168 avss.n3876 0.00406061
R30002 avss.n8227 avss.n3842 0.00406061
R30003 avss.n7750 avss.n7749 0.00406061
R30004 avss.n7761 avss.n7591 0.00406061
R30005 avss.n7751 avss.n7604 0.00406061
R30006 avss.n7674 avss.n7662 0.00406061
R30007 avss.n7713 avss.n7668 0.00406061
R30008 avss.n7816 avss.n3959 0.00406061
R30009 avss.n7781 avss.n3970 0.00406061
R30010 avss.n7815 avss.n3960 0.00406061
R30011 avss.n7874 avss.n3926 0.00406061
R30012 avss.n7397 avss.n7396 0.00406061
R30013 avss.n7408 avss.n7238 0.00406061
R30014 avss.n7398 avss.n7251 0.00406061
R30015 avss.n7321 avss.n7309 0.00406061
R30016 avss.n7360 avss.n7315 0.00406061
R30017 avss.n7463 avss.n4043 0.00406061
R30018 avss.n7428 avss.n4054 0.00406061
R30019 avss.n7462 avss.n4044 0.00406061
R30020 avss.n7521 avss.n4010 0.00406061
R30021 avss.n7044 avss.n7043 0.00406061
R30022 avss.n7055 avss.n6885 0.00406061
R30023 avss.n7045 avss.n6898 0.00406061
R30024 avss.n6968 avss.n6956 0.00406061
R30025 avss.n7007 avss.n6962 0.00406061
R30026 avss.n7110 avss.n4127 0.00406061
R30027 avss.n7075 avss.n4138 0.00406061
R30028 avss.n7109 avss.n4128 0.00406061
R30029 avss.n7168 avss.n4094 0.00406061
R30030 avss.n6691 avss.n6690 0.00406061
R30031 avss.n6702 avss.n6532 0.00406061
R30032 avss.n6692 avss.n6545 0.00406061
R30033 avss.n6615 avss.n6603 0.00406061
R30034 avss.n6654 avss.n6609 0.00406061
R30035 avss.n6757 avss.n4211 0.00406061
R30036 avss.n6722 avss.n4222 0.00406061
R30037 avss.n6756 avss.n4212 0.00406061
R30038 avss.n6815 avss.n4178 0.00406061
R30039 avss.n6338 avss.n6337 0.00406061
R30040 avss.n6349 avss.n6179 0.00406061
R30041 avss.n6339 avss.n6192 0.00406061
R30042 avss.n6262 avss.n6250 0.00406061
R30043 avss.n6301 avss.n6256 0.00406061
R30044 avss.n6404 avss.n4295 0.00406061
R30045 avss.n6369 avss.n4306 0.00406061
R30046 avss.n6403 avss.n4296 0.00406061
R30047 avss.n6462 avss.n4262 0.00406061
R30048 avss.n5985 avss.n5984 0.00406061
R30049 avss.n5996 avss.n5826 0.00406061
R30050 avss.n5986 avss.n5839 0.00406061
R30051 avss.n5909 avss.n5897 0.00406061
R30052 avss.n5948 avss.n5903 0.00406061
R30053 avss.n6051 avss.n4379 0.00406061
R30054 avss.n6016 avss.n4390 0.00406061
R30055 avss.n6050 avss.n4380 0.00406061
R30056 avss.n6109 avss.n4346 0.00406061
R30057 avss.n5632 avss.n5631 0.00406061
R30058 avss.n5643 avss.n5473 0.00406061
R30059 avss.n5633 avss.n5486 0.00406061
R30060 avss.n5556 avss.n5544 0.00406061
R30061 avss.n5595 avss.n5550 0.00406061
R30062 avss.n5698 avss.n4463 0.00406061
R30063 avss.n5663 avss.n4474 0.00406061
R30064 avss.n5697 avss.n4464 0.00406061
R30065 avss.n5756 avss.n4430 0.00406061
R30066 avss.n5287 avss.n5286 0.00406061
R30067 avss.n5094 avss.n5092 0.00406061
R30068 avss.n5288 avss.n5136 0.00406061
R30069 avss.n5216 avss.n5198 0.00406061
R30070 avss.n5345 avss.n4547 0.00406061
R30071 avss.n5310 avss.n4558 0.00406061
R30072 avss.n5344 avss.n4548 0.00406061
R30073 avss.n5403 avss.n4514 0.00406061
R30074 avss.n4933 avss.n4932 0.00406061
R30075 avss.n4740 avss.n4738 0.00406061
R30076 avss.n4934 avss.n4782 0.00406061
R30077 avss.n4862 avss.n4844 0.00406061
R30078 avss.n4991 avss.n4631 0.00406061
R30079 avss.n4956 avss.n4642 0.00406061
R30080 avss.n4990 avss.n4632 0.00406061
R30081 avss.n5049 avss.n4598 0.00406061
R30082 avss.n2385 avss.n2384 0.00406061
R30083 avss.n2480 avss.n2479 0.00406061
R30084 avss.n2459 avss.n2458 0.00406061
R30085 avss.n9158 avss.n9157 0.00406061
R30086 avss.n9116 avss.n9115 0.00406061
R30087 avss.n2583 avss.n2582 0.00406061
R30088 avss.n2537 avss.n2536 0.00406061
R30089 avss.n2516 avss.n2515 0.00406061
R30090 avss.n9047 avss.n9046 0.00406061
R30091 avss.n2169 avss.n2168 0.00406061
R30092 avss.n2264 avss.n2263 0.00406061
R30093 avss.n2243 avss.n2242 0.00406061
R30094 avss.n9379 avss.n9378 0.00406061
R30095 avss.n9337 avss.n9336 0.00406061
R30096 avss.n2367 avss.n2366 0.00406061
R30097 avss.n2321 avss.n2320 0.00406061
R30098 avss.n2300 avss.n2299 0.00406061
R30099 avss.n9268 avss.n9267 0.00406061
R30100 avss.n1953 avss.n1952 0.00406061
R30101 avss.n2048 avss.n2047 0.00406061
R30102 avss.n2027 avss.n2026 0.00406061
R30103 avss.n9600 avss.n9599 0.00406061
R30104 avss.n9558 avss.n9557 0.00406061
R30105 avss.n2151 avss.n2150 0.00406061
R30106 avss.n2105 avss.n2104 0.00406061
R30107 avss.n2084 avss.n2083 0.00406061
R30108 avss.n9489 avss.n9488 0.00406061
R30109 avss.n1737 avss.n1736 0.00406061
R30110 avss.n1832 avss.n1831 0.00406061
R30111 avss.n1811 avss.n1810 0.00406061
R30112 avss.n9821 avss.n9820 0.00406061
R30113 avss.n9779 avss.n9778 0.00406061
R30114 avss.n1935 avss.n1934 0.00406061
R30115 avss.n1889 avss.n1888 0.00406061
R30116 avss.n1868 avss.n1867 0.00406061
R30117 avss.n9710 avss.n9709 0.00406061
R30118 avss.n1521 avss.n1520 0.00406061
R30119 avss.n1616 avss.n1615 0.00406061
R30120 avss.n1595 avss.n1594 0.00406061
R30121 avss.n10042 avss.n10041 0.00406061
R30122 avss.n10000 avss.n9999 0.00406061
R30123 avss.n1719 avss.n1718 0.00406061
R30124 avss.n1673 avss.n1672 0.00406061
R30125 avss.n1652 avss.n1651 0.00406061
R30126 avss.n9931 avss.n9930 0.00406061
R30127 avss.n1305 avss.n1304 0.00406061
R30128 avss.n1400 avss.n1399 0.00406061
R30129 avss.n1379 avss.n1378 0.00406061
R30130 avss.n10263 avss.n10262 0.00406061
R30131 avss.n10221 avss.n10220 0.00406061
R30132 avss.n1503 avss.n1502 0.00406061
R30133 avss.n1457 avss.n1456 0.00406061
R30134 avss.n1436 avss.n1435 0.00406061
R30135 avss.n10152 avss.n10151 0.00406061
R30136 avss.n1089 avss.n1088 0.00406061
R30137 avss.n1184 avss.n1183 0.00406061
R30138 avss.n1163 avss.n1162 0.00406061
R30139 avss.n10484 avss.n10483 0.00406061
R30140 avss.n10442 avss.n10441 0.00406061
R30141 avss.n1287 avss.n1286 0.00406061
R30142 avss.n1241 avss.n1240 0.00406061
R30143 avss.n1220 avss.n1219 0.00406061
R30144 avss.n10373 avss.n10372 0.00406061
R30145 avss.n873 avss.n872 0.00406061
R30146 avss.n968 avss.n967 0.00406061
R30147 avss.n947 avss.n946 0.00406061
R30148 avss.n10705 avss.n10704 0.00406061
R30149 avss.n10663 avss.n10662 0.00406061
R30150 avss.n1071 avss.n1070 0.00406061
R30151 avss.n1025 avss.n1024 0.00406061
R30152 avss.n1004 avss.n1003 0.00406061
R30153 avss.n10594 avss.n10593 0.00406061
R30154 avss.n657 avss.n656 0.00406061
R30155 avss.n752 avss.n751 0.00406061
R30156 avss.n731 avss.n730 0.00406061
R30157 avss.n10926 avss.n10925 0.00406061
R30158 avss.n10884 avss.n10883 0.00406061
R30159 avss.n855 avss.n854 0.00406061
R30160 avss.n809 avss.n808 0.00406061
R30161 avss.n788 avss.n787 0.00406061
R30162 avss.n10815 avss.n10814 0.00406061
R30163 avss.n441 avss.n440 0.00406061
R30164 avss.n536 avss.n535 0.00406061
R30165 avss.n515 avss.n514 0.00406061
R30166 avss.n11147 avss.n11146 0.00406061
R30167 avss.n11105 avss.n11104 0.00406061
R30168 avss.n639 avss.n638 0.00406061
R30169 avss.n593 avss.n592 0.00406061
R30170 avss.n572 avss.n571 0.00406061
R30171 avss.n11036 avss.n11035 0.00406061
R30172 avss.n11304 avss.n11303 0.00406061
R30173 avss.n11365 avss.n11364 0.00406061
R30174 avss.n11344 avss.n11343 0.00406061
R30175 avss.n414 avss.n413 0.00406061
R30176 avss.n314 avss.n313 0.00406061
R30177 avss.n268 avss.n267 0.00406061
R30178 avss.n247 avss.n246 0.00406061
R30179 avss.n11257 avss.n11256 0.00406061
R30180 avss.n11525 avss.n11524 0.00406061
R30181 avss.n11586 avss.n11585 0.00406061
R30182 avss.n11565 avss.n11564 0.00406061
R30183 avss.n197 avss.n196 0.00406061
R30184 avss.n97 avss.n96 0.00406061
R30185 avss.n51 avss.n50 0.00406061
R30186 avss.n30 avss.n29 0.00406061
R30187 avss.n11478 avss.n11477 0.00406061
R30188 avss.n8774 avss.n8723 0.00334838
R30189 avss.n8835 avss.n8620 0.00334838
R30190 avss.n8832 avss.n8620 0.00334838
R30191 avss.n8968 avss.n3669 0.00334838
R30192 avss.n8971 avss.n3669 0.00334838
R30193 avss.n8421 avss.n8370 0.00334838
R30194 avss.n8482 avss.n8267 0.00334838
R30195 avss.n8479 avss.n8267 0.00334838
R30196 avss.n8615 avss.n3753 0.00334838
R30197 avss.n8618 avss.n3753 0.00334838
R30198 avss.n8068 avss.n8017 0.00334838
R30199 avss.n8129 avss.n7914 0.00334838
R30200 avss.n8126 avss.n7914 0.00334838
R30201 avss.n8262 avss.n3837 0.00334838
R30202 avss.n8265 avss.n3837 0.00334838
R30203 avss.n7715 avss.n7664 0.00334838
R30204 avss.n7776 avss.n7561 0.00334838
R30205 avss.n7773 avss.n7561 0.00334838
R30206 avss.n7909 avss.n3921 0.00334838
R30207 avss.n7912 avss.n3921 0.00334838
R30208 avss.n7362 avss.n7311 0.00334838
R30209 avss.n7423 avss.n7208 0.00334838
R30210 avss.n7420 avss.n7208 0.00334838
R30211 avss.n7556 avss.n4005 0.00334838
R30212 avss.n7559 avss.n4005 0.00334838
R30213 avss.n7009 avss.n6958 0.00334838
R30214 avss.n7070 avss.n6855 0.00334838
R30215 avss.n7067 avss.n6855 0.00334838
R30216 avss.n7203 avss.n4089 0.00334838
R30217 avss.n7206 avss.n4089 0.00334838
R30218 avss.n6656 avss.n6605 0.00334838
R30219 avss.n6717 avss.n6502 0.00334838
R30220 avss.n6714 avss.n6502 0.00334838
R30221 avss.n6850 avss.n4173 0.00334838
R30222 avss.n6853 avss.n4173 0.00334838
R30223 avss.n6303 avss.n6252 0.00334838
R30224 avss.n6364 avss.n6149 0.00334838
R30225 avss.n6361 avss.n6149 0.00334838
R30226 avss.n6497 avss.n4257 0.00334838
R30227 avss.n6500 avss.n4257 0.00334838
R30228 avss.n5950 avss.n5899 0.00334838
R30229 avss.n6011 avss.n5796 0.00334838
R30230 avss.n6008 avss.n5796 0.00334838
R30231 avss.n6144 avss.n4341 0.00334838
R30232 avss.n6147 avss.n4341 0.00334838
R30233 avss.n5597 avss.n5546 0.00334838
R30234 avss.n5658 avss.n5443 0.00334838
R30235 avss.n5655 avss.n5443 0.00334838
R30236 avss.n5791 avss.n4425 0.00334838
R30237 avss.n5794 avss.n4425 0.00334838
R30238 avss.n5303 avss.n5089 0.00334838
R30239 avss.n5438 avss.n4509 0.00334838
R30240 avss.n5441 avss.n4509 0.00334838
R30241 avss.n4949 avss.n4735 0.00334838
R30242 avss.n5084 avss.n4593 0.00334838
R30243 avss.n5087 avss.n4593 0.00334838
R30244 avss.n9191 avss.n9101 0.00334838
R30245 avss.n2485 avss.n2484 0.00334838
R30246 avss.n2484 avss.n2483 0.00334838
R30247 avss.n9082 avss.n9081 0.00334838
R30248 avss.n9083 avss.n9082 0.00334838
R30249 avss.n9412 avss.n9322 0.00334838
R30250 avss.n2269 avss.n2268 0.00334838
R30251 avss.n2268 avss.n2267 0.00334838
R30252 avss.n9303 avss.n9302 0.00334838
R30253 avss.n9304 avss.n9303 0.00334838
R30254 avss.n9633 avss.n9543 0.00334838
R30255 avss.n2053 avss.n2052 0.00334838
R30256 avss.n2052 avss.n2051 0.00334838
R30257 avss.n9524 avss.n9523 0.00334838
R30258 avss.n9525 avss.n9524 0.00334838
R30259 avss.n9854 avss.n9764 0.00334838
R30260 avss.n1837 avss.n1836 0.00334838
R30261 avss.n1836 avss.n1835 0.00334838
R30262 avss.n9745 avss.n9744 0.00334838
R30263 avss.n9746 avss.n9745 0.00334838
R30264 avss.n10075 avss.n9985 0.00334838
R30265 avss.n1621 avss.n1620 0.00334838
R30266 avss.n1620 avss.n1619 0.00334838
R30267 avss.n9966 avss.n9965 0.00334838
R30268 avss.n9967 avss.n9966 0.00334838
R30269 avss.n10296 avss.n10206 0.00334838
R30270 avss.n1405 avss.n1404 0.00334838
R30271 avss.n1404 avss.n1403 0.00334838
R30272 avss.n10187 avss.n10186 0.00334838
R30273 avss.n10188 avss.n10187 0.00334838
R30274 avss.n10517 avss.n10427 0.00334838
R30275 avss.n1189 avss.n1188 0.00334838
R30276 avss.n1188 avss.n1187 0.00334838
R30277 avss.n10408 avss.n10407 0.00334838
R30278 avss.n10409 avss.n10408 0.00334838
R30279 avss.n10738 avss.n10648 0.00334838
R30280 avss.n973 avss.n972 0.00334838
R30281 avss.n972 avss.n971 0.00334838
R30282 avss.n10629 avss.n10628 0.00334838
R30283 avss.n10630 avss.n10629 0.00334838
R30284 avss.n10959 avss.n10869 0.00334838
R30285 avss.n757 avss.n756 0.00334838
R30286 avss.n756 avss.n755 0.00334838
R30287 avss.n10850 avss.n10849 0.00334838
R30288 avss.n10851 avss.n10850 0.00334838
R30289 avss.n11180 avss.n11090 0.00334838
R30290 avss.n541 avss.n540 0.00334838
R30291 avss.n540 avss.n539 0.00334838
R30292 avss.n11071 avss.n11070 0.00334838
R30293 avss.n11072 avss.n11071 0.00334838
R30294 avss.n11403 avss.n11313 0.00334838
R30295 avss.n11292 avss.n11291 0.00334838
R30296 avss.n11293 avss.n11292 0.00334838
R30297 avss.n11624 avss.n11534 0.00334838
R30298 avss.n11513 avss.n11512 0.00334838
R30299 avss.n11514 avss.n11513 0.00334838
R30300 avss.n8969 avss.n3672 0.00277937
R30301 avss.n8970 avss.n8969 0.00277937
R30302 avss.n8616 avss.n3756 0.00277937
R30303 avss.n8617 avss.n8616 0.00277937
R30304 avss.n8263 avss.n3840 0.00277937
R30305 avss.n8264 avss.n8263 0.00277937
R30306 avss.n7910 avss.n3924 0.00277937
R30307 avss.n7911 avss.n7910 0.00277937
R30308 avss.n7557 avss.n4008 0.00277937
R30309 avss.n7558 avss.n7557 0.00277937
R30310 avss.n7204 avss.n4092 0.00277937
R30311 avss.n7205 avss.n7204 0.00277937
R30312 avss.n6851 avss.n4176 0.00277937
R30313 avss.n6852 avss.n6851 0.00277937
R30314 avss.n6498 avss.n4260 0.00277937
R30315 avss.n6499 avss.n6498 0.00277937
R30316 avss.n6145 avss.n4344 0.00277937
R30317 avss.n6146 avss.n6145 0.00277937
R30318 avss.n5792 avss.n4428 0.00277937
R30319 avss.n5793 avss.n5792 0.00277937
R30320 avss.n5251 avss.n5250 0.00277937
R30321 avss.n5251 avss.n5206 0.00277937
R30322 avss.n5439 avss.n4512 0.00277937
R30323 avss.n5440 avss.n5439 0.00277937
R30324 avss.n4897 avss.n4896 0.00277937
R30325 avss.n4897 avss.n4852 0.00277937
R30326 avss.n5085 avss.n4596 0.00277937
R30327 avss.n5086 avss.n5085 0.00277937
R30328 avss.n9004 avss.n9003 0.00277937
R30329 avss.n9005 avss.n9004 0.00277937
R30330 avss.n9225 avss.n9224 0.00277937
R30331 avss.n9226 avss.n9225 0.00277937
R30332 avss.n9446 avss.n9445 0.00277937
R30333 avss.n9447 avss.n9446 0.00277937
R30334 avss.n9667 avss.n9666 0.00277937
R30335 avss.n9668 avss.n9667 0.00277937
R30336 avss.n9888 avss.n9887 0.00277937
R30337 avss.n9889 avss.n9888 0.00277937
R30338 avss.n10109 avss.n10108 0.00277937
R30339 avss.n10110 avss.n10109 0.00277937
R30340 avss.n10330 avss.n10329 0.00277937
R30341 avss.n10331 avss.n10330 0.00277937
R30342 avss.n10551 avss.n10550 0.00277937
R30343 avss.n10552 avss.n10551 0.00277937
R30344 avss.n10772 avss.n10771 0.00277937
R30345 avss.n10773 avss.n10772 0.00277937
R30346 avss.n10993 avss.n10992 0.00277937
R30347 avss.n10994 avss.n10993 0.00277937
R30348 avss.n371 avss.n370 0.00277937
R30349 avss.n372 avss.n371 0.00277937
R30350 avss.n11214 avss.n11213 0.00277937
R30351 avss.n11215 avss.n11214 0.00277937
R30352 avss.n154 avss.n153 0.00277937
R30353 avss.n155 avss.n154 0.00277937
R30354 avss.n11435 avss.n11434 0.00277937
R30355 avss.n11436 avss.n11435 0.00277937
R30356 avss.n8698 avss.n8697 0.00263636
R30357 avss.n8638 avss.n8633 0.00263636
R30358 avss.n8690 avss.n8688 0.00263636
R30359 avss.n8696 avss.n8683 0.00263636
R30360 avss.n8702 avss.n8684 0.00263636
R30361 avss.n8754 avss.n8750 0.00263636
R30362 avss.n8888 avss.n3696 0.00263636
R30363 avss.n3738 avss.n3733 0.00263636
R30364 avss.n8884 avss.n8883 0.00263636
R30365 avss.n8887 avss.n3697 0.00263636
R30366 avss.n8898 avss.n3698 0.00263636
R30367 avss.n8958 avss.n8957 0.00263636
R30368 avss.n8345 avss.n8344 0.00263636
R30369 avss.n8285 avss.n8280 0.00263636
R30370 avss.n8337 avss.n8335 0.00263636
R30371 avss.n8343 avss.n8330 0.00263636
R30372 avss.n8349 avss.n8331 0.00263636
R30373 avss.n8401 avss.n8397 0.00263636
R30374 avss.n8535 avss.n3780 0.00263636
R30375 avss.n3822 avss.n3817 0.00263636
R30376 avss.n8531 avss.n8530 0.00263636
R30377 avss.n8534 avss.n3781 0.00263636
R30378 avss.n8545 avss.n3782 0.00263636
R30379 avss.n8605 avss.n8604 0.00263636
R30380 avss.n7992 avss.n7991 0.00263636
R30381 avss.n7932 avss.n7927 0.00263636
R30382 avss.n7984 avss.n7982 0.00263636
R30383 avss.n7990 avss.n7977 0.00263636
R30384 avss.n7996 avss.n7978 0.00263636
R30385 avss.n8048 avss.n8044 0.00263636
R30386 avss.n8182 avss.n3864 0.00263636
R30387 avss.n3906 avss.n3901 0.00263636
R30388 avss.n8178 avss.n8177 0.00263636
R30389 avss.n8181 avss.n3865 0.00263636
R30390 avss.n8192 avss.n3866 0.00263636
R30391 avss.n8252 avss.n8251 0.00263636
R30392 avss.n7639 avss.n7638 0.00263636
R30393 avss.n7579 avss.n7574 0.00263636
R30394 avss.n7631 avss.n7629 0.00263636
R30395 avss.n7637 avss.n7624 0.00263636
R30396 avss.n7643 avss.n7625 0.00263636
R30397 avss.n7695 avss.n7691 0.00263636
R30398 avss.n7829 avss.n3948 0.00263636
R30399 avss.n3990 avss.n3985 0.00263636
R30400 avss.n7825 avss.n7824 0.00263636
R30401 avss.n7828 avss.n3949 0.00263636
R30402 avss.n7839 avss.n3950 0.00263636
R30403 avss.n7899 avss.n7898 0.00263636
R30404 avss.n7286 avss.n7285 0.00263636
R30405 avss.n7226 avss.n7221 0.00263636
R30406 avss.n7278 avss.n7276 0.00263636
R30407 avss.n7284 avss.n7271 0.00263636
R30408 avss.n7290 avss.n7272 0.00263636
R30409 avss.n7342 avss.n7338 0.00263636
R30410 avss.n7476 avss.n4032 0.00263636
R30411 avss.n4074 avss.n4069 0.00263636
R30412 avss.n7472 avss.n7471 0.00263636
R30413 avss.n7475 avss.n4033 0.00263636
R30414 avss.n7486 avss.n4034 0.00263636
R30415 avss.n7546 avss.n7545 0.00263636
R30416 avss.n6933 avss.n6932 0.00263636
R30417 avss.n6873 avss.n6868 0.00263636
R30418 avss.n6925 avss.n6923 0.00263636
R30419 avss.n6931 avss.n6918 0.00263636
R30420 avss.n6937 avss.n6919 0.00263636
R30421 avss.n6989 avss.n6985 0.00263636
R30422 avss.n7123 avss.n4116 0.00263636
R30423 avss.n4158 avss.n4153 0.00263636
R30424 avss.n7119 avss.n7118 0.00263636
R30425 avss.n7122 avss.n4117 0.00263636
R30426 avss.n7133 avss.n4118 0.00263636
R30427 avss.n7193 avss.n7192 0.00263636
R30428 avss.n6580 avss.n6579 0.00263636
R30429 avss.n6520 avss.n6515 0.00263636
R30430 avss.n6572 avss.n6570 0.00263636
R30431 avss.n6578 avss.n6565 0.00263636
R30432 avss.n6584 avss.n6566 0.00263636
R30433 avss.n6636 avss.n6632 0.00263636
R30434 avss.n6770 avss.n4200 0.00263636
R30435 avss.n4242 avss.n4237 0.00263636
R30436 avss.n6766 avss.n6765 0.00263636
R30437 avss.n6769 avss.n4201 0.00263636
R30438 avss.n6780 avss.n4202 0.00263636
R30439 avss.n6840 avss.n6839 0.00263636
R30440 avss.n6227 avss.n6226 0.00263636
R30441 avss.n6167 avss.n6162 0.00263636
R30442 avss.n6219 avss.n6217 0.00263636
R30443 avss.n6225 avss.n6212 0.00263636
R30444 avss.n6231 avss.n6213 0.00263636
R30445 avss.n6283 avss.n6279 0.00263636
R30446 avss.n6417 avss.n4284 0.00263636
R30447 avss.n4326 avss.n4321 0.00263636
R30448 avss.n6413 avss.n6412 0.00263636
R30449 avss.n6416 avss.n4285 0.00263636
R30450 avss.n6427 avss.n4286 0.00263636
R30451 avss.n6487 avss.n6486 0.00263636
R30452 avss.n5874 avss.n5873 0.00263636
R30453 avss.n5814 avss.n5809 0.00263636
R30454 avss.n5866 avss.n5864 0.00263636
R30455 avss.n5872 avss.n5859 0.00263636
R30456 avss.n5878 avss.n5860 0.00263636
R30457 avss.n5930 avss.n5926 0.00263636
R30458 avss.n6064 avss.n4368 0.00263636
R30459 avss.n4410 avss.n4405 0.00263636
R30460 avss.n6060 avss.n6059 0.00263636
R30461 avss.n6063 avss.n4369 0.00263636
R30462 avss.n6074 avss.n4370 0.00263636
R30463 avss.n6134 avss.n6133 0.00263636
R30464 avss.n5521 avss.n5520 0.00263636
R30465 avss.n5461 avss.n5456 0.00263636
R30466 avss.n5513 avss.n5511 0.00263636
R30467 avss.n5519 avss.n5506 0.00263636
R30468 avss.n5525 avss.n5507 0.00263636
R30469 avss.n5577 avss.n5573 0.00263636
R30470 avss.n5711 avss.n4452 0.00263636
R30471 avss.n4494 avss.n4489 0.00263636
R30472 avss.n5707 avss.n5706 0.00263636
R30473 avss.n5710 avss.n4453 0.00263636
R30474 avss.n5721 avss.n4454 0.00263636
R30475 avss.n5781 avss.n5780 0.00263636
R30476 avss.n5175 avss.n5174 0.00263636
R30477 avss.n5113 avss.n5108 0.00263636
R30478 avss.n5167 avss.n5165 0.00263636
R30479 avss.n5173 avss.n5160 0.00263636
R30480 avss.n5179 avss.n5161 0.00263636
R30481 avss.n5236 avss.n5232 0.00263636
R30482 avss.n5358 avss.n4536 0.00263636
R30483 avss.n4578 avss.n4573 0.00263636
R30484 avss.n5354 avss.n5353 0.00263636
R30485 avss.n5357 avss.n4537 0.00263636
R30486 avss.n5368 avss.n4538 0.00263636
R30487 avss.n5428 avss.n5427 0.00263636
R30488 avss.n4821 avss.n4820 0.00263636
R30489 avss.n4759 avss.n4754 0.00263636
R30490 avss.n4813 avss.n4811 0.00263636
R30491 avss.n4819 avss.n4806 0.00263636
R30492 avss.n4825 avss.n4807 0.00263636
R30493 avss.n4882 avss.n4878 0.00263636
R30494 avss.n5004 avss.n4620 0.00263636
R30495 avss.n4662 avss.n4657 0.00263636
R30496 avss.n5000 avss.n4999 0.00263636
R30497 avss.n5003 avss.n4621 0.00263636
R30498 avss.n5014 avss.n4622 0.00263636
R30499 avss.n5074 avss.n5073 0.00263636
R30500 avss.n9177 avss.n9176 0.00263636
R30501 avss.n2423 avss.n2422 0.00263636
R30502 avss.n2442 avss.n2433 0.00263636
R30503 avss.n9119 avss.n9118 0.00263636
R30504 avss.n9122 avss.n9121 0.00263636
R30505 avss.n9097 avss.n9096 0.00263636
R30506 avss.n8976 avss.n8975 0.00263636
R30507 avss.n2570 avss.n2569 0.00263636
R30508 avss.n2499 avss.n2490 0.00263636
R30509 avss.n9008 avss.n9007 0.00263636
R30510 avss.n9011 avss.n9010 0.00263636
R30511 avss.n9077 avss.n9076 0.00263636
R30512 avss.n9398 avss.n9397 0.00263636
R30513 avss.n2207 avss.n2206 0.00263636
R30514 avss.n2226 avss.n2217 0.00263636
R30515 avss.n9340 avss.n9339 0.00263636
R30516 avss.n9343 avss.n9342 0.00263636
R30517 avss.n9318 avss.n9317 0.00263636
R30518 avss.n9197 avss.n9196 0.00263636
R30519 avss.n2354 avss.n2353 0.00263636
R30520 avss.n2283 avss.n2274 0.00263636
R30521 avss.n9229 avss.n9228 0.00263636
R30522 avss.n9232 avss.n9231 0.00263636
R30523 avss.n9298 avss.n9297 0.00263636
R30524 avss.n9619 avss.n9618 0.00263636
R30525 avss.n1991 avss.n1990 0.00263636
R30526 avss.n2010 avss.n2001 0.00263636
R30527 avss.n9561 avss.n9560 0.00263636
R30528 avss.n9564 avss.n9563 0.00263636
R30529 avss.n9539 avss.n9538 0.00263636
R30530 avss.n9418 avss.n9417 0.00263636
R30531 avss.n2138 avss.n2137 0.00263636
R30532 avss.n2067 avss.n2058 0.00263636
R30533 avss.n9450 avss.n9449 0.00263636
R30534 avss.n9453 avss.n9452 0.00263636
R30535 avss.n9519 avss.n9518 0.00263636
R30536 avss.n9840 avss.n9839 0.00263636
R30537 avss.n1775 avss.n1774 0.00263636
R30538 avss.n1794 avss.n1785 0.00263636
R30539 avss.n9782 avss.n9781 0.00263636
R30540 avss.n9785 avss.n9784 0.00263636
R30541 avss.n9760 avss.n9759 0.00263636
R30542 avss.n9639 avss.n9638 0.00263636
R30543 avss.n1922 avss.n1921 0.00263636
R30544 avss.n1851 avss.n1842 0.00263636
R30545 avss.n9671 avss.n9670 0.00263636
R30546 avss.n9674 avss.n9673 0.00263636
R30547 avss.n9740 avss.n9739 0.00263636
R30548 avss.n10061 avss.n10060 0.00263636
R30549 avss.n1559 avss.n1558 0.00263636
R30550 avss.n1578 avss.n1569 0.00263636
R30551 avss.n10003 avss.n10002 0.00263636
R30552 avss.n10006 avss.n10005 0.00263636
R30553 avss.n9981 avss.n9980 0.00263636
R30554 avss.n9860 avss.n9859 0.00263636
R30555 avss.n1706 avss.n1705 0.00263636
R30556 avss.n1635 avss.n1626 0.00263636
R30557 avss.n9892 avss.n9891 0.00263636
R30558 avss.n9895 avss.n9894 0.00263636
R30559 avss.n9961 avss.n9960 0.00263636
R30560 avss.n10282 avss.n10281 0.00263636
R30561 avss.n1343 avss.n1342 0.00263636
R30562 avss.n1362 avss.n1353 0.00263636
R30563 avss.n10224 avss.n10223 0.00263636
R30564 avss.n10227 avss.n10226 0.00263636
R30565 avss.n10202 avss.n10201 0.00263636
R30566 avss.n10081 avss.n10080 0.00263636
R30567 avss.n1490 avss.n1489 0.00263636
R30568 avss.n1419 avss.n1410 0.00263636
R30569 avss.n10113 avss.n10112 0.00263636
R30570 avss.n10116 avss.n10115 0.00263636
R30571 avss.n10182 avss.n10181 0.00263636
R30572 avss.n10503 avss.n10502 0.00263636
R30573 avss.n1127 avss.n1126 0.00263636
R30574 avss.n1146 avss.n1137 0.00263636
R30575 avss.n10445 avss.n10444 0.00263636
R30576 avss.n10448 avss.n10447 0.00263636
R30577 avss.n10423 avss.n10422 0.00263636
R30578 avss.n10302 avss.n10301 0.00263636
R30579 avss.n1274 avss.n1273 0.00263636
R30580 avss.n1203 avss.n1194 0.00263636
R30581 avss.n10334 avss.n10333 0.00263636
R30582 avss.n10337 avss.n10336 0.00263636
R30583 avss.n10403 avss.n10402 0.00263636
R30584 avss.n10724 avss.n10723 0.00263636
R30585 avss.n911 avss.n910 0.00263636
R30586 avss.n930 avss.n921 0.00263636
R30587 avss.n10666 avss.n10665 0.00263636
R30588 avss.n10669 avss.n10668 0.00263636
R30589 avss.n10644 avss.n10643 0.00263636
R30590 avss.n10523 avss.n10522 0.00263636
R30591 avss.n1058 avss.n1057 0.00263636
R30592 avss.n987 avss.n978 0.00263636
R30593 avss.n10555 avss.n10554 0.00263636
R30594 avss.n10558 avss.n10557 0.00263636
R30595 avss.n10624 avss.n10623 0.00263636
R30596 avss.n10945 avss.n10944 0.00263636
R30597 avss.n695 avss.n694 0.00263636
R30598 avss.n714 avss.n705 0.00263636
R30599 avss.n10887 avss.n10886 0.00263636
R30600 avss.n10890 avss.n10889 0.00263636
R30601 avss.n10865 avss.n10864 0.00263636
R30602 avss.n10744 avss.n10743 0.00263636
R30603 avss.n842 avss.n841 0.00263636
R30604 avss.n771 avss.n762 0.00263636
R30605 avss.n10776 avss.n10775 0.00263636
R30606 avss.n10779 avss.n10778 0.00263636
R30607 avss.n10845 avss.n10844 0.00263636
R30608 avss.n11166 avss.n11165 0.00263636
R30609 avss.n479 avss.n478 0.00263636
R30610 avss.n498 avss.n489 0.00263636
R30611 avss.n11108 avss.n11107 0.00263636
R30612 avss.n11111 avss.n11110 0.00263636
R30613 avss.n11086 avss.n11085 0.00263636
R30614 avss.n10965 avss.n10964 0.00263636
R30615 avss.n626 avss.n625 0.00263636
R30616 avss.n555 avss.n546 0.00263636
R30617 avss.n10997 avss.n10996 0.00263636
R30618 avss.n11000 avss.n10999 0.00263636
R30619 avss.n11066 avss.n11065 0.00263636
R30620 avss.n342 avss.n341 0.00263636
R30621 avss.n11398 avss.n11397 0.00263636
R30622 avss.n11327 avss.n11318 0.00263636
R30623 avss.n375 avss.n374 0.00263636
R30624 avss.n378 avss.n377 0.00263636
R30625 avss.n337 avss.n336 0.00263636
R30626 avss.n11186 avss.n11185 0.00263636
R30627 avss.n301 avss.n300 0.00263636
R30628 avss.n230 avss.n221 0.00263636
R30629 avss.n11218 avss.n11217 0.00263636
R30630 avss.n11221 avss.n11220 0.00263636
R30631 avss.n11287 avss.n11286 0.00263636
R30632 avss.n125 avss.n124 0.00263636
R30633 avss.n11619 avss.n11618 0.00263636
R30634 avss.n11548 avss.n11539 0.00263636
R30635 avss.n158 avss.n157 0.00263636
R30636 avss.n161 avss.n160 0.00263636
R30637 avss.n120 avss.n119 0.00263636
R30638 avss.n11407 avss.n11406 0.00263636
R30639 avss.n84 avss.n83 0.00263636
R30640 avss.n13 avss.n4 0.00263636
R30641 avss.n11439 avss.n11438 0.00263636
R30642 avss.n11442 avss.n11441 0.00263636
R30643 avss.n11508 avss.n11507 0.00263636
R30644 avss.n3352 avss.n3286 0.00258333
R30645 avss.n3456 avss.n3455 0.00258333
R30646 avss.n8769 avss.n8768 0.00239394
R30647 avss.n8737 avss.n8730 0.00239394
R30648 avss.n8672 avss.n8661 0.00239394
R30649 avss.n8659 avss.n8658 0.00239394
R30650 avss.n8851 avss.n3714 0.00239394
R30651 avss.n8873 avss.n8872 0.00239394
R30652 avss.n8940 avss.n3684 0.00239394
R30653 avss.n8946 avss.n8945 0.00239394
R30654 avss.n8416 avss.n8415 0.00239394
R30655 avss.n8384 avss.n8377 0.00239394
R30656 avss.n8319 avss.n8308 0.00239394
R30657 avss.n8306 avss.n8305 0.00239394
R30658 avss.n8498 avss.n3798 0.00239394
R30659 avss.n8520 avss.n8519 0.00239394
R30660 avss.n8587 avss.n3768 0.00239394
R30661 avss.n8593 avss.n8592 0.00239394
R30662 avss.n8063 avss.n8062 0.00239394
R30663 avss.n8031 avss.n8024 0.00239394
R30664 avss.n7966 avss.n7955 0.00239394
R30665 avss.n7953 avss.n7952 0.00239394
R30666 avss.n8145 avss.n3882 0.00239394
R30667 avss.n8167 avss.n8166 0.00239394
R30668 avss.n8234 avss.n3852 0.00239394
R30669 avss.n8240 avss.n8239 0.00239394
R30670 avss.n7710 avss.n7709 0.00239394
R30671 avss.n7678 avss.n7671 0.00239394
R30672 avss.n7613 avss.n7602 0.00239394
R30673 avss.n7600 avss.n7599 0.00239394
R30674 avss.n7792 avss.n3966 0.00239394
R30675 avss.n7814 avss.n7813 0.00239394
R30676 avss.n7881 avss.n3936 0.00239394
R30677 avss.n7887 avss.n7886 0.00239394
R30678 avss.n7357 avss.n7356 0.00239394
R30679 avss.n7325 avss.n7318 0.00239394
R30680 avss.n7260 avss.n7249 0.00239394
R30681 avss.n7247 avss.n7246 0.00239394
R30682 avss.n7439 avss.n4050 0.00239394
R30683 avss.n7461 avss.n7460 0.00239394
R30684 avss.n7528 avss.n4020 0.00239394
R30685 avss.n7534 avss.n7533 0.00239394
R30686 avss.n7004 avss.n7003 0.00239394
R30687 avss.n6972 avss.n6965 0.00239394
R30688 avss.n6907 avss.n6896 0.00239394
R30689 avss.n6894 avss.n6893 0.00239394
R30690 avss.n7086 avss.n4134 0.00239394
R30691 avss.n7108 avss.n7107 0.00239394
R30692 avss.n7175 avss.n4104 0.00239394
R30693 avss.n7181 avss.n7180 0.00239394
R30694 avss.n6651 avss.n6650 0.00239394
R30695 avss.n6619 avss.n6612 0.00239394
R30696 avss.n6554 avss.n6543 0.00239394
R30697 avss.n6541 avss.n6540 0.00239394
R30698 avss.n6733 avss.n4218 0.00239394
R30699 avss.n6755 avss.n6754 0.00239394
R30700 avss.n6822 avss.n4188 0.00239394
R30701 avss.n6828 avss.n6827 0.00239394
R30702 avss.n6298 avss.n6297 0.00239394
R30703 avss.n6266 avss.n6259 0.00239394
R30704 avss.n6201 avss.n6190 0.00239394
R30705 avss.n6188 avss.n6187 0.00239394
R30706 avss.n6380 avss.n4302 0.00239394
R30707 avss.n6402 avss.n6401 0.00239394
R30708 avss.n6469 avss.n4272 0.00239394
R30709 avss.n6475 avss.n6474 0.00239394
R30710 avss.n5945 avss.n5944 0.00239394
R30711 avss.n5913 avss.n5906 0.00239394
R30712 avss.n5848 avss.n5837 0.00239394
R30713 avss.n5835 avss.n5834 0.00239394
R30714 avss.n6027 avss.n4386 0.00239394
R30715 avss.n6049 avss.n6048 0.00239394
R30716 avss.n6116 avss.n4356 0.00239394
R30717 avss.n6122 avss.n6121 0.00239394
R30718 avss.n5592 avss.n5591 0.00239394
R30719 avss.n5560 avss.n5553 0.00239394
R30720 avss.n5495 avss.n5484 0.00239394
R30721 avss.n5482 avss.n5481 0.00239394
R30722 avss.n5674 avss.n4470 0.00239394
R30723 avss.n5696 avss.n5695 0.00239394
R30724 avss.n5763 avss.n4440 0.00239394
R30725 avss.n5769 avss.n5768 0.00239394
R30726 avss.n5249 avss.n5248 0.00239394
R30727 avss.n5220 avss.n5213 0.00239394
R30728 avss.n5149 avss.n5134 0.00239394
R30729 avss.n5294 avss.n5097 0.00239394
R30730 avss.n5321 avss.n4554 0.00239394
R30731 avss.n5343 avss.n5342 0.00239394
R30732 avss.n5410 avss.n4524 0.00239394
R30733 avss.n5416 avss.n5415 0.00239394
R30734 avss.n4895 avss.n4894 0.00239394
R30735 avss.n4866 avss.n4859 0.00239394
R30736 avss.n4795 avss.n4780 0.00239394
R30737 avss.n4940 avss.n4743 0.00239394
R30738 avss.n4967 avss.n4638 0.00239394
R30739 avss.n4989 avss.n4988 0.00239394
R30740 avss.n5056 avss.n4608 0.00239394
R30741 avss.n5062 avss.n5061 0.00239394
R30742 avss.n9113 avss.n9110 0.00239394
R30743 avss.n9167 avss.n9166 0.00239394
R30744 avss.n2456 avss.n2453 0.00239394
R30745 avss.n2475 avss.n2474 0.00239394
R30746 avss.n2532 avss.n2531 0.00239394
R30747 avss.n2513 avss.n2510 0.00239394
R30748 avss.n9056 avss.n9055 0.00239394
R30749 avss.n9001 avss.n8998 0.00239394
R30750 avss.n9334 avss.n9331 0.00239394
R30751 avss.n9388 avss.n9387 0.00239394
R30752 avss.n2240 avss.n2237 0.00239394
R30753 avss.n2259 avss.n2258 0.00239394
R30754 avss.n2316 avss.n2315 0.00239394
R30755 avss.n2297 avss.n2294 0.00239394
R30756 avss.n9277 avss.n9276 0.00239394
R30757 avss.n9222 avss.n9219 0.00239394
R30758 avss.n9555 avss.n9552 0.00239394
R30759 avss.n9609 avss.n9608 0.00239394
R30760 avss.n2024 avss.n2021 0.00239394
R30761 avss.n2043 avss.n2042 0.00239394
R30762 avss.n2100 avss.n2099 0.00239394
R30763 avss.n2081 avss.n2078 0.00239394
R30764 avss.n9498 avss.n9497 0.00239394
R30765 avss.n9443 avss.n9440 0.00239394
R30766 avss.n9776 avss.n9773 0.00239394
R30767 avss.n9830 avss.n9829 0.00239394
R30768 avss.n1808 avss.n1805 0.00239394
R30769 avss.n1827 avss.n1826 0.00239394
R30770 avss.n1884 avss.n1883 0.00239394
R30771 avss.n1865 avss.n1862 0.00239394
R30772 avss.n9719 avss.n9718 0.00239394
R30773 avss.n9664 avss.n9661 0.00239394
R30774 avss.n9997 avss.n9994 0.00239394
R30775 avss.n10051 avss.n10050 0.00239394
R30776 avss.n1592 avss.n1589 0.00239394
R30777 avss.n1611 avss.n1610 0.00239394
R30778 avss.n1668 avss.n1667 0.00239394
R30779 avss.n1649 avss.n1646 0.00239394
R30780 avss.n9940 avss.n9939 0.00239394
R30781 avss.n9885 avss.n9882 0.00239394
R30782 avss.n10218 avss.n10215 0.00239394
R30783 avss.n10272 avss.n10271 0.00239394
R30784 avss.n1376 avss.n1373 0.00239394
R30785 avss.n1395 avss.n1394 0.00239394
R30786 avss.n1452 avss.n1451 0.00239394
R30787 avss.n1433 avss.n1430 0.00239394
R30788 avss.n10161 avss.n10160 0.00239394
R30789 avss.n10106 avss.n10103 0.00239394
R30790 avss.n10439 avss.n10436 0.00239394
R30791 avss.n10493 avss.n10492 0.00239394
R30792 avss.n1160 avss.n1157 0.00239394
R30793 avss.n1179 avss.n1178 0.00239394
R30794 avss.n1236 avss.n1235 0.00239394
R30795 avss.n1217 avss.n1214 0.00239394
R30796 avss.n10382 avss.n10381 0.00239394
R30797 avss.n10327 avss.n10324 0.00239394
R30798 avss.n10660 avss.n10657 0.00239394
R30799 avss.n10714 avss.n10713 0.00239394
R30800 avss.n944 avss.n941 0.00239394
R30801 avss.n963 avss.n962 0.00239394
R30802 avss.n1020 avss.n1019 0.00239394
R30803 avss.n1001 avss.n998 0.00239394
R30804 avss.n10603 avss.n10602 0.00239394
R30805 avss.n10548 avss.n10545 0.00239394
R30806 avss.n10881 avss.n10878 0.00239394
R30807 avss.n10935 avss.n10934 0.00239394
R30808 avss.n728 avss.n725 0.00239394
R30809 avss.n747 avss.n746 0.00239394
R30810 avss.n804 avss.n803 0.00239394
R30811 avss.n785 avss.n782 0.00239394
R30812 avss.n10824 avss.n10823 0.00239394
R30813 avss.n10769 avss.n10766 0.00239394
R30814 avss.n11102 avss.n11099 0.00239394
R30815 avss.n11156 avss.n11155 0.00239394
R30816 avss.n512 avss.n509 0.00239394
R30817 avss.n531 avss.n530 0.00239394
R30818 avss.n588 avss.n587 0.00239394
R30819 avss.n569 avss.n566 0.00239394
R30820 avss.n11045 avss.n11044 0.00239394
R30821 avss.n10990 avss.n10987 0.00239394
R30822 avss.n368 avss.n365 0.00239394
R30823 avss.n423 avss.n422 0.00239394
R30824 avss.n11341 avss.n11338 0.00239394
R30825 avss.n11360 avss.n11359 0.00239394
R30826 avss.n263 avss.n262 0.00239394
R30827 avss.n244 avss.n241 0.00239394
R30828 avss.n11266 avss.n11265 0.00239394
R30829 avss.n11211 avss.n11208 0.00239394
R30830 avss.n151 avss.n148 0.00239394
R30831 avss.n206 avss.n205 0.00239394
R30832 avss.n11562 avss.n11559 0.00239394
R30833 avss.n11581 avss.n11580 0.00239394
R30834 avss.n46 avss.n45 0.00239394
R30835 avss.n27 avss.n24 0.00239394
R30836 avss.n11487 avss.n11486 0.00239394
R30837 avss.n11432 avss.n11429 0.00239394
R30838 avss.n2963 avss.n2960 0.00230459
R30839 avss.n3020 avss.n2944 0.00230459
R30840 avss.n3134 avss.n2927 0.00230459
R30841 avss.n2611 avss.n2610 0.00230459
R30842 avss.n11628 avss.n11627 0.00200055
R30843 avss.n8827 avss.n8628 0.00192424
R30844 avss.n8826 avss.n8621 0.00192424
R30845 avss.n8787 avss.n8786 0.00192424
R30846 avss.n8782 avss.n8717 0.00192424
R30847 avss.n8760 avss.n8759 0.00192424
R30848 avss.n3747 avss.n3728 0.00192424
R30849 avss.n8845 avss.n3722 0.00192424
R30850 avss.n8916 avss.n3691 0.00192424
R30851 avss.n8929 avss.n3687 0.00192424
R30852 avss.n8964 avss.n3681 0.00192424
R30853 avss.n8474 avss.n8275 0.00192424
R30854 avss.n8473 avss.n8268 0.00192424
R30855 avss.n8434 avss.n8433 0.00192424
R30856 avss.n8429 avss.n8364 0.00192424
R30857 avss.n8407 avss.n8406 0.00192424
R30858 avss.n3831 avss.n3812 0.00192424
R30859 avss.n8492 avss.n3806 0.00192424
R30860 avss.n8563 avss.n3775 0.00192424
R30861 avss.n8576 avss.n3771 0.00192424
R30862 avss.n8611 avss.n3765 0.00192424
R30863 avss.n8121 avss.n7922 0.00192424
R30864 avss.n8120 avss.n7915 0.00192424
R30865 avss.n8081 avss.n8080 0.00192424
R30866 avss.n8076 avss.n8011 0.00192424
R30867 avss.n8054 avss.n8053 0.00192424
R30868 avss.n3915 avss.n3896 0.00192424
R30869 avss.n8139 avss.n3890 0.00192424
R30870 avss.n8210 avss.n3859 0.00192424
R30871 avss.n8223 avss.n3855 0.00192424
R30872 avss.n8258 avss.n3849 0.00192424
R30873 avss.n7768 avss.n7569 0.00192424
R30874 avss.n7767 avss.n7562 0.00192424
R30875 avss.n7728 avss.n7727 0.00192424
R30876 avss.n7723 avss.n7658 0.00192424
R30877 avss.n7701 avss.n7700 0.00192424
R30878 avss.n3999 avss.n3980 0.00192424
R30879 avss.n7786 avss.n3974 0.00192424
R30880 avss.n7857 avss.n3943 0.00192424
R30881 avss.n7870 avss.n3939 0.00192424
R30882 avss.n7905 avss.n3933 0.00192424
R30883 avss.n7415 avss.n7216 0.00192424
R30884 avss.n7414 avss.n7209 0.00192424
R30885 avss.n7375 avss.n7374 0.00192424
R30886 avss.n7370 avss.n7305 0.00192424
R30887 avss.n7348 avss.n7347 0.00192424
R30888 avss.n4083 avss.n4064 0.00192424
R30889 avss.n7433 avss.n4058 0.00192424
R30890 avss.n7504 avss.n4027 0.00192424
R30891 avss.n7517 avss.n4023 0.00192424
R30892 avss.n7552 avss.n4017 0.00192424
R30893 avss.n7062 avss.n6863 0.00192424
R30894 avss.n7061 avss.n6856 0.00192424
R30895 avss.n7022 avss.n7021 0.00192424
R30896 avss.n7017 avss.n6952 0.00192424
R30897 avss.n6995 avss.n6994 0.00192424
R30898 avss.n4167 avss.n4148 0.00192424
R30899 avss.n7080 avss.n4142 0.00192424
R30900 avss.n7151 avss.n4111 0.00192424
R30901 avss.n7164 avss.n4107 0.00192424
R30902 avss.n7199 avss.n4101 0.00192424
R30903 avss.n6709 avss.n6510 0.00192424
R30904 avss.n6708 avss.n6503 0.00192424
R30905 avss.n6669 avss.n6668 0.00192424
R30906 avss.n6664 avss.n6599 0.00192424
R30907 avss.n6642 avss.n6641 0.00192424
R30908 avss.n4251 avss.n4232 0.00192424
R30909 avss.n6727 avss.n4226 0.00192424
R30910 avss.n6798 avss.n4195 0.00192424
R30911 avss.n6811 avss.n4191 0.00192424
R30912 avss.n6846 avss.n4185 0.00192424
R30913 avss.n6356 avss.n6157 0.00192424
R30914 avss.n6355 avss.n6150 0.00192424
R30915 avss.n6316 avss.n6315 0.00192424
R30916 avss.n6311 avss.n6246 0.00192424
R30917 avss.n6289 avss.n6288 0.00192424
R30918 avss.n4335 avss.n4316 0.00192424
R30919 avss.n6374 avss.n4310 0.00192424
R30920 avss.n6445 avss.n4279 0.00192424
R30921 avss.n6458 avss.n4275 0.00192424
R30922 avss.n6493 avss.n4269 0.00192424
R30923 avss.n6003 avss.n5804 0.00192424
R30924 avss.n6002 avss.n5797 0.00192424
R30925 avss.n5963 avss.n5962 0.00192424
R30926 avss.n5958 avss.n5893 0.00192424
R30927 avss.n5936 avss.n5935 0.00192424
R30928 avss.n4419 avss.n4400 0.00192424
R30929 avss.n6021 avss.n4394 0.00192424
R30930 avss.n6092 avss.n4363 0.00192424
R30931 avss.n6105 avss.n4359 0.00192424
R30932 avss.n6140 avss.n4353 0.00192424
R30933 avss.n5650 avss.n5451 0.00192424
R30934 avss.n5649 avss.n5444 0.00192424
R30935 avss.n5610 avss.n5609 0.00192424
R30936 avss.n5605 avss.n5540 0.00192424
R30937 avss.n5583 avss.n5582 0.00192424
R30938 avss.n4503 avss.n4484 0.00192424
R30939 avss.n5668 avss.n4478 0.00192424
R30940 avss.n5739 avss.n4447 0.00192424
R30941 avss.n5752 avss.n4443 0.00192424
R30942 avss.n5787 avss.n4437 0.00192424
R30943 avss.n5126 avss.n5125 0.00192424
R30944 avss.n5127 avss.n5091 0.00192424
R30945 avss.n5265 avss.n5264 0.00192424
R30946 avss.n5260 avss.n5194 0.00192424
R30947 avss.n5242 avss.n5241 0.00192424
R30948 avss.n4587 avss.n4568 0.00192424
R30949 avss.n5315 avss.n4562 0.00192424
R30950 avss.n5386 avss.n4531 0.00192424
R30951 avss.n5399 avss.n4527 0.00192424
R30952 avss.n5434 avss.n4521 0.00192424
R30953 avss.n4772 avss.n4771 0.00192424
R30954 avss.n4773 avss.n4737 0.00192424
R30955 avss.n4911 avss.n4910 0.00192424
R30956 avss.n4906 avss.n4840 0.00192424
R30957 avss.n4888 avss.n4887 0.00192424
R30958 avss.n4671 avss.n4652 0.00192424
R30959 avss.n4961 avss.n4646 0.00192424
R30960 avss.n5032 avss.n4615 0.00192424
R30961 avss.n5045 avss.n4611 0.00192424
R30962 avss.n5080 avss.n4605 0.00192424
R30963 avss.n2406 avss.n2397 0.00192424
R30964 avss.n2396 avss.n2395 0.00192424
R30965 avss.n9150 avss.n9149 0.00192424
R30966 avss.n9152 avss.n9151 0.00192424
R30967 avss.n9088 avss.n9087 0.00192424
R30968 avss.n2553 avss.n2544 0.00192424
R30969 avss.n2543 avss.n2542 0.00192424
R30970 avss.n9039 avss.n9038 0.00192424
R30971 avss.n9041 avss.n9040 0.00192424
R30972 avss.n9068 avss.n9067 0.00192424
R30973 avss.n2190 avss.n2181 0.00192424
R30974 avss.n2180 avss.n2179 0.00192424
R30975 avss.n9371 avss.n9370 0.00192424
R30976 avss.n9373 avss.n9372 0.00192424
R30977 avss.n9309 avss.n9308 0.00192424
R30978 avss.n2337 avss.n2328 0.00192424
R30979 avss.n2327 avss.n2326 0.00192424
R30980 avss.n9260 avss.n9259 0.00192424
R30981 avss.n9262 avss.n9261 0.00192424
R30982 avss.n9289 avss.n9288 0.00192424
R30983 avss.n1974 avss.n1965 0.00192424
R30984 avss.n1964 avss.n1963 0.00192424
R30985 avss.n9592 avss.n9591 0.00192424
R30986 avss.n9594 avss.n9593 0.00192424
R30987 avss.n9530 avss.n9529 0.00192424
R30988 avss.n2121 avss.n2112 0.00192424
R30989 avss.n2111 avss.n2110 0.00192424
R30990 avss.n9481 avss.n9480 0.00192424
R30991 avss.n9483 avss.n9482 0.00192424
R30992 avss.n9510 avss.n9509 0.00192424
R30993 avss.n1758 avss.n1749 0.00192424
R30994 avss.n1748 avss.n1747 0.00192424
R30995 avss.n9813 avss.n9812 0.00192424
R30996 avss.n9815 avss.n9814 0.00192424
R30997 avss.n9751 avss.n9750 0.00192424
R30998 avss.n1905 avss.n1896 0.00192424
R30999 avss.n1895 avss.n1894 0.00192424
R31000 avss.n9702 avss.n9701 0.00192424
R31001 avss.n9704 avss.n9703 0.00192424
R31002 avss.n9731 avss.n9730 0.00192424
R31003 avss.n1542 avss.n1533 0.00192424
R31004 avss.n1532 avss.n1531 0.00192424
R31005 avss.n10034 avss.n10033 0.00192424
R31006 avss.n10036 avss.n10035 0.00192424
R31007 avss.n9972 avss.n9971 0.00192424
R31008 avss.n1689 avss.n1680 0.00192424
R31009 avss.n1679 avss.n1678 0.00192424
R31010 avss.n9923 avss.n9922 0.00192424
R31011 avss.n9925 avss.n9924 0.00192424
R31012 avss.n9952 avss.n9951 0.00192424
R31013 avss.n1326 avss.n1317 0.00192424
R31014 avss.n1316 avss.n1315 0.00192424
R31015 avss.n10255 avss.n10254 0.00192424
R31016 avss.n10257 avss.n10256 0.00192424
R31017 avss.n10193 avss.n10192 0.00192424
R31018 avss.n1473 avss.n1464 0.00192424
R31019 avss.n1463 avss.n1462 0.00192424
R31020 avss.n10144 avss.n10143 0.00192424
R31021 avss.n10146 avss.n10145 0.00192424
R31022 avss.n10173 avss.n10172 0.00192424
R31023 avss.n1110 avss.n1101 0.00192424
R31024 avss.n1100 avss.n1099 0.00192424
R31025 avss.n10476 avss.n10475 0.00192424
R31026 avss.n10478 avss.n10477 0.00192424
R31027 avss.n10414 avss.n10413 0.00192424
R31028 avss.n1257 avss.n1248 0.00192424
R31029 avss.n1247 avss.n1246 0.00192424
R31030 avss.n10365 avss.n10364 0.00192424
R31031 avss.n10367 avss.n10366 0.00192424
R31032 avss.n10394 avss.n10393 0.00192424
R31033 avss.n894 avss.n885 0.00192424
R31034 avss.n884 avss.n883 0.00192424
R31035 avss.n10697 avss.n10696 0.00192424
R31036 avss.n10699 avss.n10698 0.00192424
R31037 avss.n10635 avss.n10634 0.00192424
R31038 avss.n1041 avss.n1032 0.00192424
R31039 avss.n1031 avss.n1030 0.00192424
R31040 avss.n10586 avss.n10585 0.00192424
R31041 avss.n10588 avss.n10587 0.00192424
R31042 avss.n10615 avss.n10614 0.00192424
R31043 avss.n678 avss.n669 0.00192424
R31044 avss.n668 avss.n667 0.00192424
R31045 avss.n10918 avss.n10917 0.00192424
R31046 avss.n10920 avss.n10919 0.00192424
R31047 avss.n10856 avss.n10855 0.00192424
R31048 avss.n825 avss.n816 0.00192424
R31049 avss.n815 avss.n814 0.00192424
R31050 avss.n10807 avss.n10806 0.00192424
R31051 avss.n10809 avss.n10808 0.00192424
R31052 avss.n10836 avss.n10835 0.00192424
R31053 avss.n462 avss.n453 0.00192424
R31054 avss.n452 avss.n451 0.00192424
R31055 avss.n11139 avss.n11138 0.00192424
R31056 avss.n11141 avss.n11140 0.00192424
R31057 avss.n11077 avss.n11076 0.00192424
R31058 avss.n609 avss.n600 0.00192424
R31059 avss.n599 avss.n598 0.00192424
R31060 avss.n11028 avss.n11027 0.00192424
R31061 avss.n11030 avss.n11029 0.00192424
R31062 avss.n11057 avss.n11056 0.00192424
R31063 avss.n11380 avss.n11371 0.00192424
R31064 avss.n11370 avss.n11369 0.00192424
R31065 avss.n406 avss.n405 0.00192424
R31066 avss.n408 avss.n407 0.00192424
R31067 avss.n328 avss.n327 0.00192424
R31068 avss.n284 avss.n275 0.00192424
R31069 avss.n274 avss.n273 0.00192424
R31070 avss.n11249 avss.n11248 0.00192424
R31071 avss.n11251 avss.n11250 0.00192424
R31072 avss.n11278 avss.n11277 0.00192424
R31073 avss.n11601 avss.n11592 0.00192424
R31074 avss.n11591 avss.n11590 0.00192424
R31075 avss.n189 avss.n188 0.00192424
R31076 avss.n191 avss.n190 0.00192424
R31077 avss.n111 avss.n110 0.00192424
R31078 avss.n67 avss.n58 0.00192424
R31079 avss.n57 avss.n56 0.00192424
R31080 avss.n11470 avss.n11469 0.00192424
R31081 avss.n11472 avss.n11471 0.00192424
R31082 avss.n11499 avss.n11498 0.00192424
R31083 avss.n11631 avss.n11628 0.00148276
R31084 avss.n8832 avss.n8624 0.00121212
R31085 avss.n8664 avss.n8653 0.00121212
R31086 avss.n8657 avss.n8654 0.00121212
R31087 avss.n8665 avss.n8655 0.00121212
R31088 avss.n8673 avss.n8663 0.00121212
R31089 avss.n8739 avss.n8738 0.00121212
R31090 avss.n8767 avss.n8727 0.00121212
R31091 avss.n8843 avss.n8842 0.00121212
R31092 avss.n8863 avss.n8862 0.00121212
R31093 avss.n8850 avss.n3715 0.00121212
R31094 avss.n8861 avss.n3716 0.00121212
R31095 avss.n8874 avss.n3709 0.00121212
R31096 avss.n8939 avss.n8938 0.00121212
R31097 avss.n8947 avss.n3672 0.00121212
R31098 avss.n8479 avss.n8271 0.00121212
R31099 avss.n8311 avss.n8300 0.00121212
R31100 avss.n8304 avss.n8301 0.00121212
R31101 avss.n8312 avss.n8302 0.00121212
R31102 avss.n8320 avss.n8310 0.00121212
R31103 avss.n8386 avss.n8385 0.00121212
R31104 avss.n8414 avss.n8374 0.00121212
R31105 avss.n8490 avss.n8489 0.00121212
R31106 avss.n8510 avss.n8509 0.00121212
R31107 avss.n8497 avss.n3799 0.00121212
R31108 avss.n8508 avss.n3800 0.00121212
R31109 avss.n8521 avss.n3793 0.00121212
R31110 avss.n8586 avss.n8585 0.00121212
R31111 avss.n8594 avss.n3756 0.00121212
R31112 avss.n8126 avss.n7918 0.00121212
R31113 avss.n7958 avss.n7947 0.00121212
R31114 avss.n7951 avss.n7948 0.00121212
R31115 avss.n7959 avss.n7949 0.00121212
R31116 avss.n7967 avss.n7957 0.00121212
R31117 avss.n8033 avss.n8032 0.00121212
R31118 avss.n8061 avss.n8021 0.00121212
R31119 avss.n8137 avss.n8136 0.00121212
R31120 avss.n8157 avss.n8156 0.00121212
R31121 avss.n8144 avss.n3883 0.00121212
R31122 avss.n8155 avss.n3884 0.00121212
R31123 avss.n8168 avss.n3877 0.00121212
R31124 avss.n8233 avss.n8232 0.00121212
R31125 avss.n8241 avss.n3840 0.00121212
R31126 avss.n7773 avss.n7565 0.00121212
R31127 avss.n7605 avss.n7594 0.00121212
R31128 avss.n7598 avss.n7595 0.00121212
R31129 avss.n7606 avss.n7596 0.00121212
R31130 avss.n7614 avss.n7604 0.00121212
R31131 avss.n7680 avss.n7679 0.00121212
R31132 avss.n7708 avss.n7668 0.00121212
R31133 avss.n7784 avss.n7783 0.00121212
R31134 avss.n7804 avss.n7803 0.00121212
R31135 avss.n7791 avss.n3967 0.00121212
R31136 avss.n7802 avss.n3968 0.00121212
R31137 avss.n7815 avss.n3961 0.00121212
R31138 avss.n7880 avss.n7879 0.00121212
R31139 avss.n7888 avss.n3924 0.00121212
R31140 avss.n7420 avss.n7212 0.00121212
R31141 avss.n7252 avss.n7241 0.00121212
R31142 avss.n7245 avss.n7242 0.00121212
R31143 avss.n7253 avss.n7243 0.00121212
R31144 avss.n7261 avss.n7251 0.00121212
R31145 avss.n7327 avss.n7326 0.00121212
R31146 avss.n7355 avss.n7315 0.00121212
R31147 avss.n7431 avss.n7430 0.00121212
R31148 avss.n7451 avss.n7450 0.00121212
R31149 avss.n7438 avss.n4051 0.00121212
R31150 avss.n7449 avss.n4052 0.00121212
R31151 avss.n7462 avss.n4045 0.00121212
R31152 avss.n7527 avss.n7526 0.00121212
R31153 avss.n7535 avss.n4008 0.00121212
R31154 avss.n7067 avss.n6859 0.00121212
R31155 avss.n6899 avss.n6888 0.00121212
R31156 avss.n6892 avss.n6889 0.00121212
R31157 avss.n6900 avss.n6890 0.00121212
R31158 avss.n6908 avss.n6898 0.00121212
R31159 avss.n6974 avss.n6973 0.00121212
R31160 avss.n7002 avss.n6962 0.00121212
R31161 avss.n7078 avss.n7077 0.00121212
R31162 avss.n7098 avss.n7097 0.00121212
R31163 avss.n7085 avss.n4135 0.00121212
R31164 avss.n7096 avss.n4136 0.00121212
R31165 avss.n7109 avss.n4129 0.00121212
R31166 avss.n7174 avss.n7173 0.00121212
R31167 avss.n7182 avss.n4092 0.00121212
R31168 avss.n6714 avss.n6506 0.00121212
R31169 avss.n6546 avss.n6535 0.00121212
R31170 avss.n6539 avss.n6536 0.00121212
R31171 avss.n6547 avss.n6537 0.00121212
R31172 avss.n6555 avss.n6545 0.00121212
R31173 avss.n6621 avss.n6620 0.00121212
R31174 avss.n6649 avss.n6609 0.00121212
R31175 avss.n6725 avss.n6724 0.00121212
R31176 avss.n6745 avss.n6744 0.00121212
R31177 avss.n6732 avss.n4219 0.00121212
R31178 avss.n6743 avss.n4220 0.00121212
R31179 avss.n6756 avss.n4213 0.00121212
R31180 avss.n6821 avss.n6820 0.00121212
R31181 avss.n6829 avss.n4176 0.00121212
R31182 avss.n6361 avss.n6153 0.00121212
R31183 avss.n6193 avss.n6182 0.00121212
R31184 avss.n6186 avss.n6183 0.00121212
R31185 avss.n6194 avss.n6184 0.00121212
R31186 avss.n6202 avss.n6192 0.00121212
R31187 avss.n6268 avss.n6267 0.00121212
R31188 avss.n6296 avss.n6256 0.00121212
R31189 avss.n6372 avss.n6371 0.00121212
R31190 avss.n6392 avss.n6391 0.00121212
R31191 avss.n6379 avss.n4303 0.00121212
R31192 avss.n6390 avss.n4304 0.00121212
R31193 avss.n6403 avss.n4297 0.00121212
R31194 avss.n6468 avss.n6467 0.00121212
R31195 avss.n6476 avss.n4260 0.00121212
R31196 avss.n6008 avss.n5800 0.00121212
R31197 avss.n5840 avss.n5829 0.00121212
R31198 avss.n5833 avss.n5830 0.00121212
R31199 avss.n5841 avss.n5831 0.00121212
R31200 avss.n5849 avss.n5839 0.00121212
R31201 avss.n5915 avss.n5914 0.00121212
R31202 avss.n5943 avss.n5903 0.00121212
R31203 avss.n6019 avss.n6018 0.00121212
R31204 avss.n6039 avss.n6038 0.00121212
R31205 avss.n6026 avss.n4387 0.00121212
R31206 avss.n6037 avss.n4388 0.00121212
R31207 avss.n6050 avss.n4381 0.00121212
R31208 avss.n6115 avss.n6114 0.00121212
R31209 avss.n6123 avss.n4344 0.00121212
R31210 avss.n5655 avss.n5447 0.00121212
R31211 avss.n5487 avss.n5476 0.00121212
R31212 avss.n5480 avss.n5477 0.00121212
R31213 avss.n5488 avss.n5478 0.00121212
R31214 avss.n5496 avss.n5486 0.00121212
R31215 avss.n5562 avss.n5561 0.00121212
R31216 avss.n5590 avss.n5550 0.00121212
R31217 avss.n5666 avss.n5665 0.00121212
R31218 avss.n5686 avss.n5685 0.00121212
R31219 avss.n5673 avss.n4471 0.00121212
R31220 avss.n5684 avss.n4472 0.00121212
R31221 avss.n5697 avss.n4465 0.00121212
R31222 avss.n5762 avss.n5761 0.00121212
R31223 avss.n5770 avss.n4428 0.00121212
R31224 avss.n5300 avss.n5089 0.00121212
R31225 avss.n5140 avss.n5137 0.00121212
R31226 avss.n5138 avss.n5098 0.00121212
R31227 avss.n5142 avss.n5141 0.00121212
R31228 avss.n5150 avss.n5136 0.00121212
R31229 avss.n5222 avss.n5221 0.00121212
R31230 avss.n5250 avss.n5207 0.00121212
R31231 avss.n5313 avss.n5312 0.00121212
R31232 avss.n5333 avss.n5332 0.00121212
R31233 avss.n5320 avss.n4555 0.00121212
R31234 avss.n5331 avss.n4556 0.00121212
R31235 avss.n5344 avss.n4549 0.00121212
R31236 avss.n5409 avss.n5408 0.00121212
R31237 avss.n5417 avss.n4512 0.00121212
R31238 avss.n4946 avss.n4735 0.00121212
R31239 avss.n4786 avss.n4783 0.00121212
R31240 avss.n4784 avss.n4744 0.00121212
R31241 avss.n4788 avss.n4787 0.00121212
R31242 avss.n4796 avss.n4782 0.00121212
R31243 avss.n4868 avss.n4867 0.00121212
R31244 avss.n4896 avss.n4853 0.00121212
R31245 avss.n4959 avss.n4958 0.00121212
R31246 avss.n4979 avss.n4978 0.00121212
R31247 avss.n4966 avss.n4639 0.00121212
R31248 avss.n4977 avss.n4640 0.00121212
R31249 avss.n4990 avss.n4633 0.00121212
R31250 avss.n5055 avss.n5054 0.00121212
R31251 avss.n5063 avss.n4596 0.00121212
R31252 avss.n2483 avss.n2393 0.00121212
R31253 avss.n2389 avss.n2388 0.00121212
R31254 avss.n2467 avss.n2466 0.00121212
R31255 avss.n2464 avss.n2463 0.00121212
R31256 avss.n2458 avss.n2457 0.00121212
R31257 avss.n9171 avss.n9170 0.00121212
R31258 avss.n9115 avss.n9114 0.00121212
R31259 avss.n2592 avss.n2591 0.00121212
R31260 avss.n2587 avss.n2586 0.00121212
R31261 avss.n2524 avss.n2523 0.00121212
R31262 avss.n2521 avss.n2520 0.00121212
R31263 avss.n2515 avss.n2514 0.00121212
R31264 avss.n9060 avss.n9059 0.00121212
R31265 avss.n9003 avss.n9002 0.00121212
R31266 avss.n2267 avss.n2177 0.00121212
R31267 avss.n2173 avss.n2172 0.00121212
R31268 avss.n2251 avss.n2250 0.00121212
R31269 avss.n2248 avss.n2247 0.00121212
R31270 avss.n2242 avss.n2241 0.00121212
R31271 avss.n9392 avss.n9391 0.00121212
R31272 avss.n9336 avss.n9335 0.00121212
R31273 avss.n2376 avss.n2375 0.00121212
R31274 avss.n2371 avss.n2370 0.00121212
R31275 avss.n2308 avss.n2307 0.00121212
R31276 avss.n2305 avss.n2304 0.00121212
R31277 avss.n2299 avss.n2298 0.00121212
R31278 avss.n9281 avss.n9280 0.00121212
R31279 avss.n9224 avss.n9223 0.00121212
R31280 avss.n2051 avss.n1961 0.00121212
R31281 avss.n1957 avss.n1956 0.00121212
R31282 avss.n2035 avss.n2034 0.00121212
R31283 avss.n2032 avss.n2031 0.00121212
R31284 avss.n2026 avss.n2025 0.00121212
R31285 avss.n9613 avss.n9612 0.00121212
R31286 avss.n9557 avss.n9556 0.00121212
R31287 avss.n2160 avss.n2159 0.00121212
R31288 avss.n2155 avss.n2154 0.00121212
R31289 avss.n2092 avss.n2091 0.00121212
R31290 avss.n2089 avss.n2088 0.00121212
R31291 avss.n2083 avss.n2082 0.00121212
R31292 avss.n9502 avss.n9501 0.00121212
R31293 avss.n9445 avss.n9444 0.00121212
R31294 avss.n1835 avss.n1745 0.00121212
R31295 avss.n1741 avss.n1740 0.00121212
R31296 avss.n1819 avss.n1818 0.00121212
R31297 avss.n1816 avss.n1815 0.00121212
R31298 avss.n1810 avss.n1809 0.00121212
R31299 avss.n9834 avss.n9833 0.00121212
R31300 avss.n9778 avss.n9777 0.00121212
R31301 avss.n1944 avss.n1943 0.00121212
R31302 avss.n1939 avss.n1938 0.00121212
R31303 avss.n1876 avss.n1875 0.00121212
R31304 avss.n1873 avss.n1872 0.00121212
R31305 avss.n1867 avss.n1866 0.00121212
R31306 avss.n9723 avss.n9722 0.00121212
R31307 avss.n9666 avss.n9665 0.00121212
R31308 avss.n1619 avss.n1529 0.00121212
R31309 avss.n1525 avss.n1524 0.00121212
R31310 avss.n1603 avss.n1602 0.00121212
R31311 avss.n1600 avss.n1599 0.00121212
R31312 avss.n1594 avss.n1593 0.00121212
R31313 avss.n10055 avss.n10054 0.00121212
R31314 avss.n9999 avss.n9998 0.00121212
R31315 avss.n1728 avss.n1727 0.00121212
R31316 avss.n1723 avss.n1722 0.00121212
R31317 avss.n1660 avss.n1659 0.00121212
R31318 avss.n1657 avss.n1656 0.00121212
R31319 avss.n1651 avss.n1650 0.00121212
R31320 avss.n9944 avss.n9943 0.00121212
R31321 avss.n9887 avss.n9886 0.00121212
R31322 avss.n1403 avss.n1313 0.00121212
R31323 avss.n1309 avss.n1308 0.00121212
R31324 avss.n1387 avss.n1386 0.00121212
R31325 avss.n1384 avss.n1383 0.00121212
R31326 avss.n1378 avss.n1377 0.00121212
R31327 avss.n10276 avss.n10275 0.00121212
R31328 avss.n10220 avss.n10219 0.00121212
R31329 avss.n1512 avss.n1511 0.00121212
R31330 avss.n1507 avss.n1506 0.00121212
R31331 avss.n1444 avss.n1443 0.00121212
R31332 avss.n1441 avss.n1440 0.00121212
R31333 avss.n1435 avss.n1434 0.00121212
R31334 avss.n10165 avss.n10164 0.00121212
R31335 avss.n10108 avss.n10107 0.00121212
R31336 avss.n1187 avss.n1097 0.00121212
R31337 avss.n1093 avss.n1092 0.00121212
R31338 avss.n1171 avss.n1170 0.00121212
R31339 avss.n1168 avss.n1167 0.00121212
R31340 avss.n1162 avss.n1161 0.00121212
R31341 avss.n10497 avss.n10496 0.00121212
R31342 avss.n10441 avss.n10440 0.00121212
R31343 avss.n1296 avss.n1295 0.00121212
R31344 avss.n1291 avss.n1290 0.00121212
R31345 avss.n1228 avss.n1227 0.00121212
R31346 avss.n1225 avss.n1224 0.00121212
R31347 avss.n1219 avss.n1218 0.00121212
R31348 avss.n10386 avss.n10385 0.00121212
R31349 avss.n10329 avss.n10328 0.00121212
R31350 avss.n971 avss.n881 0.00121212
R31351 avss.n877 avss.n876 0.00121212
R31352 avss.n955 avss.n954 0.00121212
R31353 avss.n952 avss.n951 0.00121212
R31354 avss.n946 avss.n945 0.00121212
R31355 avss.n10718 avss.n10717 0.00121212
R31356 avss.n10662 avss.n10661 0.00121212
R31357 avss.n1080 avss.n1079 0.00121212
R31358 avss.n1075 avss.n1074 0.00121212
R31359 avss.n1012 avss.n1011 0.00121212
R31360 avss.n1009 avss.n1008 0.00121212
R31361 avss.n1003 avss.n1002 0.00121212
R31362 avss.n10607 avss.n10606 0.00121212
R31363 avss.n10550 avss.n10549 0.00121212
R31364 avss.n755 avss.n665 0.00121212
R31365 avss.n661 avss.n660 0.00121212
R31366 avss.n739 avss.n738 0.00121212
R31367 avss.n736 avss.n735 0.00121212
R31368 avss.n730 avss.n729 0.00121212
R31369 avss.n10939 avss.n10938 0.00121212
R31370 avss.n10883 avss.n10882 0.00121212
R31371 avss.n864 avss.n863 0.00121212
R31372 avss.n859 avss.n858 0.00121212
R31373 avss.n796 avss.n795 0.00121212
R31374 avss.n793 avss.n792 0.00121212
R31375 avss.n787 avss.n786 0.00121212
R31376 avss.n10828 avss.n10827 0.00121212
R31377 avss.n10771 avss.n10770 0.00121212
R31378 avss.n539 avss.n449 0.00121212
R31379 avss.n445 avss.n444 0.00121212
R31380 avss.n523 avss.n522 0.00121212
R31381 avss.n520 avss.n519 0.00121212
R31382 avss.n514 avss.n513 0.00121212
R31383 avss.n11160 avss.n11159 0.00121212
R31384 avss.n11104 avss.n11103 0.00121212
R31385 avss.n648 avss.n647 0.00121212
R31386 avss.n643 avss.n642 0.00121212
R31387 avss.n580 avss.n579 0.00121212
R31388 avss.n577 avss.n576 0.00121212
R31389 avss.n571 avss.n570 0.00121212
R31390 avss.n11049 avss.n11048 0.00121212
R31391 avss.n10992 avss.n10991 0.00121212
R31392 avss.n11403 avss.n11312 0.00121212
R31393 avss.n11308 avss.n11307 0.00121212
R31394 avss.n11352 avss.n11351 0.00121212
R31395 avss.n11349 avss.n11348 0.00121212
R31396 avss.n11343 avss.n11342 0.00121212
R31397 avss.n427 avss.n426 0.00121212
R31398 avss.n370 avss.n369 0.00121212
R31399 avss.n323 avss.n322 0.00121212
R31400 avss.n318 avss.n317 0.00121212
R31401 avss.n255 avss.n254 0.00121212
R31402 avss.n252 avss.n251 0.00121212
R31403 avss.n246 avss.n245 0.00121212
R31404 avss.n11270 avss.n11269 0.00121212
R31405 avss.n11213 avss.n11212 0.00121212
R31406 avss.n11624 avss.n11533 0.00121212
R31407 avss.n11529 avss.n11528 0.00121212
R31408 avss.n11573 avss.n11572 0.00121212
R31409 avss.n11570 avss.n11569 0.00121212
R31410 avss.n11564 avss.n11563 0.00121212
R31411 avss.n210 avss.n209 0.00121212
R31412 avss.n153 avss.n152 0.00121212
R31413 avss.n106 avss.n105 0.00121212
R31414 avss.n101 avss.n100 0.00121212
R31415 avss.n38 avss.n37 0.00121212
R31416 avss.n35 avss.n34 0.00121212
R31417 avss.n29 avss.n28 0.00121212
R31418 avss.n11491 avss.n11490 0.00121212
R31419 avss.n11434 avss.n11433 0.00121212
R31420 avss.n2675 avss.n2621 0.00101777
R31421 avss.n2653 avss.n2648 0.00101777
R31422 avss.n2916 avss.n2625 0.00101777
R31423 avss.n2805 avss.n2796 0.00101777
R31424 avss.n3619 avss.n2613 0.00101777
R31425 avss.n3027 avss.n3022 0.00101777
R31426 avss.n2965 avss.n2620 0.00101777
R31427 avss.n3140 avss.n2919 0.00101777
R31428 avss.n4953 avss.n4952 0.000675758
R31429 avss.n5088 avss.n4592 0.000675758
R31430 avss.n5307 avss.n5306 0.000675758
R31431 avss.n5442 avss.n4508 0.000675758
R31432 avss.n11626 avss.n11517 0.000675758
R31433 avss.n11516 avss.n11515 0.000675758
R31434 avss.n11405 avss.n11296 0.000675758
R31435 avss.n11295 avss.n11294 0.000675758
R31436 avss.n5660 avss.n5659 0.000674349
R31437 avss.n5795 avss.n4424 0.000674349
R31438 avss.n6013 avss.n6012 0.000674349
R31439 avss.n6148 avss.n4340 0.000674349
R31440 avss.n6366 avss.n6365 0.000674349
R31441 avss.n6501 avss.n4256 0.000674349
R31442 avss.n6719 avss.n6718 0.000674349
R31443 avss.n6854 avss.n4172 0.000674349
R31444 avss.n11184 avss.n11183 0.000674349
R31445 avss.n11182 avss.n11073 0.000674349
R31446 avss.n10963 avss.n10962 0.000674349
R31447 avss.n10961 avss.n10852 0.000674349
R31448 avss.n10742 avss.n10741 0.000674349
R31449 avss.n10740 avss.n10631 0.000674349
R31450 avss.n10521 avss.n10520 0.000674349
R31451 avss.n10519 avss.n10410 0.000674349
R31452 avss.n7072 avss.n7071 0.000672962
R31453 avss.n7207 avss.n4088 0.000672962
R31454 avss.n7425 avss.n7424 0.000672962
R31455 avss.n7560 avss.n4004 0.000672962
R31456 avss.n7778 avss.n7777 0.000672962
R31457 avss.n7913 avss.n3920 0.000672962
R31458 avss.n8131 avss.n8130 0.000672962
R31459 avss.n8266 avss.n3836 0.000672962
R31460 avss.n10300 avss.n10299 0.000672962
R31461 avss.n10298 avss.n10189 0.000672962
R31462 avss.n10079 avss.n10078 0.000672962
R31463 avss.n10077 avss.n9968 0.000672962
R31464 avss.n9858 avss.n9857 0.000672962
R31465 avss.n9856 avss.n9747 0.000672962
R31466 avss.n9637 avss.n9636 0.000672962
R31467 avss.n9635 avss.n9526 0.000672962
R31468 avss.n8484 avss.n8483 0.000671598
R31469 avss.n8619 avss.n3752 0.000671598
R31470 avss.n8837 avss.n8836 0.000671598
R31471 avss.n8972 avss.n3668 0.000671598
R31472 avss.n9416 avss.n9415 0.000671598
R31473 avss.n9414 avss.n9305 0.000671598
R31474 avss.n9195 avss.n9194 0.000671598
R31475 avss.n9193 avss.n9084 0.000671598
R31476 comparator_0.trim_0.n4.n11 comparator_0.trim_0.n4.t13 18.7845
R31477 comparator_0.trim_0.n4 comparator_0.trim_0.n4.t8 17.4527
R31478 comparator_0.trim_0.n4.n8 comparator_0.trim_0.n4.t12 17.4005
R31479 comparator_0.trim_0.n4.n8 comparator_0.trim_0.n4.t9 17.4005
R31480 comparator_0.trim_0.n4.n9 comparator_0.trim_0.n4.t11 17.4005
R31481 comparator_0.trim_0.n4.n9 comparator_0.trim_0.n4.t15 17.4005
R31482 comparator_0.trim_0.n4.n10 comparator_0.trim_0.n4.t10 17.4005
R31483 comparator_0.trim_0.n4.n10 comparator_0.trim_0.n4.t14 17.4005
R31484 comparator_0.trim_0.n4.n0 comparator_0.trim_0.n4.t3 2.33023
R31485 comparator_0.trim_0.n4.n2 comparator_0.trim_0.n4.n1 2.24237
R31486 comparator_0.trim_0.n4.n4 comparator_0.trim_0.n4.n3 2.24237
R31487 comparator_0.trim_0.n4.n1 comparator_0.trim_0.n4.n0 2.22512
R31488 comparator_0.trim_0.n4.n5 comparator_0.trim_0.n4.n4 2.22512
R31489 comparator_0.trim_0.n4.n3 comparator_0.trim_0.n4.n2 2.19064
R31490 comparator_0.trim_0.n4 comparator_0.trim_0.n4.t7 1.31756
R31491 comparator_0.trim_0.n4.n14 comparator_0.trim_0.n4.n13 1.01343
R31492 comparator_0.trim_0.n4.n13 comparator_0.trim_0.n4.n12 1.00912
R31493 comparator_0.trim_0.n4.n12 comparator_0.trim_0.n4.n11 0.974638
R31494 comparator_0.trim_0.n4.n6 comparator_0.trim_0.n4.n5 0.950849
R31495 comparator_0.trim_0.n4.n14 comparator_0.trim_0.n4.n6 0.703086
R31496 comparator_0.trim_0.n4.n14 comparator_0.trim_0.n4 0.612569
R31497 comparator_0.trim_0.n4.n11 comparator_0.trim_0.n4.n10 0.496573
R31498 comparator_0.trim_0.n4.n13 comparator_0.trim_0.n4.n8 0.436228
R31499 comparator_0.trim_0.n4.n12 comparator_0.trim_0.n4.n9 0.436228
R31500 comparator_0.trim_0.n4.n7 comparator_0.trim_0.n4 0.280672
R31501 comparator_0.trim_0.n4.n14 comparator_0.trim_0.n4.n7 0.207397
R31502 comparator_0.trim_0.n4.n7 comparator_0.trim_0.n4 0.17713
R31503 comparator_0.trim_0.n4.n5 comparator_0.trim_0.n4.t4 0.087375
R31504 comparator_0.trim_0.n4.n4 comparator_0.trim_0.n4.t1 0.087375
R31505 comparator_0.trim_0.n4.n3 comparator_0.trim_0.n4.t6 0.087375
R31506 comparator_0.trim_0.n4.n2 comparator_0.trim_0.n4.t2 0.087375
R31507 comparator_0.trim_0.n4.n1 comparator_0.trim_0.n4.t0 0.087375
R31508 comparator_0.trim_0.n4.n0 comparator_0.trim_0.n4.t5 0.087375
R31509 comparator_0.trim_0.n4.n6 comparator_0.trim_0.n4 0.0608448
R31510 comparator_0.trim_0.n4 comparator_0.trim_0.n4.n14 0.0608448
R31511 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n1 111.322
R31512 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y.n3 50.4671
R31513 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t0 26.5955
R31514 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t2 26.5955
R31515 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t1 24.9236
R31516 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t4 24.9236
R31517 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y.n5 13.5995
R31518 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n5 dac_0.sky130_fd_sc_hd__inv_2_0.Y 12.0325
R31519 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y.n4 11.2645
R31520 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_0.Y 8.80626
R31521 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_0.Y 6.1445
R31522 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n5 dac_0.sky130_fd_sc_hd__inv_2_0.Y 5.3765
R31523 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_0.Y 4.65505
R31524 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y.n2 2.0485
R31525 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_0.Y 1.55202
R31526 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y.t3 0.127353
R31527 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_0.Y 0.0462978
R31528 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t3 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n0 0.0391355
R31529 vinn.n8 vinn.t79 29.3118
R31530 vinn.n22 vinn.t11 29.3118
R31531 vinn.n37 vinn.t44 29.3118
R31532 vinn.n52 vinn.t24 29.3118
R31533 vinn.n13 vinn.t78 29.3084
R31534 vinn.n27 vinn.t19 29.3084
R31535 vinn.n42 vinn.t47 29.3084
R31536 vinn.n57 vinn.t21 29.3084
R31537 vinn.n6 vinn.t76 28.5655
R31538 vinn.n6 vinn.t72 28.5655
R31539 vinn.n4 vinn.t73 28.5655
R31540 vinn.n4 vinn.t70 28.5655
R31541 vinn.n2 vinn.t74 28.5655
R31542 vinn.n2 vinn.t77 28.5655
R31543 vinn.n0 vinn.t75 28.5655
R31544 vinn.n0 vinn.t71 28.5655
R31545 vinn.n20 vinn.t13 28.5655
R31546 vinn.n20 vinn.t14 28.5655
R31547 vinn.n18 vinn.t12 28.5655
R31548 vinn.n18 vinn.t15 28.5655
R31549 vinn.n16 vinn.t17 28.5655
R31550 vinn.n16 vinn.t16 28.5655
R31551 vinn.n14 vinn.t18 28.5655
R31552 vinn.n14 vinn.t10 28.5655
R31553 vinn.n35 vinn.t42 28.5655
R31554 vinn.n35 vinn.t40 28.5655
R31555 vinn.n33 vinn.t48 28.5655
R31556 vinn.n33 vinn.t41 28.5655
R31557 vinn.n31 vinn.t45 28.5655
R31558 vinn.n31 vinn.t49 28.5655
R31559 vinn.n29 vinn.t46 28.5655
R31560 vinn.n29 vinn.t43 28.5655
R31561 vinn.n50 vinn.t22 28.5655
R31562 vinn.n50 vinn.t29 28.5655
R31563 vinn.n48 vinn.t26 28.5655
R31564 vinn.n48 vinn.t25 28.5655
R31565 vinn.n46 vinn.t27 28.5655
R31566 vinn.n46 vinn.t20 28.5655
R31567 vinn.n44 vinn.t28 28.5655
R31568 vinn.n44 vinn.t23 28.5655
R31569 vinn.n8 vinn.t6 18.1397
R31570 vinn.n13 vinn.t9 18.1397
R31571 vinn.n22 vinn.t53 18.1397
R31572 vinn.n27 vinn.t59 18.1397
R31573 vinn.n37 vinn.t64 18.1397
R31574 vinn.n42 vinn.t60 18.1397
R31575 vinn.n52 vinn.t32 18.1397
R31576 vinn.n57 vinn.t39 18.1397
R31577 vinn.n7 vinn.t3 17.4005
R31578 vinn.n7 vinn.t7 17.4005
R31579 vinn.n5 vinn.t8 17.4005
R31580 vinn.n5 vinn.t0 17.4005
R31581 vinn.n3 vinn.t1 17.4005
R31582 vinn.n3 vinn.t4 17.4005
R31583 vinn.n1 vinn.t2 17.4005
R31584 vinn.n1 vinn.t5 17.4005
R31585 vinn.n21 vinn.t57 17.4005
R31586 vinn.n21 vinn.t58 17.4005
R31587 vinn.n19 vinn.t54 17.4005
R31588 vinn.n19 vinn.t50 17.4005
R31589 vinn.n17 vinn.t55 17.4005
R31590 vinn.n17 vinn.t51 17.4005
R31591 vinn.n15 vinn.t56 17.4005
R31592 vinn.n15 vinn.t52 17.4005
R31593 vinn.n36 vinn.t66 17.4005
R31594 vinn.n36 vinn.t61 17.4005
R31595 vinn.n34 vinn.t68 17.4005
R31596 vinn.n34 vinn.t62 17.4005
R31597 vinn.n32 vinn.t65 17.4005
R31598 vinn.n32 vinn.t69 17.4005
R31599 vinn.n30 vinn.t63 17.4005
R31600 vinn.n30 vinn.t67 17.4005
R31601 vinn.n51 vinn.t33 17.4005
R31602 vinn.n51 vinn.t37 17.4005
R31603 vinn.n49 vinn.t34 17.4005
R31604 vinn.n49 vinn.t38 17.4005
R31605 vinn.n47 vinn.t35 17.4005
R31606 vinn.n47 vinn.t30 17.4005
R31607 vinn.n45 vinn.t36 17.4005
R31608 vinn.n45 vinn.t31 17.4005
R31609 vinn.n59 vinn.n58 8.59648
R31610 vinn.n61 vinn.n60 7.00774
R31611 vinn.n60 vinn.n59 6.6802
R31612 vinn vinn.n61 2.91369
R31613 vinn.n61 vinn 2.19494
R31614 vinn.n59 vinn.n43 1.91314
R31615 vinn.n60 vinn.n28 1.91178
R31616 vinn.n10 vinn.n9 0.811311
R31617 vinn.n24 vinn.n23 0.811311
R31618 vinn.n39 vinn.n38 0.811311
R31619 vinn.n54 vinn.n53 0.811311
R31620 vinn.n12 vinn.n11 0.799575
R31621 vinn.n26 vinn.n25 0.799575
R31622 vinn.n41 vinn.n40 0.799575
R31623 vinn.n56 vinn.n55 0.799575
R31624 vinn.n11 vinn.n10 0.794419
R31625 vinn.n25 vinn.n24 0.794419
R31626 vinn.n40 vinn.n39 0.794419
R31627 vinn.n55 vinn.n54 0.794419
R31628 vinn.n9 vinn.n8 0.787662
R31629 vinn.n23 vinn.n22 0.787662
R31630 vinn.n38 vinn.n37 0.787662
R31631 vinn.n53 vinn.n52 0.787662
R31632 vinn.n13 vinn.n12 0.773526
R31633 vinn.n27 vinn.n26 0.773526
R31634 vinn.n42 vinn.n41 0.773526
R31635 vinn.n57 vinn.n56 0.773526
R31636 vinn.n9 vinn.n6 0.746823
R31637 vinn.n10 vinn.n4 0.746823
R31638 vinn.n11 vinn.n2 0.746823
R31639 vinn.n23 vinn.n20 0.746823
R31640 vinn.n24 vinn.n18 0.746823
R31641 vinn.n25 vinn.n16 0.746823
R31642 vinn.n38 vinn.n35 0.746823
R31643 vinn.n39 vinn.n33 0.746823
R31644 vinn.n40 vinn.n31 0.746823
R31645 vinn.n53 vinn.n50 0.746823
R31646 vinn.n54 vinn.n48 0.746823
R31647 vinn.n55 vinn.n46 0.746823
R31648 vinn.n12 vinn.n0 0.743351
R31649 vinn.n26 vinn.n14 0.743351
R31650 vinn.n41 vinn.n29 0.743351
R31651 vinn.n56 vinn.n44 0.743351
R31652 vinn.n9 vinn.n7 0.739748
R31653 vinn.n10 vinn.n5 0.739748
R31654 vinn.n11 vinn.n3 0.739748
R31655 vinn.n12 vinn.n1 0.739748
R31656 vinn.n23 vinn.n21 0.739748
R31657 vinn.n24 vinn.n19 0.739748
R31658 vinn.n25 vinn.n17 0.739748
R31659 vinn.n26 vinn.n15 0.739748
R31660 vinn.n38 vinn.n36 0.739748
R31661 vinn.n39 vinn.n34 0.739748
R31662 vinn.n40 vinn.n32 0.739748
R31663 vinn.n41 vinn.n30 0.739748
R31664 vinn.n53 vinn.n51 0.739748
R31665 vinn.n54 vinn.n49 0.739748
R31666 vinn.n55 vinn.n47 0.739748
R31667 vinn.n56 vinn.n45 0.739748
R31668 vinn vinn.n13 0.627876
R31669 vinn.n28 vinn.n27 0.580651
R31670 vinn.n43 vinn.n42 0.579111
R31671 vinn.n58 vinn.n57 0.573599
R31672 vinn.n58 vinn 0.063
R31673 vinn.n43 vinn 0.0583961
R31674 vinn.n28 vinn 0.056769
R31675 dac_1.out.n20 dac_1.out.t87 130.87
R31676 dac_1.out.n74 dac_1.out.t74 28.5655
R31677 dac_1.out.n74 dac_1.out.t71 28.5655
R31678 dac_1.out.n27 dac_1.out.t17 28.5655
R31679 dac_1.out.n27 dac_1.out.t12 28.5655
R31680 dac_1.out.n30 dac_1.out.t16 28.5655
R31681 dac_1.out.n30 dac_1.out.t11 28.5655
R31682 dac_1.out.n25 dac_1.out.t15 28.5655
R31683 dac_1.out.n25 dac_1.out.t10 28.5655
R31684 dac_1.out.n24 dac_1.out.t14 28.5655
R31685 dac_1.out.n24 dac_1.out.t19 28.5655
R31686 dac_1.out.n23 dac_1.out.t18 28.5655
R31687 dac_1.out.n23 dac_1.out.t13 28.5655
R31688 dac_1.out.n39 dac_1.out.t48 28.5655
R31689 dac_1.out.n39 dac_1.out.t44 28.5655
R31690 dac_1.out.n42 dac_1.out.t40 28.5655
R31691 dac_1.out.n42 dac_1.out.t43 28.5655
R31692 dac_1.out.n37 dac_1.out.t46 28.5655
R31693 dac_1.out.n37 dac_1.out.t42 28.5655
R31694 dac_1.out.n36 dac_1.out.t45 28.5655
R31695 dac_1.out.n36 dac_1.out.t49 28.5655
R31696 dac_1.out.n35 dac_1.out.t41 28.5655
R31697 dac_1.out.n35 dac_1.out.t47 28.5655
R31698 dac_1.out.n51 dac_1.out.t23 28.5655
R31699 dac_1.out.n51 dac_1.out.t21 28.5655
R31700 dac_1.out.n54 dac_1.out.t20 28.5655
R31701 dac_1.out.n54 dac_1.out.t27 28.5655
R31702 dac_1.out.n49 dac_1.out.t29 28.5655
R31703 dac_1.out.n49 dac_1.out.t26 28.5655
R31704 dac_1.out.n48 dac_1.out.t28 28.5655
R31705 dac_1.out.n48 dac_1.out.t25 28.5655
R31706 dac_1.out.n47 dac_1.out.t24 28.5655
R31707 dac_1.out.n47 dac_1.out.t22 28.5655
R31708 dac_1.out.n64 dac_1.out.t72 28.5655
R31709 dac_1.out.n64 dac_1.out.t79 28.5655
R31710 dac_1.out.n69 dac_1.out.t75 28.5655
R31711 dac_1.out.n69 dac_1.out.t76 28.5655
R31712 dac_1.out.n71 dac_1.out.t73 28.5655
R31713 dac_1.out.n71 dac_1.out.t77 28.5655
R31714 dac_1.out.n73 dac_1.out.t70 28.5655
R31715 dac_1.out.n73 dac_1.out.t78 28.5655
R31716 dac_1.out.n28 dac_1.out.t55 17.4005
R31717 dac_1.out.n28 dac_1.out.t52 17.4005
R31718 dac_1.out.n31 dac_1.out.t54 17.4005
R31719 dac_1.out.n31 dac_1.out.t59 17.4005
R31720 dac_1.out.n26 dac_1.out.t53 17.4005
R31721 dac_1.out.n26 dac_1.out.t58 17.4005
R31722 dac_1.out.n33 dac_1.out.t51 17.4005
R31723 dac_1.out.n33 dac_1.out.t57 17.4005
R31724 dac_1.out.n34 dac_1.out.t56 17.4005
R31725 dac_1.out.n34 dac_1.out.t50 17.4005
R31726 dac_1.out.n40 dac_1.out.t66 17.4005
R31727 dac_1.out.n40 dac_1.out.t61 17.4005
R31728 dac_1.out.n43 dac_1.out.t68 17.4005
R31729 dac_1.out.n43 dac_1.out.t64 17.4005
R31730 dac_1.out.n38 dac_1.out.t63 17.4005
R31731 dac_1.out.n38 dac_1.out.t60 17.4005
R31732 dac_1.out.n45 dac_1.out.t62 17.4005
R31733 dac_1.out.n45 dac_1.out.t67 17.4005
R31734 dac_1.out.n46 dac_1.out.t69 17.4005
R31735 dac_1.out.n46 dac_1.out.t65 17.4005
R31736 dac_1.out.n52 dac_1.out.t31 17.4005
R31737 dac_1.out.n52 dac_1.out.t39 17.4005
R31738 dac_1.out.n55 dac_1.out.t30 17.4005
R31739 dac_1.out.n55 dac_1.out.t36 17.4005
R31740 dac_1.out.n50 dac_1.out.t38 17.4005
R31741 dac_1.out.n50 dac_1.out.t35 17.4005
R31742 dac_1.out.n57 dac_1.out.t37 17.4005
R31743 dac_1.out.n57 dac_1.out.t34 17.4005
R31744 dac_1.out.n58 dac_1.out.t32 17.4005
R31745 dac_1.out.n58 dac_1.out.t33 17.4005
R31746 dac_1.out.n68 dac_1.out.t2 17.4005
R31747 dac_1.out.n68 dac_1.out.t7 17.4005
R31748 dac_1.out.n70 dac_1.out.t3 17.4005
R31749 dac_1.out.n70 dac_1.out.t4 17.4005
R31750 dac_1.out.n72 dac_1.out.t0 17.4005
R31751 dac_1.out.n72 dac_1.out.t5 17.4005
R31752 dac_1.out.n77 dac_1.out.t8 17.4005
R31753 dac_1.out.n77 dac_1.out.t6 17.4005
R31754 dac_1.out.n75 dac_1.out.t1 17.4005
R31755 dac_1.out.n75 dac_1.out.t9 17.4005
R31756 dac_1.out.n21 dac_1.out.n20 9.84842
R31757 dac_1.out.n59 dac_1.out 8.6431
R31758 dac_1.out.n60 dac_1.out.n59 6.19787
R31759 dac_1.out.n66 dac_1.out.n65 4.58032
R31760 dac_1.out.n61 dac_1.out.n60 4.3755
R31761 dac_1.out.n13 dac_1.out 3.9297
R31762 dac_1.out.n12 dac_1.out 3.4597
R31763 dac_1.out.n19 dac_1.out 2.9897
R31764 dac_1.out.n1 dac_1.out.n24 2.5289
R31765 dac_1.out.n4 dac_1.out.n36 2.5289
R31766 dac_1.out.n7 dac_1.out.n48 2.5289
R31767 dac_1.out.n10 dac_1.out.n69 2.5289
R31768 dac_1.out.n0 dac_1.out.n30 2.52132
R31769 dac_1.out.n3 dac_1.out.n42 2.52132
R31770 dac_1.out.n6 dac_1.out.n54 2.52132
R31771 dac_1.out.n11 dac_1.out.n73 2.52132
R31772 dac_1.out.n18 dac_1.out 2.5197
R31773 dac_1.out dac_1.out.n62 2.47089
R31774 dac_1.out.n32 dac_1.out.n25 2.45817
R31775 dac_1.out.n44 dac_1.out.n37 2.45817
R31776 dac_1.out.n56 dac_1.out.n49 2.45817
R31777 dac_1.out.n78 dac_1.out.n71 2.45817
R31778 dac_1.out.n76 dac_1.out.n74 2.4534
R31779 dac_1.out.n29 dac_1.out.n27 2.4534
R31780 dac_1.out.n41 dac_1.out.n39 2.4534
R31781 dac_1.out.n53 dac_1.out.n51 2.4534
R31782 dac_1.out.n60 dac_1.out 2.42846
R31783 dac_1.out.n59 dac_1.out 2.29984
R31784 dac_1.out.n17 dac_1.out 2.0497
R31785 dac_1.out.n62 dac_1.out.n61 1.90839
R31786 dac_1.out.n20 dac_1.out 1.88285
R31787 dac_1.out.n16 dac_1.out 1.5797
R31788 dac_1.out.n15 dac_1.out 1.1097
R31789 dac_1.out dac_1.out.n5 1.05971
R31790 dac_1.out dac_1.out.n9 1.05971
R31791 dac_1.out dac_1.out.n2 1.05955
R31792 dac_1.out.t83 dac_1.out 0.773227
R31793 dac_1.out.n1 dac_1.out.n33 0.750533
R31794 dac_1.out.n4 dac_1.out.n45 0.750533
R31795 dac_1.out.n7 dac_1.out.n57 0.750533
R31796 dac_1.out.n10 dac_1.out.n70 0.750533
R31797 dac_1.out.n2 dac_1.out.n34 0.747922
R31798 dac_1.out.n5 dac_1.out.n46 0.747922
R31799 dac_1.out.n8 dac_1.out.n58 0.747922
R31800 dac_1.out.n9 dac_1.out.n68 0.747922
R31801 dac_1.out.n32 dac_1.out.n26 0.729365
R31802 dac_1.out.n44 dac_1.out.n38 0.729365
R31803 dac_1.out.n56 dac_1.out.n50 0.729365
R31804 dac_1.out.n78 dac_1.out.n72 0.729365
R31805 dac_1.out.n0 dac_1.out.n31 0.725192
R31806 dac_1.out.n3 dac_1.out.n43 0.725192
R31807 dac_1.out.n6 dac_1.out.n55 0.725192
R31808 dac_1.out.n11 dac_1.out.n77 0.725192
R31809 dac_1.out.n1 dac_1.out.n32 0.720895
R31810 dac_1.out.n4 dac_1.out.n44 0.720895
R31811 dac_1.out.n7 dac_1.out.n56 0.720895
R31812 dac_1.out.n10 dac_1.out.n78 0.720895
R31813 dac_1.out.n32 dac_1.out.n0 0.714316
R31814 dac_1.out.n44 dac_1.out.n3 0.714316
R31815 dac_1.out.n56 dac_1.out.n6 0.714316
R31816 dac_1.out.n78 dac_1.out.n11 0.714316
R31817 dac_1.out.t80 dac_1.out 0.685649
R31818 dac_1.out.n29 dac_1.out.n28 0.66743
R31819 dac_1.out.n41 dac_1.out.n40 0.66743
R31820 dac_1.out.n53 dac_1.out.n52 0.66743
R31821 dac_1.out.n76 dac_1.out.n75 0.665483
R31822 dac_1.out.n14 dac_1.out 0.6397
R31823 dac_1.out.t82 dac_1.out 0.598071
R31824 dac_1.out.t89 dac_1.out 0.510494
R31825 dac_1.out.n61 dac_1.out.n22 0.437652
R31826 dac_1.out.t81 dac_1.out 0.422916
R31827 dac_1.out.t88 dac_1.out 0.335339
R31828 dac_1.out.t85 dac_1.out 0.247761
R31829 dac_1.out.t82 dac_1.out.n19 0.218267
R31830 dac_1.out.t80 dac_1.out.n12 0.218267
R31831 dac_1.out.t84 dac_1.out 0.218267
R31832 dac_1.out.t86 dac_1.out.n14 0.218267
R31833 dac_1.out.t85 dac_1.out.n15 0.218267
R31834 dac_1.out.t88 dac_1.out.n16 0.218267
R31835 dac_1.out.t81 dac_1.out.n17 0.218267
R31836 dac_1.out.t89 dac_1.out.n18 0.218267
R31837 dac_1.out.t86 dac_1.out 0.160183
R31838 dac_1.out.n65 dac_1.out.n64 0.100193
R31839 dac_1.out.t84 dac_1.out 0.0726056
R31840 dac_1.out.n62 dac_1.out 0.063
R31841 dac_1.out.n66 dac_1.out.n63 0.0421667
R31842 dac_1.out.n2 dac_1.out.n23 2.52329
R31843 dac_1.out.n5 dac_1.out.n35 2.52329
R31844 dac_1.out.n8 dac_1.out.n47 2.52329
R31845 dac_1.out dac_1.out.n8 1.07616
R31846 dac_1.out.n11 dac_1.out.n76 0.711026
R31847 dac_1.out.n6 dac_1.out.n53 0.711026
R31848 dac_1.out.n3 dac_1.out.n41 0.711026
R31849 dac_1.out.n0 dac_1.out.n29 0.711026
R31850 dac_1.out.n8 dac_1.out.n7 0.658395
R31851 dac_1.out.n5 dac_1.out.n4 0.658395
R31852 dac_1.out.n2 dac_1.out.n1 0.658395
R31853 dac_1.out.n9 dac_1.out.n10 0.651816
R31854 dac_1.out.n9 dac_1.out.n67 0.585149
R31855 dac_1.out dac_1.out.t83 0.398433
R31856 dac_1.out dac_1.out.t89 0.398433
R31857 dac_1.out.t82 dac_1.out 0.398433
R31858 dac_1.out.t80 dac_1.out 0.398433
R31859 dac_1.out.t84 dac_1.out 0.398433
R31860 dac_1.out.t86 dac_1.out 0.398433
R31861 dac_1.out.t85 dac_1.out 0.398433
R31862 dac_1.out.t88 dac_1.out 0.398433
R31863 dac_1.out.t81 dac_1.out 0.398433
R31864 dac_1.out.n21 dac_1.out 0.268269
R31865 dac_1.out.n22 dac_1.out 0.240069
R31866 dac_1.out.t83 dac_1.out.n13 0.240015
R31867 dac_1.out.n22 dac_1.out 0.203383
R31868 dac_1.out dac_1.out.n21 0.175183
R31869 dac_1.out.n12 dac_1.out.t82 0.0475
R31870 dac_1.out.n18 dac_1.out.t81 0.0475
R31871 dac_1.out.n17 dac_1.out.t88 0.0475
R31872 dac_1.out.n13 dac_1.out.t80 0.0475
R31873 dac_1.out.n15 dac_1.out.t86 0.0475
R31874 dac_1.out.n14 dac_1.out.t84 0.0475
R31875 dac_1.out.n16 dac_1.out.t85 0.0475
R31876 dac_1.out.n19 dac_1.out.t89 0.0475
R31877 dac_1.out.n67 dac_1.out.n66 0.0310556
R31878 ctln1.n3 ctln1.t3 212.081
R31879 ctln1.n2 ctln1.t1 212.081
R31880 ctln1.n3 ctln1.t0 139.78
R31881 ctln1.n2 ctln1.t2 139.78
R31882 ctln1.n3 ctln1.n2 61.346
R31883 ctln1.n5 ctln1.n3 38.5428
R31884 ctln1.n5 ctln1.n0 9.30881
R31885 ctln1.n6 ctln1.n5 9.3005
R31886 ctln1.n7 ctln1.n6 9.01417
R31887 ctln1.n4 ctln1 3.09989
R31888 ctln1.n8 ctln1 1.62182
R31889 ctln1.n5 ctln1.n4 1.53719
R31890 ctln1.n7 ctln1.n0 0.0569565
R31891 ctln1.n6 ctln1.n1 0.03175
R31892 ctln1 ctln1.n8 0.0225588
R31893 ctln1.n8 ctln1 0.0149231
R31894 ctln1 ctln1.n7 0.00771154
R31895 ctln1.n4 ctln1.n1 0.00148276
R31896 ctln1.n1 ctln1.n0 0.00100057
R31897 sample.n64 sample.t16 212.081
R31898 sample.n66 sample.t0 212.081
R31899 sample.n63 sample.t22 212.081
R31900 sample.n71 sample.t6 212.081
R31901 sample.n45 sample.t36 212.081
R31902 sample.n47 sample.t2 212.081
R31903 sample.n44 sample.t39 212.081
R31904 sample.n52 sample.t19 212.081
R31905 sample.n26 sample.t10 212.081
R31906 sample.n28 sample.t18 212.081
R31907 sample.n25 sample.t1 212.081
R31908 sample.n33 sample.t23 212.081
R31909 sample.n5 sample.t11 212.081
R31910 sample.n7 sample.t57 212.081
R31911 sample.n4 sample.t15 212.081
R31912 sample.n12 sample.t42 212.081
R31913 sample.n142 sample.t38 212.081
R31914 sample.n144 sample.t17 212.081
R31915 sample.n141 sample.t43 212.081
R31916 sample.n150 sample.t9 212.081
R31917 sample.n122 sample.t5 212.081
R31918 sample.n124 sample.t28 212.081
R31919 sample.n121 sample.t7 212.081
R31920 sample.n129 sample.t49 212.081
R31921 sample.n103 sample.t45 212.081
R31922 sample.n105 sample.t25 212.081
R31923 sample.n102 sample.t52 212.081
R31924 sample.n110 sample.t29 212.081
R31925 sample.n84 sample.t35 212.081
R31926 sample.n86 sample.t46 212.081
R31927 sample.n83 sample.t27 212.081
R31928 sample.n91 sample.t54 212.081
R31929 sample.n64 sample.t53 139.78
R31930 sample.n66 sample.t30 139.78
R31931 sample.n63 sample.t60 139.78
R31932 sample.n71 sample.t34 139.78
R31933 sample.n45 sample.t8 139.78
R31934 sample.n47 sample.t32 139.78
R31935 sample.n44 sample.t12 139.78
R31936 sample.n52 sample.t58 139.78
R31937 sample.n26 sample.t41 139.78
R31938 sample.n28 sample.t56 139.78
R31939 sample.n25 sample.t31 139.78
R31940 sample.n33 sample.t61 139.78
R31941 sample.n5 sample.t44 139.78
R31942 sample.n7 sample.t24 139.78
R31943 sample.n4 sample.t51 139.78
R31944 sample.n12 sample.t14 139.78
R31945 sample.n142 sample.t63 139.78
R31946 sample.n144 sample.t47 139.78
R31947 sample.n141 sample.t50 139.78
R31948 sample.n150 sample.t62 139.78
R31949 sample.n122 sample.t21 139.78
R31950 sample.n124 sample.t26 139.78
R31951 sample.n121 sample.t13 139.78
R31952 sample.n129 sample.t3 139.78
R31953 sample.n103 sample.t4 139.78
R31954 sample.n105 sample.t55 139.78
R31955 sample.n102 sample.t59 139.78
R31956 sample.n110 sample.t40 139.78
R31957 sample.n84 sample.t20 139.78
R31958 sample.n86 sample.t48 139.78
R31959 sample.n83 sample.t33 139.78
R31960 sample.n91 sample.t37 139.78
R31961 sample.n65 sample 78.3045
R31962 sample.n46 sample 78.3045
R31963 sample.n27 sample 78.3045
R31964 sample.n6 sample 78.3045
R31965 sample.n143 sample 78.3045
R31966 sample.n123 sample 78.3045
R31967 sample.n104 sample 78.3045
R31968 sample.n85 sample 78.3045
R31969 sample.n68 sample.n67 76.0005
R31970 sample.n70 sample.n69 76.0005
R31971 sample.n49 sample.n48 76.0005
R31972 sample.n51 sample.n50 76.0005
R31973 sample.n30 sample.n29 76.0005
R31974 sample.n32 sample.n31 76.0005
R31975 sample.n9 sample.n8 76.0005
R31976 sample.n11 sample.n10 76.0005
R31977 sample.n146 sample.n145 76.0005
R31978 sample.n149 sample.n148 76.0005
R31979 sample.n126 sample.n125 76.0005
R31980 sample.n128 sample.n127 76.0005
R31981 sample.n107 sample.n106 76.0005
R31982 sample.n109 sample.n108 76.0005
R31983 sample.n88 sample.n87 76.0005
R31984 sample.n90 sample.n89 76.0005
R31985 sample.n72 sample.n71 44.8017
R31986 sample.n53 sample.n52 44.8017
R31987 sample.n34 sample.n33 44.8017
R31988 sample.n13 sample.n12 44.8017
R31989 sample.n151 sample.n150 44.8017
R31990 sample.n130 sample.n129 44.8017
R31991 sample.n111 sample.n110 44.8017
R31992 sample.n92 sample.n91 44.8017
R31993 sample.n65 sample.n64 30.6732
R31994 sample.n66 sample.n65 30.6732
R31995 sample.n67 sample.n66 30.6732
R31996 sample.n67 sample.n63 30.6732
R31997 sample.n70 sample.n63 30.6732
R31998 sample.n71 sample.n70 30.6732
R31999 sample.n46 sample.n45 30.6732
R32000 sample.n47 sample.n46 30.6732
R32001 sample.n48 sample.n47 30.6732
R32002 sample.n48 sample.n44 30.6732
R32003 sample.n51 sample.n44 30.6732
R32004 sample.n52 sample.n51 30.6732
R32005 sample.n27 sample.n26 30.6732
R32006 sample.n28 sample.n27 30.6732
R32007 sample.n29 sample.n28 30.6732
R32008 sample.n29 sample.n25 30.6732
R32009 sample.n32 sample.n25 30.6732
R32010 sample.n33 sample.n32 30.6732
R32011 sample.n6 sample.n5 30.6732
R32012 sample.n7 sample.n6 30.6732
R32013 sample.n8 sample.n7 30.6732
R32014 sample.n8 sample.n4 30.6732
R32015 sample.n11 sample.n4 30.6732
R32016 sample.n12 sample.n11 30.6732
R32017 sample.n143 sample.n142 30.6732
R32018 sample.n144 sample.n143 30.6732
R32019 sample.n145 sample.n144 30.6732
R32020 sample.n145 sample.n141 30.6732
R32021 sample.n149 sample.n141 30.6732
R32022 sample.n150 sample.n149 30.6732
R32023 sample.n123 sample.n122 30.6732
R32024 sample.n124 sample.n123 30.6732
R32025 sample.n125 sample.n124 30.6732
R32026 sample.n125 sample.n121 30.6732
R32027 sample.n128 sample.n121 30.6732
R32028 sample.n129 sample.n128 30.6732
R32029 sample.n104 sample.n103 30.6732
R32030 sample.n105 sample.n104 30.6732
R32031 sample.n106 sample.n105 30.6732
R32032 sample.n106 sample.n102 30.6732
R32033 sample.n109 sample.n102 30.6732
R32034 sample.n110 sample.n109 30.6732
R32035 sample.n85 sample.n84 30.6732
R32036 sample.n86 sample.n85 30.6732
R32037 sample.n87 sample.n86 30.6732
R32038 sample.n87 sample.n83 30.6732
R32039 sample.n90 sample.n83 30.6732
R32040 sample.n91 sample.n90 30.6732
R32041 sample.n155 sample 27.0493
R32042 sample.n68 sample 19.2005
R32043 sample.n49 sample 19.2005
R32044 sample.n30 sample 19.2005
R32045 sample.n9 sample 19.2005
R32046 sample.n146 sample 19.2005
R32047 sample.n126 sample 19.2005
R32048 sample.n107 sample 19.2005
R32049 sample.n88 sample 19.2005
R32050 sample.n69 sample 17.1525
R32051 sample.n50 sample 17.1525
R32052 sample.n31 sample 17.1525
R32053 sample.n10 sample 17.1525
R32054 sample.n148 sample 17.1525
R32055 sample.n127 sample 17.1525
R32056 sample.n108 sample 17.1525
R32057 sample.n89 sample 17.1525
R32058 sample sample.n60 12.2885
R32059 sample sample.n41 12.2885
R32060 sample sample.n22 12.2885
R32061 sample sample.n2 12.2885
R32062 sample sample.n147 12.2885
R32063 sample.n132 sample 12.2885
R32064 sample.n113 sample 12.2885
R32065 sample.n94 sample 12.2885
R32066 sample.n60 sample.n58 9.34456
R32067 sample.n41 sample.n39 9.34456
R32068 sample.n22 sample.n20 9.34456
R32069 sample.n133 sample.n132 9.34456
R32070 sample.n114 sample.n113 9.34456
R32071 sample.n95 sample.n94 9.34456
R32072 sample.n147 sample.n137 9.34405
R32073 sample.n72 sample.n59 9.3005
R32074 sample.n62 sample.n61 9.3005
R32075 sample.n53 sample.n40 9.3005
R32076 sample.n43 sample.n42 9.3005
R32077 sample.n34 sample.n21 9.3005
R32078 sample.n24 sample.n23 9.3005
R32079 sample.n140 sample.n139 9.3005
R32080 sample.n152 sample.n151 9.3005
R32081 sample.n130 sample.n120 9.3005
R32082 sample.n119 sample.n118 9.3005
R32083 sample.n111 sample.n101 9.3005
R32084 sample.n100 sample.n99 9.3005
R32085 sample.n92 sample.n82 9.3005
R32086 sample.n81 sample.n80 9.3005
R32087 sample.n61 sample.n57 9.01011
R32088 sample.n42 sample.n38 9.01011
R32089 sample.n23 sample.n19 9.01011
R32090 sample.n139 sample.n136 9.01011
R32091 sample.n134 sample.n118 9.01011
R32092 sample.n115 sample.n99 9.01011
R32093 sample.n96 sample.n80 9.01011
R32094 sample.n154 sample.n153 9.0005
R32095 sample.n69 sample 6.4005
R32096 sample.n50 sample 6.4005
R32097 sample.n31 sample 6.4005
R32098 sample.n10 sample 6.4005
R32099 sample.n148 sample 6.4005
R32100 sample.n127 sample 6.4005
R32101 sample.n108 sample 6.4005
R32102 sample.n89 sample 6.4005
R32103 sample.n76 sample 5.80233
R32104 sample.n77 sample 5.80233
R32105 sample.n78 sample 5.80233
R32106 sample sample.n155 4.85416
R32107 sample.n73 sample.n60 4.6085
R32108 sample.n72 sample.n62 4.6085
R32109 sample.n54 sample.n41 4.6085
R32110 sample.n53 sample.n43 4.6085
R32111 sample.n35 sample.n22 4.6085
R32112 sample.n34 sample.n24 4.6085
R32113 sample.n14 sample.n2 4.6085
R32114 sample.n13 sample.n3 4.6085
R32115 sample.n147 sample.n138 4.6085
R32116 sample.n151 sample.n140 4.6085
R32117 sample.n132 sample.n131 4.6085
R32118 sample.n130 sample.n119 4.6085
R32119 sample.n113 sample.n112 4.6085
R32120 sample.n111 sample.n100 4.6085
R32121 sample.n94 sample.n93 4.6085
R32122 sample.n92 sample.n81 4.6085
R32123 sample.n75 sample.n74 4.501
R32124 sample.n56 sample.n55 4.501
R32125 sample.n37 sample.n36 4.501
R32126 sample.n135 sample.n117 4.501
R32127 sample.n116 sample.n98 4.501
R32128 sample.n97 sample.n79 4.501
R32129 sample sample.n68 4.3525
R32130 sample sample.n49 4.3525
R32131 sample sample.n30 4.3525
R32132 sample sample.n9 4.3525
R32133 sample sample.n146 4.3525
R32134 sample sample.n126 4.3525
R32135 sample sample.n107 4.3525
R32136 sample sample.n88 4.3525
R32137 sample.n62 sample 1.7925
R32138 sample.n43 sample 1.7925
R32139 sample.n24 sample 1.7925
R32140 sample.n3 sample 1.7925
R32141 sample.n140 sample 1.7925
R32142 sample.n119 sample 1.7925
R32143 sample.n100 sample 1.7925
R32144 sample.n81 sample 1.7925
R32145 sample sample.n75 0.958647
R32146 sample.n76 sample.n56 0.897671
R32147 sample.n77 sample.n37 0.897671
R32148 sample.n78 sample.n18 0.897671
R32149 sample sample.n135 0.897671
R32150 sample sample.n116 0.897671
R32151 sample sample.n97 0.897671
R32152 sample sample.n154 0.869696
R32153 sample.n73 sample.n72 0.2565
R32154 sample.n54 sample.n53 0.2565
R32155 sample.n35 sample.n34 0.2565
R32156 sample.n14 sample.n13 0.2565
R32157 sample.n151 sample.n138 0.2565
R32158 sample.n131 sample.n130 0.2565
R32159 sample.n112 sample.n111 0.2565
R32160 sample.n93 sample.n92 0.2565
R32161 sample.n155 sample 0.119402
R32162 sample sample.n76 0.0614756
R32163 sample sample.n77 0.0614756
R32164 sample sample.n78 0.0614756
R32165 sample.n155 sample 0.0614756
R32166 sample.n154 sample.n136 0.0557885
R32167 sample.n61 sample.n59 0.0437692
R32168 sample.n42 sample.n40 0.0437692
R32169 sample.n23 sample.n21 0.0437692
R32170 sample.n1 sample.n0 0.0437692
R32171 sample.n152 sample.n139 0.0437692
R32172 sample.n120 sample.n118 0.0437692
R32173 sample.n101 sample.n99 0.0437692
R32174 sample.n82 sample.n80 0.0437692
R32175 sample.n75 sample.n57 0.0286442
R32176 sample.n56 sample.n38 0.0286442
R32177 sample.n37 sample.n19 0.0286442
R32178 sample.n18 sample.n17 0.0286442
R32179 sample.n135 sample.n134 0.0286442
R32180 sample.n116 sample.n115 0.0286442
R32181 sample.n97 sample.n96 0.0286442
R32182 sample.n74 sample.n59 0.00290385
R32183 sample.n55 sample.n40 0.00290385
R32184 sample.n36 sample.n21 0.00290385
R32185 sample.n15 sample.n1 0.00290385
R32186 sample.n153 sample.n152 0.00290385
R32187 sample.n120 sample.n117 0.00290385
R32188 sample.n101 sample.n98 0.00290385
R32189 sample.n82 sample.n79 0.00290385
R32190 sample.n137 sample.n136 0.00266047
R32191 sample.n58 sample.n57 0.00216539
R32192 sample.n39 sample.n38 0.00216539
R32193 sample.n20 sample.n19 0.00216539
R32194 sample.n17 sample.n16 0.00216539
R32195 sample.n134 sample.n133 0.00216539
R32196 sample.n115 sample.n114 0.00216539
R32197 sample.n96 sample.n95 0.00216539
R32198 sample.n74 sample.n58 0.0015031
R32199 sample.n55 sample.n39 0.0015031
R32200 sample.n36 sample.n20 0.0015031
R32201 sample.n16 sample.n15 0.0015031
R32202 sample.n133 sample.n117 0.0015031
R32203 sample.n114 sample.n98 0.0015031
R32204 sample.n95 sample.n79 0.0015031
R32205 sample.n74 sample.n73 0.0011688
R32206 sample.n55 sample.n54 0.0011688
R32207 sample.n36 sample.n35 0.0011688
R32208 sample.n15 sample.n14 0.0011688
R32209 sample.n153 sample.n138 0.0011688
R32210 sample.n131 sample.n117 0.0011688
R32211 sample.n112 sample.n98 0.0011688
R32212 sample.n93 sample.n79 0.0011688
R32213 sample.n153 sample.n137 0.00100797
R32214 trimb4 trimb4.n6 280.863
R32215 trimb4.n0 trimb4.t7 135.841
R32216 trimb4.n2 trimb4.t3 135.841
R32217 trimb4.n2 trimb4.t4 135.52
R32218 trimb4.n3 trimb4.t0 135.52
R32219 trimb4.n4 trimb4.t5 135.52
R32220 trimb4.n5 trimb4.t1 135.52
R32221 trimb4.n1 trimb4.t6 135.52
R32222 trimb4.n0 trimb4.t2 135.52
R32223 trimb4.n1 trimb4.n0 0.321152
R32224 trimb4.n5 trimb4.n4 0.321152
R32225 trimb4.n4 trimb4.n3 0.321152
R32226 trimb4.n3 trimb4.n2 0.321152
R32227 trimb4.n6 trimb4.n1 0.163543
R32228 trimb4.n6 trimb4.n5 0.158109
R32229 comparator_0.trim_1.n4.n10 comparator_0.trim_1.n4.t0 18.7845
R32230 comparator_0.trim_1.n4.n0 comparator_0.trim_1.n4.t4 17.6293
R32231 comparator_0.trim_1.n4.n9 comparator_0.trim_1.n4.t5 17.4005
R32232 comparator_0.trim_1.n4.n9 comparator_0.trim_1.n4.t1 17.4005
R32233 comparator_0.trim_1.n4.n8 comparator_0.trim_1.n4.t6 17.4005
R32234 comparator_0.trim_1.n4.n8 comparator_0.trim_1.n4.t2 17.4005
R32235 comparator_0.trim_1.n4.n12 comparator_0.trim_1.n4.t7 17.4005
R32236 comparator_0.trim_1.n4.n12 comparator_0.trim_1.n4.t3 17.4005
R32237 comparator_0.trim_1.n4.n1 comparator_0.trim_1.n4.t12 2.32979
R32238 comparator_0.trim_1.n4.n3 comparator_0.trim_1.n4.n2 2.24237
R32239 comparator_0.trim_1.n4.n5 comparator_0.trim_1.n4.n4 2.24237
R32240 comparator_0.trim_1.n4.n2 comparator_0.trim_1.n4.n1 2.22512
R32241 comparator_0.trim_1.n4.n6 comparator_0.trim_1.n4.n5 2.22512
R32242 comparator_0.trim_1.n4.n4 comparator_0.trim_1.n4.n3 2.19064
R32243 comparator_0.trim_1.n4 comparator_0.trim_1.n4.t8 1.31712
R32244 comparator_0.trim_1.n4.n14 comparator_0.trim_1.n4.n13 1.01343
R32245 comparator_0.trim_1.n4.n13 comparator_0.trim_1.n4.n11 1.00912
R32246 comparator_0.trim_1.n4.n11 comparator_0.trim_1.n4.n10 0.974638
R32247 comparator_0.trim_1.n4.n14 comparator_0.trim_1.n4 0.953086
R32248 comparator_0.trim_1.n4.n7 comparator_0.trim_1.n4.n6 0.950849
R32249 comparator_0.trim_1.n4.n0 comparator_0.trim_1.n4 0.731478
R32250 comparator_0.trim_1.n4.n14 comparator_0.trim_1.n4.n7 0.703086
R32251 comparator_0.trim_1.n4.n10 comparator_0.trim_1.n4.n9 0.500883
R32252 comparator_0.trim_1.n4.n13 comparator_0.trim_1.n4.n12 0.436228
R32253 comparator_0.trim_1.n4.n11 comparator_0.trim_1.n4.n8 0.436228
R32254 comparator_0.trim_1.n4.n14 comparator_0.trim_1.n4.n0 0.207397
R32255 comparator_0.trim_1.n4.n7 comparator_0.trim_1.n4 0.1255
R32256 comparator_0.trim_1.n4.n6 comparator_0.trim_1.n4.t13 0.0869357
R32257 comparator_0.trim_1.n4.n5 comparator_0.trim_1.n4.t9 0.0869357
R32258 comparator_0.trim_1.n4.n4 comparator_0.trim_1.n4.t15 0.0869357
R32259 comparator_0.trim_1.n4.n3 comparator_0.trim_1.n4.t14 0.0869357
R32260 comparator_0.trim_1.n4.n2 comparator_0.trim_1.n4.t10 0.0869357
R32261 comparator_0.trim_1.n4.n1 comparator_0.trim_1.n4.t11 0.0869357
R32262 comparator_0.trim_1.n4.n7 comparator_0.trim_1.n4 0.0608448
R32263 comparator_0.trim_1.n4 comparator_0.trim_1.n4.n14 0.0608448
R32264 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n1 111.322
R32265 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.n3 50.4671
R32266 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t3 26.5955
R32267 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t5 26.5955
R32268 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t4 24.9236
R32269 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t6 24.9236
R32270 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n5 dac_1.sky130_fd_sc_hd__inv_2_2.Y 13.5685
R32271 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.n4 11.2645
R32272 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.n5 9.41342
R32273 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_2.Y 6.1445
R32274 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_2.Y 4.65505
R32275 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n5 dac_1.sky130_fd_sc_hd__inv_2_2.Y 3.8405
R32276 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.n2 2.0485
R32277 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_2.Y 1.55202
R32278 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t2 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.197458
R32279 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.18982
R32280 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.t2 0.1012
R32281 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.n0 0.0316375
R32282 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.t1 0.00959054
R32283 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t2 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.00959054
R32284 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y.t0 0.00959054
R32285 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n0 111.322
R32286 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y.n2 50.4671
R32287 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t2 26.5955
R32288 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t3 26.5955
R32289 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t4 24.9236
R32290 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t1 24.9236
R32291 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y.n4 13.5995
R32292 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_0.Y 12.0325
R32293 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y.n3 11.2645
R32294 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n5 dac_1.sky130_fd_sc_hd__inv_2_0.Y 8.80626
R32295 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_0.Y 6.1445
R32296 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_0.Y 5.3765
R32297 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_0.Y 4.65505
R32298 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y.n1 2.0485
R32299 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_0.Y 1.55202
R32300 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y.t0 0.127353
R32301 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n5 dac_1.sky130_fd_sc_hd__inv_2_0.Y 0.0465389
R32302 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n5 0.0388945
R32303 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n1 111.322
R32304 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.n3 50.4671
R32305 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t2 26.5955
R32306 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t0 26.5955
R32307 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t1 24.9236
R32308 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t3 24.9236
R32309 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n5 dac_0.sky130_fd_sc_hd__inv_2_8.Y 12.0325
R32310 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.n5 11.5369
R32311 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.n4 11.2645
R32312 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_8.Y 6.1445
R32313 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n5 dac_0.sky130_fd_sc_hd__inv_2_8.Y 5.3765
R32314 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_8.Y 4.65505
R32315 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.n2 2.0485
R32316 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_8.Y 1.55202
R32317 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.t4 0.123153
R32318 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_8.Y 0.114063
R32319 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y.n0 0.0918889
R32320 comparator_0.in.n0 comparator_0.in.t2 29.998
R32321 comparator_0.in.n2 comparator_0.in.t1 17.4323
R32322 comparator_0.in comparator_0.in.t0 17.431
R32323 comparator_0.in.t15 comparator_0.in 16.6643
R32324 comparator_0.in.t6 comparator_0.in 14.0781
R32325 comparator_0.in.t10 comparator_0.in 11.4574
R32326 comparator_0.in.t17 comparator_0.in 10.4986
R32327 comparator_0.in.t7 comparator_0.in 8.89705
R32328 comparator_0.in.t8 comparator_0.in 6.28498
R32329 comparator_0.in.t12 comparator_0.in 4.94368
R32330 comparator_0.in.t15 comparator_0.in 4.25505
R32331 comparator_0.in.t4 comparator_0.in 3.69016
R32332 comparator_0.in.t6 comparator_0.in 3.57323
R32333 comparator_0.in.t10 comparator_0.in 2.88232
R32334 comparator_0.in.t9 comparator_0.in.t3 2.35849
R32335 comparator_0.in.t10 comparator_0.in.t6 2.23767
R32336 comparator_0.in.t18 comparator_0.in.t13 2.22905
R32337 comparator_0.in.t8 comparator_0.in.t7 2.22905
R32338 comparator_0.in.t14 comparator_0.in.t5 2.21181
R32339 comparator_0.in.t7 comparator_0.in 2.20732
R32340 comparator_0.in.t6 comparator_0.in.t15 2.20319
R32341 comparator_0.in.t16 comparator_0.in.t18 2.17733
R32342 comparator_0.in.t7 comparator_0.in.t10 2.17733
R32343 comparator_0.in.t15 comparator_0.in.t12 2.08671
R32344 comparator_0.in.t11 comparator_0.in.t4 2.08671
R32345 comparator_0.in.t4 comparator_0.in.t8 2.06947
R32346 comparator_0.in.t5 comparator_0.in.t17 2.06427
R32347 comparator_0.in.n1 comparator_0.in.t14 1.91194
R32348 comparator_0.in.n0 comparator_0.in.t9 1.75296
R32349 comparator_0.in.t8 comparator_0.in 1.66103
R32350 comparator_0.in.n3 comparator_0.in.n1 1.42291
R32351 comparator_0.in.t11 comparator_0.in 1.07809
R32352 comparator_0.in.t4 comparator_0.in 0.976935
R32353 comparator_0.in comparator_0.in.n3 0.503789
R32354 comparator_0.in comparator_0.in.t11 0.491879
R32355 comparator_0.in.n3 comparator_0.in.n2 0.470895
R32356 comparator_0.in.t13 comparator_0.in.n0 0.459352
R32357 comparator_0.in.n1 comparator_0.in.t16 0.317613
R32358 comparator_0.in.n2 comparator_0.in 0.297615
R32359 comparator_0.in.t11 comparator_0.in 0.288298
R32360 trimb2 trimb2.n0 146.279
R32361 trimb2.n0 trimb2.t0 135.803
R32362 trimb2.n0 trimb2.t1 135.52
R32363 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n0 111.322
R32364 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y.n2 50.4671
R32365 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t1 26.5955
R32366 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t2 26.5955
R32367 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t3 24.9236
R32368 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t0 24.9236
R32369 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_1.Y 13.0565
R32370 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y.n3 11.2645
R32371 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y.n4 9.31437
R32372 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_1.Y 6.1445
R32373 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_1.Y 4.65505
R32374 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_1.Y 4.3525
R32375 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y.n1 2.0485
R32376 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_1.Y 1.55202
R32377 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n6 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n5 0.122545
R32378 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n6 dac_0.sky130_fd_sc_hd__inv_2_1.Y 0.0979204
R32379 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y.n6 0.0328004
R32380 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n3 111.32
R32381 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y.n0 50.4671
R32382 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t4 26.5955
R32383 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t0 26.5955
R32384 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t1 24.9236
R32385 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t3 24.9236
R32386 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y.n2 13.5685
R32387 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y.n1 11.2645
R32388 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_5.Y 6.1445
R32389 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_5.Y 5.7129
R32390 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_5.Y 4.65505
R32391 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_5.Y 3.8405
R32392 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y.t2 3.62224
R32393 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_5.Y 2.0485
R32394 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y.n4 1.55202
R32395 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t2 dac_0.sky130_fd_sc_hd__inv_2_5.Y 0.178636
R32396 ctlp1.n1 ctlp1.t3 212.081
R32397 ctlp1.n2 ctlp1.t2 212.081
R32398 ctlp1.n4 ctlp1 152.97
R32399 ctlp1.n1 ctlp1.t1 139.78
R32400 ctlp1.n2 ctlp1.t0 139.78
R32401 ctlp1.n3 ctlp1.n0 73.5281
R32402 ctlp1.n2 ctlp1.n1 61.346
R32403 ctlp1.n3 ctlp1.n2 25.3953
R32404 ctlp1.n5 ctlp1.n4 9.3005
R32405 ctlp1.n4 ctlp1.n3 7.13769
R32406 ctlp1 ctlp1.n0 2.13383
R32407 ctlp1.n6 ctlp1 1.68065
R32408 ctlp1 ctlp1.n5 0.783662
R32409 ctlp1.n5 ctlp1.n0 0.194439
R32410 ctlp1 ctlp1.n6 0.0225588
R32411 ctlp1.n6 ctlp1 0.0149231
R32412 ctln7.n3 ctln7.t2 212.081
R32413 ctln7.n2 ctln7.t0 212.081
R32414 ctln7.n3 ctln7.t3 139.78
R32415 ctln7.n2 ctln7.t1 139.78
R32416 ctln7.n3 ctln7.n2 61.346
R32417 ctln7.n5 ctln7.n3 38.5428
R32418 ctln7.n5 ctln7.n0 9.30881
R32419 ctln7.n6 ctln7.n5 9.3005
R32420 ctln7.n7 ctln7.n6 9.01417
R32421 ctln7.n4 ctln7 3.23067
R32422 ctln7.n8 ctln7 1.67697
R32423 ctln7.n5 ctln7.n4 1.2812
R32424 ctln7.n7 ctln7.n0 0.0569565
R32425 ctln7.n6 ctln7.n1 0.03175
R32426 ctln7 ctln7.n8 0.0225588
R32427 ctln7.n8 ctln7 0.0149231
R32428 ctln7 ctln7.n7 0.00771154
R32429 ctln7.n4 ctln7.n1 0.00147336
R32430 ctln7.n1 ctln7.n0 0.00100057
R32431 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n3 111.32
R32432 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y.n0 50.4671
R32433 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t4 26.5955
R32434 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t2 26.5955
R32435 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t5 24.9236
R32436 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t3 24.9236
R32437 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y.n2 13.3125
R32438 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y.n1 11.2645
R32439 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_3.Y 11.1343
R32440 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_3.Y 6.1445
R32441 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_3.Y 4.65505
R32442 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_3.Y 4.0965
R32443 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 3.02296
R32444 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_3.Y 2.0485
R32445 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y.n4 1.55202
R32446 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t1 dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.227625
R32447 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t1 0.174201
R32448 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.158396
R32449 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n0 111.322
R32450 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.n2 50.4671
R32451 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t2 26.5955
R32452 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t3 26.5955
R32453 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t4 24.9236
R32454 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t1 24.9236
R32455 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_8.Y 12.0325
R32456 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.n4 11.5369
R32457 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.n3 11.2645
R32458 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_8.Y 6.1445
R32459 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_8.Y 5.3765
R32460 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_8.Y 4.65505
R32461 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.n1 2.0485
R32462 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_8.Y 1.55202
R32463 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.123153
R32464 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.n5 0.122835
R32465 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y.t0 0.114063
R32466 comparator_0.trim_0.n3 comparator_0.trim_0.n3.t7 18.7775
R32467 comparator_0.trim_0.n3 comparator_0.trim_0.n3.t6 17.7991
R32468 comparator_0.trim_0.n3.n0 comparator_0.trim_0.n3.t4 17.4005
R32469 comparator_0.trim_0.n3.n0 comparator_0.trim_0.n3.t5 17.4005
R32470 comparator_0.trim_0.n3.t3 comparator_0.trim_0.n3.t0 2.32781
R32471 comparator_0.trim_0.n3.t1 comparator_0.trim_0.n3.t3 2.22512
R32472 comparator_0.trim_0.n3 comparator_0.trim_0.n3.t1 1.78771
R32473 comparator_0.trim_0.n3 comparator_0.trim_0.n3.t2 0.482237
R32474 comparator_0.trim_0.n3 comparator_0.trim_0.n3.n0 0.460422
R32475 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n0 111.322
R32476 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y.n2 50.4671
R32477 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t1 26.5955
R32478 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t2 26.5955
R32479 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t3 24.9236
R32480 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t4 24.9236
R32481 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_1.Y 13.0565
R32482 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y.n3 11.2645
R32483 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y.n4 9.31437
R32484 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_1.Y 6.1445
R32485 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_1.Y 4.65505
R32486 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_1.Y 4.3525
R32487 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y.n1 2.0485
R32488 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_1.Y 1.55202
R32489 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.117746
R32490 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n6 dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.107011
R32491 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n6 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n5 0.0589115
R32492 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n6 0.0237099
R32493 ctlp7.n0 ctlp7.t0 212.081
R32494 ctlp7.n1 ctlp7.t2 212.081
R32495 ctlp7.n0 ctlp7.t1 139.78
R32496 ctlp7.n1 ctlp7.t3 139.78
R32497 ctlp7.n1 ctlp7.n0 61.346
R32498 ctlp7.n2 ctlp7.n1 37.7187
R32499 ctlp7.n2 ctlp7 2.00759
R32500 ctlp7.n3 ctlp7 1.64021
R32501 ctlp7 ctlp7.n2 0.884093
R32502 ctlp7 ctlp7.n3 0.0225588
R32503 ctlp7.n3 ctlp7 0.0149231
R32504 ctlp2.n1 ctlp2.t3 212.081
R32505 ctlp2.n2 ctlp2.t2 212.081
R32506 ctlp2.n4 ctlp2 152.97
R32507 ctlp2.n1 ctlp2.t1 139.78
R32508 ctlp2.n2 ctlp2.t0 139.78
R32509 ctlp2.n3 ctlp2.n0 73.3576
R32510 ctlp2.n2 ctlp2.n1 61.346
R32511 ctlp2.n3 ctlp2.n2 25.0059
R32512 ctlp2.n5 ctlp2.n4 9.3005
R32513 ctlp2.n4 ctlp2.n3 6.74837
R32514 ctlp2 ctlp2.n0 2.13383
R32515 ctlp2.n6 ctlp2 1.68065
R32516 ctlp2 ctlp2.n5 0.783662
R32517 ctlp2.n5 ctlp2.n0 0.194439
R32518 ctlp2 ctlp2.n6 0.0225588
R32519 ctlp2.n6 ctlp2 0.0149231
R32520 ctln3.n3 ctln3.t0 212.081
R32521 ctln3.n2 ctln3.t2 212.081
R32522 ctln3.n3 ctln3.t1 139.78
R32523 ctln3.n2 ctln3.t3 139.78
R32524 ctln3.n3 ctln3.n2 61.346
R32525 ctln3.n5 ctln3.n3 38.5428
R32526 ctln3.n5 ctln3.n0 9.30881
R32527 ctln3.n6 ctln3.n5 9.3005
R32528 ctln3.n7 ctln3.n6 9.01417
R32529 ctln3.n4 ctln3 3.09989
R32530 ctln3.n8 ctln3 1.65124
R32531 ctln3.n5 ctln3.n4 1.53719
R32532 ctln3.n7 ctln3.n0 0.0569565
R32533 ctln3.n6 ctln3.n1 0.03175
R32534 ctln3 ctln3.n8 0.0225588
R32535 ctln3.n8 ctln3 0.0149231
R32536 ctln3 ctln3.n7 0.00771154
R32537 ctln3.n4 ctln3.n1 0.00148276
R32538 ctln3.n1 ctln3.n0 0.00100057
R32539 ctlp3.n1 ctlp3.t2 212.081
R32540 ctlp3.n2 ctlp3.t1 212.081
R32541 ctlp3.n4 ctlp3 152.97
R32542 ctlp3.n1 ctlp3.t0 139.78
R32543 ctlp3.n2 ctlp3.t3 139.78
R32544 ctlp3.n3 ctlp3.n0 73.5281
R32545 ctlp3.n2 ctlp3.n1 61.346
R32546 ctlp3.n3 ctlp3.n2 25.3953
R32547 ctlp3.n5 ctlp3.n4 9.3005
R32548 ctlp3.n4 ctlp3.n3 7.13769
R32549 ctlp3 ctlp3.n0 2.13383
R32550 ctlp3.n6 ctlp3 1.68065
R32551 ctlp3 ctlp3.n5 0.783662
R32552 ctlp3.n5 ctlp3.n0 0.194439
R32553 ctlp3 ctlp3.n6 0.0225588
R32554 ctlp3.n6 ctlp3 0.0149231
R32555 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n3 111.32
R32556 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y.n0 50.4671
R32557 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t1 26.5955
R32558 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n3 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t0 26.5955
R32559 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t2 24.9236
R32560 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n0 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t3 24.9236
R32561 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y.n2 13.3125
R32562 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y.n1 11.2645
R32563 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_3.Y 11.1343
R32564 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_3.Y 6.1445
R32565 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n1 dac_0.sky130_fd_sc_hd__inv_2_3.Y 4.65505
R32566 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n2 dac_0.sky130_fd_sc_hd__inv_2_3.Y 4.0965
R32567 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y.t4 3.02296
R32568 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n4 dac_0.sky130_fd_sc_hd__inv_2_3.Y 2.0485
R32569 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y.n4 1.55202
R32570 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.123153
R32571 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t4 dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.114063
R32572 ctlp4.n0 ctlp4.t2 212.081
R32573 ctlp4.n1 ctlp4.t1 212.081
R32574 ctlp4.n0 ctlp4.t0 139.78
R32575 ctlp4.n1 ctlp4.t3 139.78
R32576 ctlp4.n1 ctlp4.n0 61.346
R32577 ctlp4.n2 ctlp4.n1 38.3778
R32578 ctlp4.n2 ctlp4 2.00798
R32579 ctlp4.n3 ctlp4 1.68432
R32580 ctlp4 ctlp4.n2 0.8837
R32581 ctlp4 ctlp4.n3 0.0225588
R32582 ctlp4.n3 ctlp4 0.0149231
R32583 trim2.n1 trim2.n0 146.195
R32584 trim2.n0 trim2.t0 135.803
R32585 trim2.n0 trim2.t1 135.52
R32586 trim2.n1 trim2 0.614724
R32587 trim2 trim2.n1 0.209739
R32588 clkc.n0 clkc.t1 144.124
R32589 clkc.n1 clkc.t4 144.066
R32590 clkc.n0 clkc.t3 142.685
R32591 clkc.n1 clkc.t0 142.679
R32592 clkc.n2 clkc.t5 135.874
R32593 clkc.n2 clkc.t2 135.452
R32594 clkc.n3 clkc.n2 10.8919
R32595 clkc.n3 clkc.n1 2.36324
R32596 clkc.n4 clkc.n0 2.36268
R32597 clkc clkc.n4 1.56717
R32598 clkc.n4 clkc.n3 1.50883
R32599 comp.n50 comp.t4 112.225
R32600 comp.n49 comp.t3 107.12
R32601 comp.n36 comp.t1 28.5655
R32602 comp.n49 comp.t0 24.7678
R32603 comp.n10 comp.t2 17.4005
R32604 comp.n16 comp.n15 13.177
R32605 comp.n42 comp.n41 13.177
R32606 comp.n1 comp.n0 9.31767
R32607 comp.n25 comp.n24 9.31767
R32608 comp.n5 comp.n4 9.3005
R32609 comp.n12 comp.n11 9.3005
R32610 comp.n17 comp.n16 9.3005
R32611 comp.n43 comp.n42 9.3005
R32612 comp.n38 comp.n37 9.3005
R32613 comp.n29 comp.n28 9.3005
R32614 comp.n37 comp.n36 9.0206
R32615 comp.n14 comp.n13 9.0005
R32616 comp.n3 comp.n2 9.0005
R32617 comp.n40 comp.n39 9.0005
R32618 comp.n27 comp.n26 9.0005
R32619 comp.n11 comp.n10 8.50005
R32620 comp.n7 comp.n6 3.0005
R32621 comp.n21 comp.n20 3.0005
R32622 comp.n31 comp.n30 3.0005
R32623 comp.n45 comp.n44 3.0005
R32624 comp.n51 comp.n48 2.77388
R32625 comp comp.n51 1.03175
R32626 comp.n48 comp.n47 0.682942
R32627 comp.n48 comp.n23 0.660969
R32628 comp.n51 comp.n50 0.462457
R32629 comp.n50 comp.n49 0.318208
R32630 comp.n19 comp.n18 0.0525833
R32631 comp.n35 comp.n34 0.0525833
R32632 comp.n20 comp.n19 0.0421667
R32633 comp.n44 comp.n35 0.0400833
R32634 comp.n9 comp.n8 0.0395625
R32635 comp.n33 comp.n32 0.0395625
R32636 comp.n14 comp.n12 0.0338333
R32637 comp.n40 comp.n38 0.0338333
R32638 comp.n21 comp.n9 0.03175
R32639 comp.n32 comp.n31 0.03175
R32640 comp.n47 comp.n46 0.03175
R32641 comp.n23 comp.n22 0.0301875
R32642 comp.n8 comp.n7 0.0301875
R32643 comp.n45 comp.n33 0.0301875
R32644 comp.n27 comp.n25 0.0176028
R32645 comp.n3 comp.n1 0.0175994
R32646 comp.n20 comp.n17 0.00675
R32647 comp.n6 comp.n5 0.00675
R32648 comp.n22 comp.n21 0.00675
R32649 comp.n30 comp.n29 0.00675
R32650 comp.n44 comp.n43 0.00675
R32651 comp.n46 comp.n45 0.00675
R32652 comp.n17 comp.n14 0.00258333
R32653 comp.n5 comp.n3 0.00258333
R32654 comp.n29 comp.n27 0.00258333
R32655 comp.n43 comp.n40 0.00258333
R32656 trim3.n0 trim3.t3 135.841
R32657 trim3.n1 trim3.t2 135.841
R32658 trim3.n1 trim3.t1 135.52
R32659 trim3.n0 trim3.t0 135.52
R32660 trim3.n3 trim3.n2 68.9103
R32661 trim3.n3 trim3 0.647821
R32662 trim3 trim3.n3 0.193682
R32663 trim3.n2 trim3.n0 0.168978
R32664 trim3.n2 trim3.n1 0.152674
R32665 ctlp0.n1 ctlp0.t0 212.081
R32666 ctlp0.n2 ctlp0.t3 212.081
R32667 ctlp0.n4 ctlp0 152.776
R32668 ctlp0.n1 ctlp0.t2 139.78
R32669 ctlp0.n2 ctlp0.t1 139.78
R32670 ctlp0.n3 ctlp0.n0 73.1879
R32671 ctlp0.n2 ctlp0.n1 61.346
R32672 ctlp0.n3 ctlp0.n2 24.6151
R32673 ctlp0.n5 ctlp0.n4 9.3005
R32674 ctlp0.n4 ctlp0.n3 6.35747
R32675 ctlp0 ctlp0.n0 2.13383
R32676 ctlp0.n6 ctlp0 1.67697
R32677 ctlp0 ctlp0.n5 1.1018
R32678 ctlp0.n5 ctlp0.n0 0.388379
R32679 ctlp0 ctlp0.n6 0.0225588
R32680 ctlp0.n6 ctlp0 0.0149231
R32681 trimb3.n0 trimb3.t1 135.841
R32682 trimb3.n1 trimb3.t2 135.841
R32683 trimb3.n1 trimb3.t0 135.52
R32684 trimb3.n0 trimb3.t3 135.52
R32685 trimb3 trimb3.n2 68.9784
R32686 trimb3.n2 trimb3.n0 0.168978
R32687 trimb3.n2 trimb3.n1 0.152674
R32688 comparator_0.trim_1.n3.n4 comparator_0.trim_1.n3.t2 18.7775
R32689 comparator_0.trim_1.n3.n5 comparator_0.trim_1.n3.t1 17.7991
R32690 comparator_0.trim_1.n3.n3 comparator_0.trim_1.n3.t0 17.4005
R32691 comparator_0.trim_1.n3.n3 comparator_0.trim_1.n3.t3 17.4005
R32692 comparator_0.trim_1.n3.n1 comparator_0.trim_1.n3.t7 2.32825
R32693 comparator_0.trim_1.n3.n2 comparator_0.trim_1.n3.n1 2.22512
R32694 comparator_0.trim_1.n3 comparator_0.trim_1.n3.n0 2.2074
R32695 comparator_0.trim_1.n3 comparator_0.trim_1.n3.n5 1.14274
R32696 comparator_0.trim_1.n3.n5 comparator_0.trim_1.n3.n4 0.966017
R32697 comparator_0.trim_1.n3.n4 comparator_0.trim_1.n3.n3 0.464714
R32698 comparator_0.trim_1.n3.n0 comparator_0.trim_1.n3.t6 0.1594
R32699 comparator_0.trim_1.n3.n0 comparator_0.trim_1.n3 0.13936
R32700 comparator_0.trim_1.n3.n2 comparator_0.trim_1.n3.t5 0.087375
R32701 comparator_0.trim_1.n3.n1 comparator_0.trim_1.n3.t4 0.087375
R32702 comparator_0.trim_1.n3.n0 comparator_0.trim_1.n3.n2 0.0757832
R32703 comparator_0.ip.n0 comparator_0.ip.t0 29.6956
R32704 comparator_0.ip.n3 comparator_0.ip.t1 17.4323
R32705 comparator_0.ip comparator_0.ip.t2 17.4118
R32706 comparator_0.ip.t4 comparator_0.ip 16.6643
R32707 comparator_0.ip.t3 comparator_0.ip 14.0781
R32708 comparator_0.ip.t16 comparator_0.ip 11.4574
R32709 comparator_0.ip.t6 comparator_0.ip 10.4986
R32710 comparator_0.ip.t14 comparator_0.ip 8.89705
R32711 comparator_0.ip.t10 comparator_0.ip 6.28498
R32712 comparator_0.ip.t17 comparator_0.ip 4.94368
R32713 comparator_0.ip.t4 comparator_0.ip 4.25505
R32714 comparator_0.ip.t18 comparator_0.ip 3.69016
R32715 comparator_0.ip.t3 comparator_0.ip 3.57323
R32716 comparator_0.ip.t16 comparator_0.ip 2.88232
R32717 comparator_0.ip.t5 comparator_0.ip.t9 2.35849
R32718 comparator_0.ip.t16 comparator_0.ip.t3 2.23767
R32719 comparator_0.ip.t12 comparator_0.ip.t8 2.22905
R32720 comparator_0.ip.t10 comparator_0.ip.t14 2.22905
R32721 comparator_0.ip.t7 comparator_0.ip.t11 2.21181
R32722 comparator_0.ip.t14 comparator_0.ip 2.20732
R32723 comparator_0.ip.t3 comparator_0.ip.t4 2.20319
R32724 comparator_0.ip.t13 comparator_0.ip.t12 2.17733
R32725 comparator_0.ip.t14 comparator_0.ip.t16 2.17733
R32726 comparator_0.ip.t4 comparator_0.ip.t17 2.08671
R32727 comparator_0.ip.t15 comparator_0.ip.t18 2.08671
R32728 comparator_0.ip.t18 comparator_0.ip.t10 2.06947
R32729 comparator_0.ip.t11 comparator_0.ip.t6 2.06427
R32730 comparator_0.ip.n1 comparator_0.ip.t7 1.89901
R32731 comparator_0.ip.n0 comparator_0.ip.t5 1.67537
R32732 comparator_0.ip.t10 comparator_0.ip 1.66103
R32733 comparator_0.ip.n2 comparator_0.ip.n1 1.17722
R32734 comparator_0.ip.t15 comparator_0.ip 1.07809
R32735 comparator_0.ip.t18 comparator_0.ip 0.976935
R32736 comparator_0.ip.n3 comparator_0.ip.n2 0.556421
R32737 comparator_0.ip.t8 comparator_0.ip.n0 0.536938
R32738 comparator_0.ip comparator_0.ip.t15 0.491879
R32739 comparator_0.ip.n2 comparator_0.ip 0.418263
R32740 comparator_0.ip.n1 comparator_0.ip.t13 0.330544
R32741 comparator_0.ip comparator_0.ip.n3 0.3005
R32742 comparator_0.ip.t15 comparator_0.ip 0.288298
R32743 trimb0 trimb0.t0 135.525
R32744 trim1.n0 trim1 155.963
R32745 trim1 trim1.t0 135.52
R32746 trim1.n0 trim1 0.550132
R32747 trim1 trim1.n0 0.2505
R32748 ctlp5.n1 ctlp5.t2 212.081
R32749 ctlp5.n2 ctlp5.t0 212.081
R32750 ctlp5.n4 ctlp5 152.97
R32751 ctlp5.n1 ctlp5.t3 139.78
R32752 ctlp5.n2 ctlp5.t1 139.78
R32753 ctlp5.n3 ctlp5.n0 73.3576
R32754 ctlp5.n2 ctlp5.n1 61.346
R32755 ctlp5.n3 ctlp5.n2 25.0059
R32756 ctlp5.n5 ctlp5.n4 9.3005
R32757 ctlp5.n4 ctlp5.n3 6.74837
R32758 ctlp5 ctlp5.n0 2.13383
R32759 ctlp5.n6 ctlp5 1.688
R32760 ctlp5 ctlp5.n5 0.783662
R32761 ctlp5.n5 ctlp5.n0 0.194439
R32762 ctlp5 ctlp5.n6 0.0225588
R32763 ctlp5.n6 ctlp5 0.0149231
R32764 ctln0.n3 ctln0.t2 212.081
R32765 ctln0.n2 ctln0.t0 212.081
R32766 ctln0.n3 ctln0.t3 139.78
R32767 ctln0.n2 ctln0.t1 139.78
R32768 ctln0.n3 ctln0.n2 61.346
R32769 ctln0.n5 ctln0.n3 37.8794
R32770 ctln0.n5 ctln0.n0 9.3127
R32771 ctln0.n6 ctln0.n5 9.3005
R32772 ctln0.n7 ctln0.n6 9.01808
R32773 ctln0.n4 ctln0 3.61245
R32774 ctln0.n8 ctln0 1.6255
R32775 ctln0.n5 ctln0.n4 1.0252
R32776 ctln0.n7 ctln0.n0 0.0569562
R32777 ctln0.n6 ctln0.n1 0.0278438
R32778 ctln0 ctln0.n8 0.0225588
R32779 ctln0.n8 ctln0 0.0149231
R32780 ctln0 ctln0.n7 0.00771154
R32781 ctln0.n4 ctln0.n1 0.00146432
R32782 ctln0.n1 ctln0.n0 0.00100086
R32783 ctln6.n3 ctln6.t1 212.081
R32784 ctln6.n2 ctln6.t0 212.081
R32785 ctln6.n3 ctln6.t3 139.78
R32786 ctln6.n2 ctln6.t2 139.78
R32787 ctln6.n3 ctln6.n2 61.346
R32788 ctln6.n5 ctln6.n3 37.8794
R32789 ctln6.n5 ctln6.n0 9.31076
R32790 ctln6.n6 ctln6.n5 9.3005
R32791 ctln6.n7 ctln6.n6 9.01612
R32792 ctln6.n4 ctln6 3.48667
R32793 ctln6.n8 ctln6 1.66594
R32794 ctln6.n5 ctln6.n4 1.2812
R32795 ctln6.n7 ctln6.n0 0.0569564
R32796 ctln6.n6 ctln6.n1 0.0297969
R32797 ctln6 ctln6.n8 0.0225588
R32798 ctln6.n8 ctln6 0.0149231
R32799 ctln6 ctln6.n7 0.00771154
R32800 ctln6.n4 ctln6.n1 0.00147336
R32801 ctln6.n1 ctln6.n0 0.00100072
R32802 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n3 111.32
R32803 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y.n0 50.4671
R32804 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t2 26.5955
R32805 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n3 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t3 26.5955
R32806 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t4 24.9236
R32807 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n0 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t1 24.9236
R32808 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y.n2 13.5685
R32809 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y.n1 11.2645
R32810 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_5.Y 6.1445
R32811 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_5.Y 5.7129
R32812 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n1 dac_1.sky130_fd_sc_hd__inv_2_5.Y 4.65505
R32813 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n2 dac_1.sky130_fd_sc_hd__inv_2_5.Y 3.8405
R32814 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y.t0 3.62224
R32815 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n4 dac_1.sky130_fd_sc_hd__inv_2_5.Y 2.0485
R32816 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y.n4 1.55202
R32817 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t0 dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.179216
R32818 trim0 trim0.t0 135.525
R32819 trimb1 trimb1.t0 135.52
R32820 ctln2.n3 ctln2.t1 212.081
R32821 ctln2.n2 ctln2.t0 212.081
R32822 ctln2.n3 ctln2.t3 139.78
R32823 ctln2.n2 ctln2.t2 139.78
R32824 ctln2.n3 ctln2.n2 61.346
R32825 ctln2.n5 ctln2.n3 37.8794
R32826 ctln2.n5 ctln2.n0 9.30881
R32827 ctln2.n6 ctln2.n5 9.3005
R32828 ctln2.n7 ctln2.n6 9.01417
R32829 ctln2.n4 ctln2 3.48667
R32830 ctln2.n8 ctln2 1.62918
R32831 ctln2.n5 ctln2.n4 1.2812
R32832 ctln2.n7 ctln2.n0 0.0569565
R32833 ctln2.n6 ctln2.n1 0.03175
R32834 ctln2 ctln2.n8 0.0225588
R32835 ctln2.n8 ctln2 0.0149231
R32836 ctln2 ctln2.n7 0.00771154
R32837 ctln2.n4 ctln2.n1 0.00147336
R32838 ctln2.n1 ctln2.n0 0.00100057
R32839 ctln5.n3 ctln5.t1 212.081
R32840 ctln5.n2 ctln5.t0 212.081
R32841 ctln5.n3 ctln5.t3 139.78
R32842 ctln5.n2 ctln5.t2 139.78
R32843 ctln5.n3 ctln5.n2 61.346
R32844 ctln5.n5 ctln5.n3 38.5428
R32845 ctln5.n5 ctln5.n0 9.30881
R32846 ctln5.n6 ctln5.n5 9.3005
R32847 ctln5.n7 ctln5.n6 9.01417
R32848 ctln5.n4 ctln5 3.23067
R32849 ctln5.n8 ctln5 1.67329
R32850 ctln5.n5 ctln5.n4 1.2812
R32851 ctln5.n7 ctln5.n0 0.0569565
R32852 ctln5.n6 ctln5.n1 0.03175
R32853 ctln5 ctln5.n8 0.0225588
R32854 ctln5.n8 ctln5 0.0149231
R32855 ctln5 ctln5.n7 0.00771154
R32856 ctln5.n4 ctln5.n1 0.00147336
R32857 ctln5.n1 ctln5.n0 0.00100057
R32858 ctlp6.n1 ctlp6.t1 212.081
R32859 ctlp6.n2 ctlp6.t0 212.081
R32860 ctlp6.n4 ctlp6 152.776
R32861 ctlp6.n1 ctlp6.t3 139.78
R32862 ctlp6.n2 ctlp6.t2 139.78
R32863 ctlp6.n3 ctlp6.n0 73.3576
R32864 ctlp6.n2 ctlp6.n1 61.346
R32865 ctlp6.n3 ctlp6.n2 25.0059
R32866 ctlp6.n5 ctlp6.n4 9.3005
R32867 ctlp6.n4 ctlp6.n3 6.74837
R32868 ctlp6 ctlp6.n0 2.13383
R32869 ctlp6.n6 ctlp6 1.65124
R32870 ctlp6 ctlp6.n5 0.945726
R32871 ctlp6.n5 ctlp6.n0 0.388379
R32872 ctlp6 ctlp6.n6 0.0225588
R32873 ctlp6.n6 ctlp6 0.0149231
R32874 ctln4.n3 ctln4.t1 212.081
R32875 ctln4.n2 ctln4.t0 212.081
R32876 ctln4.n3 ctln4.t3 139.78
R32877 ctln4.n2 ctln4.t2 139.78
R32878 ctln4.n3 ctln4.n2 61.346
R32879 ctln4.n5 ctln4.n3 38.5428
R32880 ctln4.n5 ctln4.n0 9.30881
R32881 ctln4.n6 ctln4.n5 9.3005
R32882 ctln4.n7 ctln4.n6 9.01417
R32883 ctln4.n4 ctln4 3.09989
R32884 ctln4.n8 ctln4 1.66962
R32885 ctln4.n5 ctln4.n4 1.53719
R32886 ctln4.n7 ctln4.n0 0.0569565
R32887 ctln4.n6 ctln4.n1 0.03175
R32888 ctln4 ctln4.n8 0.0225588
R32889 ctln4.n8 ctln4 0.0149231
R32890 ctln4 ctln4.n7 0.00771154
R32891 ctln4.n4 ctln4.n1 0.00148276
R32892 ctln4.n1 ctln4.n0 0.00100057
C0 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln3 0.00135f
C1 dac_0.sky130_fd_sc_hd__inv_2_7.Y avdd 0.49f
C2 comparator_0.vp dac_0.carray_0.unitcap_231.cn 0.51f
C3 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_104.cn 0.18f
C4 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_176.cn 0.18f
C5 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_334.cn 0.348f
C6 dac_1.out dac_1.sw_top_0.en_buf 0.678f
C7 avdd ctlp4 0.116f
C8 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_326.cn 0.043f
C9 dac_1.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.trim_0.n3 0.0103f
C10 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_338.cn 0.00213f
C11 ctln7 ctln4 5.84e-20
C12 ctln6 ctln5 0.106f
C13 dac_0.carray_0.unitcap_247.cn dac_0.carray_0.unitcap_239.cn 0.0902f
C14 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_330.cn 0.145f
C15 comparator_0.vp dac_1.carray_0.unitcap_151.cn 0.00925f
C16 dac_1.carray_0.unitcap_152.cn avdd 0.111f
C17 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln5 2.14e-21
C18 avdd trim3 3.8e-19
C19 dac_1.out dac_0.carray_0.unitcap_207.cn 0.00925f
C20 comparator_0.trim_0.n4 avdd 0.0529f
C21 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_199.cn 0.18f
C22 comparator_0.vp ctlp6 5.61e-19
C23 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_239.cn 0.161f
C24 dac_1.out dac_1.carray_0.unitcap_143.cn 0.51f
C25 dac_0.carray_0.unitcap_9.cn sample 0.00958f
C26 comparator_0.vp dac_0.carray_0.unitcap_200.cn 0.514f
C27 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_39.cn 0.18f
C28 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y 3.39e-19
C29 dac_1.carray_0.unitcap_183.cn dac_1.carray_0.unitcap_175.cn 0.0902f
C30 dac_1.out dac_1.sw_top_1.net1 0.302f
C31 dac_1.carray_0.unitcap_12.cn avdd 0.00155f
C32 comparator_0.trim_1.n3 trimb3 0.231f
C33 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.0139f
C34 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp2 0.16f
C35 comparator_0.vp dac_0.carray_0.unitcap_15.cn 0.501f
C36 dac_1.carray_0.unitcap_288.cn dac_1.carray_0.unitcap_256.cn 0.18f
C37 dac_1.carray_0.unitcap_208.cn dac_1.carray_0.unitcap_224.cn 0.0902f
C38 dac_0.carray_0.unitcap_337.cn dac_0.carray_0.unitcap_336.cn 0.18f
C39 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_8.Y 0.00886f
C40 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_88.cn 0.18f
C41 dac_1.carray_0.unitcap_12.cn vinn 0.00544f
C42 comparator_0.ip trimb2 0.0957f
C43 comparator_0.vp dac_0.carray_0.unitcap_215.cn 0.51f
C44 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_160.cn 0.18f
C45 comparator_0.ip dac_0.carray_0.unitcap_334.cn 0.00909f
C46 dac_0.carray_0.unitcap_39.cn dac_0.carray_0.unitcap_63.cn 0.0902f
C47 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y 0.663f
C48 comparator_0.in dac_1.carray_0.unitcap_334.cn 0.00864f
C49 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_255.cn 0.00213f
C50 comparator_0.vp dac_1.carray_0.unitcap_159.cn 0.00925f
C51 dac_1.carray_0.unitcap_324.cn ctln0 0.00176f
C52 dac_1.carray_0.unitcap_128.cn avdd 0.111f
C53 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp5 0.0515f
C54 dac_1.out dac_0.carray_0.unitcap_199.cn 0.00925f
C55 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_7.cn 0.18f
C56 dac_0.sw_top_0.en_buf comparator_0.vp 0.678f
C57 dac_0.carray_0.unitcap_208.cn dac_0.carray_0.unitcap_224.cn 0.0902f
C58 comparator_0.trim_1.n0 comparator_0.outp 0.0181f
C59 comparator_0.outp trimb3 2.12e-19
C60 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_328.cn 0.00139f
C61 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.carray_0.unitcap_328.cn 0.317f
C62 dac_0.carray_0.unitcap_191.cn dac_1.carray_0.unitcap_191.cn 0.128f
C63 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_175.cn 0.18f
C64 dac_1.out dac_1.carray_0.unitcap_119.cn 0.51f
C65 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_247.cn 0.161f
C66 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_1.Y 35.4f
C67 dac_0.carray_0.unitcap_322.cn ctlp4 1.86e-19
C68 comparator_0.vp dac_0.carray_0.unitcap_192.cn 0.514f
C69 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln5 1.78e-19
C70 avdd ctln7 0.118f
C71 comparator_0.trim_0.n2 comparator_0.trim_0.n0 1.16e-19
C72 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_47.cn 0.18f
C73 comparator_0.outp trimb0 0.0437f
C74 dac_0.carray_0.unitcap_31.cn dac_0.carray_0.unitcap_7.cn 0.0902f
C75 dac_1.carray_0.unitcap_80.cn sample 7.14e-19
C76 comparator_0.vp dac_0.carray_0.unitcap_337.cn 0.506f
C77 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_1.out 2.16e-19
C78 dac_0.sky130_fd_sc_hd__inv_2_4.Y avdd 0.223f
C79 dac_1.carray_0.unitcap_23.cn sample 0.00259f
C80 dac_0.sky130_fd_sc_hd__inv_2_5.Y comparator_0.ip 1.73e-19
C81 dac_0.sw_top_1.net1 comparator_0.vp 0.302f
C82 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_144.cn 0.18f
C83 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_64.cn 0.18f
C84 comparator_0.vp dac_0.carray_0.unitcap_191.cn 0.51f
C85 dac_1.out dac_1.sw_top_1.en_buf 0.696f
C86 dac_1.out sample 0.167f
C87 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_331.cn 0.135f
C88 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_328.cn 0.00869f
C89 dac_0.carray_0.unitcap_223.cn dac_0.carray_0.unitcap_247.cn 0.0902f
C90 comparator_0.vp dac_1.carray_0.unitcap_135.cn 0.00925f
C91 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_239.cn 0.00213f
C92 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_31.cn 0.18f
C93 dac_1.carray_0.unitcap_136.cn avdd 0.103f
C94 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_331.cn 0.0064f
C95 dac_1.out dac_0.carray_0.unitcap_175.cn 0.00925f
C96 comparator_0.trim_1.n3 ctlp6 0.00229f
C97 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_183.cn 0.18f
C98 dac_1.sky130_fd_sc_hd__inv_2_1.Y ctln6 0.159f
C99 dac_1.out dac_1.carray_0.unitcap_127.cn 0.51f
C100 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_223.cn 0.161f
C101 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 7.78e-22
C102 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.00124f
C103 comparator_0.vp dac_0.carray_0.unitcap_168.cn 0.514f
C104 dac_0.sky130_fd_sc_hd__inv_2_3.Y avdd 0.23f
C105 dac_1.carray_0.unitcap_167.cn dac_1.carray_0.unitcap_183.cn 0.0902f
C106 comparator_0.trim_1.n1 comparator_0.outp 0.0162f
C107 dac_1.carray_0.unitcap_14.cn avdd 0.00155f
C108 dac_1.carray_0.unitcap_326.cn dac_1.carray_0.unitcap_328.cn 0.18f
C109 dac_1.carray_0.unitcap_72.cn sample 0.00246f
C110 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.554f
C111 dac_0.sw_top_3.net1 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.461f
C112 dac_1.carray_0.unitcap_184.cn dac_1.carray_0.unitcap_208.cn 0.0902f
C113 comparator_0.vp dac_0.carray_0.unitcap_14.cn 0.556f
C114 comparator_0.trim_0.n2 comparator_0.trim_0.n1 0.217f
C115 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln4 0.0827f
C116 dac_1.carray_0.unitcap_15.cn sample 0.0343f
C117 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_152.cn 0.18f
C118 comparator_0.trim_1.n0 trimb0 0.117f
C119 comparator_0.vp dac_0.carray_0.unitcap_207.cn 0.51f
C120 dac_1.carray_0.unitcap_14.cn vinn 0.00135f
C121 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_80.cn 0.18f
C122 dac_0.carray_0.unitcap_47.cn dac_0.carray_0.unitcap_39.cn 0.0902f
C123 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_247.cn 0.00213f
C124 comparator_0.in dac_1.carray_0.unitcap_331.cn 0.00283f
C125 comparator_0.vp dac_1.carray_0.unitcap_143.cn 0.00925f
C126 dac_1.carray_0.unitcap_112.cn avdd 0.112f
C127 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_23.cn 0.18f
C128 comparator_0.diff comparator_0.ip 0.155f
C129 dac_1.out dac_0.carray_0.unitcap_183.cn 0.00925f
C130 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_2.Y 84.2f
C131 dac_0.sw_top_1.en_buf comparator_0.vp 0.696f
C132 dac_0.carray_0.unitcap_184.cn dac_0.carray_0.unitcap_208.cn 0.0902f
C133 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_6.Y 0.00789f
C134 dac_0.carray_0.unitcap_207.cn dac_1.carray_0.unitcap_207.cn 0.128f
C135 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_326.cn 0.00139f
C136 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_167.cn 0.18f
C137 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.carray_0.unitcap_324.cn 0.289f
C138 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.carray_0.unitcap_322.cn 0.137f
C139 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_231.cn 0.161f
C140 dac_1.out dac_1.carray_0.unitcap_103.cn 0.51f
C141 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln2 0.16f
C142 comparator_0.vp dac_0.carray_0.unitcap_176.cn 0.514f
C143 dac_1.sw_top_1.en_buf dac_1.carray_0.unitcap_48.cn 8.31e-19
C144 dac_1.carray_0.unitcap_48.cn sample 0.00246f
C145 comparator_0.vp dac_0.carray_0.unitcap_330.cn 0.502f
C146 dac_0.sky130_fd_sc_hd__inv_2_7.Y ctlp0 0.0476f
C147 dac_0.carray_0.unitcap_23.cn dac_0.carray_0.unitcap_31.cn 0.0902f
C148 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.325f
C149 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_128.cn 0.18f
C150 comparator_0.vp dac_0.carray_0.unitcap_199.cn 0.51f
C151 comparator_0.trim_1.n1 comparator_0.trim_1.n0 0.207f
C152 comparator_0.trim_1.n1 trimb3 0.00122f
C153 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_72.cn 0.18f
C154 dac_1.out dac_1.sw_top_3.en_buf 0.692f
C155 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_330.cn 0.0919f
C156 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_322.cn 0.0046f
C157 dac_1.sky130_fd_sc_hd__inv_2_6.Y ctln2 3.42e-19
C158 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_223.cn 0.181f
C159 dac_0.carray_0.unitcap_231.cn dac_0.carray_0.unitcap_223.cn 0.0902f
C160 comparator_0.vp dac_1.carray_0.unitcap_119.cn 0.00925f
C161 dac_1.carray_0.unitcap_120.cn avdd 0.111f
C162 comparator_0.vp dac_1.sky130_fd_sc_hd__inv_2_1.Y 8.01e-19
C163 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_334.cn 0.00192f
C164 dac_1.sky130_fd_sc_hd__inv_2_6.VPB avdd 0.81f
C165 dac_1.sky130_fd_sc_hd__inv_2_2.Y ctln6 0.00123f
C166 dac_1.out dac_0.carray_0.unitcap_167.cn 0.00925f
C167 comparator_0.trim_1.n4 a_33300_6679# 0.00509f
C168 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 1.29e-23
C169 comparator_0.trim_1.n1 trimb0 0.00397f
C170 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_232.cn 0.18f
C171 avdd ctlp2 0.118f
C172 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_151.cn 0.18f
C173 comparator_0.in clkc 0.372f
C174 dac_1.out dac_1.carray_0.unitcap_111.cn 0.51f
C175 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_215.cn 0.161f
C176 comparator_0.vp dac_0.carray_0.unitcap_160.cn 0.514f
C177 dac_0.sky130_fd_sc_hd__inv_2_8.Y comparator_0.vp 8.84f
C178 dac_1.carray_0.unitcap_151.cn dac_1.carray_0.unitcap_167.cn 0.0902f
C179 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_207.cn 0.18f
C180 dac_1.carray_0.unitcap_56.cn sample 0.0026f
C181 comparator_0.vp dac_0.carray_0.unitcap_12.cn 0.556f
C182 comparator_0.vp sample 0.167f
C183 dac_1.carray_0.unitcap_10.cn dac_1.carray_0.unitcap_288.cn 0.18f
C184 dac_1.carray_0.unitcap_200.cn dac_1.carray_0.unitcap_184.cn 0.0902f
C185 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_48.cn 0.18f
C186 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_0.Y 17.5f
C187 comparator_0.diff trimb4 4.81e-20
C188 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_5.Y 0.00798f
C189 comparator_0.vp dac_0.carray_0.unitcap_175.cn 0.51f
C190 comparator_0.trim_0.n3 trim2 0.00123f
C191 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y 0.357f
C192 comparator_0.in dac_1.carray_0.unitcap_330.cn 0.00277f
C193 comparator_0.vp dac_1.carray_0.unitcap_127.cn 0.00925f
C194 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_231.cn 0.18f
C195 dac_1.carray_0.unitcap_96.cn avdd 0.111f
C196 dac_1.out dac_0.carray_0.unitcap_151.cn 0.00925f
C197 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_336.cn 0.00473f
C198 dac_0.carray_0.unitcap_0.cn sample 0.00246f
C199 comparator_0.trim_1.n4 clkc 0.192f
C200 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp5 1.48e-19
C201 dac_0.sw_top_3.en_buf comparator_0.vp 0.692f
C202 dac_0.carray_0.unitcap_200.cn dac_0.carray_0.unitcap_184.cn 0.0902f
C203 dac_1.out comparator_0.trim_0.n3 0.00137f
C204 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_240.cn 0.18f
C205 dac_0.carray_0.unitcap_199.cn dac_1.carray_0.unitcap_199.cn 0.128f
C206 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_159.cn 0.18f
C207 dac_0.sw_top_0.net1 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.402f
C208 dac_1.carray_0.unitcap_8.cn sample 0.00246f
C209 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_334.cn 0.0395f
C210 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.carray_0.unitcap_324.cn 0.00391f
C211 dac_1.out dac_1.carray_0.unitcap_95.cn 0.51f
C212 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_191.cn 0.161f
C213 comparator_0.ip avdd 0.51f
C214 comparator_0.vp dac_0.carray_0.unitcap_144.cn 0.514f
C215 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp3 0.00135f
C216 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_199.cn 0.18f
C217 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.134f
C218 dac_1.carray_0.unitcap_32.cn sample 0.00246f
C219 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp0 0.00131f
C220 comparator_0.in trim3 0.102f
C221 dac_0.carray_0.unitcap_15.cn dac_0.carray_0.unitcap_23.cn 0.0902f
C222 comparator_0.vp dac_0.carray_0.unitcap_331.cn 0.501f
C223 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln7 2.79e-20
C224 comparator_0.in comparator_0.trim_0.n4 4.85f
C225 dac_0.carray_0.unitcap_322.cn ctlp2 8.69e-19
C226 comparator_0.vp dac_0.carray_0.unitcap_183.cn 0.51f
C227 dac_1.sky130_fd_sc_hd__inv_2_0.Y ctln6 0.0512f
C228 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 1.23e-21
C229 dac_1.out dac_1.sw_top_2.en_buf 0.516f
C230 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_56.cn 0.18f
C231 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_337.cn 0.0902f
C232 comparator_0.in trim0 0.0297f
C233 comparator_0.vp dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.0188f
C234 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.carray_0.unitcap_326.cn 0.00179f
C235 comparator_0.vp dac_1.carray_0.unitcap_103.cn 0.00925f
C236 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_215.cn 0.18f
C237 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_326.cn 8.52e-19
C238 dac_0.carray_0.unitcap_215.cn dac_0.carray_0.unitcap_231.cn 0.0902f
C239 dac_1.out dac_0.carray_0.unitcap_159.cn 0.00925f
C240 dac_1.carray_0.unitcap_322.cn ctln2 8.69e-19
C241 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_338.cn 0.00473f
C242 dac_1.carray_0.unitcap_104.cn avdd 0.0919f
C243 comparator_0.trim_0.n3 ctln6 0.00221f
C244 dac_0.carray_0.unitcap_24.cn sample 0.00277f
C245 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_135.cn 0.18f
C246 dac_1.out dac_1.carray_0.unitcap_71.cn 0.51f
C247 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_207.cn 0.161f
C248 comparator_0.vp dac_0.carray_0.unitcap_152.cn 0.514f
C249 dac_0.sky130_fd_sc_hd__inv_2_2.Y ctlp7 0.16f
C250 dac_0.sky130_fd_sc_hd__inv_2_8.Y comparator_0.trim_1.n3 0.00559f
C251 dac_1.carray_0.unitcap_159.cn dac_1.carray_0.unitcap_151.cn 0.0902f
C252 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_175.cn 0.18f
C253 dac_1.carray_0.unitcap_334.cn dac_1.carray_0.unitcap_326.cn 0.18f
C254 ctln3 ctln2 0.105f
C255 comparator_0.vp dac_0.carray_0.unitcap_13.cn 0.558f
C256 dac_1.carray_0.unitcap_40.cn sample 0.00329f
C257 comparator_0.trim_1.n4 comparator_0.trim_0.n4 0.12f
C258 dac_1.carray_0.unitcap_192.cn dac_1.carray_0.unitcap_200.cn 0.0902f
C259 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_239.cn 0.18f
C260 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.carray_0.unitcap_320.cn 0.00177f
C261 comparator_0.vp dac_0.carray_0.unitcap_167.cn 0.51f
C262 comparator_0.trim_0.n0 trim2 2.84e-19
C263 comparator_0.in ctln7 0.0124f
C264 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_32.cn 0.18f
C265 dac_0.sky130_fd_sc_hd__inv_2_6.Y comparator_0.vp 0.539f
C266 comparator_0.in dac_1.carray_0.unitcap_337.cn 0.00308f
C267 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_191.cn 0.18f
C268 comparator_0.vp dac_1.carray_0.unitcap_111.cn 0.00925f
C269 dac_1.carray_0.unitcap_88.cn avdd 0.111f
C270 dac_1.out dac_0.carray_0.unitcap_135.cn 0.00925f
C271 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_255.cn 0.00473f
C272 comparator_0.diff dac_1.out 0.0419f
C273 avdd trimb4 0.0756f
C274 dac_0.carray_0.unitcap_192.cn dac_0.carray_0.unitcap_200.cn 0.0902f
C275 dac_0.sw_top_2.en_buf comparator_0.vp 0.516f
C276 dac_0.carray_0.unitcap_16.cn sample 0.00246f
C277 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.105f
C278 dac_0.carray_0.unitcap_175.cn dac_1.carray_0.unitcap_175.cn 0.128f
C279 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_331.cn 0.0404f
C280 dac_1.out dac_1.carray_0.unitcap_87.cn 0.51f
C281 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_199.cn 0.161f
C282 comparator_0.vp dac_0.carray_0.unitcap_128.cn 0.514f
C283 clkc trim4 0.00154f
C284 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_183.cn 0.18f
C285 dac_1.sw_top_3.en_buf dac_1.carray_0.unitcap_32.cn 2.32e-19
C286 comparator_0.trim_1.n3 dac_0.carray_0.unitcap_331.cn 0.0174f
C287 comparator_0.vp dac_1.sky130_fd_sc_hd__inv_2_0.Y 1.97e-19
C288 comparator_0.vp dac_0.carray_0.unitcap_334.cn 0.501f
C289 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_247.cn 0.18f
C290 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_40.cn 0.18f
C291 comparator_0.vp dac_0.carray_0.unitcap_151.cn 0.51f
C292 dac_0.carray_0.unitcap_9.cn avdd 0.0125f
C293 avdd ctln1 0.12f
C294 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.carray_0.unitcap_328.cn 0.00101f
C295 dac_1.out ctln4 5.62e-19
C296 dac_0.carray_0.unitcap_191.cn dac_0.carray_0.unitcap_215.cn 0.0902f
C297 dac_1.carray_0.unitcap_64.cn avdd 0.112f
C298 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_328.cn 2e-20
C299 comparator_0.vp dac_1.carray_0.unitcap_95.cn 0.00925f
C300 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_239.cn 0.00473f
C301 comparator_0.outp latch_0.Qn 0.0168f
C302 dac_1.out dac_0.carray_0.unitcap_143.cn 0.00925f
C303 comparator_0.trim_0.n1 trim2 0.0715f
C304 comparator_0.outn clkc 0.259f
C305 dac_0.carray_0.unitcap_328.cn ctlp5 0.00202f
C306 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_175.cn 0.161f
C307 dac_1.out dac_1.carray_0.unitcap_79.cn 0.51f
C308 dac_0.sw_top_0.en_buf dac_0.sw_top_1.net1 4.9e-19
C309 comparator_0.vp dac_0.carray_0.unitcap_136.cn 0.514f
C310 dac_0.sky130_fd_sc_hd__inv_2_6.VPB avdd 0.918f
C311 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_167.cn 0.18f
C312 dac_0.sky130_fd_sc_hd__inv_2_5.Y comparator_0.vp 2.01f
C313 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.00798f
C314 dac_1.carray_0.unitcap_135.cn dac_1.carray_0.unitcap_159.cn 0.0902f
C315 comparator_0.trim_1.n2 clkc 5.88e-20
C316 dac_0.sky130_fd_sc_hd__inv_2_1.Y avdd 0.365f
C317 dac_0.carray_0.unitcap_14.cn dac_0.carray_0.unitcap_15.cn 0.18f
C318 dac_1.carray_0.unitcap_11.cn dac_1.carray_0.unitcap_10.cn 0.18f
C319 comparator_0.vp dac_0.carray_0.unitcap_11.cn 0.556f
C320 dac_1.carray_0.unitcap_168.cn dac_1.carray_0.unitcap_192.cn 0.0902f
C321 dac_0.sw_top_2.en_buf dac_0.carray_0.unitcap_24.cn 6.3e-19
C322 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_338.cn 0.18f
C323 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln2 4.16e-20
C324 trim4 trim3 0.0218f
C325 avdd ctlp5 0.116f
C326 comparator_0.vp dac_0.carray_0.unitcap_159.cn 0.51f
C327 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_338.cn 0.18f
C328 comparator_0.trim_0.n4 trim4 0.359f
C329 dac_0.carray_0.unitcap_320.cn avdd 0.0981f
C330 ctln6 ctln4 1.34e-20
C331 comparator_0.in dac_1.carray_0.unitcap_336.cn 0.00468f
C332 comparator_0.vp dac_1.carray_0.unitcap_71.cn 0.00925f
C333 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln4 5.67e-19
C334 avdd trim2 4.46e-19
C335 comparator_0.in comparator_0.trim_0.n2 1.18f
C336 dac_1.out dac_0.carray_0.unitcap_119.cn 0.00925f
C337 dac_1.carray_0.unitcap_80.cn avdd 0.0709f
C338 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_247.cn 0.00473f
C339 dac_0.sw_top_2.net1 sample 0.0371f
C340 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_6.Y 0.00789f
C341 dac_0.carray_0.unitcap_168.cn dac_0.carray_0.unitcap_192.cn 0.0902f
C342 comparator_0.vp vinp 9.61f
C343 dac_0.carray_0.unitcap_183.cn dac_1.carray_0.unitcap_183.cn 0.128f
C344 dac_1.out dac_1.carray_0.unitcap_55.cn 0.51f
C345 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_183.cn 0.161f
C346 comparator_0.vp dac_0.carray_0.unitcap_112.cn 0.514f
C347 dac_1.out avdd 6.18f
C348 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_151.cn 0.18f
C349 comparator_0.trim_1.n3 trimb2 0.00123f
C350 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp3 0.0494f
C351 comparator_0.outn trim3 9.68e-20
C352 comparator_0.trim_1.n3 dac_0.carray_0.unitcap_334.cn 0.0151f
C353 dac_1.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.in 0.0266f
C354 dac_0.carray_0.unitcap_23.cn sample 0.00259f
C355 comparator_0.vp dac_0.carray_0.unitcap_326.cn 0.501f
C356 dac_0.sw_top_3.en_buf dac_0.sw_top_2.net1 4.9e-19
C357 dac_0.sw_top_1.en_buf dac_0.sw_top_0.en_buf 0.00289f
C358 comparator_0.outn comparator_0.trim_0.n4 0.804f
C359 dac_1.out vinn 9.61f
C360 comparator_0.ip trimb1 0.0878f
C361 comparator_0.vp comparator_0.diff 0.0502f
C362 comparator_0.vp dac_0.carray_0.unitcap_135.cn 0.51f
C363 comparator_0.outn trim0 0.00216f
C364 dac_0.carray_0.unitcap_321.cn avdd 0.0672f
C365 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.carray_0.unitcap_322.cn 0.001f
C366 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.29e-23
C367 comparator_0.vp dac_1.carray_0.unitcap_87.cn 0.00925f
C368 dac_0.carray_0.unitcap_207.cn dac_0.carray_0.unitcap_191.cn 0.0902f
C369 dac_0.sky130_fd_sc_hd__inv_2_0.Y ctlp7 2.65e-19
C370 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp6 2.22e-19
C371 dac_1.out dac_0.carray_0.unitcap_127.cn 0.00925f
C372 dac_1.carray_0.unitcap_72.cn avdd 0.112f
C373 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_223.cn 0.00473f
C374 comparator_0.outp trimb2 0.0102f
C375 dac_1.carray_0.unitcap_7.cn dac_1.carray_0.unitcap_47.cn 0.0902f
C376 dac_0.sw_top_1.en_buf dac_0.sw_top_1.net1 0.585f
C377 avdd ctln6 0.116f
C378 dac_1.out dac_1.carray_0.unitcap_63.cn 0.51f
C379 dac_1.carray_0.unitcap_15.cn avdd 0.00155f
C380 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_167.cn 0.161f
C381 dac_0.carray_0.unitcap_9.cn dac_0.carray_0.unitcap_256.cn 0.18f
C382 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln4 0.0503f
C383 dac_1.sky130_fd_sc_hd__inv_2_4.Y avdd 0.226f
C384 comparator_0.vp dac_0.carray_0.unitcap_120.cn 0.514f
C385 dac_0.sky130_fd_sc_hd__inv_2_5.Y comparator_0.trim_1.n3 1.4e-19
C386 dac_1.carray_0.unitcap_143.cn dac_1.carray_0.unitcap_135.cn 0.0902f
C387 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_159.cn 0.18f
C388 comparator_0.outp comparator_0.trim_0.n3 5.99e-20
C389 comparator_0.vp dac_0.carray_0.unitcap_10.cn 0.557f
C390 dac_0.carray_0.unitcap_330.cn dac_0.carray_0.unitcap_337.cn 0.18f
C391 dac_1.sw_top_2.net1 sample 0.0371f
C392 dac_1.carray_0.unitcap_331.cn dac_1.carray_0.unitcap_334.cn 0.18f
C393 dac_0.carray_0.unitcap_15.cn sample 0.0343f
C394 dac_1.carray_0.unitcap_176.cn dac_1.carray_0.unitcap_168.cn 0.0902f
C395 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.134f
C396 comparator_0.vp dac_0.carray_0.unitcap_143.cn 0.51f
C397 dac_0.carray_0.unitcap_248.cn avdd 0.095f
C398 comparator_0.ip comparator_0.in 0.254f
C399 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln7 2.25e-19
C400 dac_1.carray_0.unitcap_48.cn avdd 0.111f
C401 comparator_0.vp dac_1.carray_0.unitcap_79.cn 0.00925f
C402 dac_1.out dac_0.carray_0.unitcap_103.cn 0.00925f
C403 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_231.cn 0.00473f
C404 dac_0.sw_top_0.en_buf sample 0.485f
C405 dac_0.carray_0.unitcap_176.cn dac_0.carray_0.unitcap_168.cn 0.0902f
C406 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.carray_0.unitcap_322.cn 0.001f
C407 dac_1.sky130_fd_sc_hd__inv_2_1.Y ctln5 0.00139f
C408 dac_0.carray_0.unitcap_167.cn dac_1.carray_0.unitcap_167.cn 0.128f
C409 dac_1.sw_top_0.en_buf dac_1.sw_top_1.net1 4.9e-19
C410 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_151.cn 0.161f
C411 dac_1.out dac_1.carray_0.unitcap_39.cn 0.51f
C412 comparator_0.vp dac_0.carray_0.unitcap_96.cn 0.514f
C413 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_135.cn 0.18f
C414 comparator_0.trim_1.n0 trimb2 2.84e-19
C415 trimb3 trimb2 0.0356f
C416 comparator_0.vp dac_0.carray_0.unitcap_328.cn 0.501f
C417 dac_0.sw_top_2.en_buf dac_0.sw_top_2.net1 0.585f
C418 dac_0.sky130_fd_sc_hd__inv_2_0.Y ctlp4 0.00127f
C419 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln3 0.0829f
C420 dac_1.sky130_fd_sc_hd__inv_2_3.Y avdd 0.233f
C421 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_336.cn 0.00473f
C422 comparator_0.trim_1.n4 comparator_0.ip 4.88f
C423 dac_0.sw_top_1.net1 sample 0.037f
C424 trimb2 trimb0 7.61e-19
C425 comparator_0.vp dac_0.carray_0.unitcap_119.cn 0.51f
C426 dac_1.sw_top_2.net1 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.358f
C427 dac_0.carray_0.unitcap_232.cn avdd 0.095f
C428 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.carray_0.unitcap_324.cn 8.63e-19
C429 dac_1.out dac_1.carray_0.unitcap_320.cn 0.496f
C430 dac_0.carray_0.unitcap_199.cn dac_0.carray_0.unitcap_207.cn 0.0902f
C431 dac_1.sky130_fd_sc_hd__inv_2_7.Y avdd 0.353f
C432 dac_1.carray_0.unitcap_56.cn avdd 0.0854f
C433 comparator_0.vp dac_1.carray_0.unitcap_55.cn 0.00925f
C434 dac_1.out dac_0.carray_0.unitcap_111.cn 0.00925f
C435 comparator_0.vp avdd 5.39f
C436 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_215.cn 0.00473f
C437 comparator_0.trim_0.n2 trim4 0.00188f
C438 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln1 0.00126f
C439 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_159.cn 0.161f
C440 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp0 0.0827f
C441 dac_1.out dac_1.carray_0.unitcap_47.cn 0.51f
C442 dac_0.carray_0.unitcap_320.cn dac_0.carray_0.unitcap_324.cn 0.18f
C443 comparator_0.vp dac_0.carray_0.unitcap_104.cn 0.514f
C444 dac_1.carray_0.unitcap_326.cn ctln7 0.00199f
C445 comparator_0.outp comparator_0.diff 0.002f
C446 dac_1.carray_0.unitcap_119.cn dac_1.carray_0.unitcap_143.cn 0.0902f
C447 dac_0.carray_0.unitcap_12.cn dac_0.carray_0.unitcap_14.cn 0.18f
C448 dac_1.carray_0.unitcap_13.cn dac_1.carray_0.unitcap_11.cn 0.18f
C449 dac_1.sw_top_1.en_buf dac_1.sw_top_0.en_buf 0.00289f
C450 dac_1.sw_top_3.en_buf dac_1.sw_top_2.net1 4.9e-19
C451 dac_0.sky130_fd_sc_hd__inv_2_7.Y ctlp1 3.56e-20
C452 dac_1.sw_top_0.en_buf sample 0.485f
C453 dac_0.carray_0.unitcap_14.cn sample 0.0343f
C454 comparator_0.vp dac_0.carray_0.unitcap_288.cn 0.558f
C455 ctlp0 ctlp5 7.15e-20
C456 dac_1.carray_0.unitcap_160.cn dac_1.carray_0.unitcap_176.cn 0.0902f
C457 dac_0.carray_0.unitcap_0.cn avdd 0.0965f
C458 dac_1.carray_0.unitcap_8.cn avdd 0.113f
C459 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_338.cn 0.00473f
C460 dac_1.sky130_fd_sc_hd__inv_2_6.VPB trim4 8.6e-19
C461 comparator_0.trim_1.n1 trimb2 0.0715f
C462 comparator_0.vp dac_0.carray_0.unitcap_127.cn 0.51f
C463 dac_0.carray_0.unitcap_240.cn avdd 0.0893f
C464 dac_1.sky130_fd_sc_hd__inv_2_6.Y ctln1 0.0498f
C465 dac_1.out dac_1.carray_0.unitcap_321.cn 0.512f
C466 comparator_0.vp dac_1.carray_0.unitcap_63.cn 0.00925f
C467 comparator_0.outn comparator_0.trim_0.n2 0.00406f
C468 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_191.cn 0.00473f
C469 dac_1.carray_0.unitcap_32.cn avdd 0.113f
C470 dac_1.out dac_0.carray_0.unitcap_95.cn 0.00925f
C471 dac_0.sw_top_1.en_buf sample 0.561f
C472 dac_0.carray_0.unitcap_160.cn dac_0.carray_0.unitcap_176.cn 0.0902f
C473 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.carray_0.unitcap_328.cn 0.00101f
C474 avdd ctlp3 0.116f
C475 dac_1.sw_top_1.en_buf dac_1.sw_top_1.net1 0.585f
C476 dac_0.carray_0.unitcap_151.cn dac_1.carray_0.unitcap_151.cn 0.128f
C477 dac_1.sw_top_1.net1 sample 0.037f
C478 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_135.cn 0.161f
C479 comparator_0.vp dac_0.carray_0.unitcap_88.cn 0.514f
C480 comparator_0.trim_1.n4 trimb4 0.359f
C481 dac_0.sky130_fd_sc_hd__inv_2_2.Y comparator_0.ip 0.095f
C482 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y 1.23e-21
C483 comparator_0.vp dac_0.carray_0.unitcap_322.cn 0.502f
C484 dac_0.carray_0.unitcap_24.cn avdd 0.0856f
C485 dac_0.sw_top_3.en_buf dac_0.sw_top_1.en_buf 0.00289f
C486 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_5.Y 2.01f
C487 dac_0.sw_top_2.net1 vinp 0.368f
C488 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_255.cn 0.00473f
C489 dac_1.carray_0.unitcap_324.cn avdd 0.0115f
C490 comparator_0.vp dac_0.carray_0.unitcap_103.cn 0.51f
C491 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.00886f
C492 dac_0.carray_0.unitcap_216.cn avdd 0.0957f
C493 comparator_0.trim_0.n3 trim1 4.9e-20
C494 dac_1.sw_top_0.en_buf dac_1.sky130_fd_sc_hd__inv_2_2.Y 1.27f
C495 dac_1.out dac_1.carray_0.unitcap_248.cn 0.514f
C496 comparator_0.vp dac_1.carray_0.unitcap_39.cn 0.00925f
C497 dac_1.carray_0.unitcap_40.cn avdd 0.111f
C498 dac_0.carray_0.unitcap_175.cn dac_0.carray_0.unitcap_199.cn 0.0902f
C499 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_207.cn 0.00473f
C500 a_33300_6679# clkc 0.0762f
C501 comparator_0.trim_1.n3 avdd 0.0396f
C502 dac_1.out dac_0.carray_0.unitcap_71.cn 0.00925f
C503 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp6 5.79e-19
C504 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y 0.105f
C505 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_143.cn 0.18f
C506 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_6.Y 0.539f
C507 comparator_0.vp dac_0.carray_0.unitcap_64.cn 0.514f
C508 dac_1.carray_0.unitcap_127.cn dac_1.carray_0.unitcap_119.cn 0.0902f
C509 dac_1.sw_top_1.net1 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.424f
C510 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp1 0.159f
C511 comparator_0.in trim2 0.0957f
C512 dac_0.carray_0.unitcap_12.cn sample 0.0343f
C513 dac_1.sky130_fd_sc_hd__inv_2_7.Y dac_1.carray_0.unitcap_320.cn 0.119f
C514 dac_1.sw_top_2.en_buf dac_1.sw_top_2.net1 0.585f
C515 comparator_0.vp dac_0.carray_0.unitcap_256.cn 0.557f
C516 dac_1.carray_0.unitcap_330.cn dac_1.carray_0.unitcap_331.cn 0.18f
C517 dac_0.carray_0.unitcap_331.cn dac_0.carray_0.unitcap_330.cn 0.18f
C518 dac_1.sw_top_1.en_buf sample 0.561f
C519 dac_1.carray_0.unitcap_144.cn dac_1.carray_0.unitcap_160.cn 0.0902f
C520 dac_0.carray_0.unitcap_322.cn ctlp3 0.00202f
C521 dac_0.carray_0.unitcap_16.cn avdd 0.0966f
C522 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln6 5.79e-19
C523 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 0.736f
C524 comparator_0.outp avdd 1.03f
C525 dac_1.sky130_fd_sc_hd__inv_2_0.Y ctln5 0.16f
C526 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_239.cn 0.00473f
C527 dac_0.carray_0.unitcap_8.cn dac_0.carray_0.unitcap_9.cn 0.18f
C528 comparator_0.vp dac_0.carray_0.unitcap_111.cn 0.51f
C529 dac_0.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.trim_1.n4 5.74e-21
C530 comparator_0.ip comparator_0.outn 0.0302f
C531 dac_1.out comparator_0.in 0.25f
C532 dac_0.carray_0.unitcap_224.cn avdd 0.095f
C533 dac_0.sky130_fd_sc_hd__inv_2_1.Y comparator_0.trim_1.n4 0.00288f
C534 dac_1.out dac_1.carray_0.unitcap_232.cn 0.514f
C535 comparator_0.vp dac_1.carray_0.unitcap_47.cn 0.00925f
C536 dac_1.out dac_0.carray_0.unitcap_87.cn 0.00925f
C537 dac_0.sw_top_2.net1 dac_0.carray_0.unitcap_10.cn 0.00207f
C538 comparator_0.trim_1.n2 comparator_0.ip 1.18f
C539 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_199.cn 0.00473f
C540 dac_0.sw_top_3.en_buf sample 0.561f
C541 dac_0.carray_0.unitcap_144.cn dac_0.carray_0.unitcap_160.cn 0.0902f
C542 comparator_0.trim_0.n3 ctln5 0.00158f
C543 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.carray_0.unitcap_326.cn 0.00179f
C544 dac_0.carray_0.unitcap_159.cn dac_1.carray_0.unitcap_159.cn 0.128f
C545 dac_0.sky130_fd_sc_hd__inv_2_2.Y trimb4 0.00591f
C546 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y 4.21f
C547 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_119.cn 0.18f
C548 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.sky130_fd_sc_hd__inv_2_6.Y 0.571f
C549 comparator_0.vp dac_0.carray_0.unitcap_80.cn 0.514f
C550 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_331.cn 0.0404f
C551 dac_1.out dac_1.carray_0.unitcap_9.cn 0.557f
C552 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_337.cn 0.0902f
C553 ctlp4 ctlp7 5.84e-20
C554 latch_0.Qn a_33300_5579# 0.0695f
C555 dac_1.sky130_fd_sc_hd__inv_2_7.Y dac_1.carray_0.unitcap_321.cn 0.18f
C556 comparator_0.vp dac_0.carray_0.unitcap_324.cn 0.505f
C557 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y 3.39e-19
C558 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_247.cn 0.00473f
C559 dac_1.out dac_1.carray_0.unitcap_0.cn 0.514f
C560 dac_0.sw_top_0.en_buf vinp 0.417f
C561 comparator_0.trim_1.n4 dac_1.out 0.00632f
C562 comparator_0.vp dac_0.carray_0.unitcap_95.cn 0.51f
C563 comparator_0.trim_0.n0 trim1 0.0594f
C564 comparator_0.in ctln6 0.00359f
C565 dac_0.carray_0.unitcap_208.cn avdd 0.0949f
C566 dac_1.sw_top_1.en_buf dac_1.sky130_fd_sc_hd__inv_2_2.Y 1.04f
C567 dac_1.sky130_fd_sc_hd__inv_2_2.Y sample 2.53f
C568 comparator_0.vp ctlp0 6.77e-19
C569 dac_1.out dac_1.carray_0.unitcap_240.cn 0.514f
C570 dac_0.carray_0.unitcap_183.cn dac_0.carray_0.unitcap_175.cn 0.0902f
C571 comparator_0.trim_1.n0 avdd 0.041f
C572 avdd trimb3 0.0585f
C573 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y 1.12f
C574 dac_1.out dac_0.carray_0.unitcap_79.cn 0.00925f
C575 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_175.cn 0.00473f
C576 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_9.cn 0.0902f
C577 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_239.cn 0.18f
C578 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_127.cn 0.18f
C579 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_248.cn 0.18f
C580 dac_1.carray_0.unitcap_324.cn dac_1.carray_0.unitcap_320.cn 0.18f
C581 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_7.Y 2.23e-21
C582 comparator_0.vp dac_0.carray_0.unitcap_72.cn 0.514f
C583 dac_0.sw_top_1.net1 vinp 0.368f
C584 clkc trim3 0.00176f
C585 avdd trimb0 0.172f
C586 dac_1.out dac_1.carray_0.unitcap_322.cn 0.502f
C587 dac_1.carray_0.unitcap_103.cn dac_1.carray_0.unitcap_127.cn 0.0902f
C588 comparator_0.trim_0.n4 clkc 0.0822f
C589 dac_1.sw_top_3.en_buf dac_1.sw_top_1.en_buf 0.00289f
C590 dac_1.carray_0.unitcap_12.cn dac_1.carray_0.unitcap_13.cn 0.18f
C591 dac_0.carray_0.unitcap_13.cn dac_0.carray_0.unitcap_12.cn 0.18f
C592 dac_0.sw_top_2.net1 avdd 0.844f
C593 dac_1.sw_top_3.en_buf sample 0.561f
C594 dac_0.carray_0.unitcap_13.cn sample 0.0343f
C595 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.0152f
C596 dac_1.carray_0.unitcap_152.cn dac_1.carray_0.unitcap_144.cn 0.0902f
C597 clkc trim0 8.72e-20
C598 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_6.Y 0.0961f
C599 dac_1.out dac_1.carray_0.unitcap_24.cn 0.514f
C600 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_223.cn 0.00473f
C601 comparator_0.vp dac_0.carray_0.unitcap_71.cn 0.51f
C602 comparator_0.trim_1.n2 trimb4 0.00188f
C603 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 4.21f
C604 dac_0.carray_0.unitcap_184.cn avdd 0.0768f
C605 avdd ctln0 0.124f
C606 dac_1.out dac_1.carray_0.unitcap_216.cn 0.514f
C607 ctlp1 ctlp2 0.106f
C608 dac_1.out ctln3 9.29e-19
C609 dac_1.sky130_fd_sc_hd__inv_2_6.Y dac_1.sky130_fd_sc_hd__inv_2_7.Y 0.543f
C610 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y 3.32f
C611 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_183.cn 0.00473f
C612 dac_1.out dac_0.carray_0.unitcap_55.cn 0.00925f
C613 dac_0.sw_top_2.en_buf sample 0.621f
C614 dac_0.carray_0.unitcap_152.cn dac_0.carray_0.unitcap_144.cn 0.0902f
C615 comparator_0.trim_0.n1 trim1 0.184f
C616 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_247.cn 0.18f
C617 dac_0.carray_0.unitcap_14.cn vinp 0.00135f
C618 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_3.Y 4.08e-19
C619 dac_0.carray_0.unitcap_328.cn ctlp6 0.00108f
C620 dac_0.carray_0.unitcap_135.cn dac_1.carray_0.unitcap_135.cn 0.128f
C621 dac_0.sky130_fd_sc_hd__inv_2_0.Y comparator_0.ip 0.0123f
C622 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_103.cn 0.18f
C623 comparator_0.trim_0.n4 dac_1.carray_0.unitcap_330.cn 0.00503f
C624 comparator_0.trim_0.n3 dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.00672f
C625 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_334.cn 0.0395f
C626 comparator_0.vp dac_0.carray_0.unitcap_48.cn 0.514f
C627 comparator_0.trim_1.n1 avdd 0.0161f
C628 dac_1.out dac_1.carray_0.unitcap_256.cn 0.557f
C629 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.carray_0.unitcap_322.cn 0.137f
C630 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp7 5.61e-22
C631 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_330.cn 0.0919f
C632 comparator_0.vp comparator_0.in 0.0157f
C633 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.out 0.0185f
C634 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln1 5.89e-21
C635 dac_0.sw_top_2.en_buf dac_0.sw_top_3.en_buf 0.00289f
C636 dac_1.out dac_1.carray_0.unitcap_16.cn 0.515f
C637 dac_0.sw_top_1.en_buf vinp 0.705f
C638 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_231.cn 0.00473f
C639 avdd ctlp6 0.116f
C640 comparator_0.vp dac_0.carray_0.unitcap_87.cn 0.51f
C641 dac_1.sw_top_3.en_buf dac_1.sky130_fd_sc_hd__inv_2_2.Y 1.15f
C642 comparator_0.trim_0.n4 trim3 0.0166f
C643 dac_0.carray_0.unitcap_200.cn avdd 0.095f
C644 ctln5 ctln4 0.106f
C645 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln3 1.86e-19
C646 dac_1.out dac_1.carray_0.unitcap_224.cn 0.514f
C647 dac_0.carray_0.unitcap_167.cn dac_0.carray_0.unitcap_183.cn 0.0902f
C648 dac_1.out trim4 0.00119f
C649 dac_1.out dac_0.carray_0.unitcap_63.cn 0.00925f
C650 dac_0.carray_0.unitcap_15.cn avdd 0.00155f
C651 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp7 1.78e-19
C652 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_167.cn 0.00473f
C653 dac_1.sw_top_2.net1 avdd 0.844f
C654 comparator_0.trim_0.n4 trim0 0.00934f
C655 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_111.cn 0.18f
C656 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y 0.246f
C657 comparator_0.vp dac_0.carray_0.unitcap_56.cn 0.514f
C658 dac_1.sw_top_2.net1 vinn 0.368f
C659 dac_1.out dac_1.carray_0.unitcap_328.cn 0.501f
C660 comparator_0.trim_1.n3 trimb1 4.9e-20
C661 dac_1.carray_0.unitcap_111.cn dac_1.carray_0.unitcap_103.cn 0.0902f
C662 comparator_0.outn trim2 0.00254f
C663 comparator_0.vp comparator_0.trim_1.n4 0.0361f
C664 dac_1.sw_top_2.en_buf sample 0.621f
C665 dac_0.carray_0.unitcap_11.cn sample 0.0348f
C666 dac_1.carray_0.unitcap_337.cn dac_1.carray_0.unitcap_330.cn 0.18f
C667 dac_0.carray_0.unitcap_334.cn dac_0.carray_0.unitcap_331.cn 0.18f
C668 dac_1.carray_0.unitcap_128.cn dac_1.carray_0.unitcap_152.cn 0.0902f
C669 dac_0.sw_top_0.en_buf avdd 1.98f
C670 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_215.cn 0.00473f
C671 dac_1.sky130_fd_sc_hd__inv_2_6.Y dac_1.carray_0.unitcap_324.cn 0.173f
C672 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_322.cn 0.0046f
C673 dac_1.out comparator_0.outn 0.0121f
C674 comparator_0.vp dac_0.carray_0.unitcap_79.cn 0.51f
C675 dac_1.carray_0.unitcap_9.cn dac_1.carray_0.unitcap_8.cn 0.18f
C676 dac_0.carray_0.unitcap_192.cn avdd 0.095f
C677 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y 0.554f
C678 dac_0.sky130_fd_sc_hd__inv_2_0.Y trimb4 7.19e-19
C679 dac_1.out dac_1.carray_0.unitcap_208.cn 0.514f
C680 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_8.Y 8.84f
C681 comparator_0.vp dac_0.carray_0.unitcap_8.cn 0.503f
C682 comparator_0.outp trimb1 0.0065f
C683 dac_1.out dac_0.carray_0.unitcap_39.cn 0.00925f
C684 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_151.cn 0.00473f
C685 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.sky130_fd_sc_hd__inv_2_4.Y 0.00132f
C686 dac_0.carray_0.unitcap_128.cn dac_0.carray_0.unitcap_152.cn 0.0902f
C687 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp4 5.67e-19
C688 dac_0.carray_0.unitcap_12.cn vinp 0.00544f
C689 sample vinp 0.0271f
C690 comparator_0.trim_0.n3 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.0576f
C691 dac_0.carray_0.unitcap_143.cn dac_1.carray_0.unitcap_143.cn 0.128f
C692 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_95.cn 0.18f
C693 comparator_0.trim_0.n4 dac_1.carray_0.unitcap_337.cn 0.0275f
C694 dac_0.sw_top_1.net1 avdd 0.849f
C695 avdd ctln5 0.116f
C696 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln3 0.161f
C697 dac_1.carray_0.unitcap_328.cn ctln6 0.00108f
C698 comparator_0.vp dac_0.carray_0.unitcap_32.cn 0.514f
C699 dac_1.out dac_1.carray_0.unitcap_288.cn 0.558f
C700 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_326.cn 0.00139f
C701 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.carray_0.unitcap_328.cn 0.317f
C702 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_331.cn 0.135f
C703 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_336.cn 0.161f
C704 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.0925f
C705 dac_0.sw_top_3.en_buf vinp 0.705f
C706 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_191.cn 0.00473f
C707 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp4 0.0503f
C708 comparator_0.vp dac_0.carray_0.unitcap_55.cn 0.51f
C709 comparator_0.trim_0.n2 clkc 5.56e-20
C710 dac_0.carray_0.unitcap_168.cn avdd 0.0611f
C711 dac_1.sw_top_2.en_buf dac_1.sky130_fd_sc_hd__inv_2_2.Y 1.16f
C712 dac_1.out dac_1.carray_0.unitcap_184.cn 0.514f
C713 dac_0.carray_0.unitcap_151.cn dac_0.carray_0.unitcap_167.cn 0.0902f
C714 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln6 2.22e-19
C715 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_159.cn 0.00473f
C716 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 3.2e-19
C717 dac_1.out dac_0.carray_0.unitcap_47.cn 0.00925f
C718 dac_1.sw_top_0.en_buf avdd 1.98f
C719 dac_0.carray_0.unitcap_14.cn avdd 0.00155f
C720 dac_1.sky130_fd_sc_hd__inv_2_1.Y ctln4 3.6e-21
C721 comparator_0.outp comparator_0.in 0.0259f
C722 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_71.cn 0.18f
C723 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_0.Y 0.0089f
C724 comparator_0.vp dac_0.sky130_fd_sc_hd__inv_2_2.Y 84.2f
C725 comparator_0.vp dac_0.carray_0.unitcap_40.cn 0.514f
C726 comparator_0.trim_1.n0 trimb1 0.0594f
C727 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y 3.32f
C728 dac_1.sw_top_0.en_buf vinn 0.417f
C729 trimb3 trimb1 7.6e-20
C730 dac_1.out dac_1.carray_0.unitcap_326.cn 0.501f
C731 comparator_0.trim_1.n4 comparator_0.trim_1.n3 0.461f
C732 dac_1.carray_0.unitcap_0.cn dac_1.carray_0.unitcap_40.cn 0.0902f
C733 dac_1.carray_0.unitcap_95.cn dac_1.carray_0.unitcap_111.cn 0.0902f
C734 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_338.cn 0.161f
C735 dac_0.carray_0.unitcap_11.cn dac_0.carray_0.unitcap_13.cn 0.18f
C736 dac_1.sw_top_2.en_buf dac_1.sw_top_3.en_buf 0.00289f
C737 dac_1.carray_0.unitcap_14.cn dac_1.carray_0.unitcap_12.cn 0.18f
C738 dac_0.sw_top_1.en_buf avdd 1.98f
C739 dac_0.carray_0.unitcap_10.cn sample 0.0376f
C740 dac_0.sky130_fd_sc_hd__inv_2_0.Y ctlp5 0.16f
C741 dac_1.carray_0.unitcap_136.cn dac_1.carray_0.unitcap_128.cn 0.0902f
C742 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln2 0.0828f
C743 dac_1.sw_top_1.net1 avdd 0.849f
C744 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y 5.1e-21
C745 a_33300_6679# comparator_0.ip 0.00843f
C746 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_328.cn 0.00869f
C747 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_207.cn 0.00473f
C748 comparator_0.vp trim4 9.93e-21
C749 trimb1 trimb0 0.0476f
C750 comparator_0.vp dac_0.carray_0.unitcap_63.cn 0.51f
C751 dac_1.carray_0.unitcap_322.cn dac_1.carray_0.unitcap_324.cn 0.18f
C752 dac_0.carray_0.unitcap_176.cn avdd 0.095f
C753 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_0.cn 0.18f
C754 dac_0.carray_0.unitcap_0.cn dac_0.carray_0.unitcap_40.cn 0.0902f
C755 dac_1.out dac_1.carray_0.unitcap_200.cn 0.514f
C756 comparator_0.trim_0.n3 dac_1.sky130_fd_sc_hd__inv_2_0.Y 0.00436f
C757 dac_1.sw_top_1.net1 vinn 0.368f
C758 comparator_0.trim_1.n4 comparator_0.outp 0.522f
C759 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_135.cn 0.00473f
C760 comparator_0.ip ctlp7 0.011f
C761 comparator_0.trim_0.n2 trim3 0.128f
C762 dac_0.sw_top_2.en_buf dac_0.carray_0.unitcap_11.cn 0.00862f
C763 dac_1.carray_0.unitcap_8.cn dac_1.carray_0.unitcap_16.cn 0.0902f
C764 dac_0.carray_0.unitcap_136.cn dac_0.carray_0.unitcap_128.cn 0.0902f
C765 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp1 0.0826f
C766 dac_0.carray_0.unitcap_119.cn dac_1.carray_0.unitcap_119.cn 0.128f
C767 dac_0.carray_0.unitcap_13.cn vinp 0.0215f
C768 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_1.out 1.97e-19
C769 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln0 1.27e-20
C770 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_87.cn 0.18f
C771 comparator_0.trim_0.n4 comparator_0.trim_0.n2 0.187f
C772 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_3.Y 1.89f
C773 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.carray_0.unitcap_328.cn 0.00139f
C774 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.carray_0.unitcap_326.cn 0.091f
C775 dac_1.out dac_1.carray_0.unitcap_10.cn 0.557f
C776 comparator_0.trim_0.n2 trim0 9.86e-19
C777 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_334.cn 0.348f
C778 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_255.cn 0.161f
C779 dac_1.sky130_fd_sc_hd__inv_2_1.Y avdd 0.404f
C780 comparator_0.vp comparator_0.outn 0.0215f
C781 ctlp2 ctlp4 3.27e-21
C782 dac_0.carray_0.unitcap_8.cn dac_0.carray_0.unitcap_16.cn 0.0902f
C783 comparator_0.ip clkc 0.121f
C784 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.251f
C785 comparator_0.trim_1.n1 trimb1 0.183f
C786 dac_0.sw_top_2.en_buf vinp 0.695f
C787 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_199.cn 0.00473f
C788 comparator_0.vp dac_0.carray_0.unitcap_39.cn 0.51f
C789 comparator_0.vp dac_1.sky130_fd_sc_hd__inv_2_8.Y 2.16e-19
C790 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_24.cn 0.18f
C791 dac_0.carray_0.unitcap_160.cn avdd 0.095f
C792 dac_0.sw_top_0.en_buf dac_0.carray_0.unitcap_80.cn 5.45e-19
C793 dac_0.sky130_fd_sc_hd__inv_2_8.Y avdd 0.26f
C794 dac_1.sky130_fd_sc_hd__inv_2_6.Y ctln0 0.16f
C795 dac_1.out dac_1.carray_0.unitcap_192.cn 0.514f
C796 dac_0.carray_0.unitcap_159.cn dac_0.carray_0.unitcap_151.cn 0.0902f
C797 dac_1.sw_top_1.en_buf avdd 1.98f
C798 dac_0.carray_0.unitcap_12.cn avdd 0.00155f
C799 avdd sample 3.12f
C800 a_33300_5579# avdd 0.381f
C801 dac_0.sky130_fd_sc_hd__inv_2_2.Y comparator_0.trim_1.n3 0.0641f
C802 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_79.cn 0.18f
C803 dac_1.sw_top_1.en_buf vinn 0.705f
C804 comparator_0.trim_1.n4 comparator_0.trim_1.n0 0.0407f
C805 comparator_0.trim_1.n4 trimb3 0.0166f
C806 sample vinn 0.027f
C807 dac_1.out dac_1.carray_0.unitcap_334.cn 0.501f
C808 dac_1.carray_0.unitcap_71.cn dac_1.carray_0.unitcap_95.cn 0.0902f
C809 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_239.cn 0.161f
C810 dac_1.carray_0.unitcap_336.cn dac_1.carray_0.unitcap_337.cn 0.18f
C811 dac_0.carray_0.unitcap_326.cn dac_0.carray_0.unitcap_334.cn 0.18f
C812 dac_0.carray_0.unitcap_288.cn sample 0.0536f
C813 dac_0.sw_top_3.en_buf avdd 1.98f
C814 dac_1.carray_0.unitcap_112.cn dac_1.carray_0.unitcap_136.cn 0.0902f
C815 comparator_0.trim_1.n4 trimb0 0.00577f
C816 dac_1.out dac_1.sw_top_3.net1 0.322f
C817 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_175.cn 0.00473f
C818 comparator_0.ip ctlp4 0.0015f
C819 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_326.cn 0.043f
C820 ctlp7 trimb4 3.66e-20
C821 comparator_0.vp dac_0.carray_0.unitcap_47.cn 0.51f
C822 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_16.cn 0.18f
C823 dac_0.carray_0.unitcap_144.cn avdd 0.0742f
C824 dac_1.out dac_1.carray_0.unitcap_168.cn 0.514f
C825 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln7 0.0932f
C826 latch_0.Qn avdd 0.551f
C827 dac_0.sw_top_2.en_buf dac_0.carray_0.unitcap_10.cn 0.0123f
C828 comparator_0.ip comparator_0.trim_0.n4 0.0147f
C829 dac_0.carray_0.unitcap_112.cn dac_0.carray_0.unitcap_136.cn 0.0902f
C830 dac_0.carray_0.unitcap_11.cn vinp 0.0736f
C831 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_336.cn 0.00213f
C832 dac_0.carray_0.unitcap_127.cn dac_1.carray_0.unitcap_127.cn 0.128f
C833 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_55.cn 0.18f
C834 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_7.cn 0.18f
C835 dac_1.sky130_fd_sc_hd__inv_2_2.Y avdd 3.53f
C836 dac_1.out dac_1.carray_0.unitcap_11.cn 0.556f
C837 trimb4 clkc 4.33e-19
C838 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.carray_0.unitcap_334.cn 2.28e-19
C839 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_326.cn 0.34f
C840 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp2 0.049f
C841 comparator_0.in trim1 0.088f
C842 comparator_0.trim_1.n3 comparator_0.outn 9.64e-20
C843 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_247.cn 0.161f
C844 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln5 1.48e-19
C845 dac_1.sky130_fd_sc_hd__inv_2_2.Y vinn 1.86f
C846 dac_1.sky130_fd_sc_hd__inv_2_0.Y ctln4 0.00127f
C847 comparator_0.trim_1.n3 comparator_0.trim_1.n2 0.264f
C848 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_183.cn 0.00473f
C849 comparator_0.trim_1.n4 comparator_0.trim_1.n1 0.0439f
C850 dac_0.carray_0.unitcap_152.cn avdd 0.0958f
C851 dac_0.sky130_fd_sc_hd__inv_2_0.Y comparator_0.vp 17.5f
C852 dac_1.out dac_1.carray_0.unitcap_176.cn 0.514f
C853 dac_0.sw_top_3.net1 comparator_0.vp 0.322f
C854 dac_0.carray_0.unitcap_135.cn dac_0.carray_0.unitcap_159.cn 0.0902f
C855 comparator_0.trim_0.n3 ctln4 0.00113f
C856 dac_0.carray_0.unitcap_13.cn avdd 0.0016f
C857 dac_1.sw_top_0.net1 dac_1.carray_0.unitcap_64.cn 1e-20
C858 dac_1.sw_top_3.en_buf avdd 1.98f
C859 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp2 0.00122f
C860 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp7 0.0932f
C861 comparator_0.outp comparator_0.outn 0.619f
C862 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_338.cn 0.00213f
C863 dac_0.sky130_fd_sc_hd__inv_2_1.Y ctlp7 0.0531f
C864 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_63.cn 0.18f
C865 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_31.cn 0.18f
C866 dac_0.sky130_fd_sc_hd__inv_2_6.Y avdd 0.234f
C867 dac_1.sw_top_3.en_buf vinn 0.705f
C868 comparator_0.trim_1.n2 comparator_0.outp 0.0319f
C869 dac_1.out dac_1.carray_0.unitcap_331.cn 0.501f
C870 dac_1.carray_0.unitcap_87.cn dac_1.carray_0.unitcap_71.cn 0.0902f
C871 ctlp5 ctlp7 1.09e-19
C872 ctln2 ctln1 0.103f
C873 ctln3 ctln0 1.18e-19
C874 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_223.cn 0.161f
C875 dac_0.carray_0.unitcap_256.cn sample 0.217f
C876 dac_0.carray_0.unitcap_10.cn dac_0.carray_0.unitcap_11.cn 0.18f
C877 dac_0.sw_top_2.en_buf avdd 1.99f
C878 dac_1.carray_0.unitcap_120.cn dac_1.carray_0.unitcap_112.cn 0.0902f
C879 comparator_0.in ctln5 0.00237f
C880 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_167.cn 0.00473f
C881 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_334.cn 0.0355f
C882 dac_0.carray_0.unitcap_128.cn avdd 0.0952f
C883 dac_0.sw_top_2.net1 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.358f
C884 comparator_0.vp ctlp1 9.29e-19
C885 dac_1.out dac_1.carray_0.unitcap_160.cn 0.514f
C886 avdd trimb2 0.0558f
C887 dac_1.sky130_fd_sc_hd__inv_2_0.Y avdd 0.303f
C888 dac_0.sw_top_2.en_buf dac_0.carray_0.unitcap_288.cn 0.00736f
C889 dac_0.carray_0.unitcap_120.cn dac_0.carray_0.unitcap_112.cn 0.0902f
C890 dac_0.carray_0.unitcap_10.cn vinp 0.0189f
C891 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_255.cn 0.00213f
C892 dac_0.carray_0.unitcap_103.cn dac_1.carray_0.unitcap_103.cn 0.128f
C893 dac_0.sky130_fd_sc_hd__inv_2_3.Y comparator_0.ip 4.53e-19
C894 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_39.cn 0.18f
C895 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_23.cn 0.18f
C896 clkc trim2 2.42e-19
C897 dac_0.carray_0.unitcap_80.cn sample 7.14e-19
C898 dac_1.out dac_1.sw_top_0.net1 0.333f
C899 comparator_0.trim_0.n3 avdd 0.00409f
C900 comparator_0.trim_1.n4 dac_0.carray_0.unitcap_337.cn 0.0265f
C901 dac_1.out dac_1.carray_0.unitcap_13.cn 0.558f
C902 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_328.cn 0.123f
C903 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_231.cn 0.161f
C904 comparator_0.outn trimb3 0.00111f
C905 dac_1.carray_0.unitcap_338.cn dac_1.carray_0.unitcap_336.cn 0.0902f
C906 dac_1.out clkc 0.0608f
C907 comparator_0.trim_1.n2 comparator_0.trim_1.n0 1.16e-19
C908 comparator_0.trim_1.n2 trimb3 0.127f
C909 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_216.cn 0.18f
C910 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_151.cn 0.00473f
C911 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_7.Y 0.00996f
C912 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.carray_0.unitcap_322.cn 0.275f
C913 dac_0.carray_0.unitcap_7.cn dac_0.carray_0.unitcap_47.cn 0.0902f
C914 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp4 0.0827f
C915 dac_0.carray_0.unitcap_136.cn avdd 0.0948f
C916 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.357f
C917 dac_0.sw_top_1.en_buf dac_0.carray_0.unitcap_48.cn 8.31e-19
C918 dac_0.sky130_fd_sc_hd__inv_2_0.Y comparator_0.trim_1.n3 0.00481f
C919 dac_0.sky130_fd_sc_hd__inv_2_1.Y ctlp4 3.6e-21
C920 dac_1.out ctln2 5.56e-19
C921 dac_0.sky130_fd_sc_hd__inv_2_2.Y ctlp6 0.00123f
C922 dac_1.out dac_1.carray_0.unitcap_144.cn 0.514f
C923 dac_0.sky130_fd_sc_hd__inv_2_5.Y avdd 0.222f
C924 dac_0.carray_0.unitcap_143.cn dac_0.carray_0.unitcap_135.cn 0.0902f
C925 comparator_0.trim_1.n2 trimb0 9.83e-19
C926 dac_1.sw_top_2.en_buf avdd 1.99f
C927 dac_0.carray_0.unitcap_11.cn avdd 0.00997f
C928 ctlp4 ctlp5 0.106f
C929 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.carray_0.unitcap_320.cn 0.119f
C930 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_239.cn 0.00213f
C931 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_47.cn 0.18f
C932 dac_0.carray_0.unitcap_72.cn sample 0.00246f
C933 dac_1.out dac_1.carray_0.unitcap_330.cn 0.502f
C934 dac_1.sw_top_2.en_buf vinn 0.695f
C935 dac_1.carray_0.unitcap_79.cn dac_1.carray_0.unitcap_87.cn 0.0902f
C936 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_215.cn 0.161f
C937 comparator_0.trim_0.n1 comparator_0.trim_0.n0 0.207f
C938 dac_0.carray_0.unitcap_328.cn dac_0.carray_0.unitcap_326.cn 0.18f
C939 trim3 trim2 0.0386f
C940 dac_1.carray_0.unitcap_96.cn dac_1.carray_0.unitcap_120.cn 0.0902f
C941 dac_0.sw_top_0.net1 comparator_0.vp 0.333f
C942 avdd vinp 3.08f
C943 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_159.cn 0.00473f
C944 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_224.cn 0.18f
C945 comparator_0.trim_0.n4 trim2 0.0233f
C946 dac_0.sw_top_0.en_buf dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.27f
C947 dac_0.carray_0.unitcap_112.cn avdd 0.0922f
C948 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln2 0.049f
C949 dac_1.out dac_1.carray_0.unitcap_152.cn 0.514f
C950 trim2 trim0 7.61e-19
C951 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.0144f
C952 comparator_0.trim_1.n2 comparator_0.trim_1.n1 0.217f
C953 dac_1.out comparator_0.trim_0.n4 0.0214f
C954 dac_0.carray_0.unitcap_326.cn avdd 5.03e-19
C955 dac_0.carray_0.unitcap_96.cn dac_0.carray_0.unitcap_120.cn 0.0902f
C956 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_247.cn 0.00213f
C957 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.carray_0.unitcap_321.cn 0.18f
C958 dac_0.carray_0.unitcap_288.cn vinp 5.91e-19
C959 dac_0.carray_0.unitcap_111.cn dac_1.carray_0.unitcap_111.cn 0.128f
C960 comparator_0.diff avdd 0.00121f
C961 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_337.cn 0.138f
C962 dac_0.carray_0.unitcap_48.cn sample 0.00246f
C963 dac_1.out dac_1.carray_0.unitcap_12.cn 0.556f
C964 comparator_0.outn trim1 0.00169f
C965 dac_0.sw_top_1.net1 dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.424f
C966 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.carray_0.unitcap_322.cn 0.00396f
C967 comparator_0.trim_1.n4 dac_0.carray_0.unitcap_330.cn 0.00649f
C968 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_191.cn 0.161f
C969 dac_1.carray_0.unitcap_255.cn dac_1.carray_0.unitcap_338.cn 0.0902f
C970 comparator_0.in a_33300_5579# 0.00575f
C971 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.134f
C972 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_135.cn 0.00473f
C973 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_4.Y 0.00883f
C974 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_208.cn 0.18f
C975 comparator_0.vp ctlp7 9.15e-19
C976 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.carray_0.unitcap_324.cn 0.173f
C977 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y 7.78e-22
C978 dac_0.carray_0.unitcap_120.cn avdd 0.0952f
C979 dac_1.out dac_1.carray_0.unitcap_128.cn 0.514f
C980 dac_0.carray_0.unitcap_119.cn dac_0.carray_0.unitcap_143.cn 0.0902f
C981 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp5 2.14e-21
C982 dac_0.carray_0.unitcap_10.cn avdd 0.021f
C983 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_223.cn 0.181f
C984 dac_1.carray_0.unitcap_9.cn sample 0.00958f
C985 dac_0.sky130_fd_sc_hd__inv_2_6.Y ctlp0 0.16f
C986 avdd ctln4 0.116f
C987 dac_1.out ctln7 9.15e-19
C988 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln2 0.00122f
C989 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_14.cn 0.0902f
C990 dac_1.carray_0.unitcap_328.cn ctln5 0.00202f
C991 comparator_0.vp clkc 0.047f
C992 dac_0.carray_0.unitcap_56.cn sample 0.0026f
C993 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.00846f
C994 dac_1.carray_0.unitcap_55.cn dac_1.carray_0.unitcap_79.cn 0.0902f
C995 dac_1.out dac_1.carray_0.unitcap_337.cn 0.506f
C996 dac_1.carray_0.unitcap_0.cn sample 0.00246f
C997 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_1.Y 0.325f
C998 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_207.cn 0.161f
C999 dac_0.sw_top_2.net1 dac_0.sw_top_3.net1 0.00267f
C1000 dac_0.carray_0.unitcap_288.cn dac_0.carray_0.unitcap_10.cn 0.18f
C1001 dac_1.carray_0.unitcap_104.cn dac_1.carray_0.unitcap_96.cn 0.0902f
C1002 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp5 1.78e-19
C1003 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_184.cn 0.18f
C1004 dac_0.sw_top_1.en_buf dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.04f
C1005 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.081f
C1006 dac_0.carray_0.unitcap_96.cn avdd 0.0948f
C1007 dac_1.out dac_1.carray_0.unitcap_136.cn 0.514f
C1008 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln5 0.0515f
C1009 dac_0.carray_0.unitcap_8.cn sample 0.00246f
C1010 dac_0.carray_0.unitcap_328.cn avdd 8.02e-19
C1011 dac_0.carray_0.unitcap_104.cn dac_0.carray_0.unitcap_96.cn 0.0902f
C1012 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_231.cn 0.18f
C1013 ctln7 ctln6 0.106f
C1014 dac_0.carray_0.unitcap_95.cn dac_1.carray_0.unitcap_95.cn 0.128f
C1015 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln7 5.61e-22
C1016 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_330.cn 7.44e-19
C1017 trimb2 trimb1 0.0771f
C1018 dac_0.carray_0.unitcap_32.cn sample 0.00246f
C1019 dac_1.out dac_1.carray_0.unitcap_14.cn 0.556f
C1020 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.108f
C1021 dac_0.sky130_fd_sc_hd__inv_2_7.Y comparator_0.vp 0.541f
C1022 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_9.cn 0.0902f
C1023 comparator_0.vp ctlp4 5.62e-19
C1024 dac_1.carray_0.unitcap_24.cn sample 0.00277f
C1025 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_199.cn 0.161f
C1026 dac_1.carray_0.unitcap_239.cn dac_1.carray_0.unitcap_255.cn 0.0902f
C1027 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln1 0.0826f
C1028 dac_0.sky130_fd_sc_hd__inv_2_0.Y ctlp6 0.0512f
C1029 comparator_0.trim_1.n3 ctlp7 0.00751f
C1030 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.00124f
C1031 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_0.cn 0.18f
C1032 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp0 1.27e-20
C1033 comparator_0.trim_0.n3 dac_1.sky130_fd_sc_hd__inv_2_5.Y 1.18e-19
C1034 comparator_0.vp comparator_0.trim_0.n4 0.002f
C1035 dac_0.carray_0.unitcap_104.cn avdd 0.0703f
C1036 dac_0.sw_top_3.en_buf dac_0.carray_0.unitcap_32.cn 2.32e-19
C1037 avdd vinn 3.08f
C1038 dac_1.out dac_1.carray_0.unitcap_112.cn 0.514f
C1039 comparator_0.outp a_33300_6679# 0.15f
C1040 dac_0.carray_0.unitcap_127.cn dac_0.carray_0.unitcap_119.cn 0.0902f
C1041 comparator_0.ip trimb4 0.104f
C1042 dac_0.carray_0.unitcap_288.cn avdd 0.119f
C1043 comparator_0.trim_0.n2 trim2 0.243f
C1044 dac_1.sw_top_2.net1 dac_1.carray_0.unitcap_10.cn 0.00207f
C1045 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.291f
C1046 dac_1.carray_0.unitcap_256.cn sample 0.217f
C1047 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_215.cn 0.18f
C1048 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp2 0.0828f
C1049 dac_1.sky130_fd_sc_hd__inv_2_1.Y trim4 1.03e-19
C1050 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_12.cn 0.0902f
C1051 dac_0.sky130_fd_sc_hd__inv_2_2.Y sample 2.53f
C1052 dac_1.carray_0.unitcap_15.cn dac_1.carray_0.unitcap_14.cn 0.18f
C1053 dac_0.carray_0.unitcap_40.cn sample 0.00329f
C1054 dac_1.out dac_1.carray_0.unitcap_336.cn 0.642f
C1055 dac_1.carray_0.unitcap_16.cn sample 0.00246f
C1056 dac_1.carray_0.unitcap_63.cn dac_1.carray_0.unitcap_55.cn 0.0902f
C1057 ctlp3 ctlp4 0.107f
C1058 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_175.cn 0.161f
C1059 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_0.Y 0.0116f
C1060 dac_0.carray_0.unitcap_322.cn dac_0.carray_0.unitcap_328.cn 0.18f
C1061 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln7 1.78e-19
C1062 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_328.cn 2e-20
C1063 dac_1.carray_0.unitcap_88.cn dac_1.carray_0.unitcap_104.cn 0.0902f
C1064 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_24.cn 0.18f
C1065 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_248.cn 0.18f
C1066 dac_0.sw_top_3.en_buf dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.15f
C1067 dac_0.carray_0.unitcap_88.cn avdd 0.0952f
C1068 comparator_0.in comparator_0.trim_0.n3 2.47f
C1069 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_337.cn 0.00682f
C1070 dac_1.out dac_1.carray_0.unitcap_120.cn 0.514f
C1071 comparator_0.outp clkc 0.129f
C1072 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.out 0.00317f
C1073 dac_0.carray_0.unitcap_322.cn avdd 0.00205f
C1074 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_191.cn 0.18f
C1075 dac_0.carray_0.unitcap_88.cn dac_0.carray_0.unitcap_104.cn 0.0902f
C1076 dac_0.sw_top_3.net1 dac_0.sw_top_1.net1 0.00267f
C1077 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.663f
C1078 dac_0.carray_0.unitcap_71.cn dac_1.carray_0.unitcap_71.cn 0.128f
C1079 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_331.cn 7.44e-19
C1080 dac_0.sky130_fd_sc_hd__inv_2_4.Y comparator_0.vp 1.03f
C1081 dac_0.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.ip 0.0265f
C1082 comparator_0.trim_1.n4 trimb2 0.0205f
C1083 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_256.cn 0.0902f
C1084 comparator_0.trim_1.n3 ctlp4 0.0012f
C1085 dac_1.out dac_1.carray_0.unitcap_338.cn 0.526f
C1086 dac_0.sky130_fd_sc_hd__inv_2_1.Y comparator_0.ip 0.0156f
C1087 dac_1.sw_top_2.net1 dac_1.sw_top_3.net1 0.00267f
C1088 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_183.cn 0.161f
C1089 dac_1.carray_0.unitcap_247.cn dac_1.carray_0.unitcap_239.cn 0.0902f
C1090 comparator_0.outn a_33300_5579# 0.197f
C1091 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.591f
C1092 comparator_0.ip ctlp5 0.00242f
C1093 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_16.cn 0.18f
C1094 dac_0.carray_0.unitcap_64.cn avdd 0.0953f
C1095 dac_1.out dac_1.carray_0.unitcap_96.cn 0.514f
C1096 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln6 0.0828f
C1097 dac_0.carray_0.unitcap_103.cn dac_0.carray_0.unitcap_127.cn 0.0902f
C1098 dac_1.sky130_fd_sc_hd__inv_2_2.Y trim4 0.00524f
C1099 dac_0.sky130_fd_sc_hd__inv_2_3.Y comparator_0.vp 4.37f
C1100 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_4.Y 0.00883f
C1101 dac_0.carray_0.unitcap_256.cn avdd 0.00523f
C1102 dac_1.carray_0.unitcap_288.cn sample 0.0536f
C1103 dac_1.carray_0.unitcap_320.cn avdd 0.111f
C1104 comparator_0.ip dac_1.out 0.0506f
C1105 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_13.cn 0.0902f
C1106 comparator_0.outp trim3 4.66e-19
C1107 comparator_0.trim_1.n0 clkc 1.59e-19
C1108 dac_0.carray_0.unitcap_336.cn dac_1.carray_0.unitcap_336.cn 0.128f
C1109 dac_1.out dac_1.carray_0.unitcap_255.cn 0.511f
C1110 comparator_0.outp comparator_0.trim_0.n4 0.00991f
C1111 dac_1.carray_0.unitcap_39.cn dac_1.carray_0.unitcap_63.cn 0.0902f
C1112 latch_0.Qn comparator_0.outn 1.66e-19
C1113 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp3 1.86e-19
C1114 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_167.cn 0.161f
C1115 dac_0.sw_top_1.en_buf dac_0.sw_top_3.net1 4.9e-19
C1116 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln4 2.49e-19
C1117 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_326.cn 8.52e-19
C1118 dac_0.carray_0.unitcap_256.cn dac_0.carray_0.unitcap_288.cn 0.18f
C1119 dac_1.carray_0.unitcap_64.cn dac_1.carray_0.unitcap_88.cn 0.0902f
C1120 trimb0 clkc 0.00269f
C1121 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_216.cn 0.18f
C1122 comparator_0.diff comparator_0.in 0.146f
C1123 dac_0.carray_0.unitcap_80.cn avdd 0.0609f
C1124 dac_0.sw_top_2.en_buf dac_0.sky130_fd_sc_hd__inv_2_2.Y 1.16f
C1125 comparator_0.in comparator_0.trim_0.n0 0.556f
C1126 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_330.cn 0.039f
C1127 dac_1.out dac_1.carray_0.unitcap_104.cn 0.514f
C1128 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.291f
C1129 dac_0.sky130_fd_sc_hd__inv_2_6.VPB trimb4 9.03e-19
C1130 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp3 0.161f
C1131 dac_0.carray_0.unitcap_324.cn avdd 0.00952f
C1132 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_200.cn 0.18f
C1133 dac_1.carray_0.unitcap_31.cn dac_1.carray_0.unitcap_7.cn 0.0902f
C1134 dac_0.carray_0.unitcap_64.cn dac_0.carray_0.unitcap_88.cn 0.0902f
C1135 dac_0.sky130_fd_sc_hd__inv_2_1.Y trimb4 5.14e-19
C1136 dac_1.carray_0.unitcap_321.cn avdd 0.0705f
C1137 dac_0.sw_top_0.en_buf dac_0.sw_top_0.net1 0.585f
C1138 comparator_0.vp dac_1.carray_0.unitcap_336.cn 0.0114f
C1139 dac_0.carray_0.unitcap_87.cn dac_1.carray_0.unitcap_87.cn 0.128f
C1140 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_255.cn 0.18f
C1141 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_1.sky130_fd_sc_hd__inv_2_0.Y 3.14e-19
C1142 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_334.cn 7.44e-19
C1143 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_3.Y 0.00846f
C1144 ctlp6 ctlp7 0.105f
C1145 avdd ctlp0 0.224f
C1146 dac_1.out dac_1.carray_0.unitcap_239.cn 0.51f
C1147 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_288.cn 0.0902f
C1148 ctln2 ctln0 1.74e-19
C1149 dac_1.sw_top_2.en_buf dac_1.carray_0.unitcap_24.cn 6.3e-19
C1150 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_151.cn 0.161f
C1151 dac_1.carray_0.unitcap_223.cn dac_1.carray_0.unitcap_247.cn 0.0902f
C1152 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_224.cn 0.18f
C1153 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_7.Y 0.00996f
C1154 comparator_0.trim_1.n4 comparator_0.diff 0.00619f
C1155 dac_1.sky130_fd_sc_hd__inv_2_0.Y trim4 2.45e-19
C1156 comparator_0.in ctln4 0.00138f
C1157 dac_0.sky130_fd_sc_hd__inv_2_8.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y 2.29f
C1158 dac_0.sw_top_1.net1 dac_0.sw_top_0.net1 0.00267f
C1159 comparator_0.vp ctlp2 5.56e-19
C1160 dac_0.carray_0.unitcap_72.cn avdd 0.0966f
C1161 dac_1.sky130_fd_sc_hd__inv_2_5.Y avdd 0.222f
C1162 dac_1.out dac_1.carray_0.unitcap_88.cn 0.514f
C1163 avdd trimb1 0.0683f
C1164 dac_0.sw_top_3.net1 sample 0.037f
C1165 dac_0.carray_0.unitcap_111.cn dac_0.carray_0.unitcap_103.cn 0.0902f
C1166 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_192.cn 0.18f
C1167 dac_1.sw_top_3.net1 dac_1.sw_top_1.net1 0.00267f
C1168 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_136.cn 0.18f
C1169 comparator_0.trim_0.n3 trim4 0.319f
C1170 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_328.cn 0.00171f
C1171 dac_1.carray_0.unitcap_10.cn sample 0.0376f
C1172 comparator_0.vp dac_1.carray_0.unitcap_338.cn 0.00925f
C1173 dac_1.carray_0.unitcap_248.cn avdd 0.111f
C1174 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_2.Y 0.134f
C1175 dac_1.out dac_1.carray_0.unitcap_7.cn 0.51f
C1176 comparator_0.in comparator_0.trim_0.n1 0.578f
C1177 comparator_0.ip dac_0.carray_0.unitcap_336.cn 0.0031f
C1178 clkc trim1 2.5e-20
C1179 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_11.cn 0.0902f
C1180 dac_0.carray_0.unitcap_338.cn dac_1.carray_0.unitcap_338.cn 0.128f
C1181 dac_1.out dac_1.carray_0.unitcap_247.cn 0.51f
C1182 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_326.cn 0.00141f
C1183 dac_1.carray_0.unitcap_47.cn dac_1.carray_0.unitcap_39.cn 0.0902f
C1184 dac_0.sw_top_3.en_buf dac_0.sw_top_3.net1 0.585f
C1185 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_159.cn 0.161f
C1186 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.sky130_fd_sc_hd__inv_2_1.Y 0.00854f
C1187 dac_1.sky130_fd_sc_hd__inv_2_6.Y avdd 0.235f
C1188 dac_0.carray_0.unitcap_324.cn dac_0.carray_0.unitcap_322.cn 0.18f
C1189 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_334.cn 0.00192f
C1190 dac_1.carray_0.unitcap_80.cn dac_1.carray_0.unitcap_64.cn 0.0902f
C1191 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_208.cn 0.18f
C1192 comparator_0.trim_1.n2 trimb2 0.243f
C1193 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp1 5.89e-21
C1194 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_8.Y 2.29f
C1195 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp5 0.0826f
C1196 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.carray_0.unitcap_255.cn 0.18f
C1197 dac_0.sky130_fd_sc_hd__inv_2_6.VPB dac_0.carray_0.unitcap_320.cn 0.00177f
C1198 dac_1.out ctln1 9.29e-19
C1199 dac_0.sky130_fd_sc_hd__inv_2_1.Y ctlp5 0.00139f
C1200 ctlp2 ctlp3 0.107f
C1201 dac_0.carray_0.unitcap_48.cn avdd 0.0948f
C1202 dac_0.sky130_fd_sc_hd__inv_2_2.Y vinp 1.86f
C1203 dac_1.out dac_1.carray_0.unitcap_64.cn 0.514f
C1204 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_331.cn 0.0439f
C1205 comparator_0.vp comparator_0.ip 0.35f
C1206 comparator_0.in avdd 0.282f
C1207 ctlp4 ctlp6 1.34e-20
C1208 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_112.cn 0.18f
C1209 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_168.cn 0.18f
C1210 dac_1.carray_0.unitcap_232.cn avdd 0.11f
C1211 comparator_0.vp dac_1.carray_0.unitcap_255.cn 0.00925f
C1212 comparator_0.trim_0.n3 dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.00508f
C1213 dac_1.carray_0.unitcap_23.cn dac_1.carray_0.unitcap_31.cn 0.0902f
C1214 dac_0.carray_0.unitcap_80.cn dac_0.carray_0.unitcap_64.cn 0.0902f
C1215 dac_1.out dac_1.carray_0.unitcap_31.cn 0.51f
C1216 dac_0.carray_0.unitcap_79.cn dac_1.carray_0.unitcap_79.cn 0.128f
C1217 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_1.sky130_fd_sc_hd__inv_2_2.Y 3.14e-19
C1218 dac_1.carray_0.unitcap_322.cn ctln4 1.86e-19
C1219 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_326.cn 0.00141f
C1220 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.carray_0.unitcap_324.cn 8.63e-19
C1221 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_10.cn 0.0902f
C1222 dac_1.out dac_1.carray_0.unitcap_223.cn 0.51f
C1223 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_1.out 8.01e-19
C1224 dac_1.sw_top_1.en_buf dac_1.sw_top_3.net1 4.9e-19
C1225 dac_1.sw_top_3.net1 sample 0.037f
C1226 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_135.cn 0.161f
C1227 dac_1.carray_0.unitcap_231.cn dac_1.carray_0.unitcap_223.cn 0.0902f
C1228 trim3 trim1 1.58e-19
C1229 dac_1.carray_0.unitcap_9.cn avdd 0.0138f
C1230 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_184.cn 0.18f
C1231 dac_1.carray_0.unitcap_321.cn dac_1.carray_0.unitcap_320.cn 0.0902f
C1232 comparator_0.trim_0.n4 trim1 0.0153f
C1233 ctln4 ctln3 0.105f
C1234 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln1 0.159f
C1235 dac_0.carray_0.unitcap_56.cn avdd 0.082f
C1236 trim1 trim0 0.0508f
C1237 comparator_0.diff trim4 4.62e-20
C1238 dac_1.carray_0.unitcap_0.cn avdd 0.112f
C1239 dac_1.out dac_1.carray_0.unitcap_80.cn 0.514f
C1240 comparator_0.trim_1.n4 avdd 0.236f
C1241 dac_0.carray_0.unitcap_95.cn dac_0.carray_0.unitcap_111.cn 0.0902f
C1242 comparator_0.ip ctlp3 5.51e-19
C1243 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_120.cn 0.18f
C1244 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_326.cn 9.72e-19
C1245 dac_1.sw_top_0.en_buf dac_1.sw_top_0.net1 0.585f
C1246 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_176.cn 0.18f
C1247 dac_1.sw_top_2.en_buf dac_1.carray_0.unitcap_288.cn 0.00736f
C1248 dac_1.carray_0.unitcap_240.cn avdd 0.094f
C1249 comparator_0.vp dac_1.carray_0.unitcap_239.cn 0.00925f
C1250 dac_1.carray_0.unitcap_11.cn sample 0.0348f
C1251 dac_1.out dac_1.carray_0.unitcap_23.cn 0.512f
C1252 dac_0.carray_0.unitcap_321.cn dac_0.carray_0.unitcap_320.cn 0.0902f
C1253 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_10.cn 0.0902f
C1254 dac_0.carray_0.unitcap_255.cn dac_1.carray_0.unitcap_255.cn 0.128f
C1255 dac_1.out dac_1.carray_0.unitcap_231.cn 0.51f
C1256 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_334.cn 7.44e-19
C1257 dac_0.carray_0.unitcap_8.cn avdd 0.102f
C1258 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_143.cn 0.18f
C1259 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_331.cn 0.0064f
C1260 dac_1.carray_0.unitcap_322.cn avdd 0.0026f
C1261 dac_1.carray_0.unitcap_72.cn dac_1.carray_0.unitcap_80.cn 0.0902f
C1262 dac_0.sw_top_0.net1 sample 0.0117f
C1263 comparator_0.vp trimb4 0.00273f
C1264 dac_1.sw_top_3.net1 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.461f
C1265 comparator_0.diff comparator_0.outn 0.00297f
C1266 dac_1.sw_top_1.net1 dac_1.sw_top_0.net1 0.00267f
C1267 dac_0.carray_0.unitcap_32.cn avdd 0.0965f
C1268 dac_0.carray_0.unitcap_324.cn ctlp0 0.00176f
C1269 comparator_0.outn comparator_0.trim_0.n0 0.00209f
C1270 comparator_0.vp dac_1.carray_0.unitcap_7.cn 0.00925f
C1271 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_334.cn 9.72e-19
C1272 dac_1.out dac_1.carray_0.unitcap_72.cn 0.514f
C1273 dac_1.carray_0.unitcap_24.cn avdd 0.11f
C1274 comparator_0.trim_1.n3 comparator_0.ip 2.47f
C1275 dac_0.sky130_fd_sc_hd__inv_2_4.Y ctlp6 1.36e-21
C1276 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_96.cn 0.18f
C1277 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_160.cn 0.18f
C1278 dac_0.sky130_fd_sc_hd__inv_2_6.Y ctlp1 0.0498f
C1279 dac_0.carray_0.unitcap_72.cn dac_0.carray_0.unitcap_80.cn 0.0902f
C1280 dac_1.carray_0.unitcap_15.cn dac_1.carray_0.unitcap_23.cn 0.0902f
C1281 dac_1.carray_0.unitcap_216.cn avdd 0.112f
C1282 comparator_0.vp dac_1.carray_0.unitcap_247.cn 0.00925f
C1283 avdd ctln3 0.116f
C1284 dac_1.out ctln6 5.61e-19
C1285 dac_0.carray_0.unitcap_55.cn dac_1.carray_0.unitcap_55.cn 0.128f
C1286 dac_1.out dac_1.carray_0.unitcap_15.cn 0.501f
C1287 dac_1.carray_0.unitcap_328.cn ctln4 6.13e-19
C1288 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_4.Y 1.03f
C1289 dac_1.out dac_1.carray_0.unitcap_215.cn 0.51f
C1290 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_11.cn 0.0902f
C1291 dac_1.sw_top_3.en_buf dac_1.sw_top_3.net1 0.585f
C1292 comparator_0.vp dac_0.carray_0.unitcap_9.cn 0.557f
C1293 dac_1.sky130_fd_sc_hd__inv_2_7.Y ctln1 3.56e-20
C1294 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_119.cn 0.18f
C1295 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp7 2.25e-19
C1296 dac_1.carray_0.unitcap_215.cn dac_1.carray_0.unitcap_231.cn 0.0902f
C1297 comparator_0.outp comparator_0.ip 0.394f
C1298 dac_1.carray_0.unitcap_256.cn avdd 0.0056f
C1299 dac_0.sky130_fd_sc_hd__inv_2_3.Y ctlp6 1.78e-19
C1300 dac_1.carray_0.unitcap_248.cn dac_1.carray_0.unitcap_321.cn 0.0902f
C1301 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_0.Y 0.108f
C1302 dac_0.sky130_fd_sc_hd__inv_2_2.Y avdd 3.48f
C1303 dac_0.carray_0.unitcap_40.cn avdd 0.095f
C1304 dac_1.sky130_fd_sc_hd__inv_2_8.Y ctln4 0.16f
C1305 dac_1.carray_0.unitcap_16.cn avdd 0.113f
C1306 dac_1.out dac_1.carray_0.unitcap_48.cn 0.514f
C1307 comparator_0.vp dac_1.carray_0.unitcap_31.cn 0.00925f
C1308 dac_0.carray_0.unitcap_71.cn dac_0.carray_0.unitcap_95.cn 0.0902f
C1309 dac_0.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.vp 0.00317f
C1310 dac_1.sw_top_0.net1 sample 0.0117f
C1311 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_144.cn 0.18f
C1312 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_104.cn 0.18f
C1313 comparator_0.vp dac_1.carray_0.unitcap_223.cn 0.00925f
C1314 ctln7 ctln5 1.09e-19
C1315 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_334.cn 9.72e-19
C1316 dac_1.carray_0.unitcap_13.cn sample 0.0343f
C1317 dac_1.sw_top_2.en_buf dac_1.carray_0.unitcap_10.cn 0.0123f
C1318 dac_1.out dac_0.carray_0.unitcap_336.cn 0.00955f
C1319 dac_0.sky130_fd_sc_hd__inv_2_1.Y comparator_0.vp 35.4f
C1320 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln6 1.36e-21
C1321 dac_1.carray_0.unitcap_224.cn avdd 0.11f
C1322 comparator_0.outn comparator_0.trim_0.n1 0.0021f
C1323 avdd trim4 0.0139f
C1324 dac_0.carray_0.unitcap_248.cn dac_0.carray_0.unitcap_321.cn 0.0902f
C1325 a_33300_6679# latch_0.Qn 0.117f
C1326 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_288.cn 0.0902f
C1327 dac_0.carray_0.unitcap_239.cn dac_1.carray_0.unitcap_239.cn 0.128f
C1328 a_33300_5579# clkc 6.73e-19
C1329 comparator_0.vp ctlp5 9.28e-19
C1330 dac_1.out dac_1.carray_0.unitcap_191.cn 0.51f
C1331 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_331.cn 7.44e-19
C1332 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_127.cn 0.18f
C1333 comparator_0.vp dac_0.carray_0.unitcap_320.cn 0.496f
C1334 comparator_0.trim_0.n3 dac_1.carray_0.unitcap_334.cn 0.0133f
C1335 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_330.cn 0.145f
C1336 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln0 0.0827f
C1337 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_3.Y 4.37f
C1338 dac_0.sw_top_3.net1 vinp 0.368f
C1339 dac_1.carray_0.unitcap_48.cn dac_1.carray_0.unitcap_72.cn 0.0902f
C1340 dac_1.carray_0.unitcap_328.cn avdd 8.02e-19
C1341 comparator_0.trim_1.n3 trimb4 0.319f
C1342 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp1 0.00126f
C1343 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_326.cn 9.72e-19
C1344 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.sky130_fd_sc_hd__inv_2_6.Y 5.1e-21
C1345 dac_1.out dac_1.sky130_fd_sc_hd__inv_2_7.Y 0.541f
C1346 comparator_0.vp dac_1.carray_0.unitcap_23.cn 0.00925f
C1347 comparator_0.trim_1.n0 comparator_0.ip 0.556f
C1348 comparator_0.ip trimb3 0.102f
C1349 dac_1.out dac_1.carray_0.unitcap_56.cn 0.514f
C1350 comparator_0.vp dac_1.out 5.43f
C1351 comparator_0.outn avdd 0.83f
C1352 comparator_0.trim_0.n2 trim1 0.0074f
C1353 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_88.cn 0.18f
C1354 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_152.cn 0.18f
C1355 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp3 0.0829f
C1356 comparator_0.vp dac_1.carray_0.unitcap_231.cn 0.00925f
C1357 dac_0.carray_0.unitcap_48.cn dac_0.carray_0.unitcap_72.cn 0.0902f
C1358 dac_1.carray_0.unitcap_208.cn avdd 0.111f
C1359 dac_1.out dac_0.carray_0.unitcap_338.cn 0.00925f
C1360 dac_0.carray_0.unitcap_63.cn dac_1.carray_0.unitcap_63.cn 0.128f
C1361 dac_1.carray_0.unitcap_324.cn ctln1 0.00202f
C1362 comparator_0.trim_0.n4 dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.0024f
C1363 latch_0.Qn clkc 6.65e-19
C1364 comparator_0.ip trimb0 0.0297f
C1365 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp4 0.16f
C1366 dac_1.sky130_fd_sc_hd__inv_2_8.Y avdd 0.266f
C1367 comparator_0.trim_1.n2 avdd 0.024f
C1368 dac_1.sw_top_0.net1 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.402f
C1369 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_5.Y 1.42e-19
C1370 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_13.cn 0.0902f
C1371 dac_1.out dac_1.carray_0.unitcap_207.cn 0.51f
C1372 comparator_0.vp dac_0.carray_0.unitcap_321.cn 0.512f
C1373 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_103.cn 0.18f
C1374 dac_1.sky130_fd_sc_hd__inv_2_3.Y ctln6 1.78e-19
C1375 dac_1.carray_0.unitcap_191.cn dac_1.carray_0.unitcap_215.cn 0.0902f
C1376 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_4.Y 0.251f
C1377 dac_1.carray_0.unitcap_288.cn avdd 0.119f
C1378 dac_1.out dac_1.carray_0.unitcap_8.cn 0.503f
C1379 dac_1.carray_0.unitcap_232.cn dac_1.carray_0.unitcap_248.cn 0.0902f
C1380 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.sky130_fd_sc_hd__inv_2_7.Y 0.00132f
C1381 dac_0.carray_0.unitcap_7.cn dac_1.carray_0.unitcap_7.cn 0.128f
C1382 comparator_0.vp dac_1.carray_0.unitcap_15.cn 0.00762f
C1383 dac_1.out dac_1.carray_0.unitcap_32.cn 0.514f
C1384 dac_1.carray_0.unitcap_288.cn vinn 5.91e-19
C1385 dac_0.sky130_fd_sc_hd__inv_2_6.VPB comparator_0.trim_1.n3 0.011f
C1386 dac_0.carray_0.unitcap_87.cn dac_0.carray_0.unitcap_71.cn 0.0902f
C1387 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_64.cn 0.18f
C1388 dac_0.sky130_fd_sc_hd__inv_2_1.Y comparator_0.trim_1.n3 0.00755f
C1389 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_331.cn 0.0439f
C1390 dac_1.sw_top_2.en_buf dac_1.carray_0.unitcap_11.cn 0.00862f
C1391 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_128.cn 0.18f
C1392 dac_1.carray_0.unitcap_12.cn sample 0.0343f
C1393 comparator_0.vp dac_1.carray_0.unitcap_215.cn 0.00925f
C1394 dac_1.carray_0.unitcap_184.cn avdd 0.0995f
C1395 dac_1.out dac_0.carray_0.unitcap_255.cn 0.00925f
C1396 dac_0.carray_0.unitcap_232.cn dac_0.carray_0.unitcap_248.cn 0.0902f
C1397 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_256.cn 0.0902f
C1398 comparator_0.trim_1.n1 comparator_0.ip 0.578f
C1399 dac_0.carray_0.unitcap_247.cn dac_1.carray_0.unitcap_247.cn 0.128f
C1400 comparator_0.trim_1.n4 trimb1 0.0143f
C1401 comparator_0.trim_1.n3 ctlp5 0.00164f
C1402 dac_1.sky130_fd_sc_hd__inv_2_1.Y ctln7 0.0531f
C1403 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_330.cn 7.44e-19
C1404 dac_1.out dac_1.carray_0.unitcap_199.cn 0.51f
C1405 comparator_0.trim_0.n3 dac_1.carray_0.unitcap_331.cn 0.0187f
C1406 comparator_0.vp dac_0.carray_0.unitcap_248.cn 0.514f
C1407 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_111.cn 0.18f
C1408 dac_1.sky130_fd_sc_hd__inv_2_1.Y dac_1.carray_0.unitcap_337.cn 0.13f
C1409 dac_1.carray_0.unitcap_56.cn dac_1.carray_0.unitcap_48.cn 0.0902f
C1410 dac_1.out dac_1.carray_0.unitcap_324.cn 0.505f
C1411 dac_1.carray_0.unitcap_326.cn avdd 5.03e-19
C1412 trimb4 trimb3 0.0194f
C1413 comparator_0.ip ctlp6 0.00368f
C1414 dac_1.sky130_fd_sc_hd__inv_2_6.VPB ctln5 0.0826f
C1415 comparator_0.vp dac_0.carray_0.unitcap_336.cn 0.64f
C1416 dac_1.out dac_1.carray_0.unitcap_40.cn 0.514f
C1417 dac_0.sky130_fd_sc_hd__inv_2_0.Y dac_0.carray_0.unitcap_328.cn 0.00171f
C1418 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_322.cn 0.00396f
C1419 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_80.cn 0.18f
C1420 dac_0.carray_0.unitcap_56.cn dac_0.carray_0.unitcap_48.cn 0.0902f
C1421 dac_0.carray_0.unitcap_338.cn dac_0.carray_0.unitcap_336.cn 0.0902f
C1422 comparator_0.vp dac_1.carray_0.unitcap_191.cn 0.00925f
C1423 comparator_0.trim_0.n4 dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.0524f
C1424 dac_1.out dac_0.carray_0.unitcap_239.cn 0.00925f
C1425 dac_1.carray_0.unitcap_200.cn avdd 0.11f
C1426 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y 3.2e-19
C1427 dac_0.sw_top_0.net1 vinp 0.368f
C1428 dac_0.carray_0.unitcap_39.cn dac_1.carray_0.unitcap_39.cn 0.128f
C1429 dac_1.sky130_fd_sc_hd__inv_2_3.Y dac_1.sky130_fd_sc_hd__inv_2_7.Y 0.0925f
C1430 trimb2 clkc 4.96e-19
C1431 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_12.cn 0.0902f
C1432 dac_1.out dac_1.carray_0.unitcap_175.cn 0.51f
C1433 dac_0.sky130_fd_sc_hd__inv_2_0.Y avdd 0.294f
C1434 comparator_0.trim_1.n4 comparator_0.in 0.0138f
C1435 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_95.cn 0.18f
C1436 dac_0.sw_top_3.net1 avdd 0.849f
C1437 comparator_0.vp dac_0.carray_0.unitcap_232.cn 0.514f
C1438 dac_1.sky130_fd_sc_hd__inv_2_5.Y ctln3 0.0494f
C1439 dac_1.carray_0.unitcap_207.cn dac_1.carray_0.unitcap_191.cn 0.0902f
C1440 comparator_0.outp dac_1.out 0.017f
C1441 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.sky130_fd_sc_hd__inv_2_6.Y 0.543f
C1442 dac_1.carray_0.unitcap_10.cn avdd 0.021f
C1443 dac_1.sky130_fd_sc_hd__inv_2_4.Y dac_1.carray_0.unitcap_324.cn 0.00391f
C1444 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp7 2.79e-20
C1445 dac_1.sky130_fd_sc_hd__inv_2_6.Y dac_1.carray_0.unitcap_322.cn 0.275f
C1446 comparator_0.trim_0.n3 clkc 6.61e-19
C1447 dac_1.carray_0.unitcap_240.cn dac_1.carray_0.unitcap_232.cn 0.0902f
C1448 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.sky130_fd_sc_hd__inv_2_8.Y 1.89f
C1449 dac_0.carray_0.unitcap_31.cn dac_1.carray_0.unitcap_31.cn 0.128f
C1450 comparator_0.vp dac_0.carray_0.unitcap_338.cn 0.526f
C1451 dac_1.out dac_0.carray_0.unitcap_7.cn 0.00925f
C1452 dac_1.carray_0.unitcap_10.cn vinn 0.0189f
C1453 comparator_0.ip dac_0.carray_0.unitcap_337.cn 0.00341f
C1454 dac_0.carray_0.unitcap_79.cn dac_0.carray_0.unitcap_87.cn 0.0902f
C1455 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_72.cn 0.18f
C1456 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_330.cn 0.039f
C1457 comparator_0.vp dac_1.carray_0.unitcap_207.cn 0.00925f
C1458 dac_1.carray_0.unitcap_14.cn sample 0.0343f
C1459 dac_1.carray_0.unitcap_192.cn avdd 0.111f
C1460 dac_1.out dac_0.carray_0.unitcap_247.cn 0.00925f
C1461 dac_1.sky130_fd_sc_hd__inv_2_2.Y ctln7 0.16f
C1462 comparator_0.vp dac_0.carray_0.unitcap_0.cn 0.514f
C1463 dac_0.carray_0.unitcap_240.cn dac_0.carray_0.unitcap_232.cn 0.0902f
C1464 avdd ctlp1 0.119f
C1465 dac_0.carray_0.unitcap_223.cn dac_1.carray_0.unitcap_223.cn 0.128f
C1466 dac_1.out dac_1.carray_0.unitcap_183.cn 0.51f
C1467 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_337.cn 0.138f
C1468 ctln1 ctln0 0.105f
C1469 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_71.cn 0.18f
C1470 comparator_0.vp dac_0.carray_0.unitcap_240.cn 0.514f
C1471 comparator_0.in ctln3 4.02e-19
C1472 dac_1.carray_0.unitcap_32.cn dac_1.carray_0.unitcap_56.cn 0.0902f
C1473 dac_0.carray_0.unitcap_326.cn ctlp7 0.00199f
C1474 comparator_0.vp ctlp3 9.29e-19
C1475 comparator_0.vp dac_0.carray_0.unitcap_255.cn 0.511f
C1476 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_136.cn 0.18f
C1477 dac_1.out dac_0.carray_0.unitcap_31.cn 0.00925f
C1478 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_328.cn 0.123f
C1479 dac_1.sw_top_3.net1 avdd 0.849f
C1480 comparator_0.trim_0.n3 trim3 0.231f
C1481 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_48.cn 0.18f
C1482 dac_0.carray_0.unitcap_32.cn dac_0.carray_0.unitcap_56.cn 0.0902f
C1483 dac_1.carray_0.unitcap_168.cn avdd 0.0728f
C1484 dac_0.carray_0.unitcap_255.cn dac_0.carray_0.unitcap_338.cn 0.0902f
C1485 comparator_0.vp dac_1.carray_0.unitcap_199.cn 0.00925f
C1486 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_1.Y 0.00854f
C1487 dac_1.out dac_0.carray_0.unitcap_223.cn 0.00925f
C1488 comparator_0.trim_0.n4 comparator_0.trim_0.n3 0.461f
C1489 dac_0.carray_0.unitcap_47.cn dac_1.carray_0.unitcap_47.cn 0.128f
C1490 dac_1.sky130_fd_sc_hd__inv_2_7.Y dac_1.carray_0.unitcap_324.cn 0.289f
C1491 comparator_0.vp dac_0.carray_0.unitcap_24.cn 0.514f
C1492 dac_0.sky130_fd_sc_hd__inv_2_7.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y 2.23e-21
C1493 dac_1.sw_top_3.net1 vinn 0.368f
C1494 dac_1.carray_0.unitcap_24.cn dac_1.carray_0.unitcap_0.cn 0.0902f
C1495 dac_0.sky130_fd_sc_hd__inv_2_5.Y ctlp4 2.49e-19
C1496 dac_1.out dac_1.carray_0.unitcap_167.cn 0.51f
C1497 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_14.cn 0.0902f
C1498 comparator_0.vp dac_0.carray_0.unitcap_216.cn 0.514f
C1499 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_87.cn 0.18f
C1500 comparator_0.diff clkc 0.104f
C1501 dac_1.carray_0.unitcap_199.cn dac_1.carray_0.unitcap_207.cn 0.0902f
C1502 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.sky130_fd_sc_hd__inv_2_5.Y 0.246f
C1503 comparator_0.trim_1.n2 trimb1 0.0074f
C1504 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.sky130_fd_sc_hd__inv_2_4.Y 0.571f
C1505 dac_0.sky130_fd_sc_hd__inv_2_8.Y ctlp2 4.16e-20
C1506 dac_1.carray_0.unitcap_11.cn avdd 0.00997f
C1507 comparator_0.vp comparator_0.trim_1.n3 0.00141f
C1508 dac_0.sky130_fd_sc_hd__inv_2_6.VPB ctlp6 0.0828f
C1509 dac_1.carray_0.unitcap_256.cn dac_1.carray_0.unitcap_9.cn 0.18f
C1510 comparator_0.in trim4 0.104f
C1511 dac_1.carray_0.unitcap_216.cn dac_1.carray_0.unitcap_240.cn 0.0902f
C1512 dac_1.out ctln0 6.77e-19
C1513 dac_0.sky130_fd_sc_hd__inv_2_1.Y ctlp6 0.159f
C1514 dac_0.carray_0.unitcap_24.cn dac_0.carray_0.unitcap_0.cn 0.0902f
C1515 dac_0.carray_0.unitcap_23.cn dac_1.carray_0.unitcap_23.cn 0.128f
C1516 comparator_0.vp dac_0.carray_0.unitcap_239.cn 0.51f
C1517 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_200.cn 0.18f
C1518 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_112.cn 0.18f
C1519 dac_1.carray_0.unitcap_11.cn vinn 0.0736f
C1520 dac_0.carray_0.unitcap_55.cn dac_0.carray_0.unitcap_79.cn 0.0902f
C1521 dac_1.sky130_fd_sc_hd__inv_2_0.Y ctln7 2.65e-19
C1522 comparator_0.ip dac_0.carray_0.unitcap_330.cn 0.00296f
C1523 dac_1.out dac_0.carray_0.unitcap_23.cn 0.00925f
C1524 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_56.cn 0.18f
C1525 ctlp5 ctlp6 0.105f
C1526 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_337.cn 0.00682f
C1527 dac_0.sw_top_0.net1 avdd 0.848f
C1528 comparator_0.vp dac_1.carray_0.unitcap_175.cn 0.00925f
C1529 dac_0.sky130_fd_sc_hd__inv_2_2.Y comparator_0.trim_1.n4 0.0583f
C1530 dac_1.carray_0.unitcap_176.cn avdd 0.11f
C1531 dac_1.carray_0.unitcap_322.cn ctln3 0.00202f
C1532 dac_1.out dac_0.carray_0.unitcap_231.cn 0.00925f
C1533 comparator_0.vp dac_0.carray_0.unitcap_16.cn 0.515f
C1534 dac_0.sky130_fd_sc_hd__inv_2_6.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y 0.0961f
C1535 dac_0.carray_0.unitcap_216.cn dac_0.carray_0.unitcap_240.cn 0.0902f
C1536 comparator_0.vp comparator_0.outp 0.0147f
C1537 dac_0.carray_0.unitcap_231.cn dac_1.carray_0.unitcap_231.cn 0.128f
C1538 comparator_0.trim_0.n3 ctln7 0.0071f
C1539 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.carray_0.unitcap_334.cn 2.28e-19
C1540 dac_1.out dac_1.carray_0.unitcap_151.cn 0.51f
C1541 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_336.cn 0.161f
C1542 comparator_0.vp dac_0.carray_0.unitcap_224.cn 0.514f
C1543 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_79.cn 0.18f
C1544 comparator_0.in comparator_0.outn 0.412f
C1545 trim2 trim1 0.0834f
C1546 dac_1.carray_0.unitcap_40.cn dac_1.carray_0.unitcap_32.cn 0.0902f
C1547 comparator_0.vp dac_0.carray_0.unitcap_7.cn 0.51f
C1548 comparator_0.in dac_1.sky130_fd_sc_hd__inv_2_8.Y 0.0133f
C1549 ctln4 ctln2 3.27e-21
C1550 dac_0.sky130_fd_sc_hd__inv_2_8.Y comparator_0.ip 0.0141f
C1551 dac_1.sky130_fd_sc_hd__inv_2_4.Y ctln0 0.00131f
C1552 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_232.cn 0.18f
C1553 a_33300_6679# avdd 0.385f
C1554 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_120.cn 0.18f
C1555 comparator_0.vp dac_0.carray_0.unitcap_247.cn 0.51f
C1556 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_192.cn 0.18f
C1557 dac_1.out dac_0.carray_0.unitcap_15.cn 0.00762f
C1558 dac_1.sky130_fd_sc_hd__inv_2_5.Y dac_1.carray_0.unitcap_326.cn 0.34f
C1559 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_2.Y 0.0152f
C1560 dac_0.sky130_fd_sc_hd__inv_2_3.Y dac_0.carray_0.unitcap_334.cn 0.0355f
C1561 dac_1.out dac_1.sw_top_2.net1 0.324f
C1562 comparator_0.diff comparator_0.trim_0.n4 0.00526f
C1563 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_32.cn 0.18f
C1564 comparator_0.vp dac_1.carray_0.unitcap_183.cn 0.00925f
C1565 dac_0.carray_0.unitcap_239.cn dac_0.carray_0.unitcap_255.cn 0.0902f
C1566 dac_0.carray_0.unitcap_40.cn dac_0.carray_0.unitcap_32.cn 0.0902f
C1567 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_337.cn 0.13f
C1568 dac_1.carray_0.unitcap_160.cn avdd 0.111f
C1569 dac_1.out dac_0.carray_0.unitcap_215.cn 0.00925f
C1570 comparator_0.trim_0.n4 comparator_0.trim_0.n0 0.0519f
C1571 avdd ctlp7 0.119f
C1572 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.sky130_fd_sc_hd__inv_2_5.Y 0.736f
C1573 comparator_0.trim_0.n0 trim0 0.117f
C1574 dac_1.carray_0.unitcap_16.cn dac_1.carray_0.unitcap_24.cn 0.0902f
C1575 dac_1.out dac_1.carray_0.unitcap_159.cn 0.51f
C1576 comparator_0.trim_1.n4 comparator_0.outn 0.011f
C1577 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_338.cn 0.161f
C1578 comparator_0.vp dac_0.carray_0.unitcap_208.cn 0.514f
C1579 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_55.cn 0.18f
C1580 dac_1.carray_0.unitcap_175.cn dac_1.carray_0.unitcap_199.cn 0.0902f
C1581 dac_1.sw_top_0.net1 avdd 0.848f
C1582 dac_1.carray_0.unitcap_13.cn avdd 0.0016f
C1583 comparator_0.trim_1.n4 comparator_0.trim_1.n2 0.178f
C1584 dac_1.carray_0.unitcap_328.cn dac_1.carray_0.unitcap_322.cn 0.18f
C1585 comparator_0.vp dac_0.carray_0.unitcap_31.cn 0.51f
C1586 dac_1.carray_0.unitcap_224.cn dac_1.carray_0.unitcap_216.cn 0.0902f
C1587 dac_0.carray_0.unitcap_324.cn ctlp1 0.00202f
C1588 dac_0.carray_0.unitcap_16.cn dac_0.carray_0.unitcap_24.cn 0.0902f
C1589 dac_1.sky130_fd_sc_hd__inv_2_8.Y dac_1.carray_0.unitcap_240.cn 0.18f
C1590 avdd clkc 1.01f
C1591 latch_0.Qn comparator_0.ip 0.00459f
C1592 comparator_0.vp dac_0.carray_0.unitcap_223.cn 0.51f
C1593 dac_1.sw_top_0.net1 vinn 0.368f
C1594 dac_0.sky130_fd_sc_hd__inv_2_5.Y dac_0.sky130_fd_sc_hd__inv_2_3.Y 1.12f
C1595 dac_0.carray_0.unitcap_15.cn dac_1.carray_0.unitcap_15.cn 0.128f
C1596 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_96.cn 0.18f
C1597 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_168.cn 0.18f
C1598 dac_1.carray_0.unitcap_13.cn vinn 0.0215f
C1599 dac_0.carray_0.unitcap_63.cn dac_0.carray_0.unitcap_55.cn 0.0902f
C1600 comparator_0.ip dac_0.carray_0.unitcap_331.cn 0.00296f
C1601 dac_0.sky130_fd_sc_hd__inv_2_6.Y ctlp2 3.42e-19
C1602 dac_1.sky130_fd_sc_hd__inv_2_0.Y dac_1.carray_0.unitcap_336.cn 0.00213f
C1603 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_40.cn 0.18f
C1604 comparator_0.vp dac_1.carray_0.unitcap_167.cn 0.00925f
C1605 avdd ctln2 0.118f
C1606 dac_1.out ctln5 9.28e-19
C1607 dac_1.carray_0.unitcap_144.cn avdd 0.077f
C1608 dac_1.out dac_0.carray_0.unitcap_191.cn 0.00925f
C1609 ctlp0 ctlp1 0.107f
C1610 dac_0.sw_top_2.net1 comparator_0.vp 0.324f
C1611 dac_0.carray_0.unitcap_224.cn dac_0.carray_0.unitcap_216.cn 0.0902f
C1612 comparator_0.trim_1.n3 comparator_0.outp 1.93e-20
C1613 comparator_0.trim_0.n1 trim3 0.00122f
C1614 dac_0.carray_0.unitcap_215.cn dac_1.carray_0.unitcap_215.cn 0.128f
C1615 dac_0.sky130_fd_sc_hd__inv_2_4.Y dac_0.carray_0.unitcap_326.cn 0.091f
C1616 dac_0.sky130_fd_sc_hd__inv_2_1.Y dac_0.carray_0.unitcap_207.cn 0.18f
C1617 dac_0.sw_top_0.net1 dac_0.carray_0.unitcap_64.cn 1e-20
C1618 dac_1.out dac_1.carray_0.unitcap_135.cn 0.51f
C1619 dac_1.sky130_fd_sc_hd__inv_2_7.Y ctln0 0.0476f
C1620 dac_1.sky130_fd_sc_hd__inv_2_2.Y dac_1.carray_0.unitcap_255.cn 0.161f
C1621 dac_0.carray_0.unitcap_328.cn ctlp4 6.13e-19
C1622 dac_0.sky130_fd_sc_hd__inv_2_2.Y dac_0.carray_0.unitcap_63.cn 0.18f
C1623 comparator_0.trim_0.n4 comparator_0.trim_0.n1 0.0526f
C1624 comparator_0.trim_0.n3 comparator_0.trim_0.n2 0.264f
C1625 comparator_0.vp dac_0.carray_0.unitcap_184.cn 0.514f
C1626 dac_0.sky130_fd_sc_hd__inv_2_8.Y trimb4 5.48e-20
C1627 comparator_0.trim_0.n1 trim0 0.00397f
C1628 dac_1.sw_top_0.en_buf dac_1.carray_0.unitcap_80.cn 5.45e-19
C1629 dac_1.sky130_fd_sc_hd__inv_2_6.VPB dac_1.sky130_fd_sc_hd__inv_2_0.Y 0.0089f
C1630 comparator_0.vp dac_0.carray_0.unitcap_23.cn 0.512f
C1631 ctln0 avss 0.429f
C1632 ctln1 avss 0.33f
C1633 ctln2 avss 0.329f
C1634 ctln3 avss 0.33f
C1635 ctln4 avss 0.33f
C1636 ctln5 avss 0.329f
C1637 ctln6 avss 0.328f
C1638 ctln7 avss 0.393f
C1639 vinn avss 5.32f
C1640 trim0 avss 0.878f
C1641 trim1 avss 0.707f
C1642 trim2 avss 0.914f
C1643 trim3 avss 1.32f
C1644 trim4 avss 2.1f
C1645 clkc avss 2.83f
C1646 trimb0 avss 0.761f
C1647 trimb1 avss 0.64f
C1648 trimb2 avss 0.864f
C1649 trimb3 avss 1.25f
C1650 trimb4 avss 2.05f
C1651 ctlp7 avss 0.392f
C1652 vinp avss 5.34f
C1653 ctlp6 avss 0.328f
C1654 ctlp5 avss 0.33f
C1655 ctlp4 avss 0.33f
C1656 sample avss 16.1f
C1657 ctlp3 avss 0.33f
C1658 ctlp2 avss 0.331f
C1659 ctlp1 avss 0.331f
C1660 ctlp0 avss 0.333f
C1661 avdd avss 8.19p
C1662 dac_1.carray_0.unitcap_320.cn avss 0.21f
C1663 dac_1.carray_0.unitcap_321.cn avss 0.185f
C1664 dac_1.carray_0.unitcap_248.cn avss 0.147f
C1665 dac_1.carray_0.unitcap_232.cn avss 0.147f
C1666 dac_1.carray_0.unitcap_240.cn avss 0.162f
C1667 dac_1.carray_0.unitcap_216.cn avss 0.146f
C1668 dac_1.carray_0.unitcap_224.cn avss 0.147f
C1669 dac_1.carray_0.unitcap_208.cn avss 0.147f
C1670 dac_1.carray_0.unitcap_184.cn avss 0.158f
C1671 dac_1.carray_0.unitcap_200.cn avss 0.147f
C1672 dac_1.carray_0.unitcap_192.cn avss 0.147f
C1673 dac_1.carray_0.unitcap_168.cn avss 0.183f
C1674 dac_1.carray_0.unitcap_176.cn avss 0.147f
C1675 dac_1.carray_0.unitcap_160.cn avss 0.147f
C1676 dac_1.carray_0.unitcap_144.cn avss 0.178f
C1677 dac_1.carray_0.unitcap_152.cn avss 0.146f
C1678 dac_1.carray_0.unitcap_128.cn avss 0.146f
C1679 dac_1.carray_0.unitcap_136.cn avss 0.154f
C1680 dac_1.carray_0.unitcap_112.cn avss 0.146f
C1681 dac_1.carray_0.unitcap_120.cn avss 0.146f
C1682 dac_1.carray_0.unitcap_96.cn avss 0.146f
C1683 dac_1.carray_0.unitcap_104.cn avss 0.165f
C1684 dac_1.carray_0.unitcap_88.cn avss 0.146f
C1685 dac_1.carray_0.unitcap_64.cn avss 0.151f
C1686 dac_1.carray_0.unitcap_80.cn avss 0.189f
C1687 dac_1.carray_0.unitcap_72.cn avss 0.151f
C1688 dac_1.carray_0.unitcap_48.cn avss 0.151f
C1689 dac_1.carray_0.unitcap_56.cn avss 0.176f
C1690 dac_1.carray_0.unitcap_32.cn avss 0.151f
C1691 dac_1.carray_0.unitcap_40.cn avss 0.151f
C1692 dac_1.carray_0.unitcap_0.cn avss 0.151f
C1693 dac_1.carray_0.unitcap_24.cn avss 0.153f
C1694 dac_1.carray_0.unitcap_16.cn avss 0.151f
C1695 dac_1.carray_0.unitcap_8.cn avss 0.234f
C1696 dac_1.carray_0.unitcap_324.cn avss 0.165f
C1697 dac_1.carray_0.unitcap_9.cn avss 0.218f
C1698 dac_1.carray_0.unitcap_322.cn avss 0.163f
C1699 dac_1.carray_0.unitcap_256.cn avss 0.252f
C1700 dac_1.carray_0.unitcap_328.cn avss 0.164f
C1701 dac_1.carray_0.unitcap_288.cn avss 0.179f
C1702 dac_1.carray_0.unitcap_326.cn avss 0.157f
C1703 dac_1.carray_0.unitcap_10.cn avss 0.199f
C1704 dac_1.carray_0.unitcap_334.cn avss 0.137f
C1705 dac_1.carray_0.unitcap_11.cn avss 0.184f
C1706 dac_1.carray_0.unitcap_331.cn avss 0.152f
C1707 dac_1.carray_0.unitcap_13.cn avss 0.199f
C1708 dac_1.carray_0.unitcap_330.cn avss 0.172f
C1709 dac_1.carray_0.unitcap_12.cn avss 0.199f
C1710 dac_1.carray_0.unitcap_337.cn avss 0.144f
C1711 dac_1.carray_0.unitcap_14.cn avss 0.199f
C1712 dac_1.carray_0.unitcap_336.cn avss 0.185f
C1713 dac_1.carray_0.unitcap_338.cn avss 0.118f
C1714 dac_1.carray_0.unitcap_255.cn avss 0.118f
C1715 dac_1.carray_0.unitcap_239.cn avss 0.118f
C1716 dac_1.carray_0.unitcap_247.cn avss 0.118f
C1717 dac_1.carray_0.unitcap_223.cn avss 0.118f
C1718 dac_1.carray_0.unitcap_231.cn avss 0.118f
C1719 dac_1.carray_0.unitcap_215.cn avss 0.118f
C1720 dac_1.carray_0.unitcap_191.cn avss 0.118f
C1721 dac_1.carray_0.unitcap_207.cn avss 0.118f
C1722 dac_1.carray_0.unitcap_199.cn avss 0.118f
C1723 dac_1.carray_0.unitcap_175.cn avss 0.118f
C1724 dac_1.carray_0.unitcap_183.cn avss 0.118f
C1725 dac_1.carray_0.unitcap_167.cn avss 0.118f
C1726 dac_1.carray_0.unitcap_151.cn avss 0.118f
C1727 dac_1.carray_0.unitcap_159.cn avss 0.118f
C1728 dac_1.carray_0.unitcap_135.cn avss 0.118f
C1729 dac_1.carray_0.unitcap_143.cn avss 0.124f
C1730 dac_1.carray_0.unitcap_119.cn avss 0.124f
C1731 dac_1.carray_0.unitcap_127.cn avss 0.124f
C1732 dac_1.carray_0.unitcap_103.cn avss 0.124f
C1733 dac_1.carray_0.unitcap_111.cn avss 0.124f
C1734 dac_1.carray_0.unitcap_95.cn avss 0.124f
C1735 dac_1.carray_0.unitcap_71.cn avss 0.124f
C1736 dac_1.carray_0.unitcap_87.cn avss 0.124f
C1737 dac_1.carray_0.unitcap_79.cn avss 0.124f
C1738 dac_1.carray_0.unitcap_55.cn avss 0.124f
C1739 dac_1.carray_0.unitcap_63.cn avss 0.124f
C1740 dac_1.carray_0.unitcap_39.cn avss 0.124f
C1741 dac_1.carray_0.unitcap_47.cn avss 0.124f
C1742 dac_1.carray_0.unitcap_7.cn avss 0.124f
C1743 dac_1.carray_0.unitcap_31.cn avss 0.124f
C1744 dac_1.carray_0.unitcap_23.cn avss 0.124f
C1745 dac_1.carray_0.unitcap_15.cn avss 0.205f
C1746 dac_0.carray_0.unitcap_336.cn avss 0.187f
C1747 dac_0.carray_0.unitcap_338.cn avss 0.118f
C1748 dac_0.carray_0.unitcap_255.cn avss 0.118f
C1749 dac_0.carray_0.unitcap_239.cn avss 0.118f
C1750 dac_0.carray_0.unitcap_247.cn avss 0.118f
C1751 dac_0.carray_0.unitcap_223.cn avss 0.118f
C1752 dac_0.carray_0.unitcap_231.cn avss 0.118f
C1753 dac_0.carray_0.unitcap_215.cn avss 0.118f
C1754 dac_0.carray_0.unitcap_191.cn avss 0.118f
C1755 dac_0.carray_0.unitcap_207.cn avss 0.118f
C1756 dac_0.carray_0.unitcap_199.cn avss 0.118f
C1757 dac_0.carray_0.unitcap_175.cn avss 0.118f
C1758 dac_0.carray_0.unitcap_183.cn avss 0.118f
C1759 dac_0.carray_0.unitcap_167.cn avss 0.118f
C1760 dac_0.carray_0.unitcap_151.cn avss 0.118f
C1761 dac_0.carray_0.unitcap_159.cn avss 0.118f
C1762 dac_0.carray_0.unitcap_135.cn avss 0.118f
C1763 dac_0.carray_0.unitcap_143.cn avss 0.124f
C1764 dac_0.carray_0.unitcap_119.cn avss 0.124f
C1765 dac_0.carray_0.unitcap_127.cn avss 0.124f
C1766 dac_0.carray_0.unitcap_103.cn avss 0.124f
C1767 dac_0.carray_0.unitcap_111.cn avss 0.124f
C1768 dac_0.carray_0.unitcap_95.cn avss 0.124f
C1769 dac_0.carray_0.unitcap_71.cn avss 0.124f
C1770 dac_0.carray_0.unitcap_87.cn avss 0.124f
C1771 dac_0.carray_0.unitcap_79.cn avss 0.124f
C1772 dac_0.carray_0.unitcap_55.cn avss 0.124f
C1773 dac_0.carray_0.unitcap_63.cn avss 0.124f
C1774 dac_0.carray_0.unitcap_39.cn avss 0.124f
C1775 dac_0.carray_0.unitcap_47.cn avss 0.124f
C1776 dac_0.carray_0.unitcap_7.cn avss 0.124f
C1777 dac_0.carray_0.unitcap_31.cn avss 0.124f
C1778 dac_0.carray_0.unitcap_23.cn avss 0.124f
C1779 dac_0.carray_0.unitcap_15.cn avss 0.205f
C1780 dac_0.carray_0.unitcap_337.cn avss 0.145f
C1781 dac_0.carray_0.unitcap_14.cn avss 0.199f
C1782 dac_0.carray_0.unitcap_330.cn avss 0.169f
C1783 dac_0.carray_0.unitcap_12.cn avss 0.199f
C1784 dac_0.carray_0.unitcap_331.cn avss 0.151f
C1785 dac_0.carray_0.unitcap_13.cn avss 0.199f
C1786 dac_0.carray_0.unitcap_334.cn avss 0.132f
C1787 dac_0.carray_0.unitcap_11.cn avss 0.184f
C1788 dac_0.carray_0.unitcap_326.cn avss 0.157f
C1789 dac_0.carray_0.unitcap_10.cn avss 0.199f
C1790 dac_0.carray_0.unitcap_328.cn avss 0.164f
C1791 dac_0.carray_0.unitcap_288.cn avss 0.179f
C1792 dac_0.carray_0.unitcap_322.cn avss 0.163f
C1793 dac_0.carray_0.unitcap_256.cn avss 0.252f
C1794 dac_0.carray_0.unitcap_324.cn avss 0.165f
C1795 dac_0.carray_0.unitcap_9.cn avss 0.219f
C1796 dac_0.carray_0.unitcap_320.cn avss 0.213f
C1797 dac_0.carray_0.unitcap_321.cn avss 0.179f
C1798 dac_0.carray_0.unitcap_248.cn avss 0.151f
C1799 dac_0.carray_0.unitcap_232.cn avss 0.151f
C1800 dac_0.carray_0.unitcap_240.cn avss 0.157f
C1801 dac_0.carray_0.unitcap_216.cn avss 0.151f
C1802 dac_0.carray_0.unitcap_224.cn avss 0.151f
C1803 dac_0.carray_0.unitcap_208.cn avss 0.151f
C1804 dac_0.carray_0.unitcap_184.cn avss 0.17f
C1805 dac_0.carray_0.unitcap_200.cn avss 0.151f
C1806 dac_0.carray_0.unitcap_192.cn avss 0.151f
C1807 dac_0.carray_0.unitcap_168.cn avss 0.186f
C1808 dac_0.carray_0.unitcap_176.cn avss 0.151f
C1809 dac_0.carray_0.unitcap_160.cn avss 0.151f
C1810 dac_0.carray_0.unitcap_144.cn avss 0.172f
C1811 dac_0.carray_0.unitcap_152.cn avss 0.151f
C1812 dac_0.carray_0.unitcap_128.cn avss 0.151f
C1813 dac_0.carray_0.unitcap_136.cn avss 0.151f
C1814 dac_0.carray_0.unitcap_112.cn avss 0.155f
C1815 dac_0.carray_0.unitcap_120.cn avss 0.151f
C1816 dac_0.carray_0.unitcap_96.cn avss 0.151f
C1817 dac_0.carray_0.unitcap_104.cn avss 0.177f
C1818 dac_0.carray_0.unitcap_88.cn avss 0.151f
C1819 dac_0.carray_0.unitcap_64.cn avss 0.157f
C1820 dac_0.carray_0.unitcap_80.cn avss 0.191f
C1821 dac_0.carray_0.unitcap_72.cn avss 0.156f
C1822 dac_0.carray_0.unitcap_48.cn avss 0.156f
C1823 dac_0.carray_0.unitcap_56.cn avss 0.17f
C1824 dac_0.carray_0.unitcap_32.cn avss 0.156f
C1825 dac_0.carray_0.unitcap_40.cn avss 0.156f
C1826 dac_0.carray_0.unitcap_0.cn avss 0.156f
C1827 dac_0.carray_0.unitcap_24.cn avss 0.166f
C1828 dac_0.carray_0.unitcap_16.cn avss 0.158f
C1829 dac_0.carray_0.unitcap_8.cn avss 0.239f
C1830 dac_1.sky130_fd_sc_hd__inv_2_7.Y avss 1.08f
C1831 dac_1.sky130_fd_sc_hd__inv_2_6.Y avss 0.841f
C1832 dac_1.sky130_fd_sc_hd__inv_2_4.Y avss 1.16f
C1833 dac_1.sky130_fd_sc_hd__inv_2_5.Y avss 2.65f
C1834 dac_1.sky130_fd_sc_hd__inv_2_3.Y avss 4.9f
C1835 dac_1.sky130_fd_sc_hd__inv_2_8.Y avss 14.8f
C1836 dac_1.sky130_fd_sc_hd__inv_2_0.Y avss 28.5f
C1837 dac_1.sky130_fd_sc_hd__inv_2_1.Y avss 55.3f
C1838 dac_1.sky130_fd_sc_hd__inv_2_2.Y avss 0.118p
C1839 dac_1.sw_top_0.net1 avss 1.99f
C1840 dac_1.sw_top_1.net1 avss 1.97f
C1841 dac_1.sw_top_3.net1 avss 1.97f
C1842 dac_1.sw_top_2.net1 avss 1.97f
C1843 dac_1.sw_top_0.en_buf avss 1.86f
C1844 dac_1.sw_top_1.en_buf avss 1.61f
C1845 dac_1.sw_top_3.en_buf avss 1.61f
C1846 dac_1.sw_top_2.en_buf avss 1.62f
C1847 comparator_0.trim_0.n0 avss 0.618f
C1848 comparator_0.trim_0.n1 avss 0.473f
C1849 comparator_0.trim_0.n2 avss 1.18f
C1850 comparator_0.trim_0.n3 avss 2.62f
C1851 comparator_0.trim_0.n4 avss 4.74f
C1852 a_33300_5579# avss 0.736f
C1853 comparator_0.outn avss 1.89f
C1854 comparator_0.in avss 5.51f
C1855 dac_1.out avss 0.18p
C1856 comparator_0.ip avss 5.2f
C1857 comparator_0.diff avss 0.562f
C1858 latch_0.Qn avss 1.11f
C1859 a_33300_6679# avss 0.701f
C1860 comparator_0.outp avss 2.12f
C1861 comparator_0.trim_1.n0 avss 0.596f
C1862 comparator_0.trim_1.n1 avss 0.463f
C1863 comparator_0.trim_1.n2 avss 1.17f
C1864 comparator_0.trim_1.n3 avss 2.15f
C1865 comparator_0.trim_1.n4 avss 4.56f
C1866 dac_0.sky130_fd_sc_hd__inv_2_2.Y avss 0.118p
C1867 comparator_0.vp avss 0.181p
C1868 dac_0.sky130_fd_sc_hd__inv_2_1.Y avss 55.7f
C1869 dac_0.sky130_fd_sc_hd__inv_2_0.Y avss 28.4f
C1870 dac_0.sky130_fd_sc_hd__inv_2_8.Y avss 14.4f
C1871 dac_0.sw_top_0.net1 avss 1.98f
C1872 dac_0.sw_top_1.net1 avss 1.96f
C1873 dac_0.sw_top_3.net1 avss 1.96f
C1874 dac_0.sw_top_2.net1 avss 1.97f
C1875 dac_0.sw_top_0.en_buf avss 1.86f
C1876 dac_0.sw_top_1.en_buf avss 1.61f
C1877 dac_0.sw_top_3.en_buf avss 1.61f
C1878 dac_0.sw_top_2.en_buf avss 1.62f
C1879 dac_0.sky130_fd_sc_hd__inv_2_3.Y avss 5.85f
C1880 dac_0.sky130_fd_sc_hd__inv_2_5.Y avss 2.65f
C1881 dac_0.sky130_fd_sc_hd__inv_2_4.Y avss 1.16f
C1882 dac_0.sky130_fd_sc_hd__inv_2_6.Y avss 0.84f
C1883 dac_0.sky130_fd_sc_hd__inv_2_7.Y avss 0.945f
C1884 dac_1.sky130_fd_sc_hd__inv_2_6.VPB avss 3.14f
C1885 dac_0.sky130_fd_sc_hd__inv_2_6.VPB avss 3.03f
C1886 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t0 avss 0.762f
C1887 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t4 avss 0.00265f
C1888 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t1 avss 0.00265f
C1889 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n0 avss 0.00626f
C1890 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n1 avss 0.00376f
C1891 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n2 avss 0.091f
C1892 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t2 avss 0.00407f
C1893 dac_1.sky130_fd_sc_hd__inv_2_5.Y.t3 avss 0.00407f
C1894 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n3 avss 0.0104f
C1895 dac_1.sky130_fd_sc_hd__inv_2_5.Y.n4 avss 0.0179f
C1896 comparator_0.ip.t15 avss 0.458f
C1897 comparator_0.ip.t18 avss 0.519f
C1898 comparator_0.ip.t10 avss 0.573f
C1899 comparator_0.ip.t14 avss 0.628f
C1900 comparator_0.ip.t16 avss 0.682f
C1901 comparator_0.ip.t3 avss 0.737f
C1902 comparator_0.ip.t4 avss 0.791f
C1903 comparator_0.ip.t13 avss 0.441f
C1904 comparator_0.ip.t12 avss 0.45f
C1905 comparator_0.ip.t8 avss 0.443f
C1906 comparator_0.ip.t0 avss 0.00501f
C1907 comparator_0.ip.t5 avss 0.453f
C1908 comparator_0.ip.t9 avss 0.437f
C1909 comparator_0.ip.n0 avss 0.047f
C1910 comparator_0.ip.t17 avss 0.752f
C1911 comparator_0.ip.t6 avss 0.489f
C1912 comparator_0.ip.t11 avss 0.451f
C1913 comparator_0.ip.t7 avss 0.449f
C1914 comparator_0.ip.n1 avss 0.0159f
C1915 comparator_0.ip.t2 avss 0.00378f
C1916 comparator_0.ip.n2 avss 0.0119f
C1917 comparator_0.ip.t1 avss 0.0038f
C1918 comparator_0.ip.n3 avss 0.0571f
C1919 comparator_0.trim_1.n3.n0 avss 0.372f
C1920 comparator_0.trim_1.n3.t7 avss 0.555f
C1921 comparator_0.trim_1.n3.t4 avss 0.436f
C1922 comparator_0.trim_1.n3.n1 avss 0.142f
C1923 comparator_0.trim_1.n3.t5 avss 0.436f
C1924 comparator_0.trim_1.n3.n2 avss 0.117f
C1925 comparator_0.trim_1.n3.t6 avss 0.483f
C1926 comparator_0.trim_1.n3.t1 avss 0.00667f
C1927 comparator_0.trim_1.n3.t0 avss 0.00574f
C1928 comparator_0.trim_1.n3.t3 avss 0.00574f
C1929 comparator_0.trim_1.n3.n3 avss 0.0366f
C1930 comparator_0.trim_1.n3.t2 avss 0.00947f
C1931 comparator_0.trim_1.n3.n4 avss 0.0705f
C1932 comparator_0.trim_1.n3.n5 avss 0.0604f
C1933 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t4 avss 0.71f
C1934 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t2 avss 0.00336f
C1935 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t3 avss 0.00336f
C1936 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n0 avss 0.00794f
C1937 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n1 avss 0.00477f
C1938 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n2 avss 0.181f
C1939 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t1 avss 0.00516f
C1940 dac_0.sky130_fd_sc_hd__inv_2_3.Y.t0 avss 0.00516f
C1941 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n3 avss 0.0132f
C1942 dac_0.sky130_fd_sc_hd__inv_2_3.Y.n4 avss 0.0228f
C1943 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t1 avss 0.00687f
C1944 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t2 avss 0.00687f
C1945 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n0 avss 0.0176f
C1946 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n1 avss 0.0303f
C1947 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t3 avss 0.00447f
C1948 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t4 avss 0.00447f
C1949 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n2 avss 0.0106f
C1950 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n3 avss 0.00634f
C1951 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n4 avss 0.23f
C1952 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n5 avss -0.374f
C1953 dac_1.sky130_fd_sc_hd__inv_2_1.Y.n6 avss 0.572f
C1954 dac_1.sky130_fd_sc_hd__inv_2_1.Y.t0 avss 0.436f
C1955 comparator_0.trim_0.n3.t2 avss 0.527f
C1956 comparator_0.trim_0.n3.t0 avss 0.555f
C1957 comparator_0.trim_0.n3.t3 avss 0.578f
C1958 comparator_0.trim_0.n3.t1 avss 0.57f
C1959 comparator_0.trim_0.n3.t6 avss 0.00667f
C1960 comparator_0.trim_0.n3.t7 avss 0.00947f
C1961 comparator_0.trim_0.n3.t4 avss 0.00574f
C1962 comparator_0.trim_0.n3.t5 avss 0.00574f
C1963 comparator_0.trim_0.n3.n0 avss 0.0366f
C1964 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t2 avss 0.00684f
C1965 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t3 avss 0.00684f
C1966 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n0 avss 0.0175f
C1967 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n1 avss 0.0301f
C1968 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t4 avss 0.00444f
C1969 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t1 avss 0.00444f
C1970 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n2 avss 0.0105f
C1971 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n3 avss 0.00631f
C1972 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n4 avss 0.28f
C1973 dac_1.sky130_fd_sc_hd__inv_2_8.Y.t0 avss 0.533f
C1974 dac_1.sky130_fd_sc_hd__inv_2_8.Y.n5 avss -0.778f
C1975 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t1 avss 0.842f
C1976 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t0 avss 0.819f
C1977 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t5 avss 0.00336f
C1978 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t3 avss 0.00336f
C1979 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n0 avss 0.00794f
C1980 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n1 avss 0.00477f
C1981 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n2 avss 0.181f
C1982 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t4 avss 0.00516f
C1983 dac_1.sky130_fd_sc_hd__inv_2_3.Y.t2 avss 0.00516f
C1984 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n3 avss 0.0132f
C1985 dac_1.sky130_fd_sc_hd__inv_2_3.Y.n4 avss 0.0228f
C1986 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t2 avss 0.763f
C1987 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t1 avss 0.00265f
C1988 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t3 avss 0.00265f
C1989 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n0 avss 0.00626f
C1990 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n1 avss 0.00376f
C1991 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n2 avss 0.091f
C1992 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t4 avss 0.00407f
C1993 dac_0.sky130_fd_sc_hd__inv_2_5.Y.t0 avss 0.00407f
C1994 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n3 avss 0.0104f
C1995 dac_0.sky130_fd_sc_hd__inv_2_5.Y.n4 avss 0.0179f
C1996 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t1 avss 0.00687f
C1997 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t2 avss 0.00687f
C1998 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n0 avss 0.0176f
C1999 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n1 avss 0.0303f
C2000 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t3 avss 0.00447f
C2001 dac_0.sky130_fd_sc_hd__inv_2_1.Y.t0 avss 0.00447f
C2002 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n2 avss 0.0106f
C2003 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n3 avss 0.00634f
C2004 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n4 avss 0.23f
C2005 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n5 avss -0.78f
C2006 dac_0.sky130_fd_sc_hd__inv_2_1.Y.n6 avss 0.957f
C2007 comparator_0.in.t11 avss 0.451f
C2008 comparator_0.in.t4 avss 0.512f
C2009 comparator_0.in.t8 avss 0.565f
C2010 comparator_0.in.t7 avss 0.619f
C2011 comparator_0.in.t10 avss 0.672f
C2012 comparator_0.in.t6 avss 0.726f
C2013 comparator_0.in.t15 avss 0.779f
C2014 comparator_0.in.t16 avss 0.435f
C2015 comparator_0.in.t18 avss 0.444f
C2016 comparator_0.in.t13 avss 0.436f
C2017 comparator_0.in.t2 avss 0.00531f
C2018 comparator_0.in.t9 avss 0.447f
C2019 comparator_0.in.t3 avss 0.43f
C2020 comparator_0.in.n0 avss 0.0486f
C2021 comparator_0.in.t12 avss 0.742f
C2022 comparator_0.in.t17 avss 0.482f
C2023 comparator_0.in.t5 avss 0.444f
C2024 comparator_0.in.t14 avss 0.443f
C2025 comparator_0.in.n1 avss 0.0168f
C2026 comparator_0.in.t1 avss 0.00375f
C2027 comparator_0.in.n2 avss 0.0554f
C2028 comparator_0.in.n3 avss 0.0133f
C2029 comparator_0.in.t0 avss 0.00375f
C2030 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t4 avss 0.533f
C2031 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n0 avss -0.376f
C2032 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t2 avss 0.00684f
C2033 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t0 avss 0.00684f
C2034 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n1 avss 0.0175f
C2035 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n2 avss 0.0301f
C2036 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t1 avss 0.00444f
C2037 dac_0.sky130_fd_sc_hd__inv_2_8.Y.t3 avss 0.00444f
C2038 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n3 avss 0.0105f
C2039 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n4 avss 0.00631f
C2040 dac_0.sky130_fd_sc_hd__inv_2_8.Y.n5 avss 0.28f
C2041 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t2 avss 0.00755f
C2042 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t3 avss 0.00755f
C2043 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n0 avss 0.0193f
C2044 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n1 avss 0.0333f
C2045 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t4 avss 0.00491f
C2046 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t1 avss 0.00491f
C2047 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n2 avss 0.0116f
C2048 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n3 avss 0.00697f
C2049 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n4 avss 0.287f
C2050 dac_1.sky130_fd_sc_hd__inv_2_0.Y.n5 avss 0.719f
C2051 dac_1.sky130_fd_sc_hd__inv_2_0.Y.t0 avss 0.552f
C2052 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t0 avss 0.349f
C2053 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t2 avss 0.459f
C2054 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t1 avss 0.36f
C2055 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n0 avss 0.211f
C2056 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t3 avss 0.00732f
C2057 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t5 avss 0.00732f
C2058 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n1 avss 0.0187f
C2059 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n2 avss 0.0323f
C2060 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t4 avss 0.00476f
C2061 dac_1.sky130_fd_sc_hd__inv_2_2.Y.t6 avss 0.00476f
C2062 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n3 avss 0.0113f
C2063 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n4 avss 0.00676f
C2064 dac_1.sky130_fd_sc_hd__inv_2_2.Y.n5 avss 0.288f
C2065 comparator_0.trim_1.n4.t4 avss 0.00627f
C2066 comparator_0.trim_1.n4.n0 avss 0.057f
C2067 comparator_0.trim_1.n4.t13 avss 0.437f
C2068 comparator_0.trim_1.n4.t9 avss 0.437f
C2069 comparator_0.trim_1.n4.t15 avss 0.437f
C2070 comparator_0.trim_1.n4.t14 avss 0.437f
C2071 comparator_0.trim_1.n4.t10 avss 0.437f
C2072 comparator_0.trim_1.n4.t11 avss 0.437f
C2073 comparator_0.trim_1.n4.t12 avss 0.557f
C2074 comparator_0.trim_1.n4.n1 avss 0.142f
C2075 comparator_0.trim_1.n4.n2 avss 0.138f
C2076 comparator_0.trim_1.n4.n3 avss 0.138f
C2077 comparator_0.trim_1.n4.n4 avss 0.138f
C2078 comparator_0.trim_1.n4.n5 avss 0.138f
C2079 comparator_0.trim_1.n4.n6 avss 0.129f
C2080 comparator_0.trim_1.n4.t8 avss 0.547f
C2081 comparator_0.trim_1.n4.n7 avss 0.0127f
C2082 comparator_0.trim_1.n4.t6 avss 0.00575f
C2083 comparator_0.trim_1.n4.t2 avss 0.00575f
C2084 comparator_0.trim_1.n4.n8 avss 0.0365f
C2085 comparator_0.trim_1.n4.t5 avss 0.00575f
C2086 comparator_0.trim_1.n4.t1 avss 0.00575f
C2087 comparator_0.trim_1.n4.n9 avss 0.0371f
C2088 comparator_0.trim_1.n4.t0 avss 0.00945f
C2089 comparator_0.trim_1.n4.n10 avss 0.0683f
C2090 comparator_0.trim_1.n4.n11 avss 0.0176f
C2091 comparator_0.trim_1.n4.t7 avss 0.00575f
C2092 comparator_0.trim_1.n4.t3 avss 0.00575f
C2093 comparator_0.trim_1.n4.n12 avss 0.0365f
C2094 comparator_0.trim_1.n4.n13 avss 0.0178f
C2095 comparator_0.trim_1.n4.n14 avss 0.0196f
C2096 sample.n0 avss 0.00529f
C2097 sample.n1 avss 0.00229f
C2098 sample.n2 avss 0.00766f
C2099 sample.n3 avss 0.00289f
C2100 sample.t42 avss 0.0194f
C2101 sample.t14 avss 0.0114f
C2102 sample.t15 avss 0.0194f
C2103 sample.t51 avss 0.0114f
C2104 sample.n4 avss 0.028f
C2105 sample.t57 avss 0.0194f
C2106 sample.t24 avss 0.0114f
C2107 sample.t11 avss 0.0194f
C2108 sample.t44 avss 0.0114f
C2109 sample.n5 avss 0.0262f
C2110 sample.n6 avss 0.0131f
C2111 sample.n7 avss 0.028f
C2112 sample.n8 avss 0.0128f
C2113 sample.n9 avss 0.0106f
C2114 sample.n10 avss 0.0106f
C2115 sample.n11 avss 0.0128f
C2116 sample.n12 avss 0.0325f
C2117 sample.n13 avss 0.0166f
C2118 sample.n14 avss 0.0022f
C2119 sample.n15 avss 0.00232f
C2120 sample.n16 avss 0.0055f
C2121 sample.n17 avss 0.0104f
C2122 sample.n18 avss 0.0297f
C2123 sample.n19 avss 0.0104f
C2124 sample.n20 avss 0.0055f
C2125 sample.n21 avss 0.00229f
C2126 sample.n22 avss 0.00766f
C2127 sample.n23 avss 0.00529f
C2128 sample.n24 avss 0.00289f
C2129 sample.t23 avss 0.0194f
C2130 sample.t61 avss 0.0114f
C2131 sample.t1 avss 0.0194f
C2132 sample.t31 avss 0.0114f
C2133 sample.n25 avss 0.028f
C2134 sample.t18 avss 0.0194f
C2135 sample.t56 avss 0.0114f
C2136 sample.t10 avss 0.0194f
C2137 sample.t41 avss 0.0114f
C2138 sample.n26 avss 0.0262f
C2139 sample.n27 avss 0.0131f
C2140 sample.n28 avss 0.028f
C2141 sample.n29 avss 0.0128f
C2142 sample.n30 avss 0.0106f
C2143 sample.n31 avss 0.0106f
C2144 sample.n32 avss 0.0128f
C2145 sample.n33 avss 0.0325f
C2146 sample.n34 avss 0.0166f
C2147 sample.n35 avss 0.0022f
C2148 sample.n36 avss 0.00232f
C2149 sample.n37 avss 0.0297f
C2150 sample.n38 avss 0.0104f
C2151 sample.n39 avss 0.0055f
C2152 sample.n40 avss 0.00229f
C2153 sample.n41 avss 0.00766f
C2154 sample.n42 avss 0.00529f
C2155 sample.n43 avss 0.00289f
C2156 sample.t19 avss 0.0194f
C2157 sample.t58 avss 0.0114f
C2158 sample.t39 avss 0.0194f
C2159 sample.t12 avss 0.0114f
C2160 sample.n44 avss 0.028f
C2161 sample.t2 avss 0.0194f
C2162 sample.t32 avss 0.0114f
C2163 sample.t36 avss 0.0194f
C2164 sample.t8 avss 0.0114f
C2165 sample.n45 avss 0.0262f
C2166 sample.n46 avss 0.0131f
C2167 sample.n47 avss 0.028f
C2168 sample.n48 avss 0.0128f
C2169 sample.n49 avss 0.0106f
C2170 sample.n50 avss 0.0106f
C2171 sample.n51 avss 0.0128f
C2172 sample.n52 avss 0.0325f
C2173 sample.n53 avss 0.0166f
C2174 sample.n54 avss 0.0022f
C2175 sample.n55 avss 0.00232f
C2176 sample.n56 avss 0.0297f
C2177 sample.n57 avss 0.0104f
C2178 sample.n58 avss 0.0055f
C2179 sample.n59 avss 0.00229f
C2180 sample.n60 avss 0.00766f
C2181 sample.n61 avss 0.00529f
C2182 sample.n62 avss 0.00289f
C2183 sample.t6 avss 0.0194f
C2184 sample.t34 avss 0.0114f
C2185 sample.t22 avss 0.0194f
C2186 sample.t60 avss 0.0114f
C2187 sample.n63 avss 0.028f
C2188 sample.t0 avss 0.0194f
C2189 sample.t30 avss 0.0114f
C2190 sample.t16 avss 0.0194f
C2191 sample.t53 avss 0.0114f
C2192 sample.n64 avss 0.0262f
C2193 sample.n65 avss 0.0131f
C2194 sample.n66 avss 0.028f
C2195 sample.n67 avss 0.0128f
C2196 sample.n68 avss 0.0106f
C2197 sample.n69 avss 0.0106f
C2198 sample.n70 avss 0.0128f
C2199 sample.n71 avss 0.0325f
C2200 sample.n72 avss 0.0166f
C2201 sample.n73 avss 0.0022f
C2202 sample.n74 avss 0.00232f
C2203 sample.n75 avss 0.0319f
C2204 sample.n76 avss 0.21f
C2205 sample.n77 avss 0.21f
C2206 sample.n78 avss 0.21f
C2207 sample.n79 avss 0.00232f
C2208 sample.n80 avss 0.00529f
C2209 sample.n81 avss 0.00289f
C2210 sample.n82 avss 0.00229f
C2211 sample.t37 avss 0.0114f
C2212 sample.t54 avss 0.0194f
C2213 sample.t33 avss 0.0114f
C2214 sample.t27 avss 0.0194f
C2215 sample.n83 avss 0.028f
C2216 sample.t48 avss 0.0114f
C2217 sample.t46 avss 0.0194f
C2218 sample.t20 avss 0.0114f
C2219 sample.t35 avss 0.0194f
C2220 sample.n84 avss 0.0262f
C2221 sample.n85 avss 0.0131f
C2222 sample.n86 avss 0.028f
C2223 sample.n87 avss 0.0128f
C2224 sample.n88 avss 0.0106f
C2225 sample.n89 avss 0.0106f
C2226 sample.n90 avss 0.0128f
C2227 sample.n91 avss 0.0325f
C2228 sample.n92 avss 0.0166f
C2229 sample.n93 avss 0.0022f
C2230 sample.n94 avss 0.00766f
C2231 sample.n95 avss 0.0055f
C2232 sample.n96 avss 0.0104f
C2233 sample.n97 avss 0.0297f
C2234 sample.n98 avss 0.00232f
C2235 sample.n99 avss 0.00529f
C2236 sample.n100 avss 0.00289f
C2237 sample.n101 avss 0.00229f
C2238 sample.t40 avss 0.0114f
C2239 sample.t29 avss 0.0194f
C2240 sample.t59 avss 0.0114f
C2241 sample.t52 avss 0.0194f
C2242 sample.n102 avss 0.028f
C2243 sample.t55 avss 0.0114f
C2244 sample.t25 avss 0.0194f
C2245 sample.t4 avss 0.0114f
C2246 sample.t45 avss 0.0194f
C2247 sample.n103 avss 0.0262f
C2248 sample.n104 avss 0.0131f
C2249 sample.n105 avss 0.028f
C2250 sample.n106 avss 0.0128f
C2251 sample.n107 avss 0.0106f
C2252 sample.n108 avss 0.0106f
C2253 sample.n109 avss 0.0128f
C2254 sample.n110 avss 0.0325f
C2255 sample.n111 avss 0.0166f
C2256 sample.n112 avss 0.0022f
C2257 sample.n113 avss 0.00766f
C2258 sample.n114 avss 0.0055f
C2259 sample.n115 avss 0.0104f
C2260 sample.n116 avss 0.0297f
C2261 sample.n117 avss 0.00232f
C2262 sample.n118 avss 0.00529f
C2263 sample.n119 avss 0.00289f
C2264 sample.n120 avss 0.00229f
C2265 sample.t3 avss 0.0114f
C2266 sample.t49 avss 0.0194f
C2267 sample.t13 avss 0.0114f
C2268 sample.t7 avss 0.0194f
C2269 sample.n121 avss 0.028f
C2270 sample.t26 avss 0.0114f
C2271 sample.t28 avss 0.0194f
C2272 sample.t21 avss 0.0114f
C2273 sample.t5 avss 0.0194f
C2274 sample.n122 avss 0.0262f
C2275 sample.n123 avss 0.0131f
C2276 sample.n124 avss 0.028f
C2277 sample.n125 avss 0.0128f
C2278 sample.n126 avss 0.0106f
C2279 sample.n127 avss 0.0106f
C2280 sample.n128 avss 0.0128f
C2281 sample.n129 avss 0.0325f
C2282 sample.n130 avss 0.0166f
C2283 sample.n131 avss 0.0022f
C2284 sample.n132 avss 0.00766f
C2285 sample.n133 avss 0.0055f
C2286 sample.n134 avss 0.0104f
C2287 sample.n135 avss 0.0297f
C2288 sample.n136 avss 0.00898f
C2289 sample.n137 avss 0.0055f
C2290 sample.n138 avss 0.0022f
C2291 sample.n139 avss 0.00529f
C2292 sample.n140 avss 0.00289f
C2293 sample.t62 avss 0.0114f
C2294 sample.t9 avss 0.0194f
C2295 sample.t50 avss 0.0114f
C2296 sample.t43 avss 0.0194f
C2297 sample.n141 avss 0.028f
C2298 sample.t47 avss 0.0114f
C2299 sample.t17 avss 0.0194f
C2300 sample.t63 avss 0.0114f
C2301 sample.t38 avss 0.0194f
C2302 sample.n142 avss 0.0262f
C2303 sample.n143 avss 0.0131f
C2304 sample.n144 avss 0.028f
C2305 sample.n145 avss 0.0128f
C2306 sample.n146 avss 0.0106f
C2307 sample.n147 avss 0.00766f
C2308 sample.n148 avss 0.0106f
C2309 sample.n149 avss 0.0128f
C2310 sample.n150 avss 0.0325f
C2311 sample.n151 avss 0.0166f
C2312 sample.n152 avss 0.00229f
C2313 sample.n153 avss 0.00377f
C2314 sample.n154 avss 0.0306f
C2315 sample.n155 avss 0.998f
C2316 dac_1.out.t83 avss 1.95f
C2317 dac_1.out.t89 avss 1.32f
C2318 dac_1.out.t85 avss 0.819f
C2319 dac_1.out.t84 avss 0.478f
C2320 dac_1.out.t86 avss 0.643f
C2321 dac_1.out.t80 avss 1.63f
C2322 dac_1.out.t88 avss 0.965f
C2323 dac_1.out.t81 avss 1.13f
C2324 dac_1.out.t82 avss 1.45f
C2325 dac_1.out.n0 avss 0.0369f
C2326 dac_1.out.n1 avss 0.0359f
C2327 dac_1.out.n2 avss 0.0393f
C2328 dac_1.out.n3 avss 0.0369f
C2329 dac_1.out.n4 avss 0.0359f
C2330 dac_1.out.n5 avss 0.0393f
C2331 dac_1.out.n6 avss 0.0369f
C2332 dac_1.out.n7 avss 0.0359f
C2333 dac_1.out.n8 avss 0.0393f
C2334 dac_1.out.n9 avss 0.031f
C2335 dac_1.out.n10 avss 0.0359f
C2336 dac_1.out.n11 avss 0.0369f
C2337 dac_1.out.n12 avss 0.41f
C2338 dac_1.out.n13 avss 0.427f
C2339 dac_1.out.n14 avss 0.205f
C2340 dac_1.out.n15 avss 0.236f
C2341 dac_1.out.n16 avss 0.255f
C2342 dac_1.out.n17 avss 0.306f
C2343 dac_1.out.n18 avss 0.337f
C2344 dac_1.out.n19 avss 0.345f
C2345 dac_1.out.t87 avss 0.0163f
C2346 dac_1.out.n20 avss 0.0858f
C2347 dac_1.out.n21 avss 0.378f
C2348 dac_1.out.n22 avss 0.0676f
C2349 dac_1.out.t18 avss 0.00496f
C2350 dac_1.out.t13 avss 0.00496f
C2351 dac_1.out.n23 avss 0.0351f
C2352 dac_1.out.t14 avss 0.00496f
C2353 dac_1.out.t19 avss 0.00496f
C2354 dac_1.out.n24 avss 0.0352f
C2355 dac_1.out.t15 avss 0.00496f
C2356 dac_1.out.t10 avss 0.00496f
C2357 dac_1.out.n25 avss 0.0348f
C2358 dac_1.out.t53 avss 0.00496f
C2359 dac_1.out.t58 avss 0.00496f
C2360 dac_1.out.n26 avss 0.0409f
C2361 dac_1.out.t17 avss 0.00496f
C2362 dac_1.out.t12 avss 0.00496f
C2363 dac_1.out.n27 avss 0.0349f
C2364 dac_1.out.t55 avss 0.00496f
C2365 dac_1.out.t52 avss 0.00496f
C2366 dac_1.out.n28 avss 0.0386f
C2367 dac_1.out.n29 avss 0.03f
C2368 dac_1.out.t16 avss 0.00496f
C2369 dac_1.out.t11 avss 0.00496f
C2370 dac_1.out.n30 avss 0.0346f
C2371 dac_1.out.t54 avss 0.00496f
C2372 dac_1.out.t59 avss 0.00496f
C2373 dac_1.out.n31 avss 0.0416f
C2374 dac_1.out.n32 avss 0.036f
C2375 dac_1.out.t51 avss 0.00496f
C2376 dac_1.out.t57 avss 0.00496f
C2377 dac_1.out.n33 avss 0.043f
C2378 dac_1.out.t56 avss 0.00496f
C2379 dac_1.out.t50 avss 0.00496f
C2380 dac_1.out.n34 avss 0.0428f
C2381 dac_1.out.t41 avss 0.00496f
C2382 dac_1.out.t47 avss 0.00496f
C2383 dac_1.out.n35 avss 0.0351f
C2384 dac_1.out.t45 avss 0.00496f
C2385 dac_1.out.t49 avss 0.00496f
C2386 dac_1.out.n36 avss 0.0352f
C2387 dac_1.out.t46 avss 0.00496f
C2388 dac_1.out.t42 avss 0.00496f
C2389 dac_1.out.n37 avss 0.0348f
C2390 dac_1.out.t63 avss 0.00496f
C2391 dac_1.out.t60 avss 0.00496f
C2392 dac_1.out.n38 avss 0.0409f
C2393 dac_1.out.t48 avss 0.00496f
C2394 dac_1.out.t44 avss 0.00496f
C2395 dac_1.out.n39 avss 0.0349f
C2396 dac_1.out.t66 avss 0.00496f
C2397 dac_1.out.t61 avss 0.00496f
C2398 dac_1.out.n40 avss 0.0386f
C2399 dac_1.out.n41 avss 0.03f
C2400 dac_1.out.t40 avss 0.00496f
C2401 dac_1.out.t43 avss 0.00496f
C2402 dac_1.out.n42 avss 0.0346f
C2403 dac_1.out.t68 avss 0.00496f
C2404 dac_1.out.t64 avss 0.00496f
C2405 dac_1.out.n43 avss 0.0416f
C2406 dac_1.out.n44 avss 0.036f
C2407 dac_1.out.t62 avss 0.00496f
C2408 dac_1.out.t67 avss 0.00496f
C2409 dac_1.out.n45 avss 0.043f
C2410 dac_1.out.t69 avss 0.00496f
C2411 dac_1.out.t65 avss 0.00496f
C2412 dac_1.out.n46 avss 0.0428f
C2413 dac_1.out.t24 avss 0.00496f
C2414 dac_1.out.t22 avss 0.00496f
C2415 dac_1.out.n47 avss 0.0351f
C2416 dac_1.out.t28 avss 0.00496f
C2417 dac_1.out.t25 avss 0.00496f
C2418 dac_1.out.n48 avss 0.0352f
C2419 dac_1.out.t29 avss 0.00496f
C2420 dac_1.out.t26 avss 0.00496f
C2421 dac_1.out.n49 avss 0.0348f
C2422 dac_1.out.t38 avss 0.00496f
C2423 dac_1.out.t35 avss 0.00496f
C2424 dac_1.out.n50 avss 0.0409f
C2425 dac_1.out.t23 avss 0.00496f
C2426 dac_1.out.t21 avss 0.00496f
C2427 dac_1.out.n51 avss 0.0349f
C2428 dac_1.out.t31 avss 0.00496f
C2429 dac_1.out.t39 avss 0.00496f
C2430 dac_1.out.n52 avss 0.0386f
C2431 dac_1.out.n53 avss 0.03f
C2432 dac_1.out.t20 avss 0.00496f
C2433 dac_1.out.t27 avss 0.00496f
C2434 dac_1.out.n54 avss 0.0346f
C2435 dac_1.out.t30 avss 0.00496f
C2436 dac_1.out.t36 avss 0.00496f
C2437 dac_1.out.n55 avss 0.0416f
C2438 dac_1.out.n56 avss 0.036f
C2439 dac_1.out.t37 avss 0.00496f
C2440 dac_1.out.t34 avss 0.00496f
C2441 dac_1.out.n57 avss 0.043f
C2442 dac_1.out.t32 avss 0.00496f
C2443 dac_1.out.t33 avss 0.00496f
C2444 dac_1.out.n58 avss 0.0428f
C2445 dac_1.out.n59 avss 0.17f
C2446 dac_1.out.n60 avss 0.129f
C2447 dac_1.out.n61 avss 0.0734f
C2448 dac_1.out.n62 avss 0.0441f
C2449 dac_1.out.n63 avss 0.0019f
C2450 dac_1.out.t72 avss 0.00496f
C2451 dac_1.out.t79 avss 0.00496f
C2452 dac_1.out.n64 avss 0.0222f
C2453 dac_1.out.n65 avss 0.011f
C2454 dac_1.out.n66 avss 0.00177f
C2455 dac_1.out.n67 avss 0.00658f
C2456 dac_1.out.t2 avss 0.00496f
C2457 dac_1.out.t7 avss 0.00496f
C2458 dac_1.out.n68 avss 0.0428f
C2459 dac_1.out.t75 avss 0.00496f
C2460 dac_1.out.t76 avss 0.00496f
C2461 dac_1.out.n69 avss 0.0352f
C2462 dac_1.out.t3 avss 0.00496f
C2463 dac_1.out.t4 avss 0.00496f
C2464 dac_1.out.n70 avss 0.043f
C2465 dac_1.out.t73 avss 0.00496f
C2466 dac_1.out.t77 avss 0.00496f
C2467 dac_1.out.n71 avss 0.0348f
C2468 dac_1.out.t0 avss 0.00496f
C2469 dac_1.out.t5 avss 0.00496f
C2470 dac_1.out.n72 avss 0.0409f
C2471 dac_1.out.t70 avss 0.00496f
C2472 dac_1.out.t78 avss 0.00496f
C2473 dac_1.out.n73 avss 0.0346f
C2474 dac_1.out.t74 avss 0.00496f
C2475 dac_1.out.t71 avss 0.00496f
C2476 dac_1.out.n74 avss 0.0349f
C2477 dac_1.out.t1 avss 0.00496f
C2478 dac_1.out.t9 avss 0.00496f
C2479 dac_1.out.n75 avss 0.0386f
C2480 dac_1.out.n76 avss 0.03f
C2481 dac_1.out.t8 avss 0.00496f
C2482 dac_1.out.t6 avss 0.00496f
C2483 dac_1.out.n77 avss 0.0416f
C2484 dac_1.out.n78 avss 0.036f
C2485 vinn.t78 avss 0.0219f
C2486 vinn.t9 avss 0.0241f
C2487 vinn.t75 avss 0.0182f
C2488 vinn.t71 avss 0.0182f
C2489 vinn.n0 avss 0.128f
C2490 vinn.t2 avss 0.0182f
C2491 vinn.t5 avss 0.0182f
C2492 vinn.n1 avss 0.128f
C2493 vinn.t74 avss 0.0182f
C2494 vinn.t77 avss 0.0182f
C2495 vinn.n2 avss 0.128f
C2496 vinn.t1 avss 0.0182f
C2497 vinn.t4 avss 0.0182f
C2498 vinn.n3 avss 0.128f
C2499 vinn.t73 avss 0.0182f
C2500 vinn.t70 avss 0.0182f
C2501 vinn.n4 avss 0.128f
C2502 vinn.t8 avss 0.0182f
C2503 vinn.t0 avss 0.0182f
C2504 vinn.n5 avss 0.128f
C2505 vinn.t76 avss 0.0182f
C2506 vinn.t72 avss 0.0182f
C2507 vinn.n6 avss 0.128f
C2508 vinn.t3 avss 0.0182f
C2509 vinn.t7 avss 0.0182f
C2510 vinn.n7 avss 0.128f
C2511 vinn.t79 avss 0.0219f
C2512 vinn.t6 avss 0.0241f
C2513 vinn.n8 avss 0.365f
C2514 vinn.n9 avss 0.107f
C2515 vinn.n10 avss 0.107f
C2516 vinn.n11 avss 0.107f
C2517 vinn.n12 avss 0.107f
C2518 vinn.n13 avss 0.383f
C2519 vinn.t19 avss 0.0219f
C2520 vinn.t59 avss 0.0241f
C2521 vinn.t18 avss 0.0182f
C2522 vinn.t10 avss 0.0182f
C2523 vinn.n14 avss 0.128f
C2524 vinn.t56 avss 0.0182f
C2525 vinn.t52 avss 0.0182f
C2526 vinn.n15 avss 0.128f
C2527 vinn.t17 avss 0.0182f
C2528 vinn.t16 avss 0.0182f
C2529 vinn.n16 avss 0.128f
C2530 vinn.t55 avss 0.0182f
C2531 vinn.t51 avss 0.0182f
C2532 vinn.n17 avss 0.128f
C2533 vinn.t12 avss 0.0182f
C2534 vinn.t15 avss 0.0182f
C2535 vinn.n18 avss 0.128f
C2536 vinn.t54 avss 0.0182f
C2537 vinn.t50 avss 0.0182f
C2538 vinn.n19 avss 0.128f
C2539 vinn.t13 avss 0.0182f
C2540 vinn.t14 avss 0.0182f
C2541 vinn.n20 avss 0.128f
C2542 vinn.t57 avss 0.0182f
C2543 vinn.t58 avss 0.0182f
C2544 vinn.n21 avss 0.128f
C2545 vinn.t11 avss 0.0219f
C2546 vinn.t53 avss 0.0241f
C2547 vinn.n22 avss 0.365f
C2548 vinn.n23 avss 0.107f
C2549 vinn.n24 avss 0.107f
C2550 vinn.n25 avss 0.107f
C2551 vinn.n26 avss 0.107f
C2552 vinn.n27 avss 0.381f
C2553 vinn.n28 avss 0.0808f
C2554 vinn.t47 avss 0.0219f
C2555 vinn.t60 avss 0.0241f
C2556 vinn.t46 avss 0.0182f
C2557 vinn.t43 avss 0.0182f
C2558 vinn.n29 avss 0.128f
C2559 vinn.t63 avss 0.0182f
C2560 vinn.t67 avss 0.0182f
C2561 vinn.n30 avss 0.128f
C2562 vinn.t45 avss 0.0182f
C2563 vinn.t49 avss 0.0182f
C2564 vinn.n31 avss 0.128f
C2565 vinn.t65 avss 0.0182f
C2566 vinn.t69 avss 0.0182f
C2567 vinn.n32 avss 0.128f
C2568 vinn.t48 avss 0.0182f
C2569 vinn.t41 avss 0.0182f
C2570 vinn.n33 avss 0.128f
C2571 vinn.t68 avss 0.0182f
C2572 vinn.t62 avss 0.0182f
C2573 vinn.n34 avss 0.128f
C2574 vinn.t42 avss 0.0182f
C2575 vinn.t40 avss 0.0182f
C2576 vinn.n35 avss 0.128f
C2577 vinn.t66 avss 0.0182f
C2578 vinn.t61 avss 0.0182f
C2579 vinn.n36 avss 0.128f
C2580 vinn.t44 avss 0.0219f
C2581 vinn.t64 avss 0.0241f
C2582 vinn.n37 avss 0.365f
C2583 vinn.n38 avss 0.107f
C2584 vinn.n39 avss 0.107f
C2585 vinn.n40 avss 0.107f
C2586 vinn.n41 avss 0.107f
C2587 vinn.n42 avss 0.381f
C2588 vinn.n43 avss 0.0818f
C2589 vinn.t21 avss 0.0219f
C2590 vinn.t39 avss 0.0241f
C2591 vinn.t28 avss 0.0182f
C2592 vinn.t23 avss 0.0182f
C2593 vinn.n44 avss 0.128f
C2594 vinn.t36 avss 0.0182f
C2595 vinn.t31 avss 0.0182f
C2596 vinn.n45 avss 0.128f
C2597 vinn.t27 avss 0.0182f
C2598 vinn.t20 avss 0.0182f
C2599 vinn.n46 avss 0.128f
C2600 vinn.t35 avss 0.0182f
C2601 vinn.t30 avss 0.0182f
C2602 vinn.n47 avss 0.128f
C2603 vinn.t26 avss 0.0182f
C2604 vinn.t25 avss 0.0182f
C2605 vinn.n48 avss 0.128f
C2606 vinn.t34 avss 0.0182f
C2607 vinn.t38 avss 0.0182f
C2608 vinn.n49 avss 0.128f
C2609 vinn.t22 avss 0.0182f
C2610 vinn.t29 avss 0.0182f
C2611 vinn.n50 avss 0.128f
C2612 vinn.t33 avss 0.0182f
C2613 vinn.t37 avss 0.0182f
C2614 vinn.n51 avss 0.128f
C2615 vinn.t24 avss 0.0219f
C2616 vinn.t32 avss 0.0241f
C2617 vinn.n52 avss 0.365f
C2618 vinn.n53 avss 0.107f
C2619 vinn.n54 avss 0.107f
C2620 vinn.n55 avss 0.107f
C2621 vinn.n56 avss 0.107f
C2622 vinn.n57 avss 0.381f
C2623 vinn.n58 avss 0.303f
C2624 vinn.n59 avss 0.559f
C2625 vinn.n60 avss 0.507f
C2626 vinn.n61 avss 0.394f
C2627 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n0 avss 0.719f
C2628 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t3 avss 0.552f
C2629 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t0 avss 0.00755f
C2630 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t2 avss 0.00755f
C2631 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n1 avss 0.0193f
C2632 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n2 avss 0.0333f
C2633 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t1 avss 0.00491f
C2634 dac_0.sky130_fd_sc_hd__inv_2_0.Y.t4 avss 0.00491f
C2635 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n3 avss 0.0116f
C2636 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n4 avss 0.00697f
C2637 dac_0.sky130_fd_sc_hd__inv_2_0.Y.n5 avss 0.287f
C2638 comparator_0.trim_0.n4.t4 avss 0.429f
C2639 comparator_0.trim_0.n4.t1 avss 0.429f
C2640 comparator_0.trim_0.n4.t6 avss 0.429f
C2641 comparator_0.trim_0.n4.t2 avss 0.429f
C2642 comparator_0.trim_0.n4.t0 avss 0.429f
C2643 comparator_0.trim_0.n4.t5 avss 0.429f
C2644 comparator_0.trim_0.n4.t3 avss 0.545f
C2645 comparator_0.trim_0.n4.n0 avss 0.139f
C2646 comparator_0.trim_0.n4.n1 avss 0.135f
C2647 comparator_0.trim_0.n4.n2 avss 0.135f
C2648 comparator_0.trim_0.n4.n3 avss 0.135f
C2649 comparator_0.trim_0.n4.n4 avss 0.135f
C2650 comparator_0.trim_0.n4.n5 avss 0.126f
C2651 comparator_0.trim_0.n4.t7 avss 0.535f
C2652 comparator_0.trim_0.n4.n6 avss 0.0116f
C2653 comparator_0.trim_0.n4.t8 avss 0.00574f
C2654 comparator_0.trim_0.n4.n7 avss 0.00609f
C2655 comparator_0.trim_0.n4.t12 avss 0.00563f
C2656 comparator_0.trim_0.n4.t9 avss 0.00563f
C2657 comparator_0.trim_0.n4.n8 avss 0.0358f
C2658 comparator_0.trim_0.n4.t11 avss 0.00563f
C2659 comparator_0.trim_0.n4.t15 avss 0.00563f
C2660 comparator_0.trim_0.n4.n9 avss 0.0358f
C2661 comparator_0.trim_0.n4.t13 avss 0.00925f
C2662 comparator_0.trim_0.n4.t10 avss 0.00563f
C2663 comparator_0.trim_0.n4.t14 avss 0.00563f
C2664 comparator_0.trim_0.n4.n10 avss 0.0363f
C2665 comparator_0.trim_0.n4.n11 avss 0.0669f
C2666 comparator_0.trim_0.n4.n12 avss 0.0172f
C2667 comparator_0.trim_0.n4.n13 avss 0.0174f
C2668 comparator_0.trim_0.n4.n14 avss 0.017f
C2669 avdd.t236 avss -0.00352f
C2670 avdd.n0 avss -0.00442f
C2671 avdd.n1 avss -0.00211f
C2672 avdd.n2 avss -7.31e-19
C2673 avdd.n3 avss -7.31e-19
C2674 avdd.n4 avss -7.31e-19
C2675 avdd.n5 avss -7.31e-19
C2676 avdd.n6 avss -7.31e-19
C2677 avdd.n7 avss -7.31e-19
C2678 avdd.n8 avss -7.31e-19
C2679 avdd.n9 avss -7.31e-19
C2680 avdd.n10 avss -0.00234f
C2681 avdd.t10 avss -0.00352f
C2682 avdd.n11 avss -0.00424f
C2683 avdd.n12 avss -0.00208f
C2684 avdd.n13 avss -0.00283f
C2685 avdd.n14 avss -0.00168f
C2686 avdd.t239 avss -0.00352f
C2687 avdd.n15 avss -0.00434f
C2688 avdd.t72 avss -0.00352f
C2689 avdd.n16 avss -0.00401f
C2690 avdd.n17 avss -0.00211f
C2691 avdd.n18 avss -0.00283f
C2692 avdd.n19 avss -0.00168f
C2693 avdd.t73 avss -0.00352f
C2694 avdd.n20 avss -0.00433f
C2695 avdd.t77 avss -0.00352f
C2696 avdd.n21 avss -0.004f
C2697 avdd.n22 avss -0.00209f
C2698 avdd.n23 avss -0.00283f
C2699 avdd.n24 avss -0.00168f
C2700 avdd.t78 avss -0.00352f
C2701 avdd.n25 avss -0.00434f
C2702 avdd.t151 avss -0.00352f
C2703 avdd.n26 avss -0.00401f
C2704 avdd.n27 avss -0.00211f
C2705 avdd.n28 avss -0.00283f
C2706 avdd.n29 avss -0.00168f
C2707 avdd.t152 avss -0.00352f
C2708 avdd.n30 avss -0.00434f
C2709 avdd.t268 avss -0.00352f
C2710 avdd.n31 avss -0.00401f
C2711 avdd.n32 avss -0.00211f
C2712 avdd.n33 avss -0.00283f
C2713 avdd.n34 avss -0.00168f
C2714 avdd.t3 avss -0.00352f
C2715 avdd.n35 avss -0.00434f
C2716 avdd.t123 avss -0.00352f
C2717 avdd.n36 avss -0.00401f
C2718 avdd.n37 avss -0.00213f
C2719 avdd.n38 avss -0.00283f
C2720 avdd.n39 avss -0.00168f
C2721 avdd.t124 avss -0.00352f
C2722 avdd.n40 avss -0.00434f
C2723 avdd.t112 avss -0.00352f
C2724 avdd.n41 avss -0.00401f
C2725 avdd.n42 avss -0.00211f
C2726 avdd.n43 avss -0.00283f
C2727 avdd.n44 avss -0.00168f
C2728 avdd.t27 avss -0.00352f
C2729 avdd.n45 avss -0.00433f
C2730 avdd.t110 avss -0.00352f
C2731 avdd.n46 avss -0.004f
C2732 avdd.n47 avss -0.00209f
C2733 avdd.n48 avss -0.00283f
C2734 avdd.n49 avss -0.00168f
C2735 avdd.t111 avss -0.00352f
C2736 avdd.n50 avss -0.00434f
C2737 avdd.t217 avss -0.00352f
C2738 avdd.n51 avss -0.00401f
C2739 avdd.n52 avss -7.31e-19
C2740 avdd.n53 avss -0.00283f
C2741 avdd.n54 avss -0.00168f
C2742 avdd.n55 avss -0.00111f
C2743 avdd.n56 avss -9.91e-19
C2744 avdd.n57 avss -0.00256f
C2745 avdd.n58 avss -8.47e-19
C2746 avdd.n59 avss -3.28e-19
C2747 avdd.n60 avss -3.28e-19
C2748 avdd.n61 avss -8.26e-19
C2749 avdd.n62 avss 0.0348f
C2750 avdd.n63 avss 0.00357f
C2751 avdd.n64 avss -8.47e-19
C2752 avdd.n65 avss -3.39e-19
C2753 avdd.n66 avss -8.47e-19
C2754 avdd.n67 avss 0.0344f
C2755 avdd.n68 avss 0.00466f
C2756 avdd.n69 avss -3.39e-19
C2757 avdd.n70 avss -6.67e-19
C2758 avdd.n71 avss -5.61e-19
C2759 avdd.n72 avss -3.39e-19
C2760 avdd.n73 avss -6.35e-19
C2761 avdd.n74 avss -0.00139f
C2762 avdd.n75 avss -6.88e-19
C2763 avdd.n76 avss -3.07e-19
C2764 avdd.n77 avss -1.8e-19
C2765 avdd.n78 avss 0.00821f
C2766 avdd.n79 avss -2.75e-19
C2767 avdd.n80 avss 0.0442f
C2768 avdd.n81 avss 0.0179f
C2769 avdd.n82 avss 0.0181f
C2770 avdd.n83 avss -2.75e-19
C2771 avdd.n84 avss -3.39e-19
C2772 avdd.n85 avss -3.6e-19
C2773 avdd.n86 avss -2.01e-19
C2774 avdd.n87 avss -0.0866f
C2775 avdd.n88 avss -0.00336f
C2776 avdd.n89 avss 0.00725f
C2777 avdd.n90 avss 0.0318f
C2778 avdd.n91 avss -0.00158f
C2779 avdd.n92 avss -8.47e-19
C2780 avdd.n93 avss -3.39e-19
C2781 avdd.n94 avss -4.23e-19
C2782 avdd.n95 avss -0.00173f
C2783 avdd.n96 avss 0.0098f
C2784 avdd.n97 avss 0.0298f
C2785 avdd.n98 avss -2.22e-19
C2786 avdd.n99 avss 0.0188f
C2787 avdd.n100 avss -2.33e-19
C2788 avdd.n101 avss -1.59e-19
C2789 avdd.n102 avss -2.22e-19
C2790 avdd.n103 avss 0.00821f
C2791 avdd.n104 avss -2.75e-19
C2792 avdd.n105 avss 0.0112f
C2793 avdd.n106 avss 0.0148f
C2794 avdd.n107 avss 0.0182f
C2795 avdd.n108 avss -1.8e-19
C2796 avdd.n109 avss -2.54e-19
C2797 avdd.n110 avss -2.54e-19
C2798 avdd.n111 avss -1.8e-19
C2799 avdd.n112 avss -1.16e-19
C2800 avdd.n113 avss -2.33e-19
C2801 avdd.n114 avss -0.00126f
C2802 avdd.n115 avss -0.00109f
C2803 avdd.n116 avss -0.00108f
C2804 avdd.n118 avss -3.07e-19
C2805 avdd.n119 avss 0.0374f
C2806 avdd.n120 avss 0.00358f
C2807 avdd.n121 avss 0.0192f
C2808 avdd.n122 avss -1.59e-19
C2809 avdd.n123 avss -1.8e-19
C2810 avdd.n124 avss 0.00875f
C2811 avdd.n125 avss 0.0111f
C2812 avdd.n126 avss 0.0154f
C2813 avdd.n127 avss 0.0183f
C2814 avdd.n128 avss -1.8e-19
C2815 avdd.n129 avss -2.22e-19
C2816 avdd.n130 avss -2.22e-19
C2817 avdd.n131 avss -1.8e-19
C2818 avdd.n132 avss -2.01e-19
C2819 avdd.n133 avss -9.61e-19
C2820 avdd.n134 avss -5.77e-19
C2821 avdd.n135 avss 0.0398f
C2822 avdd.n136 avss -3.07e-19
C2823 avdd.n137 avss -1.8e-19
C2824 avdd.n138 avss 0.0168f
C2825 avdd.n139 avss 0.0189f
C2826 avdd.n140 avss 0.0111f
C2827 avdd.n141 avss 0.00875f
C2828 avdd.n142 avss 0.0167f
C2829 avdd.n143 avss 0.0181f
C2830 avdd.n144 avss -3.6e-19
C2831 avdd.n145 avss -2.01e-19
C2832 avdd.n146 avss -3.07e-19
C2833 avdd.n147 avss -6.46e-19
C2834 avdd.n148 avss -0.00137f
C2835 avdd.n149 avss -0.0013f
C2836 avdd.n150 avss -5.19e-19
C2837 avdd.n151 avss 0.0386f
C2838 avdd.n152 avss 0.00873f
C2839 avdd.n153 avss 0.0111f
C2840 avdd.n154 avss 0.0148f
C2841 avdd.n155 avss 0.019f
C2842 avdd.n156 avss -1.8e-19
C2843 avdd.n157 avss 0.0184f
C2844 avdd.n158 avss -2.44e-19
C2845 avdd.n159 avss -2.33e-19
C2846 avdd.n160 avss 0.0022f
C2847 avdd.n161 avss -1.48e-19
C2848 avdd.n162 avss -1.27e-19
C2849 avdd.n163 avss -2.44e-19
C2850 avdd.n164 avss -8.15e-19
C2851 avdd.n165 avss -0.0014f
C2852 avdd.n166 avss -8.47e-19
C2853 avdd.n167 avss -3.39e-19
C2854 avdd.n168 avss -3.49e-19
C2855 avdd.n169 avss -1.38e-19
C2856 avdd.n170 avss -1.8e-19
C2857 avdd.n171 avss 0.00873f
C2858 avdd.n172 avss 0.0111f
C2859 avdd.n173 avss 0.0154f
C2860 avdd.n174 avss 0.0191f
C2861 avdd.n175 avss -1.8e-19
C2862 avdd.n176 avss 0.0184f
C2863 avdd.n177 avss -1.38e-19
C2864 avdd.n178 avss -1.8e-19
C2865 avdd.n179 avss -2.44e-19
C2866 avdd.n180 avss 0.0411f
C2867 avdd.n181 avss -1.8e-19
C2868 avdd.n182 avss -1.8e-19
C2869 avdd.n183 avss -2.96e-19
C2870 avdd.n184 avss -0.00139f
C2871 avdd.n185 avss -0.00106f
C2872 avdd.n186 avss -0.00357f
C2873 avdd.n187 avss 0.0382f
C2874 avdd.n188 avss -8.47e-19
C2875 avdd.n189 avss -3.28e-19
C2876 avdd.n190 avss -3.28e-19
C2877 avdd.n191 avss -8.26e-19
C2878 avdd.n192 avss 0.0348f
C2879 avdd.n193 avss 0.00357f
C2880 avdd.n194 avss -8.47e-19
C2881 avdd.n195 avss -3.39e-19
C2882 avdd.n196 avss -8.47e-19
C2883 avdd.n197 avss 0.0344f
C2884 avdd.n198 avss 0.00466f
C2885 avdd.n199 avss -3.39e-19
C2886 avdd.n200 avss -6.67e-19
C2887 avdd.n201 avss -5.61e-19
C2888 avdd.n202 avss -3.39e-19
C2889 avdd.n203 avss -6.35e-19
C2890 avdd.n204 avss -0.00139f
C2891 avdd.n205 avss -6.88e-19
C2892 avdd.n206 avss -3.07e-19
C2893 avdd.n207 avss -1.8e-19
C2894 avdd.n208 avss 0.00821f
C2895 avdd.n209 avss -2.75e-19
C2896 avdd.n210 avss 0.0442f
C2897 avdd.n211 avss 0.0179f
C2898 avdd.n212 avss 0.0181f
C2899 avdd.n213 avss -2.75e-19
C2900 avdd.n214 avss -3.39e-19
C2901 avdd.n215 avss -3.6e-19
C2902 avdd.n216 avss -2.01e-19
C2903 avdd.n217 avss -0.0866f
C2904 avdd.n218 avss -0.00336f
C2905 avdd.n219 avss 0.00725f
C2906 avdd.n220 avss 0.0318f
C2907 avdd.n221 avss -0.00158f
C2908 avdd.n222 avss -8.47e-19
C2909 avdd.n223 avss -3.39e-19
C2910 avdd.n224 avss -4.23e-19
C2911 avdd.n225 avss -0.00173f
C2912 avdd.n226 avss 0.0098f
C2913 avdd.n227 avss 0.0298f
C2914 avdd.n228 avss -2.22e-19
C2915 avdd.n229 avss 0.0188f
C2916 avdd.n230 avss -2.33e-19
C2917 avdd.n231 avss -1.59e-19
C2918 avdd.n232 avss -2.22e-19
C2919 avdd.n233 avss 0.00821f
C2920 avdd.n234 avss -2.75e-19
C2921 avdd.n235 avss 0.0112f
C2922 avdd.n236 avss 0.0148f
C2923 avdd.n237 avss 0.0182f
C2924 avdd.n238 avss -1.8e-19
C2925 avdd.n239 avss -2.54e-19
C2926 avdd.n240 avss -2.54e-19
C2927 avdd.n241 avss -1.8e-19
C2928 avdd.n242 avss -1.16e-19
C2929 avdd.n243 avss -2.33e-19
C2930 avdd.n244 avss -0.00126f
C2931 avdd.n245 avss -0.00109f
C2932 avdd.n246 avss -0.00108f
C2933 avdd.n248 avss -3.07e-19
C2934 avdd.n249 avss 0.0374f
C2935 avdd.n250 avss 0.00358f
C2936 avdd.n251 avss 0.0192f
C2937 avdd.n252 avss -1.59e-19
C2938 avdd.n253 avss -1.8e-19
C2939 avdd.n254 avss 0.00875f
C2940 avdd.n255 avss 0.0111f
C2941 avdd.n256 avss 0.0154f
C2942 avdd.n257 avss 0.0183f
C2943 avdd.n258 avss -1.8e-19
C2944 avdd.n259 avss -2.22e-19
C2945 avdd.n260 avss -2.22e-19
C2946 avdd.n261 avss -1.8e-19
C2947 avdd.n262 avss -2.01e-19
C2948 avdd.n263 avss -9.61e-19
C2949 avdd.n264 avss -5.77e-19
C2950 avdd.n265 avss 0.0398f
C2951 avdd.n266 avss -3.07e-19
C2952 avdd.n267 avss -1.8e-19
C2953 avdd.n268 avss 0.0168f
C2954 avdd.n269 avss 0.0189f
C2955 avdd.n270 avss 0.0111f
C2956 avdd.n271 avss 0.00875f
C2957 avdd.n272 avss 0.0167f
C2958 avdd.n273 avss 0.0181f
C2959 avdd.n274 avss -3.6e-19
C2960 avdd.n275 avss -2.01e-19
C2961 avdd.n276 avss -3.07e-19
C2962 avdd.n277 avss -6.46e-19
C2963 avdd.n278 avss -0.00137f
C2964 avdd.n279 avss -0.0013f
C2965 avdd.n280 avss -5.19e-19
C2966 avdd.n281 avss 0.0386f
C2967 avdd.n282 avss 0.00873f
C2968 avdd.n283 avss 0.0111f
C2969 avdd.n284 avss 0.0148f
C2970 avdd.n285 avss 0.019f
C2971 avdd.n286 avss -1.8e-19
C2972 avdd.n287 avss 0.0184f
C2973 avdd.n288 avss -2.44e-19
C2974 avdd.n289 avss -2.33e-19
C2975 avdd.n290 avss 0.0022f
C2976 avdd.n291 avss -1.48e-19
C2977 avdd.n292 avss -1.27e-19
C2978 avdd.n293 avss -2.44e-19
C2979 avdd.n294 avss -8.15e-19
C2980 avdd.n295 avss -0.0014f
C2981 avdd.n296 avss -8.47e-19
C2982 avdd.n297 avss -3.39e-19
C2983 avdd.n298 avss -3.49e-19
C2984 avdd.n299 avss -1.38e-19
C2985 avdd.n300 avss -1.8e-19
C2986 avdd.n301 avss 0.00873f
C2987 avdd.n302 avss 0.0111f
C2988 avdd.n303 avss 0.0154f
C2989 avdd.n304 avss 0.0191f
C2990 avdd.n305 avss -1.8e-19
C2991 avdd.n306 avss 0.0184f
C2992 avdd.n307 avss -1.38e-19
C2993 avdd.n308 avss -1.8e-19
C2994 avdd.n309 avss -2.44e-19
C2995 avdd.n310 avss 0.0411f
C2996 avdd.n311 avss -1.8e-19
C2997 avdd.n312 avss -1.8e-19
C2998 avdd.n313 avss -2.96e-19
C2999 avdd.n314 avss -0.00139f
C3000 avdd.n315 avss -0.00106f
C3001 avdd.n316 avss -0.00357f
C3002 avdd.n317 avss 0.0382f
C3003 avdd.n318 avss -8.47e-19
C3004 avdd.n319 avss -3.28e-19
C3005 avdd.n320 avss -3.28e-19
C3006 avdd.n321 avss -8.26e-19
C3007 avdd.n322 avss 0.0348f
C3008 avdd.n323 avss 0.00357f
C3009 avdd.n324 avss -8.47e-19
C3010 avdd.n325 avss -3.39e-19
C3011 avdd.n326 avss -8.47e-19
C3012 avdd.n327 avss 0.0344f
C3013 avdd.n328 avss 0.00466f
C3014 avdd.n329 avss -3.39e-19
C3015 avdd.n330 avss -6.67e-19
C3016 avdd.n331 avss -5.61e-19
C3017 avdd.n332 avss -3.39e-19
C3018 avdd.n333 avss -6.35e-19
C3019 avdd.n334 avss -0.00139f
C3020 avdd.n335 avss -6.88e-19
C3021 avdd.n336 avss -3.07e-19
C3022 avdd.n337 avss -1.8e-19
C3023 avdd.n338 avss 0.00821f
C3024 avdd.n339 avss -2.75e-19
C3025 avdd.n340 avss 0.0442f
C3026 avdd.n341 avss 0.0179f
C3027 avdd.n342 avss 0.0181f
C3028 avdd.n343 avss -2.75e-19
C3029 avdd.n344 avss -3.39e-19
C3030 avdd.n345 avss -3.6e-19
C3031 avdd.n346 avss -2.01e-19
C3032 avdd.n347 avss -0.0866f
C3033 avdd.n348 avss -0.00336f
C3034 avdd.n349 avss 0.00725f
C3035 avdd.n350 avss 0.0318f
C3036 avdd.n351 avss -0.00158f
C3037 avdd.n352 avss -8.47e-19
C3038 avdd.n353 avss -3.39e-19
C3039 avdd.n354 avss -4.23e-19
C3040 avdd.n355 avss -0.00173f
C3041 avdd.n356 avss 0.0098f
C3042 avdd.n357 avss 0.0298f
C3043 avdd.n358 avss -2.22e-19
C3044 avdd.n359 avss 0.0188f
C3045 avdd.n360 avss -2.33e-19
C3046 avdd.n361 avss -1.59e-19
C3047 avdd.n362 avss -2.22e-19
C3048 avdd.n363 avss 0.00821f
C3049 avdd.n364 avss -2.75e-19
C3050 avdd.n365 avss 0.0112f
C3051 avdd.n366 avss 0.0148f
C3052 avdd.n367 avss 0.0182f
C3053 avdd.n368 avss -1.8e-19
C3054 avdd.n369 avss -2.54e-19
C3055 avdd.n370 avss -2.54e-19
C3056 avdd.n371 avss -1.8e-19
C3057 avdd.n372 avss -1.16e-19
C3058 avdd.n373 avss -2.33e-19
C3059 avdd.n374 avss -0.00126f
C3060 avdd.n375 avss -0.00109f
C3061 avdd.n376 avss -0.00108f
C3062 avdd.n378 avss -3.07e-19
C3063 avdd.n379 avss 0.0374f
C3064 avdd.n380 avss 0.00358f
C3065 avdd.n381 avss 0.0192f
C3066 avdd.n382 avss -1.59e-19
C3067 avdd.n383 avss -1.8e-19
C3068 avdd.n384 avss 0.00875f
C3069 avdd.n385 avss 0.0111f
C3070 avdd.n386 avss 0.0154f
C3071 avdd.n387 avss 0.0183f
C3072 avdd.n388 avss -1.8e-19
C3073 avdd.n389 avss -2.22e-19
C3074 avdd.n390 avss -2.22e-19
C3075 avdd.n391 avss -1.8e-19
C3076 avdd.n392 avss -2.01e-19
C3077 avdd.n393 avss -9.61e-19
C3078 avdd.n394 avss -5.77e-19
C3079 avdd.n395 avss 0.0398f
C3080 avdd.n396 avss -3.07e-19
C3081 avdd.n397 avss -1.8e-19
C3082 avdd.n398 avss 0.0168f
C3083 avdd.n399 avss 0.0189f
C3084 avdd.n400 avss 0.0111f
C3085 avdd.n401 avss 0.00875f
C3086 avdd.n402 avss 0.0167f
C3087 avdd.n403 avss 0.0181f
C3088 avdd.n404 avss -3.6e-19
C3089 avdd.n405 avss -2.01e-19
C3090 avdd.n406 avss -3.07e-19
C3091 avdd.n407 avss -6.46e-19
C3092 avdd.n408 avss -0.00137f
C3093 avdd.n409 avss -0.0013f
C3094 avdd.n410 avss -5.19e-19
C3095 avdd.n411 avss 0.0386f
C3096 avdd.n412 avss 0.00873f
C3097 avdd.n413 avss 0.0111f
C3098 avdd.n414 avss 0.0148f
C3099 avdd.n415 avss 0.019f
C3100 avdd.n416 avss -1.8e-19
C3101 avdd.n417 avss 0.0184f
C3102 avdd.n418 avss -2.44e-19
C3103 avdd.n419 avss -2.33e-19
C3104 avdd.n420 avss 0.0022f
C3105 avdd.n421 avss -1.48e-19
C3106 avdd.n422 avss -1.27e-19
C3107 avdd.n423 avss -2.44e-19
C3108 avdd.n424 avss -8.15e-19
C3109 avdd.n425 avss -0.0014f
C3110 avdd.n426 avss -8.47e-19
C3111 avdd.n427 avss -3.39e-19
C3112 avdd.n428 avss -3.49e-19
C3113 avdd.n429 avss -1.38e-19
C3114 avdd.n430 avss -1.8e-19
C3115 avdd.n431 avss 0.00873f
C3116 avdd.n432 avss 0.0111f
C3117 avdd.n433 avss 0.0154f
C3118 avdd.n434 avss 0.0191f
C3119 avdd.n435 avss -1.8e-19
C3120 avdd.n436 avss 0.0184f
C3121 avdd.n437 avss -1.38e-19
C3122 avdd.n438 avss -1.8e-19
C3123 avdd.n439 avss -2.44e-19
C3124 avdd.n440 avss 0.0411f
C3125 avdd.n441 avss -1.8e-19
C3126 avdd.n442 avss -1.8e-19
C3127 avdd.n443 avss -2.96e-19
C3128 avdd.n444 avss -0.00139f
C3129 avdd.n445 avss -0.00106f
C3130 avdd.n446 avss -0.00357f
C3131 avdd.n447 avss 0.0382f
C3132 avdd.n448 avss -8.47e-19
C3133 avdd.n449 avss -3.28e-19
C3134 avdd.n450 avss -3.28e-19
C3135 avdd.n451 avss -8.26e-19
C3136 avdd.n452 avss 0.0348f
C3137 avdd.n453 avss 0.00357f
C3138 avdd.n454 avss -8.47e-19
C3139 avdd.n455 avss -3.39e-19
C3140 avdd.n456 avss -8.47e-19
C3141 avdd.n457 avss 0.0344f
C3142 avdd.n458 avss 0.00466f
C3143 avdd.n459 avss -3.39e-19
C3144 avdd.n460 avss -6.67e-19
C3145 avdd.n461 avss -5.61e-19
C3146 avdd.n462 avss -3.39e-19
C3147 avdd.n463 avss -6.35e-19
C3148 avdd.n464 avss -0.00139f
C3149 avdd.n465 avss -6.88e-19
C3150 avdd.n466 avss -3.07e-19
C3151 avdd.n467 avss -1.8e-19
C3152 avdd.n468 avss 0.00821f
C3153 avdd.n469 avss -2.75e-19
C3154 avdd.n470 avss 0.0442f
C3155 avdd.n471 avss 0.0179f
C3156 avdd.n472 avss 0.0181f
C3157 avdd.n473 avss -2.75e-19
C3158 avdd.n474 avss -3.39e-19
C3159 avdd.n475 avss -3.6e-19
C3160 avdd.n476 avss -2.01e-19
C3161 avdd.n477 avss -0.0866f
C3162 avdd.n478 avss -0.00336f
C3163 avdd.n479 avss 0.00725f
C3164 avdd.n480 avss 0.0318f
C3165 avdd.n481 avss -0.00158f
C3166 avdd.n482 avss -8.47e-19
C3167 avdd.n483 avss -3.39e-19
C3168 avdd.n484 avss -4.23e-19
C3169 avdd.n485 avss -0.00173f
C3170 avdd.n486 avss 0.0098f
C3171 avdd.n487 avss 0.0298f
C3172 avdd.n488 avss -2.22e-19
C3173 avdd.n489 avss 0.0188f
C3174 avdd.n490 avss -2.33e-19
C3175 avdd.n491 avss -1.59e-19
C3176 avdd.n492 avss -2.22e-19
C3177 avdd.n493 avss 0.00821f
C3178 avdd.n494 avss -2.75e-19
C3179 avdd.n495 avss 0.0112f
C3180 avdd.n496 avss 0.0148f
C3181 avdd.n497 avss 0.0182f
C3182 avdd.n498 avss -1.8e-19
C3183 avdd.n499 avss -2.54e-19
C3184 avdd.n500 avss -2.54e-19
C3185 avdd.n501 avss -1.8e-19
C3186 avdd.n502 avss -1.16e-19
C3187 avdd.n503 avss -2.33e-19
C3188 avdd.n504 avss -0.00126f
C3189 avdd.n505 avss -0.00109f
C3190 avdd.n506 avss -0.00108f
C3191 avdd.n508 avss -3.07e-19
C3192 avdd.n509 avss 0.0374f
C3193 avdd.n510 avss 0.00358f
C3194 avdd.n511 avss 0.0192f
C3195 avdd.n512 avss -1.59e-19
C3196 avdd.n513 avss -1.8e-19
C3197 avdd.n514 avss 0.00875f
C3198 avdd.n515 avss 0.0111f
C3199 avdd.n516 avss 0.0154f
C3200 avdd.n517 avss 0.0183f
C3201 avdd.n518 avss -1.8e-19
C3202 avdd.n519 avss -2.22e-19
C3203 avdd.n520 avss -2.22e-19
C3204 avdd.n521 avss -1.8e-19
C3205 avdd.n522 avss -2.01e-19
C3206 avdd.n523 avss -9.61e-19
C3207 avdd.n524 avss -5.77e-19
C3208 avdd.n525 avss 0.0398f
C3209 avdd.n526 avss -3.07e-19
C3210 avdd.n527 avss -1.8e-19
C3211 avdd.n528 avss 0.0168f
C3212 avdd.n529 avss 0.0189f
C3213 avdd.n530 avss 0.0111f
C3214 avdd.n531 avss 0.00875f
C3215 avdd.n532 avss 0.0167f
C3216 avdd.n533 avss 0.0181f
C3217 avdd.n534 avss -3.6e-19
C3218 avdd.n535 avss -2.01e-19
C3219 avdd.n536 avss -3.07e-19
C3220 avdd.n537 avss -6.46e-19
C3221 avdd.n538 avss -0.00137f
C3222 avdd.n539 avss -0.0013f
C3223 avdd.n540 avss -5.19e-19
C3224 avdd.n541 avss 0.0386f
C3225 avdd.n542 avss 0.00873f
C3226 avdd.n543 avss 0.0111f
C3227 avdd.n544 avss 0.0148f
C3228 avdd.n545 avss 0.019f
C3229 avdd.n546 avss -1.8e-19
C3230 avdd.n547 avss 0.0184f
C3231 avdd.n548 avss -2.44e-19
C3232 avdd.n549 avss -2.33e-19
C3233 avdd.n550 avss 0.0022f
C3234 avdd.n551 avss -1.48e-19
C3235 avdd.n552 avss -1.27e-19
C3236 avdd.n553 avss -2.44e-19
C3237 avdd.n554 avss -8.15e-19
C3238 avdd.n555 avss -0.0014f
C3239 avdd.n556 avss -8.47e-19
C3240 avdd.n557 avss -3.39e-19
C3241 avdd.n558 avss -3.49e-19
C3242 avdd.n559 avss -1.38e-19
C3243 avdd.n560 avss -1.8e-19
C3244 avdd.n561 avss 0.00873f
C3245 avdd.n562 avss 0.0111f
C3246 avdd.n563 avss 0.0154f
C3247 avdd.n564 avss 0.0191f
C3248 avdd.n565 avss -1.8e-19
C3249 avdd.n566 avss 0.0184f
C3250 avdd.n567 avss -1.38e-19
C3251 avdd.n568 avss -1.8e-19
C3252 avdd.n569 avss -2.44e-19
C3253 avdd.n570 avss 0.0411f
C3254 avdd.n571 avss -1.8e-19
C3255 avdd.n572 avss -1.8e-19
C3256 avdd.n573 avss -2.96e-19
C3257 avdd.n574 avss -0.00139f
C3258 avdd.n575 avss -0.00106f
C3259 avdd.n576 avss -0.00357f
C3260 avdd.n577 avss 0.0382f
C3261 avdd.n578 avss -8.47e-19
C3262 avdd.n579 avss -3.28e-19
C3263 avdd.n580 avss -3.28e-19
C3264 avdd.n581 avss -8.26e-19
C3265 avdd.n582 avss 0.0348f
C3266 avdd.n583 avss 0.00357f
C3267 avdd.n584 avss -8.47e-19
C3268 avdd.n585 avss -3.39e-19
C3269 avdd.n586 avss -8.47e-19
C3270 avdd.n587 avss 0.0344f
C3271 avdd.n588 avss 0.00466f
C3272 avdd.n589 avss -3.39e-19
C3273 avdd.n590 avss -6.67e-19
C3274 avdd.n591 avss -5.61e-19
C3275 avdd.n592 avss -3.39e-19
C3276 avdd.n593 avss -6.35e-19
C3277 avdd.n594 avss -0.00139f
C3278 avdd.n595 avss -6.88e-19
C3279 avdd.n596 avss -3.07e-19
C3280 avdd.n597 avss -1.8e-19
C3281 avdd.n598 avss 0.00821f
C3282 avdd.n599 avss -2.75e-19
C3283 avdd.n600 avss 0.0442f
C3284 avdd.n601 avss 0.0179f
C3285 avdd.n602 avss 0.0181f
C3286 avdd.n603 avss -2.75e-19
C3287 avdd.n604 avss -3.39e-19
C3288 avdd.n605 avss -3.6e-19
C3289 avdd.n606 avss -2.01e-19
C3290 avdd.n607 avss -0.0866f
C3291 avdd.n608 avss -0.00336f
C3292 avdd.n609 avss 0.00725f
C3293 avdd.n610 avss 0.0318f
C3294 avdd.n611 avss -0.00158f
C3295 avdd.n612 avss -8.47e-19
C3296 avdd.n613 avss -3.39e-19
C3297 avdd.n614 avss -4.23e-19
C3298 avdd.n615 avss -0.00173f
C3299 avdd.n616 avss 0.0098f
C3300 avdd.n617 avss 0.0298f
C3301 avdd.n618 avss -2.22e-19
C3302 avdd.n619 avss 0.0188f
C3303 avdd.n620 avss -2.33e-19
C3304 avdd.n621 avss -1.59e-19
C3305 avdd.n622 avss -2.22e-19
C3306 avdd.n623 avss 0.00821f
C3307 avdd.n624 avss -2.75e-19
C3308 avdd.n625 avss 0.0112f
C3309 avdd.n626 avss 0.0148f
C3310 avdd.n627 avss 0.0182f
C3311 avdd.n628 avss -1.8e-19
C3312 avdd.n629 avss -2.54e-19
C3313 avdd.n630 avss -2.54e-19
C3314 avdd.n631 avss -1.8e-19
C3315 avdd.n632 avss -1.16e-19
C3316 avdd.n633 avss -2.33e-19
C3317 avdd.n634 avss -0.00126f
C3318 avdd.n635 avss -0.00109f
C3319 avdd.n636 avss -0.00108f
C3320 avdd.n638 avss -3.07e-19
C3321 avdd.n639 avss 0.0374f
C3322 avdd.n640 avss 0.00358f
C3323 avdd.n641 avss 0.0192f
C3324 avdd.n642 avss -1.59e-19
C3325 avdd.n643 avss -1.8e-19
C3326 avdd.n644 avss 0.00875f
C3327 avdd.n645 avss 0.0111f
C3328 avdd.n646 avss 0.0154f
C3329 avdd.n647 avss 0.0183f
C3330 avdd.n648 avss -1.8e-19
C3331 avdd.n649 avss -2.22e-19
C3332 avdd.n650 avss -2.22e-19
C3333 avdd.n651 avss -1.8e-19
C3334 avdd.n652 avss -2.01e-19
C3335 avdd.n653 avss -9.61e-19
C3336 avdd.n654 avss -5.77e-19
C3337 avdd.n655 avss 0.0398f
C3338 avdd.n656 avss -3.07e-19
C3339 avdd.n657 avss -1.8e-19
C3340 avdd.n658 avss 0.0168f
C3341 avdd.n659 avss 0.0189f
C3342 avdd.n660 avss 0.0111f
C3343 avdd.n661 avss 0.00875f
C3344 avdd.n662 avss 0.0167f
C3345 avdd.n663 avss 0.0181f
C3346 avdd.n664 avss -3.6e-19
C3347 avdd.n665 avss -2.01e-19
C3348 avdd.n666 avss -3.07e-19
C3349 avdd.n667 avss -6.46e-19
C3350 avdd.n668 avss -0.00137f
C3351 avdd.n669 avss -0.0013f
C3352 avdd.n670 avss -5.19e-19
C3353 avdd.n671 avss 0.0386f
C3354 avdd.n672 avss 0.00873f
C3355 avdd.n673 avss 0.0111f
C3356 avdd.n674 avss 0.0148f
C3357 avdd.n675 avss 0.019f
C3358 avdd.n676 avss -1.8e-19
C3359 avdd.n677 avss 0.0184f
C3360 avdd.n678 avss -2.44e-19
C3361 avdd.n679 avss -2.33e-19
C3362 avdd.n680 avss 0.0022f
C3363 avdd.n681 avss -1.48e-19
C3364 avdd.n682 avss -1.27e-19
C3365 avdd.n683 avss -2.44e-19
C3366 avdd.n684 avss -8.15e-19
C3367 avdd.n685 avss -0.0014f
C3368 avdd.n686 avss -8.47e-19
C3369 avdd.n687 avss -3.39e-19
C3370 avdd.n688 avss -3.49e-19
C3371 avdd.n689 avss -1.38e-19
C3372 avdd.n690 avss -1.8e-19
C3373 avdd.n691 avss 0.00873f
C3374 avdd.n692 avss 0.0111f
C3375 avdd.n693 avss 0.0154f
C3376 avdd.n694 avss 0.0191f
C3377 avdd.n695 avss -1.8e-19
C3378 avdd.n696 avss 0.0184f
C3379 avdd.n697 avss -1.38e-19
C3380 avdd.n698 avss -1.8e-19
C3381 avdd.n699 avss -2.44e-19
C3382 avdd.n700 avss 0.0411f
C3383 avdd.n701 avss -1.8e-19
C3384 avdd.n702 avss -1.8e-19
C3385 avdd.n703 avss -2.96e-19
C3386 avdd.n704 avss -0.00139f
C3387 avdd.n705 avss -0.00106f
C3388 avdd.n706 avss -0.00357f
C3389 avdd.n707 avss 0.0382f
C3390 avdd.n708 avss -8.47e-19
C3391 avdd.n709 avss -3.28e-19
C3392 avdd.n710 avss -3.28e-19
C3393 avdd.n711 avss -8.26e-19
C3394 avdd.n712 avss 0.0348f
C3395 avdd.n713 avss 0.00357f
C3396 avdd.n714 avss -8.47e-19
C3397 avdd.n715 avss -3.39e-19
C3398 avdd.n716 avss -8.47e-19
C3399 avdd.n717 avss 0.0344f
C3400 avdd.n718 avss 0.00466f
C3401 avdd.n719 avss -3.39e-19
C3402 avdd.n720 avss -6.67e-19
C3403 avdd.n721 avss -5.61e-19
C3404 avdd.n722 avss -3.39e-19
C3405 avdd.n723 avss -6.35e-19
C3406 avdd.n724 avss -0.00139f
C3407 avdd.n725 avss -6.88e-19
C3408 avdd.n726 avss -3.07e-19
C3409 avdd.n727 avss -1.8e-19
C3410 avdd.n728 avss 0.00821f
C3411 avdd.n729 avss -2.75e-19
C3412 avdd.n730 avss 0.0442f
C3413 avdd.n731 avss 0.0179f
C3414 avdd.n732 avss 0.0181f
C3415 avdd.n733 avss -2.75e-19
C3416 avdd.n734 avss -3.39e-19
C3417 avdd.n735 avss -3.6e-19
C3418 avdd.n736 avss -2.01e-19
C3419 avdd.n737 avss -0.0866f
C3420 avdd.n738 avss -0.00336f
C3421 avdd.n739 avss 0.00725f
C3422 avdd.n740 avss 0.0318f
C3423 avdd.n741 avss -0.00158f
C3424 avdd.n742 avss -8.47e-19
C3425 avdd.n743 avss -3.39e-19
C3426 avdd.n744 avss -4.23e-19
C3427 avdd.n745 avss -0.00173f
C3428 avdd.n746 avss 0.0098f
C3429 avdd.n747 avss 0.0298f
C3430 avdd.n748 avss -2.22e-19
C3431 avdd.n749 avss 0.0188f
C3432 avdd.n750 avss -2.33e-19
C3433 avdd.n751 avss -1.59e-19
C3434 avdd.n752 avss -2.22e-19
C3435 avdd.n753 avss 0.00821f
C3436 avdd.n754 avss -2.75e-19
C3437 avdd.n755 avss 0.0112f
C3438 avdd.n756 avss 0.0148f
C3439 avdd.n757 avss 0.0182f
C3440 avdd.n758 avss -1.8e-19
C3441 avdd.n759 avss -2.54e-19
C3442 avdd.n760 avss -2.54e-19
C3443 avdd.n761 avss -1.8e-19
C3444 avdd.n762 avss -1.16e-19
C3445 avdd.n763 avss -2.33e-19
C3446 avdd.n764 avss -0.00126f
C3447 avdd.n765 avss -0.00109f
C3448 avdd.n766 avss -0.00108f
C3449 avdd.n768 avss -3.07e-19
C3450 avdd.n769 avss 0.0374f
C3451 avdd.n770 avss 0.00358f
C3452 avdd.n771 avss 0.0192f
C3453 avdd.n772 avss -1.59e-19
C3454 avdd.n773 avss -1.8e-19
C3455 avdd.n774 avss 0.00875f
C3456 avdd.n775 avss 0.0111f
C3457 avdd.n776 avss 0.0154f
C3458 avdd.n777 avss 0.0183f
C3459 avdd.n778 avss -1.8e-19
C3460 avdd.n779 avss -2.22e-19
C3461 avdd.n780 avss -2.22e-19
C3462 avdd.n781 avss -1.8e-19
C3463 avdd.n782 avss -2.01e-19
C3464 avdd.n783 avss -9.61e-19
C3465 avdd.n784 avss -5.77e-19
C3466 avdd.n785 avss 0.0398f
C3467 avdd.n786 avss -3.07e-19
C3468 avdd.n787 avss -1.8e-19
C3469 avdd.n788 avss 0.0168f
C3470 avdd.n789 avss 0.0189f
C3471 avdd.n790 avss 0.0111f
C3472 avdd.n791 avss 0.00875f
C3473 avdd.n792 avss 0.0167f
C3474 avdd.n793 avss 0.0181f
C3475 avdd.n794 avss -3.6e-19
C3476 avdd.n795 avss -2.01e-19
C3477 avdd.n796 avss -3.07e-19
C3478 avdd.n797 avss -6.46e-19
C3479 avdd.n798 avss -0.00137f
C3480 avdd.n799 avss -0.0013f
C3481 avdd.n800 avss -5.19e-19
C3482 avdd.n801 avss 0.0386f
C3483 avdd.n802 avss 0.00873f
C3484 avdd.n803 avss 0.0111f
C3485 avdd.n804 avss 0.0148f
C3486 avdd.n805 avss 0.019f
C3487 avdd.n806 avss -1.8e-19
C3488 avdd.n807 avss 0.0184f
C3489 avdd.n808 avss -2.44e-19
C3490 avdd.n809 avss -2.33e-19
C3491 avdd.n810 avss 0.0022f
C3492 avdd.n811 avss -1.48e-19
C3493 avdd.n812 avss -1.27e-19
C3494 avdd.n813 avss -2.44e-19
C3495 avdd.n814 avss -8.15e-19
C3496 avdd.n815 avss -0.0014f
C3497 avdd.n816 avss -8.47e-19
C3498 avdd.n817 avss -3.39e-19
C3499 avdd.n818 avss -3.49e-19
C3500 avdd.n819 avss -1.38e-19
C3501 avdd.n820 avss -1.8e-19
C3502 avdd.n821 avss 0.00873f
C3503 avdd.n822 avss 0.0111f
C3504 avdd.n823 avss 0.0154f
C3505 avdd.n824 avss 0.0191f
C3506 avdd.n825 avss -1.8e-19
C3507 avdd.n826 avss 0.0184f
C3508 avdd.n827 avss -1.38e-19
C3509 avdd.n828 avss -1.8e-19
C3510 avdd.n829 avss -2.44e-19
C3511 avdd.n830 avss 0.0411f
C3512 avdd.n831 avss -1.8e-19
C3513 avdd.n832 avss -1.8e-19
C3514 avdd.n833 avss -2.96e-19
C3515 avdd.n834 avss -0.00139f
C3516 avdd.n835 avss -0.00106f
C3517 avdd.n836 avss -0.00357f
C3518 avdd.n837 avss 0.0382f
C3519 avdd.n838 avss -8.47e-19
C3520 avdd.n839 avss -3.28e-19
C3521 avdd.n840 avss -3.28e-19
C3522 avdd.n841 avss -8.26e-19
C3523 avdd.n842 avss 0.0348f
C3524 avdd.n843 avss 0.00357f
C3525 avdd.n844 avss -8.47e-19
C3526 avdd.n845 avss -3.39e-19
C3527 avdd.n846 avss -8.47e-19
C3528 avdd.n847 avss 0.0344f
C3529 avdd.n848 avss 0.00466f
C3530 avdd.n849 avss -3.39e-19
C3531 avdd.n850 avss -6.67e-19
C3532 avdd.n851 avss -5.61e-19
C3533 avdd.n852 avss -3.39e-19
C3534 avdd.n853 avss -6.35e-19
C3535 avdd.n854 avss -0.00139f
C3536 avdd.n855 avss -6.88e-19
C3537 avdd.n856 avss -3.07e-19
C3538 avdd.n857 avss -1.8e-19
C3539 avdd.n858 avss 0.00821f
C3540 avdd.n859 avss -2.75e-19
C3541 avdd.n860 avss 0.0442f
C3542 avdd.n861 avss 0.0179f
C3543 avdd.n862 avss 0.0181f
C3544 avdd.n863 avss -2.75e-19
C3545 avdd.n864 avss -3.39e-19
C3546 avdd.n865 avss -3.6e-19
C3547 avdd.n866 avss -2.01e-19
C3548 avdd.n867 avss -0.0866f
C3549 avdd.n868 avss -0.00336f
C3550 avdd.n869 avss 0.00725f
C3551 avdd.n870 avss 0.0318f
C3552 avdd.n871 avss -0.00158f
C3553 avdd.n872 avss -8.47e-19
C3554 avdd.n873 avss -3.39e-19
C3555 avdd.n874 avss -4.23e-19
C3556 avdd.n875 avss -0.00173f
C3557 avdd.n876 avss 0.0098f
C3558 avdd.n877 avss 0.0298f
C3559 avdd.n878 avss -2.22e-19
C3560 avdd.n879 avss 0.0188f
C3561 avdd.n880 avss -2.33e-19
C3562 avdd.n881 avss -1.59e-19
C3563 avdd.n882 avss -2.22e-19
C3564 avdd.n883 avss 0.00821f
C3565 avdd.n884 avss -2.75e-19
C3566 avdd.n885 avss 0.0112f
C3567 avdd.n886 avss 0.0148f
C3568 avdd.n887 avss 0.0182f
C3569 avdd.n888 avss -1.8e-19
C3570 avdd.n889 avss -2.54e-19
C3571 avdd.n890 avss -2.54e-19
C3572 avdd.n891 avss -1.8e-19
C3573 avdd.n892 avss -1.16e-19
C3574 avdd.n893 avss -2.33e-19
C3575 avdd.n894 avss -0.00126f
C3576 avdd.n895 avss -0.00109f
C3577 avdd.n896 avss -0.00108f
C3578 avdd.n898 avss -3.07e-19
C3579 avdd.n899 avss 0.0374f
C3580 avdd.n900 avss 0.00358f
C3581 avdd.n901 avss 0.0192f
C3582 avdd.n902 avss -1.59e-19
C3583 avdd.n903 avss -1.8e-19
C3584 avdd.n904 avss 0.00875f
C3585 avdd.n905 avss 0.0111f
C3586 avdd.n906 avss 0.0154f
C3587 avdd.n907 avss 0.0183f
C3588 avdd.n908 avss -1.8e-19
C3589 avdd.n909 avss -2.22e-19
C3590 avdd.n910 avss -2.22e-19
C3591 avdd.n911 avss -1.8e-19
C3592 avdd.n912 avss -2.01e-19
C3593 avdd.n913 avss -9.61e-19
C3594 avdd.n914 avss -5.77e-19
C3595 avdd.n915 avss 0.0398f
C3596 avdd.n916 avss -3.07e-19
C3597 avdd.n917 avss -1.8e-19
C3598 avdd.n918 avss 0.0168f
C3599 avdd.n919 avss 0.0189f
C3600 avdd.n920 avss 0.0111f
C3601 avdd.n921 avss 0.00875f
C3602 avdd.n922 avss 0.0167f
C3603 avdd.n923 avss 0.0181f
C3604 avdd.n924 avss -3.6e-19
C3605 avdd.n925 avss -2.01e-19
C3606 avdd.n926 avss -3.07e-19
C3607 avdd.n927 avss -6.46e-19
C3608 avdd.n928 avss -0.00137f
C3609 avdd.n929 avss -0.0013f
C3610 avdd.n930 avss -5.19e-19
C3611 avdd.n931 avss 0.0386f
C3612 avdd.n932 avss 0.00873f
C3613 avdd.n933 avss 0.0111f
C3614 avdd.n934 avss 0.0148f
C3615 avdd.n935 avss 0.019f
C3616 avdd.n936 avss -1.8e-19
C3617 avdd.n937 avss 0.0184f
C3618 avdd.n938 avss -2.44e-19
C3619 avdd.n939 avss -2.33e-19
C3620 avdd.n940 avss 0.0022f
C3621 avdd.n941 avss -1.48e-19
C3622 avdd.n942 avss -1.27e-19
C3623 avdd.n943 avss -2.44e-19
C3624 avdd.n944 avss -8.15e-19
C3625 avdd.n945 avss -0.0014f
C3626 avdd.n946 avss -8.47e-19
C3627 avdd.n947 avss -3.39e-19
C3628 avdd.n948 avss -3.49e-19
C3629 avdd.n949 avss -1.38e-19
C3630 avdd.n950 avss -1.8e-19
C3631 avdd.n951 avss 0.00873f
C3632 avdd.n952 avss 0.0111f
C3633 avdd.n953 avss 0.0154f
C3634 avdd.n954 avss 0.0191f
C3635 avdd.n955 avss -1.8e-19
C3636 avdd.n956 avss 0.0184f
C3637 avdd.n957 avss -1.38e-19
C3638 avdd.n958 avss -1.8e-19
C3639 avdd.n959 avss -2.44e-19
C3640 avdd.n960 avss 0.0411f
C3641 avdd.n961 avss -1.8e-19
C3642 avdd.n962 avss -1.8e-19
C3643 avdd.n963 avss -2.96e-19
C3644 avdd.n964 avss -0.00139f
C3645 avdd.n965 avss -0.00106f
C3646 avdd.n966 avss -0.00357f
C3647 avdd.n967 avss 0.0382f
C3648 avdd.n968 avss -8.47e-19
C3649 avdd.n969 avss -3.28e-19
C3650 avdd.n970 avss -3.28e-19
C3651 avdd.n971 avss -8.26e-19
C3652 avdd.n972 avss 0.0348f
C3653 avdd.n973 avss 0.00357f
C3654 avdd.n974 avss -8.47e-19
C3655 avdd.n975 avss -3.39e-19
C3656 avdd.n976 avss -8.47e-19
C3657 avdd.n977 avss 0.0344f
C3658 avdd.n978 avss 0.00466f
C3659 avdd.n979 avss -3.39e-19
C3660 avdd.n980 avss -6.67e-19
C3661 avdd.n981 avss -5.61e-19
C3662 avdd.n982 avss -3.39e-19
C3663 avdd.n983 avss -6.35e-19
C3664 avdd.n984 avss -0.00139f
C3665 avdd.n985 avss -6.88e-19
C3666 avdd.n986 avss -3.07e-19
C3667 avdd.n987 avss -1.8e-19
C3668 avdd.n988 avss 0.00821f
C3669 avdd.n989 avss -2.75e-19
C3670 avdd.n990 avss 0.0442f
C3671 avdd.n991 avss 0.0179f
C3672 avdd.n992 avss 0.0181f
C3673 avdd.n993 avss -2.75e-19
C3674 avdd.n994 avss -3.39e-19
C3675 avdd.n995 avss -3.6e-19
C3676 avdd.n996 avss -2.01e-19
C3677 avdd.n997 avss -0.0866f
C3678 avdd.n998 avss -0.00336f
C3679 avdd.n999 avss 0.00725f
C3680 avdd.n1000 avss 0.0318f
C3681 avdd.n1001 avss -0.00158f
C3682 avdd.n1002 avss -8.47e-19
C3683 avdd.n1003 avss -3.39e-19
C3684 avdd.n1004 avss -4.23e-19
C3685 avdd.n1005 avss -0.00173f
C3686 avdd.n1006 avss 0.0098f
C3687 avdd.n1007 avss 0.0298f
C3688 avdd.n1008 avss -2.22e-19
C3689 avdd.n1009 avss 0.0188f
C3690 avdd.n1010 avss -2.33e-19
C3691 avdd.n1011 avss -1.59e-19
C3692 avdd.n1012 avss -2.22e-19
C3693 avdd.n1013 avss 0.00821f
C3694 avdd.n1014 avss -2.75e-19
C3695 avdd.n1015 avss 0.0112f
C3696 avdd.n1016 avss 0.0148f
C3697 avdd.n1017 avss 0.0182f
C3698 avdd.n1018 avss -1.8e-19
C3699 avdd.n1019 avss -2.54e-19
C3700 avdd.n1020 avss -2.54e-19
C3701 avdd.n1021 avss -1.8e-19
C3702 avdd.n1022 avss -1.16e-19
C3703 avdd.n1023 avss -2.33e-19
C3704 avdd.n1024 avss -0.00126f
C3705 avdd.n1025 avss -0.00109f
C3706 avdd.n1026 avss -0.00108f
C3707 avdd.n1028 avss -3.07e-19
C3708 avdd.n1029 avss 0.0374f
C3709 avdd.n1030 avss 0.00358f
C3710 avdd.n1031 avss 0.0192f
C3711 avdd.n1032 avss -1.59e-19
C3712 avdd.n1033 avss -1.8e-19
C3713 avdd.n1034 avss 0.00875f
C3714 avdd.n1035 avss 0.0111f
C3715 avdd.n1036 avss 0.0154f
C3716 avdd.n1037 avss 0.0183f
C3717 avdd.n1038 avss -1.8e-19
C3718 avdd.n1039 avss -2.22e-19
C3719 avdd.n1040 avss -2.22e-19
C3720 avdd.n1041 avss -1.8e-19
C3721 avdd.n1042 avss -2.01e-19
C3722 avdd.n1043 avss -9.61e-19
C3723 avdd.n1044 avss -5.77e-19
C3724 avdd.n1045 avss 0.0398f
C3725 avdd.n1046 avss -3.07e-19
C3726 avdd.n1047 avss -1.8e-19
C3727 avdd.n1048 avss 0.0168f
C3728 avdd.n1049 avss 0.0189f
C3729 avdd.n1050 avss 0.0111f
C3730 avdd.n1051 avss 0.00875f
C3731 avdd.n1052 avss 0.0167f
C3732 avdd.n1053 avss 0.0181f
C3733 avdd.n1054 avss -3.6e-19
C3734 avdd.n1055 avss -2.01e-19
C3735 avdd.n1056 avss -3.07e-19
C3736 avdd.n1057 avss -6.46e-19
C3737 avdd.n1058 avss -0.00137f
C3738 avdd.n1059 avss -0.0013f
C3739 avdd.n1060 avss -5.19e-19
C3740 avdd.n1061 avss 0.0386f
C3741 avdd.n1062 avss 0.00873f
C3742 avdd.n1063 avss 0.0111f
C3743 avdd.n1064 avss 0.0148f
C3744 avdd.n1065 avss 0.019f
C3745 avdd.n1066 avss -1.8e-19
C3746 avdd.n1067 avss 0.0184f
C3747 avdd.n1068 avss -2.44e-19
C3748 avdd.n1069 avss -2.33e-19
C3749 avdd.n1070 avss 0.0022f
C3750 avdd.n1071 avss -1.48e-19
C3751 avdd.n1072 avss -1.27e-19
C3752 avdd.n1073 avss -2.44e-19
C3753 avdd.n1074 avss -8.15e-19
C3754 avdd.n1075 avss -0.0014f
C3755 avdd.n1076 avss -8.47e-19
C3756 avdd.n1077 avss -3.39e-19
C3757 avdd.n1078 avss -3.49e-19
C3758 avdd.n1079 avss -1.38e-19
C3759 avdd.n1080 avss -1.8e-19
C3760 avdd.n1081 avss 0.00873f
C3761 avdd.n1082 avss 0.0111f
C3762 avdd.n1083 avss 0.0154f
C3763 avdd.n1084 avss 0.0191f
C3764 avdd.n1085 avss -1.8e-19
C3765 avdd.n1086 avss 0.0184f
C3766 avdd.n1087 avss -1.38e-19
C3767 avdd.n1088 avss -1.8e-19
C3768 avdd.n1089 avss -2.44e-19
C3769 avdd.n1090 avss 0.0411f
C3770 avdd.n1091 avss -1.8e-19
C3771 avdd.n1092 avss -1.8e-19
C3772 avdd.n1093 avss -2.96e-19
C3773 avdd.n1094 avss -0.00139f
C3774 avdd.n1095 avss -0.00106f
C3775 avdd.n1096 avss -0.00357f
C3776 avdd.n1097 avss 0.0382f
C3777 avdd.n1098 avss -8.47e-19
C3778 avdd.n1099 avss -3.28e-19
C3779 avdd.n1100 avss -3.28e-19
C3780 avdd.n1101 avss -8.26e-19
C3781 avdd.n1102 avss 0.0348f
C3782 avdd.n1103 avss 0.00357f
C3783 avdd.n1104 avss -8.47e-19
C3784 avdd.n1105 avss -3.39e-19
C3785 avdd.n1106 avss -8.47e-19
C3786 avdd.n1107 avss 0.0344f
C3787 avdd.n1108 avss 0.00466f
C3788 avdd.n1109 avss -3.39e-19
C3789 avdd.n1110 avss -6.67e-19
C3790 avdd.n1111 avss -5.61e-19
C3791 avdd.n1112 avss -3.39e-19
C3792 avdd.n1113 avss -6.35e-19
C3793 avdd.n1114 avss -0.00139f
C3794 avdd.n1115 avss -6.88e-19
C3795 avdd.n1116 avss -3.07e-19
C3796 avdd.n1117 avss -1.8e-19
C3797 avdd.n1118 avss 0.00821f
C3798 avdd.n1119 avss -2.75e-19
C3799 avdd.n1120 avss 0.0442f
C3800 avdd.n1121 avss 0.0179f
C3801 avdd.n1122 avss 0.0181f
C3802 avdd.n1123 avss -2.75e-19
C3803 avdd.n1124 avss -3.39e-19
C3804 avdd.n1125 avss -3.6e-19
C3805 avdd.n1126 avss -2.01e-19
C3806 avdd.n1127 avss -0.0866f
C3807 avdd.n1128 avss -0.00336f
C3808 avdd.n1129 avss 0.00725f
C3809 avdd.n1130 avss 0.0318f
C3810 avdd.n1131 avss -0.00158f
C3811 avdd.n1132 avss -8.47e-19
C3812 avdd.n1133 avss -3.39e-19
C3813 avdd.n1134 avss -4.23e-19
C3814 avdd.n1135 avss -0.00173f
C3815 avdd.n1136 avss 0.0098f
C3816 avdd.n1137 avss 0.0298f
C3817 avdd.n1138 avss -2.22e-19
C3818 avdd.n1139 avss 0.0188f
C3819 avdd.n1140 avss -2.33e-19
C3820 avdd.n1141 avss -1.59e-19
C3821 avdd.n1142 avss -2.22e-19
C3822 avdd.n1143 avss 0.00821f
C3823 avdd.n1144 avss -2.75e-19
C3824 avdd.n1145 avss 0.0112f
C3825 avdd.n1146 avss 0.0148f
C3826 avdd.n1147 avss 0.0182f
C3827 avdd.n1148 avss -1.8e-19
C3828 avdd.n1149 avss -2.54e-19
C3829 avdd.n1150 avss -2.54e-19
C3830 avdd.n1151 avss -1.8e-19
C3831 avdd.n1152 avss -1.16e-19
C3832 avdd.n1153 avss -2.33e-19
C3833 avdd.n1154 avss -0.00126f
C3834 avdd.n1155 avss -0.00109f
C3835 avdd.n1156 avss -0.00108f
C3836 avdd.n1158 avss -3.07e-19
C3837 avdd.n1159 avss 0.0374f
C3838 avdd.n1160 avss 0.00358f
C3839 avdd.n1161 avss 0.0192f
C3840 avdd.n1162 avss -1.59e-19
C3841 avdd.n1163 avss -1.8e-19
C3842 avdd.n1164 avss 0.00875f
C3843 avdd.n1165 avss 0.0111f
C3844 avdd.n1166 avss 0.0154f
C3845 avdd.n1167 avss 0.0183f
C3846 avdd.n1168 avss -1.8e-19
C3847 avdd.n1169 avss -2.22e-19
C3848 avdd.n1170 avss -2.22e-19
C3849 avdd.n1171 avss -1.8e-19
C3850 avdd.n1172 avss -2.01e-19
C3851 avdd.n1173 avss -9.61e-19
C3852 avdd.n1174 avss -5.77e-19
C3853 avdd.n1175 avss 0.0398f
C3854 avdd.n1176 avss -3.07e-19
C3855 avdd.n1177 avss -1.8e-19
C3856 avdd.n1178 avss 0.0168f
C3857 avdd.n1179 avss 0.0189f
C3858 avdd.n1180 avss 0.0111f
C3859 avdd.n1181 avss 0.00875f
C3860 avdd.n1182 avss 0.0167f
C3861 avdd.n1183 avss 0.0181f
C3862 avdd.n1184 avss -3.6e-19
C3863 avdd.n1185 avss -2.01e-19
C3864 avdd.n1186 avss -3.07e-19
C3865 avdd.n1187 avss -6.46e-19
C3866 avdd.n1188 avss -0.00137f
C3867 avdd.n1189 avss -0.0013f
C3868 avdd.n1190 avss -5.19e-19
C3869 avdd.n1191 avss 0.0386f
C3870 avdd.n1192 avss 0.00873f
C3871 avdd.n1193 avss 0.0111f
C3872 avdd.n1194 avss 0.0148f
C3873 avdd.n1195 avss 0.019f
C3874 avdd.n1196 avss -1.8e-19
C3875 avdd.n1197 avss 0.0184f
C3876 avdd.n1198 avss -2.44e-19
C3877 avdd.n1199 avss -2.33e-19
C3878 avdd.n1200 avss 0.0022f
C3879 avdd.n1201 avss -1.48e-19
C3880 avdd.n1202 avss -1.27e-19
C3881 avdd.n1203 avss -2.44e-19
C3882 avdd.n1204 avss -8.15e-19
C3883 avdd.n1205 avss -0.0014f
C3884 avdd.n1206 avss -8.47e-19
C3885 avdd.n1207 avss -3.39e-19
C3886 avdd.n1208 avss -3.49e-19
C3887 avdd.n1209 avss -1.38e-19
C3888 avdd.n1210 avss -1.8e-19
C3889 avdd.n1211 avss 0.00873f
C3890 avdd.n1212 avss 0.0111f
C3891 avdd.n1213 avss 0.0154f
C3892 avdd.n1214 avss 0.0191f
C3893 avdd.n1215 avss -1.8e-19
C3894 avdd.n1216 avss 0.0184f
C3895 avdd.n1217 avss -1.38e-19
C3896 avdd.n1218 avss -1.8e-19
C3897 avdd.n1219 avss -2.44e-19
C3898 avdd.n1220 avss 0.0411f
C3899 avdd.n1221 avss -1.8e-19
C3900 avdd.n1222 avss -1.8e-19
C3901 avdd.n1223 avss -2.96e-19
C3902 avdd.n1224 avss -0.00139f
C3903 avdd.n1225 avss -0.00106f
C3904 avdd.n1226 avss -0.00357f
C3905 avdd.n1227 avss 0.0382f
C3906 avdd.n1228 avss -8.47e-19
C3907 avdd.n1229 avss -3.28e-19
C3908 avdd.n1230 avss -3.28e-19
C3909 avdd.n1231 avss -8.26e-19
C3910 avdd.n1232 avss 0.0348f
C3911 avdd.n1233 avss 0.00357f
C3912 avdd.n1234 avss -8.47e-19
C3913 avdd.n1235 avss -3.39e-19
C3914 avdd.n1236 avss -8.47e-19
C3915 avdd.n1237 avss 0.0344f
C3916 avdd.n1238 avss 0.00466f
C3917 avdd.n1239 avss -3.39e-19
C3918 avdd.n1240 avss -6.67e-19
C3919 avdd.n1241 avss -5.61e-19
C3920 avdd.n1242 avss -3.39e-19
C3921 avdd.n1243 avss -6.35e-19
C3922 avdd.n1244 avss -0.00139f
C3923 avdd.n1245 avss -6.88e-19
C3924 avdd.n1246 avss -3.07e-19
C3925 avdd.n1247 avss -1.8e-19
C3926 avdd.n1248 avss 0.00821f
C3927 avdd.n1249 avss -2.75e-19
C3928 avdd.n1250 avss 0.0442f
C3929 avdd.n1251 avss 0.0179f
C3930 avdd.n1252 avss 0.0181f
C3931 avdd.n1253 avss -2.75e-19
C3932 avdd.n1254 avss -3.39e-19
C3933 avdd.n1255 avss -3.6e-19
C3934 avdd.n1256 avss -2.01e-19
C3935 avdd.n1257 avss -0.0866f
C3936 avdd.n1258 avss -0.00336f
C3937 avdd.n1259 avss 0.00725f
C3938 avdd.n1260 avss 0.0318f
C3939 avdd.n1261 avss -0.00158f
C3940 avdd.n1262 avss -8.47e-19
C3941 avdd.n1263 avss -3.39e-19
C3942 avdd.n1264 avss -4.23e-19
C3943 avdd.n1265 avss -0.00173f
C3944 avdd.n1266 avss 0.0098f
C3945 avdd.n1267 avss 0.0298f
C3946 avdd.n1268 avss -2.22e-19
C3947 avdd.n1269 avss 0.0188f
C3948 avdd.n1270 avss -2.33e-19
C3949 avdd.n1271 avss -1.59e-19
C3950 avdd.n1272 avss -2.22e-19
C3951 avdd.n1273 avss 0.00821f
C3952 avdd.n1274 avss -2.75e-19
C3953 avdd.n1275 avss 0.0112f
C3954 avdd.n1276 avss 0.0148f
C3955 avdd.n1277 avss 0.0182f
C3956 avdd.n1278 avss -1.8e-19
C3957 avdd.n1279 avss -2.54e-19
C3958 avdd.n1280 avss -2.54e-19
C3959 avdd.n1281 avss -1.8e-19
C3960 avdd.n1282 avss -1.16e-19
C3961 avdd.n1283 avss -2.33e-19
C3962 avdd.n1284 avss -0.00126f
C3963 avdd.n1285 avss -0.00109f
C3964 avdd.n1286 avss -0.00108f
C3965 avdd.n1288 avss -3.07e-19
C3966 avdd.n1289 avss 0.0374f
C3967 avdd.n1290 avss 0.00358f
C3968 avdd.n1291 avss 0.0192f
C3969 avdd.n1292 avss -1.59e-19
C3970 avdd.n1293 avss -1.8e-19
C3971 avdd.n1294 avss 0.00875f
C3972 avdd.n1295 avss 0.0111f
C3973 avdd.n1296 avss 0.0154f
C3974 avdd.n1297 avss 0.0183f
C3975 avdd.n1298 avss -1.8e-19
C3976 avdd.n1299 avss -2.22e-19
C3977 avdd.n1300 avss -2.22e-19
C3978 avdd.n1301 avss -1.8e-19
C3979 avdd.n1302 avss -2.01e-19
C3980 avdd.n1303 avss -9.61e-19
C3981 avdd.n1304 avss -5.77e-19
C3982 avdd.n1305 avss 0.0398f
C3983 avdd.n1306 avss -3.07e-19
C3984 avdd.n1307 avss -1.8e-19
C3985 avdd.n1308 avss 0.0168f
C3986 avdd.n1309 avss 0.0189f
C3987 avdd.n1310 avss 0.0111f
C3988 avdd.n1311 avss 0.00875f
C3989 avdd.n1312 avss 0.0167f
C3990 avdd.n1313 avss 0.0181f
C3991 avdd.n1314 avss -3.6e-19
C3992 avdd.n1315 avss -2.01e-19
C3993 avdd.n1316 avss -3.07e-19
C3994 avdd.n1317 avss -6.46e-19
C3995 avdd.n1318 avss -0.00137f
C3996 avdd.n1319 avss -0.0013f
C3997 avdd.n1320 avss -5.19e-19
C3998 avdd.n1321 avss 0.0386f
C3999 avdd.n1322 avss 0.00873f
C4000 avdd.n1323 avss 0.0111f
C4001 avdd.n1324 avss 0.0148f
C4002 avdd.n1325 avss 0.019f
C4003 avdd.n1326 avss -1.8e-19
C4004 avdd.n1327 avss 0.0184f
C4005 avdd.n1328 avss -2.44e-19
C4006 avdd.n1329 avss -2.33e-19
C4007 avdd.n1330 avss 0.0022f
C4008 avdd.n1331 avss -1.48e-19
C4009 avdd.n1332 avss -1.27e-19
C4010 avdd.n1333 avss -2.44e-19
C4011 avdd.n1334 avss -8.15e-19
C4012 avdd.n1335 avss -0.0014f
C4013 avdd.n1336 avss -8.47e-19
C4014 avdd.n1337 avss -3.39e-19
C4015 avdd.n1338 avss -3.49e-19
C4016 avdd.n1339 avss -1.38e-19
C4017 avdd.n1340 avss -1.8e-19
C4018 avdd.n1341 avss 0.00873f
C4019 avdd.n1342 avss 0.0111f
C4020 avdd.n1343 avss 0.0154f
C4021 avdd.n1344 avss 0.0191f
C4022 avdd.n1345 avss -1.8e-19
C4023 avdd.n1346 avss 0.0184f
C4024 avdd.n1347 avss -1.38e-19
C4025 avdd.n1348 avss -1.8e-19
C4026 avdd.n1349 avss -2.44e-19
C4027 avdd.n1350 avss 0.0411f
C4028 avdd.n1351 avss -1.8e-19
C4029 avdd.n1352 avss -1.8e-19
C4030 avdd.n1353 avss -2.96e-19
C4031 avdd.n1354 avss -0.00139f
C4032 avdd.n1355 avss -0.00106f
C4033 avdd.n1356 avss -0.00357f
C4034 avdd.n1357 avss 0.0382f
C4035 avdd.n1358 avss -8.47e-19
C4036 avdd.n1359 avss -3.28e-19
C4037 avdd.n1360 avss -3.28e-19
C4038 avdd.n1361 avss -8.26e-19
C4039 avdd.n1362 avss 0.0348f
C4040 avdd.n1363 avss 0.00357f
C4041 avdd.n1364 avss -8.47e-19
C4042 avdd.n1365 avss -3.39e-19
C4043 avdd.n1366 avss -8.47e-19
C4044 avdd.n1367 avss 0.0344f
C4045 avdd.n1368 avss 0.00466f
C4046 avdd.n1369 avss -3.39e-19
C4047 avdd.n1370 avss -6.67e-19
C4048 avdd.n1371 avss -5.61e-19
C4049 avdd.n1372 avss -3.39e-19
C4050 avdd.n1373 avss -6.35e-19
C4051 avdd.n1374 avss -0.00139f
C4052 avdd.n1375 avss -6.88e-19
C4053 avdd.n1376 avss -3.07e-19
C4054 avdd.n1377 avss -1.8e-19
C4055 avdd.n1378 avss 0.00821f
C4056 avdd.n1379 avss -2.75e-19
C4057 avdd.n1380 avss 0.0442f
C4058 avdd.n1381 avss 0.0179f
C4059 avdd.n1382 avss 0.0181f
C4060 avdd.n1383 avss -2.75e-19
C4061 avdd.n1384 avss -3.39e-19
C4062 avdd.n1385 avss -3.6e-19
C4063 avdd.n1386 avss -2.01e-19
C4064 avdd.n1387 avss -0.0866f
C4065 avdd.n1388 avss -0.00336f
C4066 avdd.n1389 avss 0.00725f
C4067 avdd.n1390 avss 0.0318f
C4068 avdd.n1391 avss -0.00158f
C4069 avdd.n1392 avss -8.47e-19
C4070 avdd.n1393 avss -3.39e-19
C4071 avdd.n1394 avss -4.23e-19
C4072 avdd.n1395 avss -0.00173f
C4073 avdd.n1396 avss 0.0098f
C4074 avdd.n1397 avss 0.0298f
C4075 avdd.n1398 avss -2.22e-19
C4076 avdd.n1399 avss 0.0188f
C4077 avdd.n1400 avss -2.33e-19
C4078 avdd.n1401 avss -1.59e-19
C4079 avdd.n1402 avss -2.22e-19
C4080 avdd.n1403 avss 0.00821f
C4081 avdd.n1404 avss -2.75e-19
C4082 avdd.n1405 avss 0.0112f
C4083 avdd.n1406 avss 0.0148f
C4084 avdd.n1407 avss 0.0182f
C4085 avdd.n1408 avss -1.8e-19
C4086 avdd.n1409 avss -2.54e-19
C4087 avdd.n1410 avss -2.54e-19
C4088 avdd.n1411 avss -1.8e-19
C4089 avdd.n1412 avss -1.16e-19
C4090 avdd.n1413 avss -2.33e-19
C4091 avdd.n1414 avss -0.00126f
C4092 avdd.n1415 avss -0.00109f
C4093 avdd.n1416 avss -0.00108f
C4094 avdd.n1418 avss -3.07e-19
C4095 avdd.n1419 avss 0.0374f
C4096 avdd.n1420 avss 0.00358f
C4097 avdd.n1421 avss 0.0192f
C4098 avdd.n1422 avss -1.59e-19
C4099 avdd.n1423 avss -1.8e-19
C4100 avdd.n1424 avss 0.00875f
C4101 avdd.n1425 avss 0.0111f
C4102 avdd.n1426 avss 0.0154f
C4103 avdd.n1427 avss 0.0183f
C4104 avdd.n1428 avss -1.8e-19
C4105 avdd.n1429 avss -2.22e-19
C4106 avdd.n1430 avss -2.22e-19
C4107 avdd.n1431 avss -1.8e-19
C4108 avdd.n1432 avss -2.01e-19
C4109 avdd.n1433 avss -9.61e-19
C4110 avdd.n1434 avss -5.77e-19
C4111 avdd.n1435 avss 0.0398f
C4112 avdd.n1436 avss -3.07e-19
C4113 avdd.n1437 avss -1.8e-19
C4114 avdd.n1438 avss 0.0168f
C4115 avdd.n1439 avss 0.0189f
C4116 avdd.n1440 avss 0.0111f
C4117 avdd.n1441 avss 0.00875f
C4118 avdd.n1442 avss 0.0167f
C4119 avdd.n1443 avss 0.0181f
C4120 avdd.n1444 avss -3.6e-19
C4121 avdd.n1445 avss -2.01e-19
C4122 avdd.n1446 avss -3.07e-19
C4123 avdd.n1447 avss -6.46e-19
C4124 avdd.n1448 avss -0.00137f
C4125 avdd.n1449 avss -0.0013f
C4126 avdd.n1450 avss -5.19e-19
C4127 avdd.n1451 avss 0.0386f
C4128 avdd.n1452 avss 0.00873f
C4129 avdd.n1453 avss 0.0111f
C4130 avdd.n1454 avss 0.0148f
C4131 avdd.n1455 avss 0.019f
C4132 avdd.n1456 avss -1.8e-19
C4133 avdd.n1457 avss 0.0184f
C4134 avdd.n1458 avss -2.44e-19
C4135 avdd.n1459 avss -2.33e-19
C4136 avdd.n1460 avss 0.0022f
C4137 avdd.n1461 avss -1.48e-19
C4138 avdd.n1462 avss -1.27e-19
C4139 avdd.n1463 avss -2.44e-19
C4140 avdd.n1464 avss -8.15e-19
C4141 avdd.n1465 avss -0.0014f
C4142 avdd.n1466 avss -8.47e-19
C4143 avdd.n1467 avss -3.39e-19
C4144 avdd.n1468 avss -3.49e-19
C4145 avdd.n1469 avss -1.38e-19
C4146 avdd.n1470 avss -1.8e-19
C4147 avdd.n1471 avss 0.00873f
C4148 avdd.n1472 avss 0.0111f
C4149 avdd.n1473 avss 0.0154f
C4150 avdd.n1474 avss 0.0191f
C4151 avdd.n1475 avss -1.8e-19
C4152 avdd.n1476 avss 0.0184f
C4153 avdd.n1477 avss -1.38e-19
C4154 avdd.n1478 avss -1.8e-19
C4155 avdd.n1479 avss -2.44e-19
C4156 avdd.n1480 avss 0.0411f
C4157 avdd.n1481 avss -1.8e-19
C4158 avdd.n1482 avss -1.8e-19
C4159 avdd.n1483 avss -2.96e-19
C4160 avdd.n1484 avss -0.00139f
C4161 avdd.n1485 avss -0.00106f
C4162 avdd.n1486 avss -0.00357f
C4163 avdd.n1487 avss 0.0382f
C4164 avdd.n1488 avss -8.47e-19
C4165 avdd.n1489 avss -3.28e-19
C4166 avdd.n1490 avss -3.28e-19
C4167 avdd.n1491 avss -8.26e-19
C4168 avdd.n1492 avss 0.0348f
C4169 avdd.n1493 avss 0.00357f
C4170 avdd.n1494 avss -8.47e-19
C4171 avdd.n1495 avss -3.39e-19
C4172 avdd.n1496 avss -8.47e-19
C4173 avdd.n1497 avss 0.0344f
C4174 avdd.n1498 avss 0.00466f
C4175 avdd.n1499 avss -3.39e-19
C4176 avdd.n1500 avss -6.67e-19
C4177 avdd.n1501 avss -5.61e-19
C4178 avdd.n1502 avss -3.39e-19
C4179 avdd.n1503 avss -6.35e-19
C4180 avdd.n1504 avss -0.00139f
C4181 avdd.n1505 avss -6.88e-19
C4182 avdd.n1506 avss -3.07e-19
C4183 avdd.n1507 avss -1.8e-19
C4184 avdd.n1508 avss 0.00821f
C4185 avdd.n1509 avss -2.75e-19
C4186 avdd.n1510 avss 0.0442f
C4187 avdd.n1511 avss 0.0179f
C4188 avdd.n1512 avss 0.0181f
C4189 avdd.n1513 avss -2.75e-19
C4190 avdd.n1514 avss -3.39e-19
C4191 avdd.n1515 avss -3.6e-19
C4192 avdd.n1516 avss -2.01e-19
C4193 avdd.n1517 avss -0.0866f
C4194 avdd.n1518 avss -0.00336f
C4195 avdd.n1519 avss 0.00725f
C4196 avdd.n1520 avss 0.0318f
C4197 avdd.n1521 avss -0.00158f
C4198 avdd.n1522 avss -8.47e-19
C4199 avdd.n1523 avss -3.39e-19
C4200 avdd.n1524 avss -4.23e-19
C4201 avdd.n1525 avss -0.00173f
C4202 avdd.n1526 avss 0.0098f
C4203 avdd.n1527 avss 0.0298f
C4204 avdd.n1528 avss -2.22e-19
C4205 avdd.n1529 avss 0.0188f
C4206 avdd.n1530 avss -2.33e-19
C4207 avdd.n1531 avss -1.59e-19
C4208 avdd.n1532 avss -2.22e-19
C4209 avdd.n1533 avss 0.00821f
C4210 avdd.n1534 avss -2.75e-19
C4211 avdd.n1535 avss 0.0112f
C4212 avdd.n1536 avss 0.0148f
C4213 avdd.n1537 avss 0.0182f
C4214 avdd.n1538 avss -1.8e-19
C4215 avdd.n1539 avss -2.54e-19
C4216 avdd.n1540 avss -2.54e-19
C4217 avdd.n1541 avss -1.8e-19
C4218 avdd.n1542 avss -1.16e-19
C4219 avdd.n1543 avss -2.33e-19
C4220 avdd.n1544 avss -0.00126f
C4221 avdd.n1545 avss -0.00109f
C4222 avdd.n1546 avss -0.00108f
C4223 avdd.n1548 avss -3.07e-19
C4224 avdd.n1549 avss 0.0374f
C4225 avdd.n1550 avss 0.00358f
C4226 avdd.n1551 avss 0.0192f
C4227 avdd.n1552 avss -1.59e-19
C4228 avdd.n1553 avss -1.8e-19
C4229 avdd.n1554 avss 0.00875f
C4230 avdd.n1555 avss 0.0111f
C4231 avdd.n1556 avss 0.0154f
C4232 avdd.n1557 avss 0.0183f
C4233 avdd.n1558 avss -1.8e-19
C4234 avdd.n1559 avss -2.22e-19
C4235 avdd.n1560 avss -2.22e-19
C4236 avdd.n1561 avss -1.8e-19
C4237 avdd.n1562 avss -2.01e-19
C4238 avdd.n1563 avss -9.61e-19
C4239 avdd.n1564 avss -5.77e-19
C4240 avdd.n1565 avss 0.0398f
C4241 avdd.n1566 avss -3.07e-19
C4242 avdd.n1567 avss -1.8e-19
C4243 avdd.n1568 avss 0.0168f
C4244 avdd.n1569 avss 0.0189f
C4245 avdd.n1570 avss 0.0111f
C4246 avdd.n1571 avss 0.00875f
C4247 avdd.n1572 avss 0.0167f
C4248 avdd.n1573 avss 0.0181f
C4249 avdd.n1574 avss -3.6e-19
C4250 avdd.n1575 avss -2.01e-19
C4251 avdd.n1576 avss -3.07e-19
C4252 avdd.n1577 avss -6.46e-19
C4253 avdd.n1578 avss -0.00137f
C4254 avdd.n1579 avss -0.0013f
C4255 avdd.n1580 avss -5.19e-19
C4256 avdd.n1581 avss 0.0386f
C4257 avdd.n1582 avss 0.00873f
C4258 avdd.n1583 avss 0.0111f
C4259 avdd.n1584 avss 0.0148f
C4260 avdd.n1585 avss 0.019f
C4261 avdd.n1586 avss -1.8e-19
C4262 avdd.n1587 avss 0.0184f
C4263 avdd.n1588 avss -2.44e-19
C4264 avdd.n1589 avss -2.33e-19
C4265 avdd.n1590 avss 0.0022f
C4266 avdd.n1591 avss -1.48e-19
C4267 avdd.n1592 avss -1.27e-19
C4268 avdd.n1593 avss -2.44e-19
C4269 avdd.n1594 avss -8.15e-19
C4270 avdd.n1595 avss -0.0014f
C4271 avdd.n1596 avss -8.47e-19
C4272 avdd.n1597 avss -3.39e-19
C4273 avdd.n1598 avss -3.49e-19
C4274 avdd.n1599 avss -1.38e-19
C4275 avdd.n1600 avss -1.8e-19
C4276 avdd.n1601 avss 0.00873f
C4277 avdd.n1602 avss 0.0111f
C4278 avdd.n1603 avss 0.0154f
C4279 avdd.n1604 avss 0.0191f
C4280 avdd.n1605 avss -1.8e-19
C4281 avdd.n1606 avss 0.0184f
C4282 avdd.n1607 avss -1.38e-19
C4283 avdd.n1608 avss -1.8e-19
C4284 avdd.n1609 avss -2.44e-19
C4285 avdd.n1610 avss 0.0411f
C4286 avdd.n1611 avss -1.8e-19
C4287 avdd.n1612 avss -1.8e-19
C4288 avdd.n1613 avss -2.96e-19
C4289 avdd.n1614 avss -0.00139f
C4290 avdd.n1615 avss -0.00106f
C4291 avdd.n1616 avss -0.00357f
C4292 avdd.n1617 avss 0.0382f
C4293 avdd.n1618 avss -0.0038f
C4294 avdd.n1619 avss -0.00562f
C4295 avdd.n1620 avss -0.00797f
C4296 avdd.t190 avss -0.0366f
C4297 avdd.n1621 avss -0.00549f
C4298 avdd.n1622 avss -0.00263f
C4299 avdd.n1623 avss -0.00484f
C4300 avdd.t317 avss -0.0156f
C4301 avdd.n1624 avss -0.0327f
C4302 avdd.t191 avss -0.0021f
C4303 avdd.n1625 avss -8.24e-19
C4304 avdd.t1 avss -0.00353f
C4305 avdd.n1626 avss -0.00283f
C4306 avdd.t164 avss -8.66e-19
C4307 avdd.t22 avss -8.66e-19
C4308 avdd.n1627 avss -0.00196f
C4309 avdd.t254 avss -0.00353f
C4310 avdd.n1628 avss -0.00489f
C4311 avdd.t80 avss -0.00288f
C4312 avdd.n1629 avss -0.00283f
C4313 avdd.t241 avss -8.66e-19
C4314 avdd.t246 avss -8.66e-19
C4315 avdd.n1630 avss -0.00196f
C4316 avdd.t249 avss -0.00288f
C4317 avdd.n1631 avss -0.00287f
C4318 avdd.n1633 avss -0.00514f
C4319 avdd.n1634 avss -0.00151f
C4320 avdd.n1635 avss -0.0158f
C4321 avdd.t252 avss -0.0265f
C4322 avdd.t244 avss -0.0264f
C4323 avdd.t255 avss -0.0215f
C4324 avdd.t256 avss -0.0215f
C4325 avdd.t247 avss -0.0215f
C4326 avdd.t257 avss -0.0161f
C4327 avdd.t243 avss -0.0215f
C4328 avdd.t251 avss -0.0215f
C4329 avdd.t242 avss -0.0215f
C4330 avdd.t250 avss -0.0161f
C4331 avdd.n1636 avss -0.0108f
C4332 avdd.n1637 avss -0.0211f
C4333 avdd.n1638 avss -0.0433f
C4334 avdd.n1639 avss -0.0109f
C4335 avdd.n1640 avss -0.00871f
C4336 avdd.n1642 avss -4.69e-19
C4337 avdd.n1643 avss -4.83e-19
C4338 avdd.n1644 avss -5.62e-19
C4339 avdd.n1645 avss -0.00521f
C4340 avdd.n1646 avss -0.00283f
C4341 avdd.t324 avss -0.00479f
C4342 avdd.n1647 avss -0.00364f
C4343 avdd.n1648 avss -0.00562f
C4344 avdd.n1649 avss -0.00797f
C4345 avdd.t210 avss -0.00215f
C4346 avdd.n1650 avss -0.00826f
C4347 avdd.n1651 avss -0.015f
C4348 avdd.n1653 avss -0.0026f
C4349 avdd.n1654 avss -0.00441f
C4350 avdd.n1655 avss -0.00365f
C4351 avdd.n1656 avss -0.0187f
C4352 avdd.t199 avss -0.0198f
C4353 avdd.t56 avss -0.0146f
C4354 avdd.t64 avss -0.0113f
C4355 avdd.t53 avss -0.0113f
C4356 avdd.t68 avss -0.0107f
C4357 avdd.t161 avss -0.0141f
C4358 avdd.t237 avss -0.0113f
C4359 avdd.t309 avss -0.0113f
C4360 avdd.t25 avss -0.0107f
C4361 avdd.t205 avss -0.0366f
C4362 avdd.n1657 avss -0.00549f
C4363 avdd.n1658 avss -0.00263f
C4364 avdd.n1659 avss -0.00484f
C4365 avdd.t325 avss -0.0156f
C4366 avdd.n1660 avss -0.0327f
C4367 avdd.t206 avss -0.0021f
C4368 avdd.n1661 avss -8.24e-19
C4369 avdd.t26 avss -0.00353f
C4370 avdd.n1662 avss -0.00283f
C4371 avdd.t238 avss -8.66e-19
C4372 avdd.t310 avss -8.66e-19
C4373 avdd.n1663 avss -0.00196f
C4374 avdd.t69 avss -0.00353f
C4375 avdd.n1664 avss -0.00489f
C4376 avdd.t162 avss -0.00288f
C4377 avdd.n1665 avss -0.00283f
C4378 avdd.t65 avss -8.66e-19
C4379 avdd.t54 avss -8.66e-19
C4380 avdd.n1666 avss -0.00196f
C4381 avdd.t57 avss -0.00288f
C4382 avdd.n1667 avss -0.00287f
C4383 avdd.n1669 avss -0.00514f
C4384 avdd.n1670 avss -0.00151f
C4385 avdd.n1671 avss -0.0158f
C4386 avdd.t63 avss -0.0265f
C4387 avdd.t70 avss -0.0264f
C4388 avdd.t66 avss -0.0215f
C4389 avdd.t60 avss -0.0215f
C4390 avdd.t55 avss -0.0215f
C4391 avdd.t61 avss -0.0161f
C4392 avdd.t67 avss -0.0215f
C4393 avdd.t59 avss -0.0215f
C4394 avdd.t62 avss -0.0215f
C4395 avdd.t58 avss -0.0161f
C4396 avdd.n1672 avss -0.0108f
C4397 avdd.n1673 avss -0.0211f
C4398 avdd.n1674 avss -0.0433f
C4399 avdd.n1675 avss -0.0109f
C4400 avdd.n1676 avss -0.00871f
C4401 avdd.n1678 avss -4.69e-19
C4402 avdd.n1679 avss -4.83e-19
C4403 avdd.n1680 avss -5.62e-19
C4404 avdd.n1681 avss -0.00521f
C4405 avdd.n1682 avss -0.00283f
C4406 avdd.t311 avss -0.00479f
C4407 avdd.n1683 avss -0.00213f
C4408 avdd.n1684 avss -0.003f
C4409 avdd.t200 avss -0.00212f
C4410 avdd.n1685 avss -0.00172f
C4411 avdd.n1686 avss -0.00788f
C4412 avdd.n1687 avss -0.00627f
C4413 avdd.t201 avss -0.00212f
C4414 avdd.n1688 avss -0.0045f
C4415 avdd.n1689 avss -0.00278f
C4416 avdd.n1690 avss -0.00145f
C4417 avdd.n1691 avss -0.00506f
C4418 avdd.n1692 avss -0.00213f
C4419 avdd.n1693 avss -0.00283f
C4420 avdd.n1694 avss -8.24e-19
C4421 avdd.n1695 avss -0.00252f
C4422 avdd.n1696 avss -8.24e-19
C4423 avdd.n1697 avss -0.00283f
C4424 avdd.n1698 avss -0.00168f
C4425 avdd.n1699 avss -0.00202f
C4426 avdd.n1700 avss -0.00278f
C4427 avdd.n1701 avss -8.24e-19
C4428 avdd.n1702 avss -0.00252f
C4429 avdd.n1703 avss -0.00283f
C4430 avdd.n1704 avss -0.00283f
C4431 avdd.n1705 avss -0.00168f
C4432 avdd.n1706 avss -0.00481f
C4433 avdd.n1707 avss -0.00653f
C4434 avdd.n1708 avss -0.00632f
C4435 avdd.n1709 avss -0.0101f
C4436 avdd.n1710 avss -0.00797f
C4437 avdd.n1711 avss -0.00562f
C4438 avdd.n1712 avss -0.00378f
C4439 avdd.n1713 avss -0.00145f
C4440 avdd.t319 avss -0.00479f
C4441 avdd.t215 avss -0.00212f
C4442 avdd.n1714 avss -0.00172f
C4443 avdd.n1715 avss -0.00788f
C4444 avdd.t216 avss -0.00212f
C4445 avdd.t180 avss -0.00288f
C4446 avdd.n1717 avss -0.00514f
C4447 avdd.n1718 avss -0.00151f
C4448 avdd.n1719 avss -0.0158f
C4449 avdd.t165 avss -0.0265f
C4450 avdd.t176 avss -0.0264f
C4451 avdd.t172 avss -0.0215f
C4452 avdd.t166 avss -0.0215f
C4453 avdd.t174 avss -0.0215f
C4454 avdd.t169 avss -0.0161f
C4455 avdd.t173 avss -0.0215f
C4456 avdd.t182 avss -0.0215f
C4457 avdd.t175 avss -0.0215f
C4458 avdd.t181 avss -0.0161f
C4459 avdd.n1720 avss -0.0108f
C4460 avdd.n1721 avss -0.0211f
C4461 avdd.n1722 avss -0.0433f
C4462 avdd.n1723 avss -0.0109f
C4463 avdd.n1724 avss -0.00871f
C4464 avdd.n1726 avss -4.69e-19
C4465 avdd.n1727 avss -4.83e-19
C4466 avdd.n1728 avss -5.62e-19
C4467 avdd.n1729 avss -0.00521f
C4468 avdd.n1730 avss -0.00506f
C4469 avdd.n1731 avss -0.00213f
C4470 avdd.t168 avss -8.66e-19
C4471 avdd.t178 avss -8.66e-19
C4472 avdd.n1732 avss -0.00196f
C4473 avdd.n1733 avss -0.00252f
C4474 avdd.n1734 avss -0.00168f
C4475 avdd.t171 avss -0.00353f
C4476 avdd.t126 avss -0.00288f
C4477 avdd.n1735 avss -0.00202f
C4478 avdd.t24 avss -8.66e-19
C4479 avdd.t106 avss -8.66e-19
C4480 avdd.n1736 avss -0.00196f
C4481 avdd.n1737 avss -0.00252f
C4482 avdd.n1738 avss -0.00168f
C4483 avdd.t209 avss -0.0021f
C4484 avdd.t318 avss -0.0156f
C4485 avdd.n1739 avss -0.0327f
C4486 avdd.n1740 avss -0.0101f
C4487 avdd.n1741 avss -0.00632f
C4488 avdd.n1742 avss -0.00484f
C4489 avdd.n1743 avss -0.00653f
C4490 avdd.t259 avss -0.00353f
C4491 avdd.n1744 avss -0.00481f
C4492 avdd.n1745 avss -8.24e-19
C4493 avdd.n1746 avss -0.00283f
C4494 avdd.n1747 avss -0.00283f
C4495 avdd.n1748 avss -0.00283f
C4496 avdd.n1749 avss -8.24e-19
C4497 avdd.n1750 avss -0.00278f
C4498 avdd.n1751 avss -0.00489f
C4499 avdd.n1752 avss -8.24e-19
C4500 avdd.n1753 avss -0.00283f
C4501 avdd.n1754 avss -0.00283f
C4502 avdd.n1755 avss -0.00283f
C4503 avdd.n1756 avss -8.24e-19
C4504 avdd.n1757 avss -0.00287f
C4505 avdd.n1758 avss -0.00278f
C4506 avdd.n1759 avss -0.0045f
C4507 avdd.n1760 avss -0.00627f
C4508 avdd.n1761 avss -0.00283f
C4509 avdd.n1762 avss -0.00213f
C4510 avdd.n1763 avss -0.00234f
C4511 avdd.n1764 avss -0.00364f
C4512 avdd.t207 avss -0.00215f
C4513 avdd.n1765 avss -0.00826f
C4514 avdd.n1766 avss -0.00924f
C4515 avdd.n1767 avss -0.0248f
C4516 avdd.t214 avss -0.0186f
C4517 avdd.t179 avss -0.0146f
C4518 avdd.t167 avss -0.0113f
C4519 avdd.t177 avss -0.0113f
C4520 avdd.t170 avss -0.0107f
C4521 avdd.t125 avss -0.0141f
C4522 avdd.t23 avss -0.0113f
C4523 avdd.t105 avss -0.0113f
C4524 avdd.t258 avss -0.0107f
C4525 avdd.t208 avss -0.0366f
C4526 avdd.t0 avss -0.0107f
C4527 avdd.t21 avss -0.0113f
C4528 avdd.t163 avss -0.0113f
C4529 avdd.t79 avss -0.0141f
C4530 avdd.t253 avss -0.0107f
C4531 avdd.t245 avss -0.0113f
C4532 avdd.t240 avss -0.0113f
C4533 avdd.t248 avss -0.0146f
C4534 avdd.t230 avss -0.0186f
C4535 avdd.n1768 avss -0.0248f
C4536 avdd.n1769 avss -0.00924f
C4537 avdd.n1770 avss -0.00549f
C4538 avdd.n1771 avss -0.00378f
C4539 avdd.n1772 avss -0.00234f
C4540 avdd.n1773 avss -0.00213f
C4541 avdd.n1774 avss -0.00263f
C4542 avdd.t231 avss -0.00212f
C4543 avdd.n1775 avss -0.00172f
C4544 avdd.n1776 avss -0.00788f
C4545 avdd.n1777 avss -0.00627f
C4546 avdd.t232 avss -0.00212f
C4547 avdd.n1778 avss -0.0045f
C4548 avdd.n1779 avss -0.00278f
C4549 avdd.n1780 avss -0.00145f
C4550 avdd.n1781 avss -0.00506f
C4551 avdd.n1782 avss -0.00213f
C4552 avdd.n1783 avss -0.00283f
C4553 avdd.n1784 avss -8.24e-19
C4554 avdd.n1785 avss -0.00252f
C4555 avdd.n1786 avss -8.24e-19
C4556 avdd.n1787 avss -0.00283f
C4557 avdd.n1788 avss -0.00168f
C4558 avdd.n1789 avss -0.00202f
C4559 avdd.n1790 avss -0.00278f
C4560 avdd.n1791 avss -8.24e-19
C4561 avdd.n1792 avss -0.00252f
C4562 avdd.n1793 avss -0.00283f
C4563 avdd.n1794 avss -0.00283f
C4564 avdd.n1795 avss -0.00168f
C4565 avdd.n1796 avss -0.00481f
C4566 avdd.n1797 avss -0.00653f
C4567 avdd.n1798 avss -0.00632f
C4568 avdd.n1799 avss -0.0101f
C4569 avdd.n1800 avss -0.00797f
C4570 avdd.n1801 avss -0.00562f
C4571 avdd.n1802 avss -0.00378f
C4572 avdd.n1803 avss -0.00145f
C4573 avdd.t315 avss -0.00479f
C4574 avdd.t234 avss -0.00212f
C4575 avdd.n1804 avss -0.00172f
C4576 avdd.n1805 avss -0.00788f
C4577 avdd.t235 avss -0.00212f
C4578 avdd.t275 avss -0.00288f
C4579 avdd.n1807 avss -0.00514f
C4580 avdd.n1808 avss -0.00151f
C4581 avdd.n1809 avss -0.0158f
C4582 avdd.t280 avss -0.0265f
C4583 avdd.t285 avss -0.0264f
C4584 avdd.t278 avss -0.0215f
C4585 avdd.t272 avss -0.0215f
C4586 avdd.t273 avss -0.0215f
C4587 avdd.t286 avss -0.0161f
C4588 avdd.t269 avss -0.0215f
C4589 avdd.t277 avss -0.0215f
C4590 avdd.t279 avss -0.0215f
C4591 avdd.t276 avss -0.0161f
C4592 avdd.n1810 avss -0.0108f
C4593 avdd.n1811 avss -0.0211f
C4594 avdd.n1812 avss -0.0433f
C4595 avdd.n1813 avss -0.0109f
C4596 avdd.n1814 avss -0.00871f
C4597 avdd.n1816 avss -4.69e-19
C4598 avdd.n1817 avss -4.83e-19
C4599 avdd.n1818 avss -5.62e-19
C4600 avdd.n1819 avss -0.00521f
C4601 avdd.n1820 avss -0.00506f
C4602 avdd.n1821 avss -0.00213f
C4603 avdd.t284 avss -8.66e-19
C4604 avdd.t271 avss -8.66e-19
C4605 avdd.n1822 avss -0.00196f
C4606 avdd.n1823 avss -0.00252f
C4607 avdd.n1824 avss -0.00168f
C4608 avdd.t282 avss -0.00353f
C4609 avdd.t84 avss -0.00288f
C4610 avdd.n1825 avss -0.00202f
C4611 avdd.t16 avss -8.66e-19
C4612 avdd.t263 avss -8.66e-19
C4613 avdd.n1826 avss -0.00196f
C4614 avdd.n1827 avss -0.00252f
C4615 avdd.n1828 avss -0.00168f
C4616 avdd.t219 avss -0.0021f
C4617 avdd.t326 avss -0.0156f
C4618 avdd.n1829 avss -0.0327f
C4619 avdd.n1830 avss -0.0101f
C4620 avdd.n1831 avss -0.00632f
C4621 avdd.n1832 avss -0.00484f
C4622 avdd.n1833 avss -0.00653f
C4623 avdd.t146 avss -0.00353f
C4624 avdd.n1834 avss -0.00481f
C4625 avdd.n1835 avss -8.24e-19
C4626 avdd.n1836 avss -0.00283f
C4627 avdd.n1837 avss -0.00283f
C4628 avdd.n1838 avss -0.00283f
C4629 avdd.n1839 avss -8.24e-19
C4630 avdd.n1840 avss -0.00278f
C4631 avdd.n1841 avss -0.00489f
C4632 avdd.n1842 avss -8.24e-19
C4633 avdd.n1843 avss -0.00283f
C4634 avdd.n1844 avss -0.00283f
C4635 avdd.n1845 avss -0.00283f
C4636 avdd.n1846 avss -8.24e-19
C4637 avdd.n1847 avss -0.00287f
C4638 avdd.n1848 avss -0.00278f
C4639 avdd.n1849 avss -0.0045f
C4640 avdd.n1850 avss -0.00627f
C4641 avdd.n1851 avss -0.00283f
C4642 avdd.n1852 avss -0.00213f
C4643 avdd.n1853 avss -0.00234f
C4644 avdd.n1854 avss -0.00364f
C4645 avdd.t192 avss -0.00215f
C4646 avdd.n1855 avss -0.00826f
C4647 avdd.n1856 avss -0.00924f
C4648 avdd.n1857 avss -0.0248f
C4649 avdd.t233 avss -0.0186f
C4650 avdd.t274 avss -0.0146f
C4651 avdd.t283 avss -0.0113f
C4652 avdd.t270 avss -0.0113f
C4653 avdd.t281 avss -0.0107f
C4654 avdd.t83 avss -0.0141f
C4655 avdd.t15 avss -0.0113f
C4656 avdd.t262 avss -0.0113f
C4657 avdd.t145 avss -0.0107f
C4658 avdd.t218 avss -0.0366f
C4659 avdd.n1858 avss -0.0151f
C4660 avdd.n1860 avss -0.0026f
C4661 avdd.n1861 avss -0.00441f
C4662 avdd.n1862 avss -0.00354f
C4663 avdd.n1863 avss -0.0113f
C4664 avdd.n1864 avss -0.0248f
C4665 avdd.t220 avss -0.00215f
C4666 avdd.n1865 avss -0.00826f
C4667 avdd.n1866 avss -0.00924f
C4668 avdd.n1867 avss -0.00549f
C4669 avdd.n1868 avss -0.00378f
C4670 avdd.n1869 avss -0.00235f
C4671 avdd.n1870 avss -6.67e-19
C4672 avdd.n1871 avss -0.00323f
C4673 avdd.n1872 avss -0.545f
C4674 avdd.n1873 avss 0.0382f
C4675 avdd.n1874 avss 0.0382f
C4676 avdd.n1875 avss 0.0382f
C4677 avdd.n1876 avss 0.0382f
C4678 avdd.n1877 avss 0.0382f
C4679 avdd.n1878 avss -0.00357f
C4680 avdd.n1879 avss -0.00108f
C4681 avdd.n1880 avss -2.01e-19
C4682 avdd.n1881 avss -0.00173f
C4683 avdd.n1882 avss -2.96e-19
C4684 avdd.n1883 avss -6.67e-19
C4685 avdd.n1884 avss -1.8e-19
C4686 avdd.n1885 avss 0.0411f
C4687 avdd.n1886 avss 0.0191f
C4688 avdd.n1887 avss -1.38e-19
C4689 avdd.n1888 avss -3.39e-19
C4690 avdd.n1889 avss 0.0111f
C4691 avdd.n1890 avss -2.22e-19
C4692 avdd.n1891 avss 0.0374f
C4693 avdd.n1892 avss 0.0112f
C4694 avdd.n1893 avss -1.8e-19
C4695 avdd.n1894 avss -1.8e-19
C4696 avdd.n1895 avss -0.00109f
C4697 avdd.n1896 avss -0.00126f
C4698 avdd.n1897 avss 0.0318f
C4699 avdd.n1898 avss -0.00139f
C4700 avdd.n1899 avss -2.22e-19
C4701 avdd.n1900 avss 0.0188f
C4702 avdd.n1901 avss -2.75e-19
C4703 avdd.n1902 avss -3.6e-19
C4704 avdd.n1903 avss -3.07e-19
C4705 avdd.n1904 avss -6.88e-19
C4706 avdd.n1905 avss 0.00725f
C4707 avdd.n1906 avss -0.00336f
C4708 avdd.n1907 avss -1.8e-19
C4709 avdd.n1908 avss -2.01e-19
C4710 avdd.n1909 avss -0.0866f
C4711 avdd.n1910 avss 0.0179f
C4712 avdd.n1911 avss 0.0442f
C4713 avdd.n1912 avss -3.39e-19
C4714 avdd.n1913 avss -2.75e-19
C4715 avdd.n1914 avss 0.0181f
C4716 avdd.n1915 avss 0.00821f
C4717 avdd.n1916 avss 0.00821f
C4718 avdd.n1917 avss -2.75e-19
C4719 avdd.n1918 avss -2.33e-19
C4720 avdd.n1919 avss -2.54e-19
C4721 avdd.n1920 avss -2.54e-19
C4722 avdd.n1921 avss -2.22e-19
C4723 avdd.n1922 avss -1.59e-19
C4724 avdd.n1923 avss 0.0298f
C4725 avdd.n1924 avss 0.0098f
C4726 avdd.n1925 avss -0.00158f
C4727 avdd.n1926 avss -8.47e-19
C4728 avdd.n1927 avss -4.23e-19
C4729 avdd.n1928 avss -3.39e-19
C4730 avdd.n1929 avss -2.33e-19
C4731 avdd.n1930 avss -1.16e-19
C4732 avdd.n1931 avss 0.0182f
C4733 avdd.n1932 avss 0.0148f
C4734 avdd.n1933 avss 0.00875f
C4735 avdd.n1935 avss -3.07e-19
C4736 avdd.n1936 avss 0.0192f
C4737 avdd.n1937 avss -1.59e-19
C4738 avdd.n1938 avss -1.8e-19
C4739 avdd.n1939 avss 0.00358f
C4740 avdd.n1940 avss -2.22e-19
C4741 avdd.n1941 avss -1.8e-19
C4742 avdd.n1942 avss -1.8e-19
C4743 avdd.n1943 avss 0.0183f
C4744 avdd.n1944 avss 0.0154f
C4745 avdd.n1945 avss 0.0154f
C4746 avdd.n1946 avss 0.0111f
C4747 avdd.n1947 avss 0.0111f
C4748 avdd.n1948 avss -1.8e-19
C4749 avdd.n1949 avss -8.15e-19
C4750 avdd.n1950 avss -1.48e-19
C4751 avdd.n1951 avss -3.39e-19
C4752 avdd.n1952 avss 0.00466f
C4753 avdd.n1953 avss -8.47e-19
C4754 avdd.n1954 avss -0.0014f
C4755 avdd.n1955 avss 0.0344f
C4756 avdd.n1956 avss -8.47e-19
C4757 avdd.n1957 avss 0.0348f
C4758 avdd.n1958 avss -5.19e-19
C4759 avdd.n1959 avss -3.07e-19
C4760 avdd.n1960 avss -3.28e-19
C4761 avdd.n1961 avss -1.8e-19
C4762 avdd.n1962 avss 0.0189f
C4763 avdd.n1963 avss -2.33e-19
C4764 avdd.n1964 avss 0.0022f
C4765 avdd.n1965 avss 0.0386f
C4766 avdd.n1966 avss -2.44e-19
C4767 avdd.n1967 avss 0.0184f
C4768 avdd.n1968 avss 0.00873f
C4769 avdd.n1969 avss 0.0168f
C4770 avdd.n1970 avss 0.0167f
C4771 avdd.n1971 avss -5.77e-19
C4772 avdd.n1972 avss -8.47e-19
C4773 avdd.n1973 avss -2.22e-19
C4774 avdd.n1974 avss 0.00875f
C4775 avdd.n1975 avss -2.54e-19
C4776 avdd.n1976 avss 0.0182f
C4777 avdd.n1977 avss 0.0111f
C4778 avdd.n1978 avss -1.59e-19
C4779 avdd.n1979 avss -3.39e-19
C4780 avdd.n1980 avss -1.59e-19
C4781 avdd.n1981 avss 3e-19
C4782 avdd.n1982 avss -2.54e-19
C4783 avdd.n1983 avss -1.8e-19
C4784 avdd.n1984 avss -1.8e-19
C4785 avdd.n1985 avss -1.16e-19
C4786 avdd.n1986 avss -2.33e-19
C4787 avdd.n1987 avss -3.39e-19
C4788 avdd.n1988 avss -8.47e-19
C4789 avdd.n1989 avss 0.0342f
C4790 avdd.n1990 avss 0.0049f
C4791 avdd.n1991 avss -8.47e-19
C4792 avdd.n1992 avss 0.0388f
C4793 avdd.n1993 avss -3.39e-19
C4794 avdd.n1994 avss -3.39e-19
C4795 avdd.n1995 avss -2.22e-19
C4796 avdd.n1996 avss -2.01e-19
C4797 avdd.n1997 avss -1.8e-19
C4798 avdd.n1998 avss -1.8e-19
C4799 avdd.n1999 avss -2.22e-19
C4800 avdd.n2000 avss 0.0111f
C4801 avdd.n2001 avss -1.8e-19
C4802 avdd.n2002 avss -2.96e-19
C4803 avdd.n2003 avss -2.44e-19
C4804 avdd.n2004 avss 0.0384f
C4805 avdd.n2006 avss -7.52e-19
C4806 avdd.n2008 avss 0.00869f
C4807 avdd.n2009 avss -1.48e-19
C4808 avdd.n2010 avss -0.00173f
C4809 avdd.n2011 avss 0.0269f
C4810 avdd.n2012 avss -1.38e-19
C4811 avdd.n2013 avss -2.44e-19
C4812 avdd.n2014 avss -1.8e-19
C4813 avdd.n2015 avss -1.8e-19
C4814 avdd.n2016 avss -1.38e-19
C4815 avdd.n2017 avss -3.49e-19
C4816 avdd.n2018 avss 0.0184f
C4817 avdd.n2019 avss 0.00873f
C4818 avdd.n2020 avss 0.0422f
C4819 avdd.n2021 avss 0.0197f
C4820 avdd.n2022 avss -2.44e-19
C4821 avdd.n2023 avss -2.44e-19
C4822 avdd.n2024 avss -2.33e-19
C4823 avdd.n2025 avss -2.33e-19
C4824 avdd.n2026 avss -1.8e-19
C4825 avdd.n2027 avss 0.019f
C4826 avdd.n2028 avss 0.00203f
C4827 avdd.n2029 avss -1.27e-19
C4828 avdd.n2030 avss 0.0382f
C4829 avdd.n2031 avss -8.47e-19
C4830 avdd.n2032 avss -3.18e-19
C4831 avdd.n2033 avss 0.03f
C4832 avdd.n2034 avss 0.00899f
C4833 avdd.n2035 avss -0.00113f
C4834 avdd.n2036 avss -0.00512f
C4835 avdd.n2037 avss -1.8e-19
C4836 avdd.n2038 avss -1.8e-19
C4837 avdd.n2039 avss 0.0191f
C4838 avdd.n2040 avss 0.0154f
C4839 avdd.n2041 avss 0.0154f
C4840 avdd.n2042 avss 0.0183f
C4841 avdd.n2043 avss -1.8e-19
C4842 avdd.n2044 avss -1.8e-19
C4843 avdd.n2045 avss -5.82e-19
C4844 avdd.n2046 avss -6.46e-19
C4845 avdd.n2047 avss -3.07e-19
C4846 avdd.n2048 avss 0.0192f
C4847 avdd.n2049 avss 0.00875f
C4848 avdd.n2050 avss 0.0148f
C4849 avdd.n2051 avss 0.0111f
C4850 avdd.n2052 avss -2.22e-19
C4851 avdd.n2053 avss 0.0192f
C4852 avdd.n2054 avss -4.76e-19
C4853 avdd.n2055 avss -0.00128f
C4854 avdd.n2056 avss 0.0346f
C4855 avdd.n2057 avss 0.00378f
C4856 avdd.n2058 avss -8.47e-19
C4857 avdd.n2059 avss 0.0398f
C4858 avdd.n2060 avss -3.07e-19
C4859 avdd.n2061 avss 0.0181f
C4860 avdd.n2062 avss -3.6e-19
C4861 avdd.n2063 avss -2.01e-19
C4862 avdd.n2064 avss -3.28e-19
C4863 avdd.n2065 avss -8.26e-19
C4864 avdd.n2066 avss -6.46e-19
C4865 avdd.n2067 avss -0.00137f
C4866 avdd.n2068 avss -0.0013f
C4867 avdd.n2069 avss 0.00357f
C4868 avdd.n2070 avss -8.47e-19
C4869 avdd.n2071 avss -3.39e-19
C4870 avdd.n2072 avss -1.27e-19
C4871 avdd.n2073 avss -2.44e-19
C4872 avdd.n2074 avss 0.019f
C4873 avdd.n2075 avss 0.0148f
C4874 avdd.n2076 avss 0.00873f
C4875 avdd.n2077 avss 0.0184f
C4876 avdd.n2078 avss -3.49e-19
C4877 avdd.n2079 avss -1.38e-19
C4878 avdd.n2080 avss -1.8e-19
C4879 avdd.n2081 avss -1.8e-19
C4880 avdd.n2082 avss -2.44e-19
C4881 avdd.n2083 avss -1.8e-19
C4882 avdd.n2084 avss -1.8e-19
C4883 avdd.n2085 avss -5.61e-19
C4884 avdd.n2086 avss -3.39e-19
C4885 avdd.n2087 avss -6.35e-19
C4886 avdd.n2088 avss -0.00139f
C4887 avdd.n2089 avss -0.00106f
C4888 avdd.n2090 avss -9.61e-19
C4889 avdd.n2091 avss 0.0382f
C4890 avdd.n2092 avss -0.193f
C4891 avdd.n2093 avss -0.00512f
C4892 avdd.n2094 avss 0.0269f
C4893 avdd.n2095 avss -2.96e-19
C4894 avdd.n2096 avss 0.00869f
C4895 avdd.n2097 avss 0.00203f
C4896 avdd.n2098 avss -2.33e-19
C4897 avdd.n2099 avss 0.019f
C4898 avdd.n2100 avss 0.0111f
C4899 avdd.n2101 avss -1.38e-19
C4900 avdd.n2102 avss -2.44e-19
C4901 avdd.n2103 avss 0.0111f
C4902 avdd.n2104 avss -1.8e-19
C4903 avdd.n2105 avss -1.8e-19
C4904 avdd.n2106 avss 0.03f
C4905 avdd.n2107 avss -3.39e-19
C4906 avdd.n2108 avss -3.39e-19
C4907 avdd.n2109 avss -1.59e-19
C4908 avdd.n2110 avss 0.0111f
C4909 avdd.n2111 avss -1.8e-19
C4910 avdd.n2112 avss -1.8e-19
C4911 avdd.n2113 avss 0.0342f
C4912 avdd.n2114 avss 0.00378f
C4913 avdd.n2115 avss -5.77e-19
C4914 avdd.n2116 avss -2.22e-19
C4915 avdd.n2117 avss 0.0168f
C4916 avdd.n2118 avss -3.6e-19
C4917 avdd.n2119 avss -1.8e-19
C4918 avdd.n2120 avss -8.26e-19
C4919 avdd.n2121 avss -0.0013f
C4920 avdd.n2122 avss -3.39e-19
C4921 avdd.n2123 avss -1.27e-19
C4922 avdd.n2124 avss 0.0022f
C4923 avdd.n2125 avss 0.019f
C4924 avdd.n2126 avss 0.0184f
C4925 avdd.n2127 avss -5.19e-19
C4926 avdd.n2128 avss 0.0386f
C4927 avdd.n2129 avss 0.0111f
C4928 avdd.n2130 avss -1.38e-19
C4929 avdd.n2131 avss -1.38e-19
C4930 avdd.n2132 avss -3.39e-19
C4931 avdd.n2133 avss -3.39e-19
C4932 avdd.n2134 avss -1.8e-19
C4933 avdd.n2135 avss 0.0411f
C4934 avdd.n2136 avss 0.0111f
C4935 avdd.n2137 avss -1.8e-19
C4936 avdd.n2138 avss -1.8e-19
C4937 avdd.n2139 avss -0.00173f
C4938 avdd.n2140 avss -2.96e-19
C4939 avdd.n2141 avss -0.00139f
C4940 avdd.n2142 avss -6.35e-19
C4941 avdd.n2143 avss -4.23e-19
C4942 avdd.n2144 avss -0.00109f
C4943 avdd.n2145 avss -0.00108f
C4944 avdd.n2146 avss 0.0374f
C4945 avdd.n2147 avss 0.0112f
C4946 avdd.n2148 avss -1.8e-19
C4947 avdd.n2149 avss -1.8e-19
C4948 avdd.n2150 avss -0.00126f
C4949 avdd.n2151 avss 0.0318f
C4950 avdd.n2152 avss -0.00139f
C4951 avdd.n2153 avss -2.22e-19
C4952 avdd.n2154 avss 0.0188f
C4953 avdd.n2155 avss -2.75e-19
C4954 avdd.n2156 avss -3.6e-19
C4955 avdd.n2157 avss -3.07e-19
C4956 avdd.n2158 avss -6.88e-19
C4957 avdd.n2159 avss 0.00725f
C4958 avdd.n2160 avss -0.00336f
C4959 avdd.n2161 avss -1.8e-19
C4960 avdd.n2162 avss -2.01e-19
C4961 avdd.n2163 avss -0.0866f
C4962 avdd.n2164 avss 0.0179f
C4963 avdd.n2165 avss 0.0442f
C4964 avdd.n2166 avss -3.39e-19
C4965 avdd.n2167 avss -2.75e-19
C4966 avdd.n2168 avss 0.0181f
C4967 avdd.n2169 avss 0.00821f
C4968 avdd.n2170 avss 0.00821f
C4969 avdd.n2171 avss -2.75e-19
C4970 avdd.n2172 avss -2.33e-19
C4971 avdd.n2173 avss -2.54e-19
C4972 avdd.n2174 avss -2.54e-19
C4973 avdd.n2175 avss -2.22e-19
C4974 avdd.n2176 avss -1.59e-19
C4975 avdd.n2177 avss 0.0298f
C4976 avdd.n2178 avss 0.0098f
C4977 avdd.n2179 avss -0.00158f
C4978 avdd.n2180 avss -8.47e-19
C4979 avdd.n2181 avss -3.39e-19
C4980 avdd.n2182 avss -2.33e-19
C4981 avdd.n2183 avss -1.16e-19
C4982 avdd.n2184 avss 0.0182f
C4983 avdd.n2185 avss 0.0148f
C4984 avdd.n2186 avss 0.00875f
C4985 avdd.n2187 avss -2.22e-19
C4986 avdd.n2188 avss -2.22e-19
C4987 avdd.n2189 avss 0.00358f
C4988 avdd.n2190 avss -1.8e-19
C4989 avdd.n2191 avss -1.59e-19
C4990 avdd.n2192 avss 0.0192f
C4991 avdd.n2193 avss -3.07e-19
C4992 avdd.n2195 avss -0.00357f
C4993 avdd.n2196 avss -0.00106f
C4994 avdd.n2197 avss -9.61e-19
C4995 avdd.n2198 avss -2.01e-19
C4996 avdd.n2199 avss 0.0183f
C4997 avdd.n2200 avss 0.0154f
C4998 avdd.n2201 avss 0.0154f
C4999 avdd.n2202 avss 0.0191f
C5000 avdd.n2203 avss -1.8e-19
C5001 avdd.n2204 avss -1.8e-19
C5002 avdd.n2205 avss -2.44e-19
C5003 avdd.n2206 avss -1.8e-19
C5004 avdd.n2207 avss -1.8e-19
C5005 avdd.n2208 avss -5.61e-19
C5006 avdd.n2209 avss 0.0344f
C5007 avdd.n2210 avss -2.44e-19
C5008 avdd.n2211 avss -8.47e-19
C5009 avdd.n2212 avss -8.15e-19
C5010 avdd.n2213 avss -0.0014f
C5011 avdd.n2214 avss -8.47e-19
C5012 avdd.n2215 avss 0.00466f
C5013 avdd.n2216 avss -3.39e-19
C5014 avdd.n2217 avss -6.67e-19
C5015 avdd.n2218 avss -3.49e-19
C5016 avdd.n2219 avss 0.0184f
C5017 avdd.n2220 avss 0.00873f
C5018 avdd.n2221 avss 0.0148f
C5019 avdd.n2222 avss 0.00873f
C5020 avdd.n2223 avss 0.0111f
C5021 avdd.n2224 avss -2.44e-19
C5022 avdd.n2225 avss -2.33e-19
C5023 avdd.n2226 avss -1.8e-19
C5024 avdd.n2227 avss -1.48e-19
C5025 avdd.n2228 avss -8.47e-19
C5026 avdd.n2229 avss 0.00357f
C5027 avdd.n2230 avss 0.0348f
C5028 avdd.n2231 avss -0.00137f
C5029 avdd.n2232 avss -6.46e-19
C5030 avdd.n2233 avss 0.0189f
C5031 avdd.n2234 avss -3.07e-19
C5032 avdd.n2235 avss -2.01e-19
C5033 avdd.n2236 avss -3.28e-19
C5034 avdd.n2237 avss -3.28e-19
C5035 avdd.n2238 avss -8.47e-19
C5036 avdd.n2239 avss 0.0398f
C5037 avdd.n2240 avss -3.07e-19
C5038 avdd.n2241 avss 0.0181f
C5039 avdd.n2242 avss 0.0167f
C5040 avdd.n2243 avss 0.00875f
C5041 avdd.n2244 avss -2.54e-19
C5042 avdd.n2245 avss -2.54e-19
C5043 avdd.n2246 avss -2.22e-19
C5044 avdd.n2247 avss 0.0192f
C5045 avdd.n2248 avss -4.76e-19
C5046 avdd.n2249 avss -0.00128f
C5047 avdd.n2250 avss 0.0346f
C5048 avdd.n2251 avss -8.47e-19
C5049 avdd.n2252 avss 0.0388f
C5050 avdd.n2253 avss -8.47e-19
C5051 avdd.n2254 avss 0.0049f
C5052 avdd.n2255 avss 3e-19
C5053 avdd.n2256 avss -8.47e-19
C5054 avdd.n2257 avss -3.39e-19
C5055 avdd.n2258 avss -2.33e-19
C5056 avdd.n2259 avss -1.16e-19
C5057 avdd.n2260 avss 0.0182f
C5058 avdd.n2261 avss 0.0148f
C5059 avdd.n2262 avss 0.00875f
C5060 avdd.n2263 avss -2.22e-19
C5061 avdd.n2264 avss -2.22e-19
C5062 avdd.n2265 avss -1.8e-19
C5063 avdd.n2266 avss -1.8e-19
C5064 avdd.n2267 avss -1.59e-19
C5065 avdd.n2268 avss 0.0192f
C5066 avdd.n2269 avss -3.07e-19
C5067 avdd.n2270 avss -6.46e-19
C5068 avdd.n2271 avss -5.82e-19
C5069 avdd.n2272 avss -7.52e-19
C5070 avdd.n2273 avss 0.00899f
C5071 avdd.n2274 avss -0.00113f
C5072 avdd.n2275 avss -8.47e-19
C5073 avdd.n2276 avss -3.39e-19
C5074 avdd.n2277 avss -3.18e-19
C5075 avdd.n2278 avss -2.01e-19
C5076 avdd.n2279 avss 0.0183f
C5077 avdd.n2280 avss 0.0154f
C5078 avdd.n2281 avss 0.0154f
C5079 avdd.n2282 avss 0.0191f
C5080 avdd.n2283 avss -1.8e-19
C5081 avdd.n2284 avss -1.8e-19
C5082 avdd.n2285 avss -1.8e-19
C5083 avdd.n2286 avss -2.44e-19
C5084 avdd.n2287 avss -1.8e-19
C5085 avdd.n2288 avss -1.8e-19
C5086 avdd.n2289 avss -1.38e-19
C5087 avdd.n2291 avss -3.49e-19
C5088 avdd.n2292 avss 0.0184f
C5089 avdd.n2293 avss 0.00873f
C5090 avdd.n2294 avss 0.0422f
C5091 avdd.n2295 avss 0.0197f
C5092 avdd.n2296 avss 0.0384f
C5093 avdd.n2297 avss -2.44e-19
C5094 avdd.n2298 avss -2.44e-19
C5095 avdd.n2299 avss -2.33e-19
C5096 avdd.n2300 avss -1.8e-19
C5097 avdd.n2301 avss -1.48e-19
C5098 avdd.n2302 avss -0.00173f
C5099 avdd.n2304 avss -1.27e-19
C5100 avdd.n2305 avss 0.0382f
C5101 avdd.n2306 avss -0.159f
C5102 avdd.n2307 avss -0.193f
C5103 avdd.n2308 avss -0.00512f
C5104 avdd.n2309 avss 0.0269f
C5105 avdd.n2310 avss -2.96e-19
C5106 avdd.n2311 avss 0.00869f
C5107 avdd.n2312 avss 0.00203f
C5108 avdd.n2313 avss -2.33e-19
C5109 avdd.n2314 avss 0.019f
C5110 avdd.n2315 avss 0.0111f
C5111 avdd.n2316 avss -1.38e-19
C5112 avdd.n2317 avss -2.44e-19
C5113 avdd.n2318 avss 0.0111f
C5114 avdd.n2319 avss -1.8e-19
C5115 avdd.n2320 avss -1.8e-19
C5116 avdd.n2321 avss 0.03f
C5117 avdd.n2322 avss -3.39e-19
C5118 avdd.n2323 avss -3.39e-19
C5119 avdd.n2324 avss -1.59e-19
C5120 avdd.n2325 avss 0.0111f
C5121 avdd.n2326 avss -1.8e-19
C5122 avdd.n2327 avss -1.8e-19
C5123 avdd.n2328 avss 0.0342f
C5124 avdd.n2329 avss 0.00378f
C5125 avdd.n2330 avss -5.77e-19
C5126 avdd.n2331 avss -2.22e-19
C5127 avdd.n2332 avss 0.0168f
C5128 avdd.n2333 avss -3.6e-19
C5129 avdd.n2334 avss -1.8e-19
C5130 avdd.n2335 avss -8.26e-19
C5131 avdd.n2336 avss -0.0013f
C5132 avdd.n2337 avss -3.39e-19
C5133 avdd.n2338 avss -1.27e-19
C5134 avdd.n2339 avss 0.0022f
C5135 avdd.n2340 avss 0.019f
C5136 avdd.n2341 avss 0.0184f
C5137 avdd.n2342 avss -5.19e-19
C5138 avdd.n2343 avss 0.0386f
C5139 avdd.n2344 avss 0.0111f
C5140 avdd.n2345 avss -1.38e-19
C5141 avdd.n2346 avss -1.38e-19
C5142 avdd.n2347 avss -3.39e-19
C5143 avdd.n2348 avss -3.39e-19
C5144 avdd.n2349 avss -1.8e-19
C5145 avdd.n2350 avss 0.0411f
C5146 avdd.n2351 avss 0.0111f
C5147 avdd.n2352 avss -1.8e-19
C5148 avdd.n2353 avss -1.8e-19
C5149 avdd.n2354 avss -0.00173f
C5150 avdd.n2355 avss -2.96e-19
C5151 avdd.n2356 avss -0.00139f
C5152 avdd.n2357 avss -6.35e-19
C5153 avdd.n2358 avss -4.23e-19
C5154 avdd.n2359 avss -0.00109f
C5155 avdd.n2360 avss -0.00108f
C5156 avdd.n2361 avss 0.0374f
C5157 avdd.n2362 avss 0.0112f
C5158 avdd.n2363 avss -1.8e-19
C5159 avdd.n2364 avss -1.8e-19
C5160 avdd.n2365 avss -0.00126f
C5161 avdd.n2366 avss 0.0318f
C5162 avdd.n2367 avss -0.00139f
C5163 avdd.n2368 avss -2.22e-19
C5164 avdd.n2369 avss 0.0188f
C5165 avdd.n2370 avss -2.75e-19
C5166 avdd.n2371 avss -3.6e-19
C5167 avdd.n2372 avss -3.07e-19
C5168 avdd.n2373 avss -6.88e-19
C5169 avdd.n2374 avss 0.00725f
C5170 avdd.n2375 avss -0.00336f
C5171 avdd.n2376 avss -1.8e-19
C5172 avdd.n2377 avss -2.01e-19
C5173 avdd.n2378 avss -0.0866f
C5174 avdd.n2379 avss 0.0179f
C5175 avdd.n2380 avss 0.0442f
C5176 avdd.n2381 avss -3.39e-19
C5177 avdd.n2382 avss -2.75e-19
C5178 avdd.n2383 avss 0.0181f
C5179 avdd.n2384 avss 0.00821f
C5180 avdd.n2385 avss 0.00821f
C5181 avdd.n2386 avss -2.75e-19
C5182 avdd.n2387 avss -2.33e-19
C5183 avdd.n2388 avss -2.54e-19
C5184 avdd.n2389 avss -2.54e-19
C5185 avdd.n2390 avss -2.22e-19
C5186 avdd.n2391 avss -1.59e-19
C5187 avdd.n2392 avss 0.0298f
C5188 avdd.n2393 avss 0.0098f
C5189 avdd.n2394 avss -0.00158f
C5190 avdd.n2395 avss -8.47e-19
C5191 avdd.n2396 avss -3.39e-19
C5192 avdd.n2397 avss -2.33e-19
C5193 avdd.n2398 avss -1.16e-19
C5194 avdd.n2399 avss 0.0182f
C5195 avdd.n2400 avss 0.0148f
C5196 avdd.n2401 avss 0.00875f
C5197 avdd.n2402 avss -2.22e-19
C5198 avdd.n2403 avss -2.22e-19
C5199 avdd.n2404 avss 0.00358f
C5200 avdd.n2405 avss -1.8e-19
C5201 avdd.n2406 avss -1.59e-19
C5202 avdd.n2407 avss 0.0192f
C5203 avdd.n2408 avss -3.07e-19
C5204 avdd.n2410 avss -0.00357f
C5205 avdd.n2411 avss -0.00106f
C5206 avdd.n2412 avss -9.61e-19
C5207 avdd.n2413 avss -2.01e-19
C5208 avdd.n2414 avss 0.0183f
C5209 avdd.n2415 avss 0.0154f
C5210 avdd.n2416 avss 0.0154f
C5211 avdd.n2417 avss 0.0191f
C5212 avdd.n2418 avss -1.8e-19
C5213 avdd.n2419 avss -1.8e-19
C5214 avdd.n2420 avss -2.44e-19
C5215 avdd.n2421 avss -1.8e-19
C5216 avdd.n2422 avss -1.8e-19
C5217 avdd.n2423 avss -5.61e-19
C5218 avdd.n2424 avss 0.0344f
C5219 avdd.n2425 avss -2.44e-19
C5220 avdd.n2426 avss -8.47e-19
C5221 avdd.n2427 avss -8.15e-19
C5222 avdd.n2428 avss -0.0014f
C5223 avdd.n2429 avss -8.47e-19
C5224 avdd.n2430 avss 0.00466f
C5225 avdd.n2431 avss -3.39e-19
C5226 avdd.n2432 avss -6.67e-19
C5227 avdd.n2433 avss -3.49e-19
C5228 avdd.n2434 avss 0.0184f
C5229 avdd.n2435 avss 0.00873f
C5230 avdd.n2436 avss 0.0148f
C5231 avdd.n2437 avss 0.00873f
C5232 avdd.n2438 avss 0.0111f
C5233 avdd.n2439 avss -2.44e-19
C5234 avdd.n2440 avss -2.33e-19
C5235 avdd.n2441 avss -1.8e-19
C5236 avdd.n2442 avss -1.48e-19
C5237 avdd.n2443 avss -8.47e-19
C5238 avdd.n2444 avss 0.00357f
C5239 avdd.n2445 avss 0.0348f
C5240 avdd.n2446 avss -0.00137f
C5241 avdd.n2447 avss -6.46e-19
C5242 avdd.n2448 avss 0.0189f
C5243 avdd.n2449 avss -3.07e-19
C5244 avdd.n2450 avss -2.01e-19
C5245 avdd.n2451 avss -3.28e-19
C5246 avdd.n2452 avss -3.28e-19
C5247 avdd.n2453 avss -8.47e-19
C5248 avdd.n2454 avss 0.0398f
C5249 avdd.n2455 avss -3.07e-19
C5250 avdd.n2456 avss 0.0181f
C5251 avdd.n2457 avss 0.0167f
C5252 avdd.n2458 avss 0.00875f
C5253 avdd.n2459 avss -2.54e-19
C5254 avdd.n2460 avss -2.54e-19
C5255 avdd.n2461 avss -2.22e-19
C5256 avdd.n2462 avss 0.0192f
C5257 avdd.n2463 avss -4.76e-19
C5258 avdd.n2464 avss -0.00128f
C5259 avdd.n2465 avss 0.0346f
C5260 avdd.n2466 avss -8.47e-19
C5261 avdd.n2467 avss 0.0388f
C5262 avdd.n2468 avss -8.47e-19
C5263 avdd.n2469 avss 0.0049f
C5264 avdd.n2470 avss 3e-19
C5265 avdd.n2471 avss -8.47e-19
C5266 avdd.n2472 avss -3.39e-19
C5267 avdd.n2473 avss -2.33e-19
C5268 avdd.n2474 avss -1.16e-19
C5269 avdd.n2475 avss 0.0182f
C5270 avdd.n2476 avss 0.0148f
C5271 avdd.n2477 avss 0.00875f
C5272 avdd.n2478 avss -2.22e-19
C5273 avdd.n2479 avss -2.22e-19
C5274 avdd.n2480 avss -1.8e-19
C5275 avdd.n2481 avss -1.8e-19
C5276 avdd.n2482 avss -1.59e-19
C5277 avdd.n2483 avss 0.0192f
C5278 avdd.n2484 avss -3.07e-19
C5279 avdd.n2485 avss -6.46e-19
C5280 avdd.n2486 avss -5.82e-19
C5281 avdd.n2487 avss -7.52e-19
C5282 avdd.n2488 avss 0.00899f
C5283 avdd.n2489 avss -0.00113f
C5284 avdd.n2490 avss -8.47e-19
C5285 avdd.n2491 avss -3.39e-19
C5286 avdd.n2492 avss -3.18e-19
C5287 avdd.n2493 avss -2.01e-19
C5288 avdd.n2494 avss 0.0183f
C5289 avdd.n2495 avss 0.0154f
C5290 avdd.n2496 avss 0.0154f
C5291 avdd.n2497 avss 0.0191f
C5292 avdd.n2498 avss -1.8e-19
C5293 avdd.n2499 avss -1.8e-19
C5294 avdd.n2500 avss -1.8e-19
C5295 avdd.n2501 avss -2.44e-19
C5296 avdd.n2502 avss -1.8e-19
C5297 avdd.n2503 avss -1.8e-19
C5298 avdd.n2504 avss -1.38e-19
C5299 avdd.n2506 avss -3.49e-19
C5300 avdd.n2507 avss 0.0184f
C5301 avdd.n2508 avss 0.00873f
C5302 avdd.n2509 avss 0.0422f
C5303 avdd.n2510 avss 0.0197f
C5304 avdd.n2511 avss 0.0384f
C5305 avdd.n2512 avss -2.44e-19
C5306 avdd.n2513 avss -2.44e-19
C5307 avdd.n2514 avss -2.33e-19
C5308 avdd.n2515 avss -1.8e-19
C5309 avdd.n2516 avss -1.48e-19
C5310 avdd.n2517 avss -0.00173f
C5311 avdd.n2519 avss -1.27e-19
C5312 avdd.n2520 avss 0.0382f
C5313 avdd.n2521 avss -0.161f
C5314 avdd.n2522 avss -0.195f
C5315 avdd.n2523 avss -0.00512f
C5316 avdd.n2524 avss 0.0269f
C5317 avdd.n2525 avss -2.96e-19
C5318 avdd.n2526 avss 0.00869f
C5319 avdd.n2527 avss 0.00203f
C5320 avdd.n2528 avss -2.33e-19
C5321 avdd.n2529 avss 0.019f
C5322 avdd.n2530 avss 0.0111f
C5323 avdd.n2531 avss -1.38e-19
C5324 avdd.n2532 avss -2.44e-19
C5325 avdd.n2533 avss 0.0111f
C5326 avdd.n2534 avss -1.8e-19
C5327 avdd.n2535 avss -1.8e-19
C5328 avdd.n2536 avss 0.03f
C5329 avdd.n2537 avss -3.39e-19
C5330 avdd.n2538 avss -3.39e-19
C5331 avdd.n2539 avss -1.59e-19
C5332 avdd.n2540 avss 0.0111f
C5333 avdd.n2541 avss -1.8e-19
C5334 avdd.n2542 avss -1.8e-19
C5335 avdd.n2543 avss 0.0342f
C5336 avdd.n2544 avss 0.00378f
C5337 avdd.n2545 avss -5.77e-19
C5338 avdd.n2546 avss -2.22e-19
C5339 avdd.n2547 avss 0.0168f
C5340 avdd.n2548 avss -3.6e-19
C5341 avdd.n2549 avss -1.8e-19
C5342 avdd.n2550 avss -8.26e-19
C5343 avdd.n2551 avss -0.0013f
C5344 avdd.n2552 avss -3.39e-19
C5345 avdd.n2553 avss -1.27e-19
C5346 avdd.n2554 avss 0.0022f
C5347 avdd.n2555 avss 0.019f
C5348 avdd.n2556 avss 0.0184f
C5349 avdd.n2557 avss -5.19e-19
C5350 avdd.n2558 avss 0.0386f
C5351 avdd.n2559 avss 0.0111f
C5352 avdd.n2560 avss -1.38e-19
C5353 avdd.n2561 avss -1.38e-19
C5354 avdd.n2562 avss -3.39e-19
C5355 avdd.n2563 avss -3.39e-19
C5356 avdd.n2564 avss -1.8e-19
C5357 avdd.n2565 avss 0.0411f
C5358 avdd.n2566 avss 0.0111f
C5359 avdd.n2567 avss -1.8e-19
C5360 avdd.n2568 avss -1.8e-19
C5361 avdd.n2569 avss -0.00173f
C5362 avdd.n2570 avss -2.96e-19
C5363 avdd.n2571 avss -0.00139f
C5364 avdd.n2572 avss -6.35e-19
C5365 avdd.n2573 avss -4.23e-19
C5366 avdd.n2574 avss -0.00109f
C5367 avdd.n2575 avss -0.00108f
C5368 avdd.n2576 avss 0.0374f
C5369 avdd.n2577 avss 0.0112f
C5370 avdd.n2578 avss -1.8e-19
C5371 avdd.n2579 avss -1.8e-19
C5372 avdd.n2580 avss -0.00126f
C5373 avdd.n2581 avss 0.0318f
C5374 avdd.n2582 avss -0.00139f
C5375 avdd.n2583 avss -2.22e-19
C5376 avdd.n2584 avss 0.0188f
C5377 avdd.n2585 avss -2.75e-19
C5378 avdd.n2586 avss -3.6e-19
C5379 avdd.n2587 avss -3.07e-19
C5380 avdd.n2588 avss -6.88e-19
C5381 avdd.n2589 avss 0.00725f
C5382 avdd.n2590 avss -0.00336f
C5383 avdd.n2591 avss -1.8e-19
C5384 avdd.n2592 avss -2.01e-19
C5385 avdd.n2593 avss -0.0866f
C5386 avdd.n2594 avss 0.0179f
C5387 avdd.n2595 avss 0.0442f
C5388 avdd.n2596 avss -3.39e-19
C5389 avdd.n2597 avss -2.75e-19
C5390 avdd.n2598 avss 0.0181f
C5391 avdd.n2599 avss 0.00821f
C5392 avdd.n2600 avss 0.00821f
C5393 avdd.n2601 avss -2.75e-19
C5394 avdd.n2602 avss -2.33e-19
C5395 avdd.n2603 avss -2.54e-19
C5396 avdd.n2604 avss -2.54e-19
C5397 avdd.n2605 avss -2.22e-19
C5398 avdd.n2606 avss -1.59e-19
C5399 avdd.n2607 avss 0.0298f
C5400 avdd.n2608 avss 0.0098f
C5401 avdd.n2609 avss -0.00158f
C5402 avdd.n2610 avss -8.47e-19
C5403 avdd.n2611 avss -3.39e-19
C5404 avdd.n2612 avss -2.33e-19
C5405 avdd.n2613 avss -1.16e-19
C5406 avdd.n2614 avss 0.0182f
C5407 avdd.n2615 avss 0.0148f
C5408 avdd.n2616 avss 0.00875f
C5409 avdd.n2617 avss -2.22e-19
C5410 avdd.n2618 avss -2.22e-19
C5411 avdd.n2619 avss 0.00358f
C5412 avdd.n2620 avss -1.8e-19
C5413 avdd.n2621 avss -1.59e-19
C5414 avdd.n2622 avss 0.0192f
C5415 avdd.n2623 avss -3.07e-19
C5416 avdd.n2625 avss -0.00357f
C5417 avdd.n2626 avss -0.00106f
C5418 avdd.n2627 avss -9.61e-19
C5419 avdd.n2628 avss -2.01e-19
C5420 avdd.n2629 avss 0.0183f
C5421 avdd.n2630 avss 0.0154f
C5422 avdd.n2631 avss 0.0154f
C5423 avdd.n2632 avss 0.0191f
C5424 avdd.n2633 avss -1.8e-19
C5425 avdd.n2634 avss -1.8e-19
C5426 avdd.n2635 avss -2.44e-19
C5427 avdd.n2636 avss -1.8e-19
C5428 avdd.n2637 avss -1.8e-19
C5429 avdd.n2638 avss -5.61e-19
C5430 avdd.n2639 avss 0.0344f
C5431 avdd.n2640 avss -2.44e-19
C5432 avdd.n2641 avss -8.47e-19
C5433 avdd.n2642 avss -8.15e-19
C5434 avdd.n2643 avss -0.0014f
C5435 avdd.n2644 avss -8.47e-19
C5436 avdd.n2645 avss 0.00466f
C5437 avdd.n2646 avss -3.39e-19
C5438 avdd.n2647 avss -6.67e-19
C5439 avdd.n2648 avss -3.49e-19
C5440 avdd.n2649 avss 0.0184f
C5441 avdd.n2650 avss 0.00873f
C5442 avdd.n2651 avss 0.0148f
C5443 avdd.n2652 avss 0.00873f
C5444 avdd.n2653 avss 0.0111f
C5445 avdd.n2654 avss -2.44e-19
C5446 avdd.n2655 avss -2.33e-19
C5447 avdd.n2656 avss -1.8e-19
C5448 avdd.n2657 avss -1.48e-19
C5449 avdd.n2658 avss -8.47e-19
C5450 avdd.n2659 avss 0.00357f
C5451 avdd.n2660 avss 0.0348f
C5452 avdd.n2661 avss -0.00137f
C5453 avdd.n2662 avss -6.46e-19
C5454 avdd.n2663 avss 0.0189f
C5455 avdd.n2664 avss -3.07e-19
C5456 avdd.n2665 avss -2.01e-19
C5457 avdd.n2666 avss -3.28e-19
C5458 avdd.n2667 avss -3.28e-19
C5459 avdd.n2668 avss -8.47e-19
C5460 avdd.n2669 avss 0.0398f
C5461 avdd.n2670 avss -3.07e-19
C5462 avdd.n2671 avss 0.0181f
C5463 avdd.n2672 avss 0.0167f
C5464 avdd.n2673 avss 0.00875f
C5465 avdd.n2674 avss -2.54e-19
C5466 avdd.n2675 avss -2.54e-19
C5467 avdd.n2676 avss -2.22e-19
C5468 avdd.n2677 avss 0.0192f
C5469 avdd.n2678 avss -4.76e-19
C5470 avdd.n2679 avss -0.00128f
C5471 avdd.n2680 avss 0.0346f
C5472 avdd.n2681 avss -8.47e-19
C5473 avdd.n2682 avss 0.0388f
C5474 avdd.n2683 avss -8.47e-19
C5475 avdd.n2684 avss 0.0049f
C5476 avdd.n2685 avss 3e-19
C5477 avdd.n2686 avss -8.47e-19
C5478 avdd.n2687 avss -3.39e-19
C5479 avdd.n2688 avss -2.33e-19
C5480 avdd.n2689 avss -1.16e-19
C5481 avdd.n2690 avss 0.0182f
C5482 avdd.n2691 avss 0.0148f
C5483 avdd.n2692 avss 0.00875f
C5484 avdd.n2693 avss -2.22e-19
C5485 avdd.n2694 avss -2.22e-19
C5486 avdd.n2695 avss -1.8e-19
C5487 avdd.n2696 avss -1.8e-19
C5488 avdd.n2697 avss -1.59e-19
C5489 avdd.n2698 avss 0.0192f
C5490 avdd.n2699 avss -3.07e-19
C5491 avdd.n2700 avss -6.46e-19
C5492 avdd.n2701 avss -5.82e-19
C5493 avdd.n2702 avss -7.52e-19
C5494 avdd.n2703 avss 0.00899f
C5495 avdd.n2704 avss -0.00113f
C5496 avdd.n2705 avss -8.47e-19
C5497 avdd.n2706 avss -3.39e-19
C5498 avdd.n2707 avss -3.18e-19
C5499 avdd.n2708 avss -2.01e-19
C5500 avdd.n2709 avss 0.0183f
C5501 avdd.n2710 avss 0.0154f
C5502 avdd.n2711 avss 0.0154f
C5503 avdd.n2712 avss 0.0191f
C5504 avdd.n2713 avss -1.8e-19
C5505 avdd.n2714 avss -1.8e-19
C5506 avdd.n2715 avss -1.8e-19
C5507 avdd.n2716 avss -2.44e-19
C5508 avdd.n2717 avss -1.8e-19
C5509 avdd.n2718 avss -1.8e-19
C5510 avdd.n2719 avss -1.38e-19
C5511 avdd.n2721 avss -3.49e-19
C5512 avdd.n2722 avss 0.0184f
C5513 avdd.n2723 avss 0.00873f
C5514 avdd.n2724 avss 0.0422f
C5515 avdd.n2725 avss 0.0197f
C5516 avdd.n2726 avss 0.0384f
C5517 avdd.n2727 avss -2.44e-19
C5518 avdd.n2728 avss -2.44e-19
C5519 avdd.n2729 avss -2.33e-19
C5520 avdd.n2730 avss -1.8e-19
C5521 avdd.n2731 avss -1.48e-19
C5522 avdd.n2732 avss -0.00173f
C5523 avdd.n2734 avss -1.27e-19
C5524 avdd.n2735 avss 0.0382f
C5525 avdd.n2736 avss -0.161f
C5526 avdd.n2737 avss -0.194f
C5527 avdd.n2738 avss -0.00512f
C5528 avdd.n2739 avss 0.0269f
C5529 avdd.n2740 avss -2.96e-19
C5530 avdd.n2741 avss 0.00869f
C5531 avdd.n2742 avss 0.00203f
C5532 avdd.n2743 avss -2.33e-19
C5533 avdd.n2744 avss 0.019f
C5534 avdd.n2745 avss 0.0111f
C5535 avdd.n2746 avss -1.38e-19
C5536 avdd.n2747 avss -2.44e-19
C5537 avdd.n2748 avss 0.0111f
C5538 avdd.n2749 avss -1.8e-19
C5539 avdd.n2750 avss -1.8e-19
C5540 avdd.n2751 avss 0.03f
C5541 avdd.n2752 avss -3.39e-19
C5542 avdd.n2753 avss -3.39e-19
C5543 avdd.n2754 avss -1.59e-19
C5544 avdd.n2755 avss 0.0111f
C5545 avdd.n2756 avss -1.8e-19
C5546 avdd.n2757 avss -1.8e-19
C5547 avdd.n2758 avss 0.0342f
C5548 avdd.n2759 avss 0.00378f
C5549 avdd.n2760 avss -5.77e-19
C5550 avdd.n2761 avss -2.22e-19
C5551 avdd.n2762 avss 0.0168f
C5552 avdd.n2763 avss -3.6e-19
C5553 avdd.n2764 avss -1.8e-19
C5554 avdd.n2765 avss -8.26e-19
C5555 avdd.n2766 avss -0.0013f
C5556 avdd.n2767 avss -3.39e-19
C5557 avdd.n2768 avss -1.27e-19
C5558 avdd.n2769 avss 0.0022f
C5559 avdd.n2770 avss 0.019f
C5560 avdd.n2771 avss 0.0184f
C5561 avdd.n2772 avss -5.19e-19
C5562 avdd.n2773 avss 0.0386f
C5563 avdd.n2774 avss 0.0111f
C5564 avdd.n2775 avss -1.38e-19
C5565 avdd.n2776 avss -1.38e-19
C5566 avdd.n2777 avss -3.39e-19
C5567 avdd.n2778 avss -3.39e-19
C5568 avdd.n2779 avss -1.8e-19
C5569 avdd.n2780 avss 0.0411f
C5570 avdd.n2781 avss 0.0111f
C5571 avdd.n2782 avss -1.8e-19
C5572 avdd.n2783 avss -1.8e-19
C5573 avdd.n2784 avss -0.00173f
C5574 avdd.n2785 avss -2.96e-19
C5575 avdd.n2786 avss -0.00139f
C5576 avdd.n2787 avss -6.35e-19
C5577 avdd.n2788 avss -4.23e-19
C5578 avdd.n2789 avss -0.00109f
C5579 avdd.n2790 avss -0.00108f
C5580 avdd.n2791 avss 0.0374f
C5581 avdd.n2792 avss 0.0112f
C5582 avdd.n2793 avss -1.8e-19
C5583 avdd.n2794 avss -1.8e-19
C5584 avdd.n2795 avss -0.00126f
C5585 avdd.n2796 avss 0.0318f
C5586 avdd.n2797 avss -0.00139f
C5587 avdd.n2798 avss -2.22e-19
C5588 avdd.n2799 avss 0.0188f
C5589 avdd.n2800 avss -2.75e-19
C5590 avdd.n2801 avss -3.6e-19
C5591 avdd.n2802 avss -3.07e-19
C5592 avdd.n2803 avss -6.88e-19
C5593 avdd.n2804 avss 0.00725f
C5594 avdd.n2805 avss -0.00336f
C5595 avdd.n2806 avss -1.8e-19
C5596 avdd.n2807 avss -2.01e-19
C5597 avdd.n2808 avss -0.0866f
C5598 avdd.n2809 avss 0.0179f
C5599 avdd.n2810 avss 0.0442f
C5600 avdd.n2811 avss -3.39e-19
C5601 avdd.n2812 avss -2.75e-19
C5602 avdd.n2813 avss 0.0181f
C5603 avdd.n2814 avss 0.00821f
C5604 avdd.n2815 avss 0.00821f
C5605 avdd.n2816 avss -2.75e-19
C5606 avdd.n2817 avss -2.33e-19
C5607 avdd.n2818 avss -2.54e-19
C5608 avdd.n2819 avss -2.54e-19
C5609 avdd.n2820 avss -2.22e-19
C5610 avdd.n2821 avss -1.59e-19
C5611 avdd.n2822 avss 0.0298f
C5612 avdd.n2823 avss 0.0098f
C5613 avdd.n2824 avss -0.00158f
C5614 avdd.n2825 avss -8.47e-19
C5615 avdd.n2826 avss -3.39e-19
C5616 avdd.n2827 avss -2.33e-19
C5617 avdd.n2828 avss -1.16e-19
C5618 avdd.n2829 avss 0.0182f
C5619 avdd.n2830 avss 0.0148f
C5620 avdd.n2831 avss 0.00875f
C5621 avdd.n2832 avss -2.22e-19
C5622 avdd.n2833 avss -2.22e-19
C5623 avdd.n2834 avss 0.00358f
C5624 avdd.n2835 avss -1.8e-19
C5625 avdd.n2836 avss -1.59e-19
C5626 avdd.n2837 avss 0.0192f
C5627 avdd.n2838 avss -3.07e-19
C5628 avdd.n2840 avss -0.00357f
C5629 avdd.n2841 avss -0.00106f
C5630 avdd.n2842 avss -9.61e-19
C5631 avdd.n2843 avss -2.01e-19
C5632 avdd.n2844 avss 0.0183f
C5633 avdd.n2845 avss 0.0154f
C5634 avdd.n2846 avss 0.0154f
C5635 avdd.n2847 avss 0.0191f
C5636 avdd.n2848 avss -1.8e-19
C5637 avdd.n2849 avss -1.8e-19
C5638 avdd.n2850 avss -2.44e-19
C5639 avdd.n2851 avss -1.8e-19
C5640 avdd.n2852 avss -1.8e-19
C5641 avdd.n2853 avss -5.61e-19
C5642 avdd.n2854 avss 0.0344f
C5643 avdd.n2855 avss -2.44e-19
C5644 avdd.n2856 avss -8.47e-19
C5645 avdd.n2857 avss -8.15e-19
C5646 avdd.n2858 avss -0.0014f
C5647 avdd.n2859 avss -8.47e-19
C5648 avdd.n2860 avss 0.00466f
C5649 avdd.n2861 avss -3.39e-19
C5650 avdd.n2862 avss -6.67e-19
C5651 avdd.n2863 avss -3.49e-19
C5652 avdd.n2864 avss 0.0184f
C5653 avdd.n2865 avss 0.00873f
C5654 avdd.n2866 avss 0.0148f
C5655 avdd.n2867 avss 0.00873f
C5656 avdd.n2868 avss 0.0111f
C5657 avdd.n2869 avss -2.44e-19
C5658 avdd.n2870 avss -2.33e-19
C5659 avdd.n2871 avss -1.8e-19
C5660 avdd.n2872 avss -1.48e-19
C5661 avdd.n2873 avss -8.47e-19
C5662 avdd.n2874 avss 0.00357f
C5663 avdd.n2875 avss 0.0348f
C5664 avdd.n2876 avss -0.00137f
C5665 avdd.n2877 avss -6.46e-19
C5666 avdd.n2878 avss 0.0189f
C5667 avdd.n2879 avss -3.07e-19
C5668 avdd.n2880 avss -2.01e-19
C5669 avdd.n2881 avss -3.28e-19
C5670 avdd.n2882 avss -3.28e-19
C5671 avdd.n2883 avss -8.47e-19
C5672 avdd.n2884 avss 0.0398f
C5673 avdd.n2885 avss -3.07e-19
C5674 avdd.n2886 avss 0.0181f
C5675 avdd.n2887 avss 0.0167f
C5676 avdd.n2888 avss 0.00875f
C5677 avdd.n2889 avss -2.54e-19
C5678 avdd.n2890 avss -2.54e-19
C5679 avdd.n2891 avss -2.22e-19
C5680 avdd.n2892 avss 0.0192f
C5681 avdd.n2893 avss -4.76e-19
C5682 avdd.n2894 avss -0.00128f
C5683 avdd.n2895 avss 0.0346f
C5684 avdd.n2896 avss -8.47e-19
C5685 avdd.n2897 avss 0.0388f
C5686 avdd.n2898 avss -8.47e-19
C5687 avdd.n2899 avss 0.0049f
C5688 avdd.n2900 avss 3e-19
C5689 avdd.n2901 avss -8.47e-19
C5690 avdd.n2902 avss -3.39e-19
C5691 avdd.n2903 avss -2.33e-19
C5692 avdd.n2904 avss -1.16e-19
C5693 avdd.n2905 avss 0.0182f
C5694 avdd.n2906 avss 0.0148f
C5695 avdd.n2907 avss 0.00875f
C5696 avdd.n2908 avss -2.22e-19
C5697 avdd.n2909 avss -2.22e-19
C5698 avdd.n2910 avss -1.8e-19
C5699 avdd.n2911 avss -1.8e-19
C5700 avdd.n2912 avss -1.59e-19
C5701 avdd.n2913 avss 0.0192f
C5702 avdd.n2914 avss -3.07e-19
C5703 avdd.n2915 avss -6.46e-19
C5704 avdd.n2916 avss -5.82e-19
C5705 avdd.n2917 avss -7.52e-19
C5706 avdd.n2918 avss 0.00899f
C5707 avdd.n2919 avss -0.00113f
C5708 avdd.n2920 avss -8.47e-19
C5709 avdd.n2921 avss -3.39e-19
C5710 avdd.n2922 avss -3.18e-19
C5711 avdd.n2923 avss -2.01e-19
C5712 avdd.n2924 avss 0.0183f
C5713 avdd.n2925 avss 0.0154f
C5714 avdd.n2926 avss 0.0154f
C5715 avdd.n2927 avss 0.0191f
C5716 avdd.n2928 avss -1.8e-19
C5717 avdd.n2929 avss -1.8e-19
C5718 avdd.n2930 avss -1.8e-19
C5719 avdd.n2931 avss -2.44e-19
C5720 avdd.n2932 avss -1.8e-19
C5721 avdd.n2933 avss -1.8e-19
C5722 avdd.n2934 avss -1.38e-19
C5723 avdd.n2936 avss -3.49e-19
C5724 avdd.n2937 avss 0.0184f
C5725 avdd.n2938 avss 0.00873f
C5726 avdd.n2939 avss 0.0422f
C5727 avdd.n2940 avss 0.0197f
C5728 avdd.n2941 avss 0.0384f
C5729 avdd.n2942 avss -2.44e-19
C5730 avdd.n2943 avss -2.44e-19
C5731 avdd.n2944 avss -2.33e-19
C5732 avdd.n2945 avss -1.8e-19
C5733 avdd.n2946 avss -1.48e-19
C5734 avdd.n2947 avss -0.00173f
C5735 avdd.n2949 avss -1.27e-19
C5736 avdd.n2950 avss 0.0382f
C5737 avdd.n2951 avss -0.16f
C5738 avdd.n2952 avss -0.195f
C5739 avdd.n2953 avss -0.00512f
C5740 avdd.n2954 avss 0.0269f
C5741 avdd.n2955 avss -2.96e-19
C5742 avdd.n2956 avss 0.00869f
C5743 avdd.n2957 avss 0.00203f
C5744 avdd.n2958 avss -2.33e-19
C5745 avdd.n2959 avss 0.019f
C5746 avdd.n2960 avss 0.0111f
C5747 avdd.n2961 avss -1.38e-19
C5748 avdd.n2962 avss -2.44e-19
C5749 avdd.n2963 avss 0.0111f
C5750 avdd.n2964 avss -1.8e-19
C5751 avdd.n2965 avss -1.8e-19
C5752 avdd.n2966 avss 0.03f
C5753 avdd.n2967 avss -3.39e-19
C5754 avdd.n2968 avss -3.39e-19
C5755 avdd.n2969 avss -1.59e-19
C5756 avdd.n2970 avss 0.0111f
C5757 avdd.n2971 avss -1.8e-19
C5758 avdd.n2972 avss -1.8e-19
C5759 avdd.n2973 avss 0.0342f
C5760 avdd.n2974 avss 0.00378f
C5761 avdd.n2975 avss -5.77e-19
C5762 avdd.n2976 avss -2.22e-19
C5763 avdd.n2977 avss 0.0168f
C5764 avdd.n2978 avss -3.6e-19
C5765 avdd.n2979 avss -1.8e-19
C5766 avdd.n2980 avss -8.26e-19
C5767 avdd.n2981 avss -0.0013f
C5768 avdd.n2982 avss -3.39e-19
C5769 avdd.n2983 avss -1.27e-19
C5770 avdd.n2984 avss 0.0022f
C5771 avdd.n2985 avss 0.019f
C5772 avdd.n2986 avss 0.0184f
C5773 avdd.n2987 avss -5.19e-19
C5774 avdd.n2988 avss 0.0386f
C5775 avdd.n2989 avss 0.0111f
C5776 avdd.n2990 avss -1.38e-19
C5777 avdd.n2991 avss -1.38e-19
C5778 avdd.n2992 avss -3.39e-19
C5779 avdd.n2993 avss -3.39e-19
C5780 avdd.n2994 avss -1.8e-19
C5781 avdd.n2995 avss 0.0411f
C5782 avdd.n2996 avss 0.0111f
C5783 avdd.n2997 avss -1.8e-19
C5784 avdd.n2998 avss -1.8e-19
C5785 avdd.n2999 avss -0.00173f
C5786 avdd.n3000 avss -2.96e-19
C5787 avdd.n3001 avss -0.00139f
C5788 avdd.n3002 avss -6.35e-19
C5789 avdd.n3003 avss -4.23e-19
C5790 avdd.n3004 avss -0.00109f
C5791 avdd.n3005 avss -0.00108f
C5792 avdd.n3006 avss 0.0374f
C5793 avdd.n3007 avss 0.0112f
C5794 avdd.n3008 avss -1.8e-19
C5795 avdd.n3009 avss -1.8e-19
C5796 avdd.n3010 avss -0.00126f
C5797 avdd.n3011 avss 0.0318f
C5798 avdd.n3012 avss -0.00139f
C5799 avdd.n3013 avss -2.22e-19
C5800 avdd.n3014 avss 0.0188f
C5801 avdd.n3015 avss -2.75e-19
C5802 avdd.n3016 avss -3.6e-19
C5803 avdd.n3017 avss -3.07e-19
C5804 avdd.n3018 avss -6.88e-19
C5805 avdd.n3019 avss 0.00725f
C5806 avdd.n3020 avss -0.00336f
C5807 avdd.n3021 avss -1.8e-19
C5808 avdd.n3022 avss -2.01e-19
C5809 avdd.n3023 avss -0.0866f
C5810 avdd.n3024 avss 0.0179f
C5811 avdd.n3025 avss 0.0442f
C5812 avdd.n3026 avss -3.39e-19
C5813 avdd.n3027 avss -2.75e-19
C5814 avdd.n3028 avss 0.0181f
C5815 avdd.n3029 avss 0.00821f
C5816 avdd.n3030 avss 0.00821f
C5817 avdd.n3031 avss -2.75e-19
C5818 avdd.n3032 avss -2.33e-19
C5819 avdd.n3033 avss -2.54e-19
C5820 avdd.n3034 avss -2.54e-19
C5821 avdd.n3035 avss -2.22e-19
C5822 avdd.n3036 avss -1.59e-19
C5823 avdd.n3037 avss 0.0298f
C5824 avdd.n3038 avss 0.0098f
C5825 avdd.n3039 avss -0.00158f
C5826 avdd.n3040 avss -8.47e-19
C5827 avdd.n3041 avss -3.39e-19
C5828 avdd.n3042 avss -2.33e-19
C5829 avdd.n3043 avss -1.16e-19
C5830 avdd.n3044 avss 0.0182f
C5831 avdd.n3045 avss 0.0148f
C5832 avdd.n3046 avss 0.00875f
C5833 avdd.n3047 avss -2.22e-19
C5834 avdd.n3048 avss -2.22e-19
C5835 avdd.n3049 avss 0.00358f
C5836 avdd.n3050 avss -1.8e-19
C5837 avdd.n3051 avss -1.59e-19
C5838 avdd.n3052 avss 0.0192f
C5839 avdd.n3053 avss -3.07e-19
C5840 avdd.n3055 avss -0.00357f
C5841 avdd.n3056 avss -0.00106f
C5842 avdd.n3057 avss -9.61e-19
C5843 avdd.n3058 avss -2.01e-19
C5844 avdd.n3059 avss 0.0183f
C5845 avdd.n3060 avss 0.0154f
C5846 avdd.n3061 avss 0.0154f
C5847 avdd.n3062 avss 0.0191f
C5848 avdd.n3063 avss -1.8e-19
C5849 avdd.n3064 avss -1.8e-19
C5850 avdd.n3065 avss -2.44e-19
C5851 avdd.n3066 avss -1.8e-19
C5852 avdd.n3067 avss -1.8e-19
C5853 avdd.n3068 avss -5.61e-19
C5854 avdd.n3069 avss 0.0344f
C5855 avdd.n3070 avss -2.44e-19
C5856 avdd.n3071 avss -8.47e-19
C5857 avdd.n3072 avss -8.15e-19
C5858 avdd.n3073 avss -0.0014f
C5859 avdd.n3074 avss -8.47e-19
C5860 avdd.n3075 avss 0.00466f
C5861 avdd.n3076 avss -3.39e-19
C5862 avdd.n3077 avss -6.67e-19
C5863 avdd.n3078 avss -3.49e-19
C5864 avdd.n3079 avss 0.0184f
C5865 avdd.n3080 avss 0.00873f
C5866 avdd.n3081 avss 0.0148f
C5867 avdd.n3082 avss 0.00873f
C5868 avdd.n3083 avss 0.0111f
C5869 avdd.n3084 avss -2.44e-19
C5870 avdd.n3085 avss -2.33e-19
C5871 avdd.n3086 avss -1.8e-19
C5872 avdd.n3087 avss -1.48e-19
C5873 avdd.n3088 avss -8.47e-19
C5874 avdd.n3089 avss 0.00357f
C5875 avdd.n3090 avss 0.0348f
C5876 avdd.n3091 avss -0.00137f
C5877 avdd.n3092 avss -6.46e-19
C5878 avdd.n3093 avss 0.0189f
C5879 avdd.n3094 avss -3.07e-19
C5880 avdd.n3095 avss -2.01e-19
C5881 avdd.n3096 avss -3.28e-19
C5882 avdd.n3097 avss -3.28e-19
C5883 avdd.n3098 avss -8.47e-19
C5884 avdd.n3099 avss 0.0398f
C5885 avdd.n3100 avss -3.07e-19
C5886 avdd.n3101 avss 0.0181f
C5887 avdd.n3102 avss 0.0167f
C5888 avdd.n3103 avss 0.00875f
C5889 avdd.n3104 avss -2.54e-19
C5890 avdd.n3105 avss -2.54e-19
C5891 avdd.n3106 avss -2.22e-19
C5892 avdd.n3107 avss 0.0192f
C5893 avdd.n3108 avss -4.76e-19
C5894 avdd.n3109 avss -0.00128f
C5895 avdd.n3110 avss 0.0346f
C5896 avdd.n3111 avss -8.47e-19
C5897 avdd.n3112 avss 0.0388f
C5898 avdd.n3113 avss -8.47e-19
C5899 avdd.n3114 avss 0.0049f
C5900 avdd.n3115 avss 3e-19
C5901 avdd.n3116 avss -8.47e-19
C5902 avdd.n3117 avss -3.39e-19
C5903 avdd.n3118 avss -2.33e-19
C5904 avdd.n3119 avss -1.16e-19
C5905 avdd.n3120 avss 0.0182f
C5906 avdd.n3121 avss 0.0148f
C5907 avdd.n3122 avss 0.00875f
C5908 avdd.n3123 avss -2.22e-19
C5909 avdd.n3124 avss -2.22e-19
C5910 avdd.n3125 avss -1.8e-19
C5911 avdd.n3126 avss -1.8e-19
C5912 avdd.n3127 avss -1.59e-19
C5913 avdd.n3128 avss 0.0192f
C5914 avdd.n3129 avss -3.07e-19
C5915 avdd.n3130 avss -6.46e-19
C5916 avdd.n3131 avss -5.82e-19
C5917 avdd.n3132 avss -7.52e-19
C5918 avdd.n3133 avss 0.00899f
C5919 avdd.n3134 avss -0.00113f
C5920 avdd.n3135 avss -8.47e-19
C5921 avdd.n3136 avss -3.39e-19
C5922 avdd.n3137 avss -3.18e-19
C5923 avdd.n3138 avss -2.01e-19
C5924 avdd.n3139 avss 0.0183f
C5925 avdd.n3140 avss 0.0154f
C5926 avdd.n3141 avss 0.0154f
C5927 avdd.n3142 avss 0.0191f
C5928 avdd.n3143 avss -1.8e-19
C5929 avdd.n3144 avss -1.8e-19
C5930 avdd.n3145 avss -1.8e-19
C5931 avdd.n3146 avss -2.44e-19
C5932 avdd.n3147 avss -1.8e-19
C5933 avdd.n3148 avss -1.8e-19
C5934 avdd.n3149 avss -1.38e-19
C5935 avdd.n3151 avss -3.49e-19
C5936 avdd.n3152 avss 0.0184f
C5937 avdd.n3153 avss 0.00873f
C5938 avdd.n3154 avss 0.0422f
C5939 avdd.n3155 avss 0.0197f
C5940 avdd.n3156 avss 0.0384f
C5941 avdd.n3157 avss -2.44e-19
C5942 avdd.n3158 avss -2.44e-19
C5943 avdd.n3159 avss -2.33e-19
C5944 avdd.n3160 avss -1.8e-19
C5945 avdd.n3161 avss -1.48e-19
C5946 avdd.n3162 avss -0.00173f
C5947 avdd.n3164 avss -1.27e-19
C5948 avdd.n3165 avss 0.0382f
C5949 avdd.n3166 avss -0.161f
C5950 avdd.n3167 avss -0.194f
C5951 avdd.n3168 avss -0.162f
C5952 avdd.n3169 avss -0.00357f
C5953 avdd.n3170 avss -0.00108f
C5954 avdd.n3171 avss -2.01e-19
C5955 avdd.n3172 avss -2.96e-19
C5956 avdd.n3173 avss -6.67e-19
C5957 avdd.n3174 avss -1.8e-19
C5958 avdd.n3175 avss 0.0411f
C5959 avdd.n3176 avss 0.0191f
C5960 avdd.n3177 avss -1.38e-19
C5961 avdd.n3178 avss -3.39e-19
C5962 avdd.n3179 avss 0.0111f
C5963 avdd.n3180 avss -2.22e-19
C5964 avdd.n3181 avss 0.0374f
C5965 avdd.n3182 avss 0.0112f
C5966 avdd.n3183 avss -1.8e-19
C5967 avdd.n3184 avss -1.8e-19
C5968 avdd.n3185 avss -0.00109f
C5969 avdd.n3186 avss -0.00126f
C5970 avdd.n3187 avss 0.0318f
C5971 avdd.n3188 avss -0.00139f
C5972 avdd.n3189 avss -2.22e-19
C5973 avdd.n3190 avss 0.0188f
C5974 avdd.n3191 avss -2.75e-19
C5975 avdd.n3192 avss -3.6e-19
C5976 avdd.n3193 avss -3.07e-19
C5977 avdd.n3194 avss -6.88e-19
C5978 avdd.n3195 avss 0.00725f
C5979 avdd.n3196 avss -0.00336f
C5980 avdd.n3197 avss -1.8e-19
C5981 avdd.n3198 avss -2.01e-19
C5982 avdd.n3199 avss -0.0866f
C5983 avdd.n3200 avss 0.0179f
C5984 avdd.n3201 avss 0.0442f
C5985 avdd.n3202 avss -3.39e-19
C5986 avdd.n3203 avss -2.75e-19
C5987 avdd.n3204 avss 0.0181f
C5988 avdd.n3205 avss 0.00821f
C5989 avdd.n3206 avss 0.00821f
C5990 avdd.n3207 avss -2.75e-19
C5991 avdd.n3208 avss -2.33e-19
C5992 avdd.n3209 avss -2.54e-19
C5993 avdd.n3210 avss -2.54e-19
C5994 avdd.n3211 avss -2.22e-19
C5995 avdd.n3212 avss -1.59e-19
C5996 avdd.n3213 avss 0.0298f
C5997 avdd.n3214 avss 0.0098f
C5998 avdd.n3215 avss -0.00158f
C5999 avdd.n3216 avss -8.47e-19
C6000 avdd.n3217 avss -4.23e-19
C6001 avdd.n3218 avss -3.39e-19
C6002 avdd.n3219 avss -2.33e-19
C6003 avdd.n3220 avss -1.16e-19
C6004 avdd.n3221 avss 0.0182f
C6005 avdd.n3222 avss 0.0148f
C6006 avdd.n3223 avss 0.00875f
C6007 avdd.n3225 avss -3.07e-19
C6008 avdd.n3226 avss 0.0192f
C6009 avdd.n3227 avss -1.59e-19
C6010 avdd.n3228 avss -1.8e-19
C6011 avdd.n3229 avss 0.00358f
C6012 avdd.n3230 avss -2.22e-19
C6013 avdd.n3231 avss -1.8e-19
C6014 avdd.n3232 avss -1.8e-19
C6015 avdd.n3233 avss 0.0183f
C6016 avdd.n3234 avss 0.0154f
C6017 avdd.n3235 avss 0.0154f
C6018 avdd.n3236 avss 0.0111f
C6019 avdd.n3237 avss 0.0111f
C6020 avdd.n3238 avss -1.8e-19
C6021 avdd.n3239 avss -8.15e-19
C6022 avdd.n3240 avss -1.48e-19
C6023 avdd.n3241 avss -3.39e-19
C6024 avdd.n3242 avss 0.00466f
C6025 avdd.n3243 avss -8.47e-19
C6026 avdd.n3244 avss -0.0014f
C6027 avdd.n3245 avss 0.0344f
C6028 avdd.n3246 avss -8.47e-19
C6029 avdd.n3247 avss 0.0348f
C6030 avdd.n3248 avss -5.19e-19
C6031 avdd.n3249 avss -3.07e-19
C6032 avdd.n3250 avss -3.28e-19
C6033 avdd.n3251 avss -1.8e-19
C6034 avdd.n3252 avss 0.0189f
C6035 avdd.n3253 avss -2.33e-19
C6036 avdd.n3254 avss 0.0022f
C6037 avdd.n3255 avss 0.0386f
C6038 avdd.n3256 avss -2.44e-19
C6039 avdd.n3257 avss 0.0184f
C6040 avdd.n3258 avss 0.00873f
C6041 avdd.n3259 avss 0.0168f
C6042 avdd.n3260 avss 0.0167f
C6043 avdd.n3261 avss -5.77e-19
C6044 avdd.n3262 avss -8.47e-19
C6045 avdd.n3263 avss -2.22e-19
C6046 avdd.n3264 avss 0.00875f
C6047 avdd.n3265 avss -2.54e-19
C6048 avdd.n3266 avss 0.0182f
C6049 avdd.n3267 avss 0.0111f
C6050 avdd.n3268 avss -1.59e-19
C6051 avdd.n3269 avss -3.39e-19
C6052 avdd.n3270 avss -1.59e-19
C6053 avdd.n3271 avss 3e-19
C6054 avdd.n3272 avss -2.54e-19
C6055 avdd.n3273 avss -1.8e-19
C6056 avdd.n3274 avss -1.8e-19
C6057 avdd.n3275 avss -1.16e-19
C6058 avdd.n3276 avss -2.33e-19
C6059 avdd.n3277 avss -3.39e-19
C6060 avdd.n3278 avss -8.47e-19
C6061 avdd.n3279 avss 0.0342f
C6062 avdd.n3280 avss 0.0049f
C6063 avdd.n3281 avss -8.47e-19
C6064 avdd.n3282 avss 0.0388f
C6065 avdd.n3283 avss -3.39e-19
C6066 avdd.n3284 avss -3.39e-19
C6067 avdd.n3285 avss -2.22e-19
C6068 avdd.n3286 avss -2.01e-19
C6069 avdd.n3287 avss -1.8e-19
C6070 avdd.n3288 avss -1.8e-19
C6071 avdd.n3289 avss -2.22e-19
C6072 avdd.n3290 avss 0.0111f
C6073 avdd.n3291 avss -1.8e-19
C6074 avdd.n3292 avss -2.96e-19
C6075 avdd.n3293 avss -2.44e-19
C6076 avdd.n3294 avss 0.0384f
C6077 avdd.n3295 avss -0.00113f
C6078 avdd.n3296 avss -0.00173f
C6079 avdd.n3297 avss -3.49e-19
C6080 avdd.n3299 avss 0.0382f
C6081 avdd.n3300 avss -3.18e-19
C6082 avdd.n3301 avss -8.47e-19
C6083 avdd.n3302 avss 0.03f
C6084 avdd.n3303 avss 0.00899f
C6085 avdd.n3304 avss -7.52e-19
C6086 avdd.n3305 avss -1.27e-19
C6087 avdd.n3306 avss -2.44e-19
C6088 avdd.n3307 avss -1.8e-19
C6089 avdd.n3308 avss -1.8e-19
C6090 avdd.n3309 avss -1.38e-19
C6091 avdd.n3310 avss -1.38e-19
C6092 avdd.n3311 avss 0.0184f
C6093 avdd.n3312 avss 0.00873f
C6094 avdd.n3313 avss 0.0422f
C6095 avdd.n3314 avss -2.33e-19
C6096 avdd.n3315 avss 0.0197f
C6097 avdd.n3316 avss -2.44e-19
C6098 avdd.n3317 avss -2.44e-19
C6099 avdd.n3318 avss -2.33e-19
C6100 avdd.n3319 avss -1.48e-19
C6101 avdd.n3320 avss -1.8e-19
C6102 avdd.n3321 avss 0.019f
C6103 avdd.n3322 avss 0.00335f
C6104 avdd.n3323 avss 0.0265f
C6105 avdd.n3324 avss 0.00778f
C6106 avdd.n3325 avss -0.00512f
C6107 avdd.n3326 avss -1.8e-19
C6108 avdd.n3327 avss -1.8e-19
C6109 avdd.n3328 avss 0.0191f
C6110 avdd.n3329 avss 0.0154f
C6111 avdd.n3330 avss 0.0154f
C6112 avdd.n3331 avss 0.0183f
C6113 avdd.n3332 avss -1.8e-19
C6114 avdd.n3333 avss -1.8e-19
C6115 avdd.n3334 avss -5.82e-19
C6116 avdd.n3335 avss -6.46e-19
C6117 avdd.n3336 avss -3.07e-19
C6118 avdd.n3337 avss 0.0192f
C6119 avdd.n3338 avss 0.00875f
C6120 avdd.n3339 avss 0.0148f
C6121 avdd.n3340 avss 0.0111f
C6122 avdd.n3341 avss -2.22e-19
C6123 avdd.n3342 avss 0.0192f
C6124 avdd.n3343 avss -4.76e-19
C6125 avdd.n3344 avss -0.00128f
C6126 avdd.n3345 avss 0.0346f
C6127 avdd.n3346 avss 0.00378f
C6128 avdd.n3347 avss -8.47e-19
C6129 avdd.n3348 avss 0.0398f
C6130 avdd.n3349 avss -3.07e-19
C6131 avdd.n3350 avss 0.0181f
C6132 avdd.n3351 avss -3.6e-19
C6133 avdd.n3352 avss -2.01e-19
C6134 avdd.n3353 avss -3.28e-19
C6135 avdd.n3354 avss -8.26e-19
C6136 avdd.n3355 avss -6.46e-19
C6137 avdd.n3356 avss -0.00137f
C6138 avdd.n3357 avss -0.0013f
C6139 avdd.n3358 avss 0.00357f
C6140 avdd.n3359 avss -8.47e-19
C6141 avdd.n3360 avss -3.39e-19
C6142 avdd.n3361 avss -1.27e-19
C6143 avdd.n3362 avss -2.44e-19
C6144 avdd.n3363 avss 0.019f
C6145 avdd.n3364 avss 0.0148f
C6146 avdd.n3365 avss 0.00873f
C6147 avdd.n3366 avss 0.0184f
C6148 avdd.n3367 avss -3.49e-19
C6149 avdd.n3368 avss -1.38e-19
C6150 avdd.n3369 avss -1.8e-19
C6151 avdd.n3370 avss -1.8e-19
C6152 avdd.n3371 avss -2.44e-19
C6153 avdd.n3372 avss -1.8e-19
C6154 avdd.n3373 avss -1.8e-19
C6155 avdd.n3374 avss -5.61e-19
C6156 avdd.n3375 avss -3.39e-19
C6157 avdd.n3376 avss -6.35e-19
C6158 avdd.n3377 avss -0.00121f
C6159 avdd.n3378 avss -0.00122f
C6160 avdd.n3379 avss -0.00173f
C6161 avdd.n3380 avss -9.75e-19
C6162 avdd.n3381 avss 0.0382f
C6163 avdd.n3382 avss -0.196f
C6164 avdd.n3383 avss -0.162f
C6165 avdd.n3384 avss -0.00357f
C6166 avdd.n3385 avss -0.00108f
C6167 avdd.n3386 avss -2.01e-19
C6168 avdd.n3387 avss -2.96e-19
C6169 avdd.n3388 avss -6.67e-19
C6170 avdd.n3389 avss -1.8e-19
C6171 avdd.n3390 avss 0.0411f
C6172 avdd.n3391 avss 0.0191f
C6173 avdd.n3392 avss -1.38e-19
C6174 avdd.n3393 avss -3.39e-19
C6175 avdd.n3394 avss 0.0111f
C6176 avdd.n3395 avss -2.22e-19
C6177 avdd.n3396 avss 0.0374f
C6178 avdd.n3397 avss 0.0112f
C6179 avdd.n3398 avss -1.8e-19
C6180 avdd.n3399 avss -1.8e-19
C6181 avdd.n3400 avss -0.00109f
C6182 avdd.n3401 avss -0.00126f
C6183 avdd.n3402 avss 0.0318f
C6184 avdd.n3403 avss -0.00139f
C6185 avdd.n3404 avss -2.22e-19
C6186 avdd.n3405 avss 0.0188f
C6187 avdd.n3406 avss -2.75e-19
C6188 avdd.n3407 avss -3.6e-19
C6189 avdd.n3408 avss -3.07e-19
C6190 avdd.n3409 avss -6.88e-19
C6191 avdd.n3410 avss 0.00725f
C6192 avdd.n3411 avss -0.00336f
C6193 avdd.n3412 avss -1.8e-19
C6194 avdd.n3413 avss -2.01e-19
C6195 avdd.n3414 avss -0.0866f
C6196 avdd.n3415 avss 0.0179f
C6197 avdd.n3416 avss 0.0442f
C6198 avdd.n3417 avss -3.39e-19
C6199 avdd.n3418 avss -2.75e-19
C6200 avdd.n3419 avss 0.0181f
C6201 avdd.n3420 avss 0.00821f
C6202 avdd.n3421 avss 0.00821f
C6203 avdd.n3422 avss -2.75e-19
C6204 avdd.n3423 avss -2.33e-19
C6205 avdd.n3424 avss -2.54e-19
C6206 avdd.n3425 avss -2.54e-19
C6207 avdd.n3426 avss -2.22e-19
C6208 avdd.n3427 avss -1.59e-19
C6209 avdd.n3428 avss 0.0298f
C6210 avdd.n3429 avss 0.0098f
C6211 avdd.n3430 avss -0.00158f
C6212 avdd.n3431 avss -8.47e-19
C6213 avdd.n3432 avss -4.23e-19
C6214 avdd.n3433 avss -3.39e-19
C6215 avdd.n3434 avss -2.33e-19
C6216 avdd.n3435 avss -1.16e-19
C6217 avdd.n3436 avss 0.0182f
C6218 avdd.n3437 avss 0.0148f
C6219 avdd.n3438 avss 0.00875f
C6220 avdd.n3440 avss -3.07e-19
C6221 avdd.n3441 avss 0.0192f
C6222 avdd.n3442 avss -1.59e-19
C6223 avdd.n3443 avss -1.8e-19
C6224 avdd.n3444 avss 0.00358f
C6225 avdd.n3445 avss -2.22e-19
C6226 avdd.n3446 avss -1.8e-19
C6227 avdd.n3447 avss -1.8e-19
C6228 avdd.n3448 avss 0.0183f
C6229 avdd.n3449 avss 0.0154f
C6230 avdd.n3450 avss 0.0154f
C6231 avdd.n3451 avss 0.0111f
C6232 avdd.n3452 avss 0.0111f
C6233 avdd.n3453 avss -1.8e-19
C6234 avdd.n3454 avss -8.15e-19
C6235 avdd.n3455 avss -1.48e-19
C6236 avdd.n3456 avss -3.39e-19
C6237 avdd.n3457 avss 0.00466f
C6238 avdd.n3458 avss -8.47e-19
C6239 avdd.n3459 avss -0.0014f
C6240 avdd.n3460 avss 0.0344f
C6241 avdd.n3461 avss -8.47e-19
C6242 avdd.n3462 avss 0.0348f
C6243 avdd.n3463 avss -5.19e-19
C6244 avdd.n3464 avss -3.07e-19
C6245 avdd.n3465 avss -3.28e-19
C6246 avdd.n3466 avss -1.8e-19
C6247 avdd.n3467 avss 0.0189f
C6248 avdd.n3468 avss -2.33e-19
C6249 avdd.n3469 avss 0.0022f
C6250 avdd.n3470 avss 0.0386f
C6251 avdd.n3471 avss -2.44e-19
C6252 avdd.n3472 avss 0.0184f
C6253 avdd.n3473 avss 0.00873f
C6254 avdd.n3474 avss 0.0168f
C6255 avdd.n3475 avss 0.0167f
C6256 avdd.n3476 avss -5.77e-19
C6257 avdd.n3477 avss -8.47e-19
C6258 avdd.n3478 avss -2.22e-19
C6259 avdd.n3479 avss 0.00875f
C6260 avdd.n3480 avss -2.54e-19
C6261 avdd.n3481 avss 0.0182f
C6262 avdd.n3482 avss 0.0111f
C6263 avdd.n3483 avss -1.59e-19
C6264 avdd.n3484 avss -3.39e-19
C6265 avdd.n3485 avss -1.59e-19
C6266 avdd.n3486 avss 3e-19
C6267 avdd.n3487 avss -2.54e-19
C6268 avdd.n3488 avss -1.8e-19
C6269 avdd.n3489 avss -1.8e-19
C6270 avdd.n3490 avss -1.16e-19
C6271 avdd.n3491 avss -2.33e-19
C6272 avdd.n3492 avss -3.39e-19
C6273 avdd.n3493 avss -8.47e-19
C6274 avdd.n3494 avss 0.0342f
C6275 avdd.n3495 avss 0.0049f
C6276 avdd.n3496 avss -8.47e-19
C6277 avdd.n3497 avss 0.0388f
C6278 avdd.n3498 avss -3.39e-19
C6279 avdd.n3499 avss -3.39e-19
C6280 avdd.n3500 avss -2.22e-19
C6281 avdd.n3501 avss -2.01e-19
C6282 avdd.n3502 avss -1.8e-19
C6283 avdd.n3503 avss -1.8e-19
C6284 avdd.n3504 avss -2.22e-19
C6285 avdd.n3505 avss 0.0111f
C6286 avdd.n3506 avss -1.8e-19
C6287 avdd.n3507 avss -2.96e-19
C6288 avdd.n3508 avss -2.44e-19
C6289 avdd.n3509 avss 0.0384f
C6290 avdd.n3510 avss -0.00113f
C6291 avdd.n3511 avss -0.00173f
C6292 avdd.n3512 avss -3.49e-19
C6293 avdd.n3514 avss 0.0382f
C6294 avdd.n3515 avss -3.18e-19
C6295 avdd.n3516 avss -8.47e-19
C6296 avdd.n3517 avss 0.03f
C6297 avdd.n3518 avss 0.00899f
C6298 avdd.n3519 avss -7.52e-19
C6299 avdd.n3520 avss -1.27e-19
C6300 avdd.n3521 avss -2.44e-19
C6301 avdd.n3522 avss -1.8e-19
C6302 avdd.n3523 avss -1.8e-19
C6303 avdd.n3524 avss -1.38e-19
C6304 avdd.n3525 avss -1.38e-19
C6305 avdd.n3526 avss 0.0184f
C6306 avdd.n3527 avss 0.00873f
C6307 avdd.n3528 avss 0.0422f
C6308 avdd.n3529 avss -2.33e-19
C6309 avdd.n3530 avss 0.0197f
C6310 avdd.n3531 avss -2.44e-19
C6311 avdd.n3532 avss -2.44e-19
C6312 avdd.n3533 avss -2.33e-19
C6313 avdd.n3534 avss -1.48e-19
C6314 avdd.n3535 avss -1.8e-19
C6315 avdd.n3536 avss 0.019f
C6316 avdd.n3537 avss 0.00335f
C6317 avdd.n3538 avss 0.0265f
C6318 avdd.n3539 avss 0.00778f
C6319 avdd.n3540 avss -0.00512f
C6320 avdd.n3541 avss -1.8e-19
C6321 avdd.n3542 avss -1.8e-19
C6322 avdd.n3543 avss 0.0191f
C6323 avdd.n3544 avss 0.0154f
C6324 avdd.n3545 avss 0.0154f
C6325 avdd.n3546 avss 0.0183f
C6326 avdd.n3547 avss -1.8e-19
C6327 avdd.n3548 avss -1.8e-19
C6328 avdd.n3549 avss -5.82e-19
C6329 avdd.n3550 avss -6.46e-19
C6330 avdd.n3551 avss -3.07e-19
C6331 avdd.n3552 avss 0.0192f
C6332 avdd.n3553 avss 0.00875f
C6333 avdd.n3554 avss 0.0148f
C6334 avdd.n3555 avss 0.0111f
C6335 avdd.n3556 avss -2.22e-19
C6336 avdd.n3557 avss 0.0192f
C6337 avdd.n3558 avss -4.76e-19
C6338 avdd.n3559 avss -0.00128f
C6339 avdd.n3560 avss 0.0346f
C6340 avdd.n3561 avss 0.00378f
C6341 avdd.n3562 avss -8.47e-19
C6342 avdd.n3563 avss 0.0398f
C6343 avdd.n3564 avss -3.07e-19
C6344 avdd.n3565 avss 0.0181f
C6345 avdd.n3566 avss -3.6e-19
C6346 avdd.n3567 avss -2.01e-19
C6347 avdd.n3568 avss -3.28e-19
C6348 avdd.n3569 avss -8.26e-19
C6349 avdd.n3570 avss -6.46e-19
C6350 avdd.n3571 avss -0.00137f
C6351 avdd.n3572 avss -0.0013f
C6352 avdd.n3573 avss 0.00357f
C6353 avdd.n3574 avss -8.47e-19
C6354 avdd.n3575 avss -3.39e-19
C6355 avdd.n3576 avss -1.27e-19
C6356 avdd.n3577 avss -2.44e-19
C6357 avdd.n3578 avss 0.019f
C6358 avdd.n3579 avss 0.0148f
C6359 avdd.n3580 avss 0.00873f
C6360 avdd.n3581 avss 0.0184f
C6361 avdd.n3582 avss -3.49e-19
C6362 avdd.n3583 avss -1.38e-19
C6363 avdd.n3584 avss -1.8e-19
C6364 avdd.n3585 avss -1.8e-19
C6365 avdd.n3586 avss -2.44e-19
C6366 avdd.n3587 avss -1.8e-19
C6367 avdd.n3588 avss -1.8e-19
C6368 avdd.n3589 avss -5.61e-19
C6369 avdd.n3590 avss -3.39e-19
C6370 avdd.n3591 avss -6.35e-19
C6371 avdd.n3592 avss -0.00121f
C6372 avdd.n3593 avss -0.00122f
C6373 avdd.n3594 avss -0.00173f
C6374 avdd.n3595 avss -9.75e-19
C6375 avdd.n3596 avss 0.0382f
C6376 avdd.n3597 avss -0.196f
C6377 avdd.n3598 avss -0.162f
C6378 avdd.n3599 avss -0.00357f
C6379 avdd.n3600 avss -0.00108f
C6380 avdd.n3601 avss -2.01e-19
C6381 avdd.n3602 avss -2.96e-19
C6382 avdd.n3603 avss -6.67e-19
C6383 avdd.n3604 avss -1.8e-19
C6384 avdd.n3605 avss 0.0411f
C6385 avdd.n3606 avss 0.0191f
C6386 avdd.n3607 avss -1.38e-19
C6387 avdd.n3608 avss -3.39e-19
C6388 avdd.n3609 avss 0.0111f
C6389 avdd.n3610 avss -2.22e-19
C6390 avdd.n3611 avss 0.0374f
C6391 avdd.n3612 avss 0.0112f
C6392 avdd.n3613 avss -1.8e-19
C6393 avdd.n3614 avss -1.8e-19
C6394 avdd.n3615 avss -0.00109f
C6395 avdd.n3616 avss -0.00126f
C6396 avdd.n3617 avss 0.0318f
C6397 avdd.n3618 avss -0.00139f
C6398 avdd.n3619 avss -2.22e-19
C6399 avdd.n3620 avss 0.0188f
C6400 avdd.n3621 avss -2.75e-19
C6401 avdd.n3622 avss -3.6e-19
C6402 avdd.n3623 avss -3.07e-19
C6403 avdd.n3624 avss -6.88e-19
C6404 avdd.n3625 avss 0.00725f
C6405 avdd.n3626 avss -0.00336f
C6406 avdd.n3627 avss -1.8e-19
C6407 avdd.n3628 avss -2.01e-19
C6408 avdd.n3629 avss -0.0866f
C6409 avdd.n3630 avss 0.0179f
C6410 avdd.n3631 avss 0.0442f
C6411 avdd.n3632 avss -3.39e-19
C6412 avdd.n3633 avss -2.75e-19
C6413 avdd.n3634 avss 0.0181f
C6414 avdd.n3635 avss 0.00821f
C6415 avdd.n3636 avss 0.00821f
C6416 avdd.n3637 avss -2.75e-19
C6417 avdd.n3638 avss -2.33e-19
C6418 avdd.n3639 avss -2.54e-19
C6419 avdd.n3640 avss -2.54e-19
C6420 avdd.n3641 avss -2.22e-19
C6421 avdd.n3642 avss -1.59e-19
C6422 avdd.n3643 avss 0.0298f
C6423 avdd.n3644 avss 0.0098f
C6424 avdd.n3645 avss -0.00158f
C6425 avdd.n3646 avss -8.47e-19
C6426 avdd.n3647 avss -4.23e-19
C6427 avdd.n3648 avss -3.39e-19
C6428 avdd.n3649 avss -2.33e-19
C6429 avdd.n3650 avss -1.16e-19
C6430 avdd.n3651 avss 0.0182f
C6431 avdd.n3652 avss 0.0148f
C6432 avdd.n3653 avss 0.00875f
C6433 avdd.n3655 avss -3.07e-19
C6434 avdd.n3656 avss 0.0192f
C6435 avdd.n3657 avss -1.59e-19
C6436 avdd.n3658 avss -1.8e-19
C6437 avdd.n3659 avss 0.00358f
C6438 avdd.n3660 avss -2.22e-19
C6439 avdd.n3661 avss -1.8e-19
C6440 avdd.n3662 avss -1.8e-19
C6441 avdd.n3663 avss 0.0183f
C6442 avdd.n3664 avss 0.0154f
C6443 avdd.n3665 avss 0.0154f
C6444 avdd.n3666 avss 0.0111f
C6445 avdd.n3667 avss 0.0111f
C6446 avdd.n3668 avss -1.8e-19
C6447 avdd.n3669 avss -8.15e-19
C6448 avdd.n3670 avss -1.48e-19
C6449 avdd.n3671 avss -3.39e-19
C6450 avdd.n3672 avss 0.00466f
C6451 avdd.n3673 avss -8.47e-19
C6452 avdd.n3674 avss -0.0014f
C6453 avdd.n3675 avss 0.0344f
C6454 avdd.n3676 avss -8.47e-19
C6455 avdd.n3677 avss 0.0348f
C6456 avdd.n3678 avss -5.19e-19
C6457 avdd.n3679 avss -3.07e-19
C6458 avdd.n3680 avss -3.28e-19
C6459 avdd.n3681 avss -1.8e-19
C6460 avdd.n3682 avss 0.0189f
C6461 avdd.n3683 avss -2.33e-19
C6462 avdd.n3684 avss 0.0022f
C6463 avdd.n3685 avss 0.0386f
C6464 avdd.n3686 avss -2.44e-19
C6465 avdd.n3687 avss 0.0184f
C6466 avdd.n3688 avss 0.00873f
C6467 avdd.n3689 avss 0.0168f
C6468 avdd.n3690 avss 0.0167f
C6469 avdd.n3691 avss -5.77e-19
C6470 avdd.n3692 avss -8.47e-19
C6471 avdd.n3693 avss -2.22e-19
C6472 avdd.n3694 avss 0.00875f
C6473 avdd.n3695 avss -2.54e-19
C6474 avdd.n3696 avss 0.0182f
C6475 avdd.n3697 avss 0.0111f
C6476 avdd.n3698 avss -1.59e-19
C6477 avdd.n3699 avss -3.39e-19
C6478 avdd.n3700 avss -1.59e-19
C6479 avdd.n3701 avss 3e-19
C6480 avdd.n3702 avss -2.54e-19
C6481 avdd.n3703 avss -1.8e-19
C6482 avdd.n3704 avss -1.8e-19
C6483 avdd.n3705 avss -1.16e-19
C6484 avdd.n3706 avss -2.33e-19
C6485 avdd.n3707 avss -3.39e-19
C6486 avdd.n3708 avss -8.47e-19
C6487 avdd.n3709 avss 0.0342f
C6488 avdd.n3710 avss 0.0049f
C6489 avdd.n3711 avss -8.47e-19
C6490 avdd.n3712 avss 0.0388f
C6491 avdd.n3713 avss -3.39e-19
C6492 avdd.n3714 avss -3.39e-19
C6493 avdd.n3715 avss -2.22e-19
C6494 avdd.n3716 avss -2.01e-19
C6495 avdd.n3717 avss -1.8e-19
C6496 avdd.n3718 avss -1.8e-19
C6497 avdd.n3719 avss -2.22e-19
C6498 avdd.n3720 avss 0.0111f
C6499 avdd.n3721 avss -1.8e-19
C6500 avdd.n3722 avss -2.96e-19
C6501 avdd.n3723 avss -2.44e-19
C6502 avdd.n3724 avss 0.0384f
C6503 avdd.n3725 avss -0.00113f
C6504 avdd.n3726 avss -0.00173f
C6505 avdd.n3727 avss -3.49e-19
C6506 avdd.n3729 avss 0.0382f
C6507 avdd.n3730 avss -3.18e-19
C6508 avdd.n3731 avss -8.47e-19
C6509 avdd.n3732 avss 0.03f
C6510 avdd.n3733 avss 0.00899f
C6511 avdd.n3734 avss -7.52e-19
C6512 avdd.n3735 avss -1.27e-19
C6513 avdd.n3736 avss -2.44e-19
C6514 avdd.n3737 avss -1.8e-19
C6515 avdd.n3738 avss -1.8e-19
C6516 avdd.n3739 avss -1.38e-19
C6517 avdd.n3740 avss -1.38e-19
C6518 avdd.n3741 avss 0.0184f
C6519 avdd.n3742 avss 0.00873f
C6520 avdd.n3743 avss 0.0422f
C6521 avdd.n3744 avss -2.33e-19
C6522 avdd.n3745 avss 0.0197f
C6523 avdd.n3746 avss -2.44e-19
C6524 avdd.n3747 avss -2.44e-19
C6525 avdd.n3748 avss -2.33e-19
C6526 avdd.n3749 avss -1.48e-19
C6527 avdd.n3750 avss -1.8e-19
C6528 avdd.n3751 avss 0.019f
C6529 avdd.n3752 avss 0.00335f
C6530 avdd.n3753 avss 0.0265f
C6531 avdd.n3754 avss 0.00778f
C6532 avdd.n3755 avss -0.00512f
C6533 avdd.n3756 avss -1.8e-19
C6534 avdd.n3757 avss -1.8e-19
C6535 avdd.n3758 avss 0.0191f
C6536 avdd.n3759 avss 0.0154f
C6537 avdd.n3760 avss 0.0154f
C6538 avdd.n3761 avss 0.0183f
C6539 avdd.n3762 avss -1.8e-19
C6540 avdd.n3763 avss -1.8e-19
C6541 avdd.n3764 avss -5.82e-19
C6542 avdd.n3765 avss -6.46e-19
C6543 avdd.n3766 avss -3.07e-19
C6544 avdd.n3767 avss 0.0192f
C6545 avdd.n3768 avss 0.00875f
C6546 avdd.n3769 avss 0.0148f
C6547 avdd.n3770 avss 0.0111f
C6548 avdd.n3771 avss -2.22e-19
C6549 avdd.n3772 avss 0.0192f
C6550 avdd.n3773 avss -4.76e-19
C6551 avdd.n3774 avss -0.00128f
C6552 avdd.n3775 avss 0.0346f
C6553 avdd.n3776 avss 0.00378f
C6554 avdd.n3777 avss -8.47e-19
C6555 avdd.n3778 avss 0.0398f
C6556 avdd.n3779 avss -3.07e-19
C6557 avdd.n3780 avss 0.0181f
C6558 avdd.n3781 avss -3.6e-19
C6559 avdd.n3782 avss -2.01e-19
C6560 avdd.n3783 avss -3.28e-19
C6561 avdd.n3784 avss -8.26e-19
C6562 avdd.n3785 avss -6.46e-19
C6563 avdd.n3786 avss -0.00137f
C6564 avdd.n3787 avss -0.0013f
C6565 avdd.n3788 avss 0.00357f
C6566 avdd.n3789 avss -8.47e-19
C6567 avdd.n3790 avss -3.39e-19
C6568 avdd.n3791 avss -1.27e-19
C6569 avdd.n3792 avss -2.44e-19
C6570 avdd.n3793 avss 0.019f
C6571 avdd.n3794 avss 0.0148f
C6572 avdd.n3795 avss 0.00873f
C6573 avdd.n3796 avss 0.0184f
C6574 avdd.n3797 avss -3.49e-19
C6575 avdd.n3798 avss -1.38e-19
C6576 avdd.n3799 avss -1.8e-19
C6577 avdd.n3800 avss -1.8e-19
C6578 avdd.n3801 avss -2.44e-19
C6579 avdd.n3802 avss -1.8e-19
C6580 avdd.n3803 avss -1.8e-19
C6581 avdd.n3804 avss -5.61e-19
C6582 avdd.n3805 avss -3.39e-19
C6583 avdd.n3806 avss -6.35e-19
C6584 avdd.n3807 avss -0.00121f
C6585 avdd.n3808 avss -0.00122f
C6586 avdd.n3809 avss -0.00173f
C6587 avdd.n3810 avss -9.75e-19
C6588 avdd.n3811 avss 0.0382f
C6589 avdd.n3812 avss -0.196f
C6590 avdd.n3813 avss -0.162f
C6591 avdd.n3814 avss -0.00357f
C6592 avdd.n3815 avss -0.00108f
C6593 avdd.n3816 avss -2.01e-19
C6594 avdd.n3817 avss -2.96e-19
C6595 avdd.n3818 avss -6.67e-19
C6596 avdd.n3819 avss -1.8e-19
C6597 avdd.n3820 avss 0.0411f
C6598 avdd.n3821 avss 0.0191f
C6599 avdd.n3822 avss -1.38e-19
C6600 avdd.n3823 avss -3.39e-19
C6601 avdd.n3824 avss 0.0111f
C6602 avdd.n3825 avss -2.22e-19
C6603 avdd.n3826 avss 0.0374f
C6604 avdd.n3827 avss 0.0112f
C6605 avdd.n3828 avss -1.8e-19
C6606 avdd.n3829 avss -1.8e-19
C6607 avdd.n3830 avss -0.00109f
C6608 avdd.n3831 avss -0.00126f
C6609 avdd.n3832 avss 0.0318f
C6610 avdd.n3833 avss -0.00139f
C6611 avdd.n3834 avss -2.22e-19
C6612 avdd.n3835 avss 0.0188f
C6613 avdd.n3836 avss -2.75e-19
C6614 avdd.n3837 avss -3.6e-19
C6615 avdd.n3838 avss -3.07e-19
C6616 avdd.n3839 avss -6.88e-19
C6617 avdd.n3840 avss 0.00725f
C6618 avdd.n3841 avss -0.00336f
C6619 avdd.n3842 avss -1.8e-19
C6620 avdd.n3843 avss -2.01e-19
C6621 avdd.n3844 avss -0.0866f
C6622 avdd.n3845 avss 0.0179f
C6623 avdd.n3846 avss 0.0442f
C6624 avdd.n3847 avss -3.39e-19
C6625 avdd.n3848 avss -2.75e-19
C6626 avdd.n3849 avss 0.0181f
C6627 avdd.n3850 avss 0.00821f
C6628 avdd.n3851 avss 0.00821f
C6629 avdd.n3852 avss -2.75e-19
C6630 avdd.n3853 avss -2.33e-19
C6631 avdd.n3854 avss -2.54e-19
C6632 avdd.n3855 avss -2.54e-19
C6633 avdd.n3856 avss -2.22e-19
C6634 avdd.n3857 avss -1.59e-19
C6635 avdd.n3858 avss 0.0298f
C6636 avdd.n3859 avss 0.0098f
C6637 avdd.n3860 avss -0.00158f
C6638 avdd.n3861 avss -8.47e-19
C6639 avdd.n3862 avss -4.23e-19
C6640 avdd.n3863 avss -3.39e-19
C6641 avdd.n3864 avss -2.33e-19
C6642 avdd.n3865 avss -1.16e-19
C6643 avdd.n3866 avss 0.0182f
C6644 avdd.n3867 avss 0.0148f
C6645 avdd.n3868 avss 0.00875f
C6646 avdd.n3870 avss -3.07e-19
C6647 avdd.n3871 avss 0.0192f
C6648 avdd.n3872 avss -1.59e-19
C6649 avdd.n3873 avss -1.8e-19
C6650 avdd.n3874 avss 0.00358f
C6651 avdd.n3875 avss -2.22e-19
C6652 avdd.n3876 avss -1.8e-19
C6653 avdd.n3877 avss -1.8e-19
C6654 avdd.n3878 avss 0.0183f
C6655 avdd.n3879 avss 0.0154f
C6656 avdd.n3880 avss 0.0154f
C6657 avdd.n3881 avss 0.0111f
C6658 avdd.n3882 avss 0.0111f
C6659 avdd.n3883 avss -1.8e-19
C6660 avdd.n3884 avss -8.15e-19
C6661 avdd.n3885 avss -1.48e-19
C6662 avdd.n3886 avss -3.39e-19
C6663 avdd.n3887 avss 0.00466f
C6664 avdd.n3888 avss -8.47e-19
C6665 avdd.n3889 avss -0.0014f
C6666 avdd.n3890 avss 0.0344f
C6667 avdd.n3891 avss -8.47e-19
C6668 avdd.n3892 avss 0.0348f
C6669 avdd.n3893 avss -5.19e-19
C6670 avdd.n3894 avss -3.07e-19
C6671 avdd.n3895 avss -3.28e-19
C6672 avdd.n3896 avss -1.8e-19
C6673 avdd.n3897 avss 0.0189f
C6674 avdd.n3898 avss -2.33e-19
C6675 avdd.n3899 avss 0.0022f
C6676 avdd.n3900 avss 0.0386f
C6677 avdd.n3901 avss -2.44e-19
C6678 avdd.n3902 avss 0.0184f
C6679 avdd.n3903 avss 0.00873f
C6680 avdd.n3904 avss 0.0168f
C6681 avdd.n3905 avss 0.0167f
C6682 avdd.n3906 avss -5.77e-19
C6683 avdd.n3907 avss -8.47e-19
C6684 avdd.n3908 avss -2.22e-19
C6685 avdd.n3909 avss 0.00875f
C6686 avdd.n3910 avss -2.54e-19
C6687 avdd.n3911 avss 0.0182f
C6688 avdd.n3912 avss 0.0111f
C6689 avdd.n3913 avss -1.59e-19
C6690 avdd.n3914 avss -3.39e-19
C6691 avdd.n3915 avss -1.59e-19
C6692 avdd.n3916 avss 3e-19
C6693 avdd.n3917 avss -2.54e-19
C6694 avdd.n3918 avss -1.8e-19
C6695 avdd.n3919 avss -1.8e-19
C6696 avdd.n3920 avss -1.16e-19
C6697 avdd.n3921 avss -2.33e-19
C6698 avdd.n3922 avss -3.39e-19
C6699 avdd.n3923 avss -8.47e-19
C6700 avdd.n3924 avss 0.0342f
C6701 avdd.n3925 avss 0.0049f
C6702 avdd.n3926 avss -8.47e-19
C6703 avdd.n3927 avss 0.0388f
C6704 avdd.n3928 avss -3.39e-19
C6705 avdd.n3929 avss -3.39e-19
C6706 avdd.n3930 avss -2.22e-19
C6707 avdd.n3931 avss -2.01e-19
C6708 avdd.n3932 avss -1.8e-19
C6709 avdd.n3933 avss -1.8e-19
C6710 avdd.n3934 avss -2.22e-19
C6711 avdd.n3935 avss 0.0111f
C6712 avdd.n3936 avss -1.8e-19
C6713 avdd.n3937 avss -2.96e-19
C6714 avdd.n3938 avss -2.44e-19
C6715 avdd.n3939 avss 0.0384f
C6716 avdd.n3940 avss -0.00113f
C6717 avdd.n3941 avss -0.00173f
C6718 avdd.n3942 avss -3.49e-19
C6719 avdd.n3944 avss 0.0382f
C6720 avdd.n3945 avss -3.18e-19
C6721 avdd.n3946 avss -8.47e-19
C6722 avdd.n3947 avss 0.03f
C6723 avdd.n3948 avss 0.00899f
C6724 avdd.n3949 avss -7.52e-19
C6725 avdd.n3950 avss -1.27e-19
C6726 avdd.n3951 avss -2.44e-19
C6727 avdd.n3952 avss -1.8e-19
C6728 avdd.n3953 avss -1.8e-19
C6729 avdd.n3954 avss -1.38e-19
C6730 avdd.n3955 avss -1.38e-19
C6731 avdd.n3956 avss 0.0184f
C6732 avdd.n3957 avss 0.00873f
C6733 avdd.n3958 avss 0.0422f
C6734 avdd.n3959 avss -2.33e-19
C6735 avdd.n3960 avss 0.0197f
C6736 avdd.n3961 avss -2.44e-19
C6737 avdd.n3962 avss -2.44e-19
C6738 avdd.n3963 avss -2.33e-19
C6739 avdd.n3964 avss -1.48e-19
C6740 avdd.n3965 avss -1.8e-19
C6741 avdd.n3966 avss 0.019f
C6742 avdd.n3967 avss 0.00335f
C6743 avdd.n3968 avss 0.0265f
C6744 avdd.n3969 avss 0.00778f
C6745 avdd.n3970 avss -0.00512f
C6746 avdd.n3971 avss -1.8e-19
C6747 avdd.n3972 avss -1.8e-19
C6748 avdd.n3973 avss 0.0191f
C6749 avdd.n3974 avss 0.0154f
C6750 avdd.n3975 avss 0.0154f
C6751 avdd.n3976 avss 0.0183f
C6752 avdd.n3977 avss -1.8e-19
C6753 avdd.n3978 avss -1.8e-19
C6754 avdd.n3979 avss -5.82e-19
C6755 avdd.n3980 avss -6.46e-19
C6756 avdd.n3981 avss -3.07e-19
C6757 avdd.n3982 avss 0.0192f
C6758 avdd.n3983 avss 0.00875f
C6759 avdd.n3984 avss 0.0148f
C6760 avdd.n3985 avss 0.0111f
C6761 avdd.n3986 avss -2.22e-19
C6762 avdd.n3987 avss 0.0192f
C6763 avdd.n3988 avss -4.76e-19
C6764 avdd.n3989 avss -0.00128f
C6765 avdd.n3990 avss 0.0346f
C6766 avdd.n3991 avss 0.00378f
C6767 avdd.n3992 avss -8.47e-19
C6768 avdd.n3993 avss 0.0398f
C6769 avdd.n3994 avss -3.07e-19
C6770 avdd.n3995 avss 0.0181f
C6771 avdd.n3996 avss -3.6e-19
C6772 avdd.n3997 avss -2.01e-19
C6773 avdd.n3998 avss -3.28e-19
C6774 avdd.n3999 avss -8.26e-19
C6775 avdd.n4000 avss -6.46e-19
C6776 avdd.n4001 avss -0.00137f
C6777 avdd.n4002 avss -0.0013f
C6778 avdd.n4003 avss 0.00357f
C6779 avdd.n4004 avss -8.47e-19
C6780 avdd.n4005 avss -3.39e-19
C6781 avdd.n4006 avss -1.27e-19
C6782 avdd.n4007 avss -2.44e-19
C6783 avdd.n4008 avss 0.019f
C6784 avdd.n4009 avss 0.0148f
C6785 avdd.n4010 avss 0.00873f
C6786 avdd.n4011 avss 0.0184f
C6787 avdd.n4012 avss -3.49e-19
C6788 avdd.n4013 avss -1.38e-19
C6789 avdd.n4014 avss -1.8e-19
C6790 avdd.n4015 avss -1.8e-19
C6791 avdd.n4016 avss -2.44e-19
C6792 avdd.n4017 avss -1.8e-19
C6793 avdd.n4018 avss -1.8e-19
C6794 avdd.n4019 avss -5.61e-19
C6795 avdd.n4020 avss -3.39e-19
C6796 avdd.n4021 avss -6.35e-19
C6797 avdd.n4022 avss -0.00121f
C6798 avdd.n4023 avss -0.00122f
C6799 avdd.n4024 avss -0.00173f
C6800 avdd.n4025 avss -9.75e-19
C6801 avdd.n4026 avss 0.0382f
C6802 avdd.n4027 avss -0.196f
C6803 avdd.n4028 avss -0.163f
C6804 avdd.n4029 avss -0.00357f
C6805 avdd.n4030 avss -0.00108f
C6806 avdd.n4031 avss -2.01e-19
C6807 avdd.n4032 avss -2.96e-19
C6808 avdd.n4033 avss -6.67e-19
C6809 avdd.n4034 avss -1.8e-19
C6810 avdd.n4035 avss 0.0411f
C6811 avdd.n4036 avss 0.0191f
C6812 avdd.n4037 avss -1.38e-19
C6813 avdd.n4038 avss -3.39e-19
C6814 avdd.n4039 avss 0.0111f
C6815 avdd.n4040 avss -2.22e-19
C6816 avdd.n4041 avss 0.0374f
C6817 avdd.n4042 avss 0.0112f
C6818 avdd.n4043 avss -1.8e-19
C6819 avdd.n4044 avss -1.8e-19
C6820 avdd.n4045 avss -0.00109f
C6821 avdd.n4046 avss -0.00126f
C6822 avdd.n4047 avss 0.0318f
C6823 avdd.n4048 avss -0.00139f
C6824 avdd.n4049 avss -2.22e-19
C6825 avdd.n4050 avss 0.0188f
C6826 avdd.n4051 avss -2.75e-19
C6827 avdd.n4052 avss -3.6e-19
C6828 avdd.n4053 avss -3.07e-19
C6829 avdd.n4054 avss -6.88e-19
C6830 avdd.n4055 avss 0.00725f
C6831 avdd.n4056 avss -0.00336f
C6832 avdd.n4057 avss -1.8e-19
C6833 avdd.n4058 avss -2.01e-19
C6834 avdd.n4059 avss -0.0866f
C6835 avdd.n4060 avss 0.0179f
C6836 avdd.n4061 avss 0.0442f
C6837 avdd.n4062 avss -3.39e-19
C6838 avdd.n4063 avss -2.75e-19
C6839 avdd.n4064 avss 0.0181f
C6840 avdd.n4065 avss 0.00821f
C6841 avdd.n4066 avss 0.00821f
C6842 avdd.n4067 avss -2.75e-19
C6843 avdd.n4068 avss -2.33e-19
C6844 avdd.n4069 avss -2.54e-19
C6845 avdd.n4070 avss -2.54e-19
C6846 avdd.n4071 avss -2.22e-19
C6847 avdd.n4072 avss -1.59e-19
C6848 avdd.n4073 avss 0.0298f
C6849 avdd.n4074 avss 0.0098f
C6850 avdd.n4075 avss -0.00158f
C6851 avdd.n4076 avss -8.47e-19
C6852 avdd.n4077 avss -4.23e-19
C6853 avdd.n4078 avss -3.39e-19
C6854 avdd.n4079 avss -2.33e-19
C6855 avdd.n4080 avss -1.16e-19
C6856 avdd.n4081 avss 0.0182f
C6857 avdd.n4082 avss 0.0148f
C6858 avdd.n4083 avss 0.00875f
C6859 avdd.n4085 avss -3.07e-19
C6860 avdd.n4086 avss 0.0192f
C6861 avdd.n4087 avss -1.59e-19
C6862 avdd.n4088 avss -1.8e-19
C6863 avdd.n4089 avss 0.00358f
C6864 avdd.n4090 avss -2.22e-19
C6865 avdd.n4091 avss -1.8e-19
C6866 avdd.n4092 avss -1.8e-19
C6867 avdd.n4093 avss 0.0183f
C6868 avdd.n4094 avss 0.0154f
C6869 avdd.n4095 avss 0.0154f
C6870 avdd.n4096 avss 0.0111f
C6871 avdd.n4097 avss 0.0111f
C6872 avdd.n4098 avss -1.8e-19
C6873 avdd.n4099 avss -8.15e-19
C6874 avdd.n4100 avss -1.48e-19
C6875 avdd.n4101 avss -3.39e-19
C6876 avdd.n4102 avss 0.00466f
C6877 avdd.n4103 avss -8.47e-19
C6878 avdd.n4104 avss -0.0014f
C6879 avdd.n4105 avss 0.0344f
C6880 avdd.n4106 avss -8.47e-19
C6881 avdd.n4107 avss 0.0348f
C6882 avdd.n4108 avss -5.19e-19
C6883 avdd.n4109 avss -3.07e-19
C6884 avdd.n4110 avss -3.28e-19
C6885 avdd.n4111 avss -1.8e-19
C6886 avdd.n4112 avss 0.0189f
C6887 avdd.n4113 avss -2.33e-19
C6888 avdd.n4114 avss 0.0022f
C6889 avdd.n4115 avss 0.0386f
C6890 avdd.n4116 avss -2.44e-19
C6891 avdd.n4117 avss 0.0184f
C6892 avdd.n4118 avss 0.00873f
C6893 avdd.n4119 avss 0.0168f
C6894 avdd.n4120 avss 0.0167f
C6895 avdd.n4121 avss -5.77e-19
C6896 avdd.n4122 avss -8.47e-19
C6897 avdd.n4123 avss -2.22e-19
C6898 avdd.n4124 avss 0.00875f
C6899 avdd.n4125 avss -2.54e-19
C6900 avdd.n4126 avss 0.0182f
C6901 avdd.n4127 avss 0.0111f
C6902 avdd.n4128 avss -1.59e-19
C6903 avdd.n4129 avss -3.39e-19
C6904 avdd.n4130 avss -1.59e-19
C6905 avdd.n4131 avss 3e-19
C6906 avdd.n4132 avss -2.54e-19
C6907 avdd.n4133 avss -1.8e-19
C6908 avdd.n4134 avss -1.8e-19
C6909 avdd.n4135 avss -1.16e-19
C6910 avdd.n4136 avss -2.33e-19
C6911 avdd.n4137 avss -3.39e-19
C6912 avdd.n4138 avss -8.47e-19
C6913 avdd.n4139 avss 0.0342f
C6914 avdd.n4140 avss 0.0049f
C6915 avdd.n4141 avss -8.47e-19
C6916 avdd.n4142 avss 0.0388f
C6917 avdd.n4143 avss -3.39e-19
C6918 avdd.n4144 avss -3.39e-19
C6919 avdd.n4145 avss -2.22e-19
C6920 avdd.n4146 avss -2.01e-19
C6921 avdd.n4147 avss -1.8e-19
C6922 avdd.n4148 avss -1.8e-19
C6923 avdd.n4149 avss -2.22e-19
C6924 avdd.n4150 avss 0.0111f
C6925 avdd.n4151 avss -1.8e-19
C6926 avdd.n4152 avss -2.96e-19
C6927 avdd.n4153 avss -2.44e-19
C6928 avdd.n4154 avss 0.0384f
C6929 avdd.n4155 avss -0.00113f
C6930 avdd.n4156 avss -0.00173f
C6931 avdd.n4157 avss -3.49e-19
C6932 avdd.n4159 avss 0.0382f
C6933 avdd.n4160 avss -3.18e-19
C6934 avdd.n4161 avss -8.47e-19
C6935 avdd.n4162 avss 0.03f
C6936 avdd.n4163 avss 0.00899f
C6937 avdd.n4164 avss -7.52e-19
C6938 avdd.n4165 avss -1.27e-19
C6939 avdd.n4166 avss -2.44e-19
C6940 avdd.n4167 avss -1.8e-19
C6941 avdd.n4168 avss -1.8e-19
C6942 avdd.n4169 avss -1.38e-19
C6943 avdd.n4170 avss -1.38e-19
C6944 avdd.n4171 avss 0.0184f
C6945 avdd.n4172 avss 0.00873f
C6946 avdd.n4173 avss 0.0422f
C6947 avdd.n4174 avss -2.33e-19
C6948 avdd.n4175 avss 0.0197f
C6949 avdd.n4176 avss -2.44e-19
C6950 avdd.n4177 avss -2.44e-19
C6951 avdd.n4178 avss -2.33e-19
C6952 avdd.n4179 avss -1.48e-19
C6953 avdd.n4180 avss -1.8e-19
C6954 avdd.n4181 avss 0.019f
C6955 avdd.n4182 avss 0.00335f
C6956 avdd.n4183 avss 0.0265f
C6957 avdd.n4184 avss 0.00778f
C6958 avdd.n4185 avss -0.00512f
C6959 avdd.n4186 avss -1.8e-19
C6960 avdd.n4187 avss -1.8e-19
C6961 avdd.n4188 avss 0.0191f
C6962 avdd.n4189 avss 0.0154f
C6963 avdd.n4190 avss 0.0154f
C6964 avdd.n4191 avss 0.0183f
C6965 avdd.n4192 avss -1.8e-19
C6966 avdd.n4193 avss -1.8e-19
C6967 avdd.n4194 avss -5.82e-19
C6968 avdd.n4195 avss -6.46e-19
C6969 avdd.n4196 avss -3.07e-19
C6970 avdd.n4197 avss 0.0192f
C6971 avdd.n4198 avss 0.00875f
C6972 avdd.n4199 avss 0.0148f
C6973 avdd.n4200 avss 0.0111f
C6974 avdd.n4201 avss -2.22e-19
C6975 avdd.n4202 avss 0.0192f
C6976 avdd.n4203 avss -4.76e-19
C6977 avdd.n4204 avss -0.00128f
C6978 avdd.n4205 avss 0.0346f
C6979 avdd.n4206 avss 0.00378f
C6980 avdd.n4207 avss -8.47e-19
C6981 avdd.n4208 avss 0.0398f
C6982 avdd.n4209 avss -3.07e-19
C6983 avdd.n4210 avss 0.0181f
C6984 avdd.n4211 avss -3.6e-19
C6985 avdd.n4212 avss -2.01e-19
C6986 avdd.n4213 avss -3.28e-19
C6987 avdd.n4214 avss -8.26e-19
C6988 avdd.n4215 avss -6.46e-19
C6989 avdd.n4216 avss -0.00137f
C6990 avdd.n4217 avss -0.0013f
C6991 avdd.n4218 avss 0.00357f
C6992 avdd.n4219 avss -8.47e-19
C6993 avdd.n4220 avss -3.39e-19
C6994 avdd.n4221 avss -1.27e-19
C6995 avdd.n4222 avss -2.44e-19
C6996 avdd.n4223 avss 0.019f
C6997 avdd.n4224 avss 0.0148f
C6998 avdd.n4225 avss 0.00873f
C6999 avdd.n4226 avss 0.0184f
C7000 avdd.n4227 avss -3.49e-19
C7001 avdd.n4228 avss -1.38e-19
C7002 avdd.n4229 avss -1.8e-19
C7003 avdd.n4230 avss -1.8e-19
C7004 avdd.n4231 avss -2.44e-19
C7005 avdd.n4232 avss -1.8e-19
C7006 avdd.n4233 avss -1.8e-19
C7007 avdd.n4234 avss -5.61e-19
C7008 avdd.n4235 avss -3.39e-19
C7009 avdd.n4236 avss -6.35e-19
C7010 avdd.n4237 avss -0.00121f
C7011 avdd.n4238 avss -0.00122f
C7012 avdd.n4239 avss -0.00173f
C7013 avdd.n4240 avss -9.75e-19
C7014 avdd.n4241 avss 0.0382f
C7015 avdd.n4242 avss -0.198f
C7016 avdd.n4243 avss -0.163f
C7017 avdd.n4244 avss -0.00357f
C7018 avdd.n4245 avss -0.00108f
C7019 avdd.n4246 avss -2.01e-19
C7020 avdd.n4247 avss -2.96e-19
C7021 avdd.n4248 avss -6.67e-19
C7022 avdd.n4249 avss -1.8e-19
C7023 avdd.n4250 avss 0.0411f
C7024 avdd.n4251 avss 0.0191f
C7025 avdd.n4252 avss -1.38e-19
C7026 avdd.n4253 avss -3.39e-19
C7027 avdd.n4254 avss 0.0111f
C7028 avdd.n4255 avss -2.22e-19
C7029 avdd.n4256 avss 0.0374f
C7030 avdd.n4257 avss 0.0112f
C7031 avdd.n4258 avss -1.8e-19
C7032 avdd.n4259 avss -1.8e-19
C7033 avdd.n4260 avss -0.00109f
C7034 avdd.n4261 avss -0.00126f
C7035 avdd.n4262 avss 0.0318f
C7036 avdd.n4263 avss -0.00139f
C7037 avdd.n4264 avss -2.22e-19
C7038 avdd.n4265 avss 0.0188f
C7039 avdd.n4266 avss -2.75e-19
C7040 avdd.n4267 avss -3.6e-19
C7041 avdd.n4268 avss -3.07e-19
C7042 avdd.n4269 avss -6.88e-19
C7043 avdd.n4270 avss 0.00725f
C7044 avdd.n4271 avss -0.00336f
C7045 avdd.n4272 avss -1.8e-19
C7046 avdd.n4273 avss -2.01e-19
C7047 avdd.n4274 avss -0.0866f
C7048 avdd.n4275 avss 0.0179f
C7049 avdd.n4276 avss 0.0442f
C7050 avdd.n4277 avss -3.39e-19
C7051 avdd.n4278 avss -2.75e-19
C7052 avdd.n4279 avss 0.0181f
C7053 avdd.n4280 avss 0.00821f
C7054 avdd.n4281 avss 0.00821f
C7055 avdd.n4282 avss -2.75e-19
C7056 avdd.n4283 avss -2.33e-19
C7057 avdd.n4284 avss -2.54e-19
C7058 avdd.n4285 avss -2.54e-19
C7059 avdd.n4286 avss -2.22e-19
C7060 avdd.n4287 avss -1.59e-19
C7061 avdd.n4288 avss 0.0298f
C7062 avdd.n4289 avss 0.0098f
C7063 avdd.n4290 avss -0.00158f
C7064 avdd.n4291 avss -8.47e-19
C7065 avdd.n4292 avss -4.23e-19
C7066 avdd.n4293 avss -3.39e-19
C7067 avdd.n4294 avss -2.33e-19
C7068 avdd.n4295 avss -1.16e-19
C7069 avdd.n4296 avss 0.0182f
C7070 avdd.n4297 avss 0.0148f
C7071 avdd.n4298 avss 0.00875f
C7072 avdd.n4300 avss -3.07e-19
C7073 avdd.n4301 avss 0.0192f
C7074 avdd.n4302 avss -1.59e-19
C7075 avdd.n4303 avss -1.8e-19
C7076 avdd.n4304 avss 0.00358f
C7077 avdd.n4305 avss -2.22e-19
C7078 avdd.n4306 avss -1.8e-19
C7079 avdd.n4307 avss -1.8e-19
C7080 avdd.n4308 avss 0.0183f
C7081 avdd.n4309 avss 0.0154f
C7082 avdd.n4310 avss 0.0154f
C7083 avdd.n4311 avss 0.0111f
C7084 avdd.n4312 avss 0.0111f
C7085 avdd.n4313 avss -1.8e-19
C7086 avdd.n4314 avss -8.15e-19
C7087 avdd.n4315 avss -1.48e-19
C7088 avdd.n4316 avss -3.39e-19
C7089 avdd.n4317 avss 0.00466f
C7090 avdd.n4318 avss -8.47e-19
C7091 avdd.n4319 avss -0.0014f
C7092 avdd.n4320 avss 0.0344f
C7093 avdd.n4321 avss -8.47e-19
C7094 avdd.n4322 avss 0.0348f
C7095 avdd.n4323 avss -5.19e-19
C7096 avdd.n4324 avss -3.07e-19
C7097 avdd.n4325 avss -3.28e-19
C7098 avdd.n4326 avss -1.8e-19
C7099 avdd.n4327 avss 0.0189f
C7100 avdd.n4328 avss -2.33e-19
C7101 avdd.n4329 avss 0.0022f
C7102 avdd.n4330 avss 0.0386f
C7103 avdd.n4331 avss -2.44e-19
C7104 avdd.n4332 avss 0.0184f
C7105 avdd.n4333 avss 0.00873f
C7106 avdd.n4334 avss 0.0168f
C7107 avdd.n4335 avss 0.0167f
C7108 avdd.n4336 avss -5.77e-19
C7109 avdd.n4337 avss -8.47e-19
C7110 avdd.n4338 avss -2.22e-19
C7111 avdd.n4339 avss 0.00875f
C7112 avdd.n4340 avss -2.54e-19
C7113 avdd.n4341 avss 0.0182f
C7114 avdd.n4342 avss 0.0111f
C7115 avdd.n4343 avss -1.59e-19
C7116 avdd.n4344 avss -3.39e-19
C7117 avdd.n4345 avss -1.59e-19
C7118 avdd.n4346 avss 3e-19
C7119 avdd.n4347 avss -2.54e-19
C7120 avdd.n4348 avss -1.8e-19
C7121 avdd.n4349 avss -1.8e-19
C7122 avdd.n4350 avss -1.16e-19
C7123 avdd.n4351 avss -2.33e-19
C7124 avdd.n4352 avss -3.39e-19
C7125 avdd.n4353 avss -8.47e-19
C7126 avdd.n4354 avss 0.0342f
C7127 avdd.n4355 avss 0.0049f
C7128 avdd.n4356 avss -8.47e-19
C7129 avdd.n4357 avss 0.0388f
C7130 avdd.n4358 avss -3.39e-19
C7131 avdd.n4359 avss -3.39e-19
C7132 avdd.n4360 avss -2.22e-19
C7133 avdd.n4361 avss -2.01e-19
C7134 avdd.n4362 avss -1.8e-19
C7135 avdd.n4363 avss -1.8e-19
C7136 avdd.n4364 avss -2.22e-19
C7137 avdd.n4365 avss 0.0111f
C7138 avdd.n4366 avss -1.8e-19
C7139 avdd.n4367 avss -2.96e-19
C7140 avdd.n4368 avss -2.44e-19
C7141 avdd.n4369 avss 0.0384f
C7142 avdd.n4370 avss -0.00113f
C7143 avdd.n4371 avss -0.00173f
C7144 avdd.n4372 avss -3.49e-19
C7145 avdd.n4374 avss 0.0382f
C7146 avdd.n4375 avss -3.18e-19
C7147 avdd.n4376 avss -8.47e-19
C7148 avdd.n4377 avss 0.03f
C7149 avdd.n4378 avss 0.00899f
C7150 avdd.n4379 avss -7.52e-19
C7151 avdd.n4380 avss -1.27e-19
C7152 avdd.n4381 avss -2.44e-19
C7153 avdd.n4382 avss -1.8e-19
C7154 avdd.n4383 avss -1.8e-19
C7155 avdd.n4384 avss -1.38e-19
C7156 avdd.n4385 avss -1.38e-19
C7157 avdd.n4386 avss 0.0184f
C7158 avdd.n4387 avss 0.00873f
C7159 avdd.n4388 avss 0.0422f
C7160 avdd.n4389 avss -2.33e-19
C7161 avdd.n4390 avss 0.0197f
C7162 avdd.n4391 avss -2.44e-19
C7163 avdd.n4392 avss -2.44e-19
C7164 avdd.n4393 avss -2.33e-19
C7165 avdd.n4394 avss -1.48e-19
C7166 avdd.n4395 avss -1.8e-19
C7167 avdd.n4396 avss 0.019f
C7168 avdd.n4397 avss 0.00335f
C7169 avdd.n4398 avss 0.0265f
C7170 avdd.n4399 avss 0.00778f
C7171 avdd.n4400 avss -0.00512f
C7172 avdd.n4401 avss -1.8e-19
C7173 avdd.n4402 avss -1.8e-19
C7174 avdd.n4403 avss 0.0191f
C7175 avdd.n4404 avss 0.0154f
C7176 avdd.n4405 avss 0.0154f
C7177 avdd.n4406 avss 0.0183f
C7178 avdd.n4407 avss -1.8e-19
C7179 avdd.n4408 avss -1.8e-19
C7180 avdd.n4409 avss -5.82e-19
C7181 avdd.n4410 avss -6.46e-19
C7182 avdd.n4411 avss -3.07e-19
C7183 avdd.n4412 avss 0.0192f
C7184 avdd.n4413 avss 0.00875f
C7185 avdd.n4414 avss 0.0148f
C7186 avdd.n4415 avss 0.0111f
C7187 avdd.n4416 avss -2.22e-19
C7188 avdd.n4417 avss 0.0192f
C7189 avdd.n4418 avss -4.76e-19
C7190 avdd.n4419 avss -0.00128f
C7191 avdd.n4420 avss 0.0346f
C7192 avdd.n4421 avss 0.00378f
C7193 avdd.n4422 avss -8.47e-19
C7194 avdd.n4423 avss 0.0398f
C7195 avdd.n4424 avss -3.07e-19
C7196 avdd.n4425 avss 0.0181f
C7197 avdd.n4426 avss -3.6e-19
C7198 avdd.n4427 avss -2.01e-19
C7199 avdd.n4428 avss -3.28e-19
C7200 avdd.n4429 avss -8.26e-19
C7201 avdd.n4430 avss -6.46e-19
C7202 avdd.n4431 avss -0.00137f
C7203 avdd.n4432 avss -0.0013f
C7204 avdd.n4433 avss 0.00357f
C7205 avdd.n4434 avss -8.47e-19
C7206 avdd.n4435 avss -3.39e-19
C7207 avdd.n4436 avss -1.27e-19
C7208 avdd.n4437 avss -2.44e-19
C7209 avdd.n4438 avss 0.019f
C7210 avdd.n4439 avss 0.0148f
C7211 avdd.n4440 avss 0.00873f
C7212 avdd.n4441 avss 0.0184f
C7213 avdd.n4442 avss -3.49e-19
C7214 avdd.n4443 avss -1.38e-19
C7215 avdd.n4444 avss -1.8e-19
C7216 avdd.n4445 avss -1.8e-19
C7217 avdd.n4446 avss -2.44e-19
C7218 avdd.n4447 avss -1.8e-19
C7219 avdd.n4448 avss -1.8e-19
C7220 avdd.n4449 avss -5.61e-19
C7221 avdd.n4450 avss -3.39e-19
C7222 avdd.n4451 avss -6.35e-19
C7223 avdd.n4452 avss -0.00121f
C7224 avdd.n4453 avss -0.00122f
C7225 avdd.n4454 avss -0.00173f
C7226 avdd.n4455 avss -9.75e-19
C7227 avdd.n4456 avss 0.0382f
C7228 avdd.n4457 avss -0.722f
C7229 avdd.n4458 avss -1.38e-19
C7230 avdd.t316 avss -7.94e-19
C7231 avdd.t4 avss -0.00135f
C7232 avdd.t323 avss -7.94e-19
C7233 avdd.t6 avss -0.00135f
C7234 avdd.n4459 avss -0.00226f
C7235 avdd.n4460 avss -0.00233f
C7236 avdd.n4461 avss -4.13e-19
C7237 avdd.n4462 avss -7.92e-19
C7238 avdd.n4463 avss -2.26e-19
C7239 avdd.n4464 avss -0.00675f
C7240 avdd.n4465 avss -9.91e-19
C7241 avdd.t5 avss -0.00352f
C7242 avdd.n4466 avss -0.00442f
C7243 avdd.n4467 avss -0.00213f
C7244 avdd.n4468 avss -7.31e-19
C7245 avdd.t2 avss -0.00352f
C7246 avdd.n4469 avss -0.004f
C7247 avdd.t8 avss -0.00352f
C7248 avdd.n4470 avss -0.00433f
C7249 avdd.n4471 avss -0.00213f
C7250 avdd.n4472 avss -7.31e-19
C7251 avdd.t74 avss -0.00352f
C7252 avdd.n4473 avss -0.00401f
C7253 avdd.t155 avss -0.00352f
C7254 avdd.n4474 avss -0.00434f
C7255 avdd.n4475 avss -0.00213f
C7256 avdd.n4476 avss -7.31e-19
C7257 avdd.t157 avss -0.00352f
C7258 avdd.n4477 avss -0.00401f
C7259 avdd.t159 avss -0.00352f
C7260 avdd.n4478 avss -0.00434f
C7261 avdd.n4479 avss -0.00213f
C7262 avdd.n4480 avss -7.31e-19
C7263 avdd.t186 avss -0.00352f
C7264 avdd.n4481 avss -0.00401f
C7265 avdd.t71 avss -0.00352f
C7266 avdd.n4482 avss -0.00434f
C7267 avdd.n4483 avss -0.00213f
C7268 avdd.n4484 avss -0.00106f
C7269 avdd.n4485 avss -7.42e-19
C7270 avdd.n4486 avss -0.00207f
C7271 avdd.n4487 avss -7.42e-19
C7272 avdd.n4488 avss -0.0169f
C7273 avdd.n4489 avss -0.00865f
C7274 avdd.n4490 avss -0.00164f
C7275 avdd.n4491 avss -7.42e-19
C7276 avdd.n4492 avss -0.00158f
C7277 avdd.n4493 avss -7.42e-19
C7278 avdd.n4494 avss -7.42e-19
C7279 avdd.n4495 avss -7.42e-19
C7280 avdd.n4496 avss -7.42e-19
C7281 avdd.n4498 avss -0.021f
C7282 avdd.n4500 avss -7.42e-19
C7283 avdd.n4501 avss -7.42e-19
C7284 avdd.n4502 avss -0.00158f
C7285 avdd.n4503 avss -0.00164f
C7286 avdd.n4504 avss -2.13e-19
C7287 avdd.n4505 avss -3.71e-19
C7288 avdd.t33 avss -0.00735f
C7289 avdd.n4506 avss -0.00735f
C7290 avdd.n4507 avss -7.42e-19
C7291 avdd.n4508 avss -7.42e-19
C7292 avdd.n4509 avss -0.00184f
C7293 avdd.n4510 avss -7.42e-19
C7294 avdd.n4511 avss -0.00735f
C7295 avdd.n4512 avss -0.00735f
C7296 avdd.n4513 avss -3.71e-19
C7297 avdd.n4514 avss -3.71e-19
C7298 avdd.n4515 avss -3.71e-19
C7299 avdd.n4516 avss -1.8e-19
C7300 avdd.n4517 avss -0.00123f
C7301 avdd.n4518 avss -1.64e-19
C7302 avdd.n4519 avss -2.02e-19
C7303 avdd.n4520 avss -9.27e-20
C7304 avdd.n4521 avss -0.00154f
C7305 avdd.n4522 avss -2.95e-19
C7306 avdd.n4523 avss -9.27e-20
C7307 avdd.n4524 avss -9.27e-20
C7308 avdd.n4525 avss -9.27e-20
C7309 avdd.n4526 avss -0.00184f
C7310 avdd.n4527 avss -0.00584f
C7311 avdd.n4528 avss -0.00735f
C7312 avdd.n4529 avss -7.42e-19
C7313 avdd.n4530 avss -7.42e-19
C7314 avdd.n4531 avss -7.42e-19
C7315 avdd.n4532 avss -7.42e-19
C7316 avdd.n4533 avss -0.0144f
C7317 avdd.n4534 avss -0.0104f
C7318 avdd.n4535 avss -7.25e-19
C7319 avdd.n4536 avss -7.42e-19
C7320 avdd.n4537 avss -3.71e-19
C7321 avdd.n4538 avss -3.71e-19
C7322 avdd.n4539 avss -7.25e-19
C7323 avdd.n4540 avss -7.42e-19
C7324 avdd.n4541 avss -7.42e-19
C7325 avdd.t289 avss -0.00735f
C7326 avdd.n4542 avss -0.0147f
C7327 avdd.n4543 avss -7.42e-19
C7328 avdd.n4544 avss -7.42e-19
C7329 avdd.n4545 avss -7.42e-19
C7330 avdd.n4546 avss -0.0147f
C7331 avdd.n4547 avss -7.42e-19
C7332 avdd.n4548 avss -7.42e-19
C7333 avdd.n4549 avss -7.42e-19
C7334 avdd.n4550 avss -0.0147f
C7335 avdd.n4551 avss -7.42e-19
C7336 avdd.n4552 avss -7.42e-19
C7337 avdd.n4553 avss -7.42e-19
C7338 avdd.t108 avss -0.00735f
C7339 avdd.n4554 avss -7.42e-19
C7340 avdd.n4555 avss -3.71e-19
C7341 avdd.n4556 avss -3.71e-19
C7342 avdd.n4557 avss -0.0121f
C7343 avdd.n4558 avss -0.00735f
C7344 avdd.n4559 avss -7.42e-19
C7345 avdd.n4560 avss -7.42e-19
C7346 avdd.n4561 avss -0.00184f
C7347 avdd.n4562 avss -7.42e-19
C7348 avdd.n4563 avss -0.00735f
C7349 avdd.n4564 avss -0.00735f
C7350 avdd.n4565 avss -3.71e-19
C7351 avdd.n4566 avss -3.71e-19
C7352 avdd.n4567 avss -2.67e-19
C7353 avdd.n4568 avss -6e-20
C7354 avdd.n4569 avss -3.22e-19
C7355 avdd.n4570 avss -0.00184f
C7356 avdd.n4571 avss -9.27e-20
C7357 avdd.n4572 avss -2.62e-19
C7358 avdd.n4573 avss -9.27e-20
C7359 avdd.n4574 avss -5.77e-19
C7360 avdd.n4575 avss -6.98e-19
C7361 avdd.n4576 avss -0.0117f
C7362 avdd.n4577 avss -7.42e-19
C7363 avdd.n4578 avss -7.42e-19
C7364 avdd.n4579 avss -7.42e-19
C7365 avdd.n4580 avss -7.42e-19
C7366 avdd.n4581 avss -0.002f
C7367 avdd.n4582 avss -0.002f
C7368 avdd.t30 avss -0.00735f
C7369 avdd.n4583 avss -0.0225f
C7370 avdd.n4584 avss -7.42e-19
C7371 avdd.n4585 avss -0.0019f
C7372 avdd.n4586 avss -1.64e-19
C7373 avdd.t34 avss -0.00173f
C7374 avdd.n4587 avss -0.011f
C7375 avdd.n4588 avss -6.54e-19
C7376 avdd.n4589 avss -2.13e-19
C7377 avdd.n4590 avss -3.05e-19
C7378 avdd.n4591 avss -9.27e-20
C7379 avdd.n4592 avss -2.18e-19
C7380 avdd.n4593 avss -5.49e-19
C7381 avdd.n4594 avss -1.64e-19
C7382 avdd.n4595 avss -9.27e-20
C7383 avdd.n4596 avss -9.27e-20
C7384 avdd.n4597 avss -1.36e-19
C7385 avdd.n4598 avss -3.55e-19
C7386 avdd.n4599 avss -0.00703f
C7387 avdd.n4600 avss -0.00605f
C7388 avdd.n4601 avss -0.00184f
C7389 avdd.n4602 avss -9.27e-20
C7390 avdd.n4603 avss -9.27e-20
C7391 avdd.n4604 avss -1.58e-19
C7392 avdd.n4605 avss -9.27e-20
C7393 avdd.n4606 avss -1.64e-19
C7394 avdd.n4607 avss -0.00127f
C7395 avdd.n4608 avss -0.00156f
C7396 avdd.n4609 avss -0.00787f
C7397 avdd.n4610 avss -0.00806f
C7398 avdd.t290 avss -0.00173f
C7399 avdd.n4611 avss -0.0017f
C7400 avdd.n4612 avss -0.011f
C7401 avdd.n4613 avss -0.00784f
C7402 avdd.n4614 avss -0.00785f
C7403 avdd.t109 avss -0.00173f
C7404 avdd.n4615 avss -0.0115f
C7405 avdd.n4616 avss -1.64e-19
C7406 avdd.n4617 avss -9.27e-20
C7407 avdd.n4618 avss -9.27e-20
C7408 avdd.n4619 avss -9.27e-20
C7409 avdd.n4620 avss -9.27e-20
C7410 avdd.n4621 avss -2.51e-19
C7411 avdd.n4622 avss -9.27e-20
C7412 avdd.n4623 avss -6.06e-19
C7413 avdd.n4624 avss -6.26e-19
C7414 avdd.n4625 avss -9.27e-20
C7415 avdd.n4626 avss -1.64e-19
C7416 avdd.n4627 avss -0.00115f
C7417 avdd.n4628 avss -0.00118f
C7418 avdd.n4629 avss -1.64e-19
C7419 avdd.n4630 avss -5.97e-19
C7420 avdd.n4631 avss -1.04e-19
C7421 avdd.n4632 avss -9.27e-20
C7422 avdd.n4633 avss -2.35e-19
C7423 avdd.n4634 avss -3.27e-19
C7424 avdd.n4635 avss -0.00184f
C7425 avdd.n4636 avss -0.00649f
C7426 avdd.n4637 avss -0.0066f
C7427 avdd.n4638 avss -3.33e-19
C7428 avdd.n4639 avss -8.18e-20
C7429 avdd.n4640 avss -9.05e-19
C7430 avdd.n4641 avss -0.00115f
C7431 avdd.n4642 avss -0.015f
C7432 avdd.t31 avss -0.00174f
C7433 avdd.n4643 avss -0.0157f
C7434 avdd.n4644 avss -0.00207f
C7435 avdd.n4645 avss -2.89e-19
C7436 avdd.n4646 avss -6.05e-19
C7437 avdd.n4647 avss -7.42e-19
C7438 avdd.n4648 avss -7.42e-19
C7439 avdd.n4649 avss -7.42e-19
C7440 avdd.n4652 avss -0.00197f
C7441 avdd.n4653 avss -0.00197f
C7442 avdd.n4654 avss -7.42e-19
C7443 avdd.n4655 avss -7.42e-19
C7444 avdd.n4656 avss -7.42e-19
C7445 avdd.n4657 avss -7.42e-19
C7446 avdd.n4659 avss -0.0266f
C7447 avdd.n4661 avss -0.00189f
C7448 avdd.n4662 avss -0.00189f
C7449 avdd.n4663 avss -0.0019f
C7450 avdd.n4664 avss -7.42e-19
C7451 avdd.n4665 avss -7.42e-19
C7452 avdd.n4666 avss -0.0104f
C7453 avdd.n4667 avss -7.42e-19
C7454 avdd.n4668 avss -7.42e-19
C7455 avdd.n4669 avss -7.42e-19
C7456 avdd.n4670 avss -7.42e-19
C7457 avdd.n4671 avss -7.42e-19
C7458 avdd.n4672 avss -0.0138f
C7459 avdd.n4673 avss -0.00735f
C7460 avdd.n4674 avss -3.71e-19
C7461 avdd.n4675 avss -8.18e-20
C7462 avdd.n4676 avss -9.27e-20
C7463 avdd.n4677 avss -2.45e-19
C7464 avdd.n4678 avss -3.38e-19
C7465 avdd.n4679 avss -0.0067f
C7466 avdd.n4680 avss -0.00638f
C7467 avdd.n4681 avss -0.00184f
C7468 avdd.n4682 avss -9.27e-20
C7469 avdd.n4683 avss -9.27e-20
C7470 avdd.n4684 avss -3.71e-19
C7471 avdd.n4685 avss -5.35e-19
C7472 avdd.n4686 avss -6.27e-19
C7473 avdd.n4687 avss -0.0124f
C7474 avdd.n4688 avss -7.42e-19
C7475 avdd.n4689 avss -7.42e-19
C7476 avdd.n4690 avss -7.42e-19
C7477 avdd.n4691 avss -7.42e-19
C7478 avdd.n4692 avss -7.42e-19
C7479 avdd.n4693 avss -7.42e-19
C7480 avdd.n4694 avss -0.0137f
C7481 avdd.n4695 avss -6.93e-19
C7482 avdd.n4696 avss -6.93e-19
C7483 avdd.n4697 avss -7.42e-19
C7484 avdd.n4698 avss -7.42e-19
C7485 avdd.n4699 avss -7.42e-19
C7486 avdd.n4700 avss -0.00995f
C7487 avdd.n4701 avss -7.42e-19
C7488 avdd.n4702 avss -7.42e-19
C7489 avdd.n4703 avss -7.42e-19
C7490 avdd.n4704 avss -7.42e-19
C7491 avdd.n4705 avss -7.42e-19
C7492 avdd.n4706 avss -0.0147f
C7493 avdd.n4707 avss -7.42e-19
C7494 avdd.n4708 avss -7.42e-19
C7495 avdd.n4709 avss -7.42e-19
C7496 avdd.n4710 avss -7.42e-19
C7497 avdd.n4711 avss -7.42e-19
C7498 avdd.n4712 avss -0.0147f
C7499 avdd.n4713 avss -7.42e-19
C7500 avdd.n4714 avss -7.42e-19
C7501 avdd.n4715 avss -7.42e-19
C7502 avdd.n4716 avss -7.42e-19
C7503 avdd.n4717 avss -7.42e-19
C7504 avdd.n4718 avss -0.0117f
C7505 avdd.n4719 avss -7.42e-19
C7506 avdd.n4720 avss -7.42e-19
C7507 avdd.n4721 avss -7.42e-19
C7508 avdd.n4722 avss -7.42e-19
C7509 avdd.n4723 avss -7.42e-19
C7510 avdd.n4724 avss -0.0147f
C7511 avdd.n4725 avss -7.42e-19
C7512 avdd.n4726 avss -7.42e-19
C7513 avdd.n4727 avss -7.42e-19
C7514 avdd.n4728 avss -7.42e-19
C7515 avdd.n4729 avss -7.42e-19
C7516 avdd.n4730 avss -0.00184f
C7517 avdd.n4731 avss -0.00724f
C7518 avdd.n4732 avss -3.65e-19
C7519 avdd.n4733 avss -1.58e-19
C7520 avdd.n4734 avss -9.27e-20
C7521 avdd.n4735 avss -2.07e-19
C7522 avdd.n4736 avss -5.29e-19
C7523 avdd.n4737 avss -6.74e-19
C7524 avdd.n4738 avss -0.00127f
C7525 avdd.n4739 avss -2.84e-19
C7526 avdd.n4740 avss -5.35e-19
C7527 avdd.n4741 avss -6.27e-19
C7528 avdd.n4742 avss -0.0124f
C7529 avdd.n4743 avss -7.42e-19
C7530 avdd.n4744 avss -7.42e-19
C7531 avdd.n4745 avss -7.42e-19
C7532 avdd.n4746 avss -7.42e-19
C7533 avdd.n4747 avss -7.42e-19
C7534 avdd.n4748 avss -7.42e-19
C7535 avdd.n4749 avss -0.0119f
C7536 avdd.n4750 avss -6.65e-19
C7537 avdd.n4751 avss -5.73e-19
C7538 avdd.n4752 avss -7.42e-19
C7539 avdd.n4753 avss -7.42e-19
C7540 avdd.n4754 avss -7.42e-19
C7541 avdd.n4755 avss -0.0147f
C7542 avdd.n4756 avss -0.00208f
C7543 avdd.n4757 avss -0.0012f
C7544 avdd.n4758 avss -0.00766f
C7545 avdd.t20 avss -0.00412f
C7546 avdd.t153 avss -0.00397f
C7547 avdd.t19 avss -0.127f
C7548 avdd.t28 avss -0.123f
C7549 avdd.t17 avss -0.0473f
C7550 avdd.n4759 avss -0.082f
C7551 avdd.t154 avss -0.00412f
C7552 avdd.t18 avss -0.00397f
C7553 avdd.t29 avss -0.00412f
C7554 avdd.t32 avss -0.00406f
C7555 avdd.n4760 avss -0.0114f
C7556 avdd.n4761 avss -0.0125f
C7557 avdd.n4762 avss -0.0368f
C7558 avdd.n4763 avss -0.0152f
C7559 avdd.n4764 avss -0.0683f
C7560 avdd.n4765 avss -0.0447f
C7561 avdd.n4766 avss -0.0018f
C7562 avdd.n4767 avss -0.00208f
C7563 avdd.n4768 avss -8.51e-19
C7564 avdd.t156 avss -0.00352f
C7565 avdd.n4769 avss -0.00411f
C7566 avdd.n4770 avss -7.31e-19
C7567 avdd.n4771 avss -0.00257f
C7568 avdd.n4772 avss -9.55e-19
C7569 avdd.n4773 avss -0.00213f
C7570 avdd.n4774 avss -0.00257f
C7571 avdd.n4775 avss -9.39e-19
C7572 avdd.t185 avss -0.00352f
C7573 avdd.n4776 avss -0.00433f
C7574 avdd.t160 avss -0.00352f
C7575 avdd.n4777 avss -0.004f
C7576 avdd.n4778 avss -7.31e-19
C7577 avdd.n4779 avss -0.00257f
C7578 avdd.n4780 avss -9.55e-19
C7579 avdd.n4781 avss -0.00213f
C7580 avdd.n4782 avss -0.00257f
C7581 avdd.n4783 avss -9.55e-19
C7582 avdd.t158 avss -0.00352f
C7583 avdd.n4784 avss -0.00434f
C7584 avdd.t288 avss -0.00352f
C7585 avdd.n4785 avss -0.00401f
C7586 avdd.n4786 avss -7.31e-19
C7587 avdd.n4787 avss -0.00257f
C7588 avdd.n4788 avss -9.7e-19
C7589 avdd.n4789 avss -0.00213f
C7590 avdd.n4790 avss -0.00257f
C7591 avdd.n4791 avss -9.55e-19
C7592 avdd.t287 avss -0.00352f
C7593 avdd.n4792 avss -0.00434f
C7594 avdd.t9 avss -0.00352f
C7595 avdd.n4793 avss -0.00401f
C7596 avdd.n4794 avss -7.31e-19
C7597 avdd.n4795 avss -0.00257f
C7598 avdd.n4796 avss -9.39e-19
C7599 avdd.n4797 avss -0.00213f
C7600 avdd.n4798 avss -0.00257f
C7601 avdd.n4799 avss -9.55e-19
C7602 avdd.t107 avss -0.00352f
C7603 avdd.n4800 avss -0.00434f
C7604 avdd.t7 avss -0.00352f
C7605 avdd.n4801 avss -0.00401f
C7606 avdd.n4802 avss -7.31e-19
C7607 avdd.n4803 avss -0.00257f
C7608 avdd.n4804 avss -9.24e-19
C7609 avdd.n4805 avss -0.00159f
C7610 avdd.n4806 avss -0.00543f
C7611 avdd.n4807 avss -0.0574f
C7612 avdd.n4808 avss -0.613f
C7613 avdd.n4809 avss -0.286f
C7614 avdd.n4810 avss 0.0269f
C7615 avdd.n4811 avss -1.27e-19
C7616 avdd.n4812 avss -2.96e-19
C7617 avdd.n4813 avss -0.00113f
C7618 avdd.n4815 avss -1.8e-19
C7619 avdd.n4816 avss -8.47e-19
C7620 avdd.n4817 avss 0.00869f
C7621 avdd.n4819 avss -0.00173f
C7622 avdd.n4820 avss -2.44e-19
C7623 avdd.n4821 avss 0.0111f
C7624 avdd.n4822 avss -1.38e-19
C7625 avdd.n4823 avss -2.44e-19
C7626 avdd.n4824 avss 0.0111f
C7627 avdd.n4825 avss -1.8e-19
C7628 avdd.n4826 avss -1.8e-19
C7629 avdd.n4827 avss 0.00908f
C7630 avdd.n4828 avss 0.03f
C7631 avdd.n4829 avss -3.39e-19
C7632 avdd.n4830 avss -3.39e-19
C7633 avdd.n4831 avss -1.59e-19
C7634 avdd.n4832 avss 0.0111f
C7635 avdd.n4833 avss -1.8e-19
C7636 avdd.n4834 avss -1.8e-19
C7637 avdd.n4835 avss 0.0342f
C7638 avdd.n4836 avss 0.00378f
C7639 avdd.n4837 avss -5.77e-19
C7640 avdd.n4838 avss -2.22e-19
C7641 avdd.n4839 avss 0.0168f
C7642 avdd.n4840 avss -3.6e-19
C7643 avdd.n4841 avss -1.8e-19
C7644 avdd.n4842 avss -8.26e-19
C7645 avdd.n4843 avss -0.0013f
C7646 avdd.n4844 avss -3.39e-19
C7647 avdd.n4845 avss -1.27e-19
C7648 avdd.n4846 avss 0.0022f
C7649 avdd.n4847 avss 0.019f
C7650 avdd.n4848 avss 0.0184f
C7651 avdd.n4849 avss -5.19e-19
C7652 avdd.n4850 avss 0.0386f
C7653 avdd.n4851 avss 0.0111f
C7654 avdd.n4852 avss -1.38e-19
C7655 avdd.n4853 avss -1.38e-19
C7656 avdd.n4854 avss -3.39e-19
C7657 avdd.n4855 avss -3.39e-19
C7658 avdd.n4856 avss -1.8e-19
C7659 avdd.n4857 avss 0.0411f
C7660 avdd.n4858 avss 0.0111f
C7661 avdd.n4859 avss -1.8e-19
C7662 avdd.n4860 avss -1.8e-19
C7663 avdd.n4861 avss -0.00173f
C7664 avdd.n4862 avss -0.00122f
C7665 avdd.n4863 avss -2.96e-19
C7666 avdd.n4864 avss -0.00121f
C7667 avdd.n4865 avss -6.35e-19
C7668 avdd.n4866 avss -0.00357f
C7669 avdd.n4867 avss -0.00109f
C7670 avdd.n4868 avss 0.0374f
C7671 avdd.n4869 avss 0.0112f
C7672 avdd.n4870 avss -1.8e-19
C7673 avdd.n4871 avss -1.8e-19
C7674 avdd.n4872 avss -0.00126f
C7675 avdd.n4873 avss 0.0318f
C7676 avdd.n4874 avss -0.00139f
C7677 avdd.n4875 avss -2.22e-19
C7678 avdd.n4876 avss 0.0188f
C7679 avdd.n4877 avss -2.75e-19
C7680 avdd.n4878 avss -3.6e-19
C7681 avdd.n4879 avss -3.07e-19
C7682 avdd.n4880 avss -6.88e-19
C7683 avdd.n4881 avss 0.00725f
C7684 avdd.n4882 avss -0.00336f
C7685 avdd.n4883 avss -1.8e-19
C7686 avdd.n4884 avss -2.01e-19
C7687 avdd.n4885 avss -0.0866f
C7688 avdd.n4886 avss 0.0179f
C7689 avdd.n4887 avss 0.0442f
C7690 avdd.n4888 avss -3.39e-19
C7691 avdd.n4889 avss -2.75e-19
C7692 avdd.n4890 avss 0.0181f
C7693 avdd.n4891 avss 0.00821f
C7694 avdd.n4892 avss 0.00821f
C7695 avdd.n4893 avss -2.75e-19
C7696 avdd.n4894 avss -2.33e-19
C7697 avdd.n4895 avss -2.54e-19
C7698 avdd.n4896 avss -2.54e-19
C7699 avdd.n4897 avss -2.22e-19
C7700 avdd.n4898 avss -1.59e-19
C7701 avdd.n4899 avss 0.0298f
C7702 avdd.n4900 avss 0.0098f
C7703 avdd.n4901 avss -0.00158f
C7704 avdd.n4902 avss -8.47e-19
C7705 avdd.n4903 avss -4.23e-19
C7706 avdd.n4904 avss -3.39e-19
C7707 avdd.n4905 avss -2.33e-19
C7708 avdd.n4906 avss -1.16e-19
C7709 avdd.n4907 avss 0.0182f
C7710 avdd.n4908 avss 0.0148f
C7711 avdd.n4909 avss 0.00875f
C7712 avdd.n4910 avss -2.22e-19
C7713 avdd.n4911 avss -2.22e-19
C7714 avdd.n4912 avss 0.00358f
C7715 avdd.n4913 avss -1.8e-19
C7716 avdd.n4914 avss -1.59e-19
C7717 avdd.n4915 avss 0.0192f
C7718 avdd.n4916 avss -3.07e-19
C7719 avdd.n4917 avss -0.00108f
C7720 avdd.n4918 avss 0.0382f
C7721 avdd.n4919 avss -9.76e-19
C7722 avdd.n4920 avss -2.01e-19
C7723 avdd.n4921 avss 0.0183f
C7724 avdd.n4922 avss 0.0154f
C7725 avdd.n4923 avss 0.0154f
C7726 avdd.n4924 avss 0.0191f
C7727 avdd.n4925 avss -1.8e-19
C7728 avdd.n4926 avss -1.8e-19
C7729 avdd.n4927 avss -2.44e-19
C7730 avdd.n4928 avss -1.8e-19
C7731 avdd.n4929 avss -1.8e-19
C7732 avdd.n4930 avss -5.61e-19
C7733 avdd.n4931 avss 0.0344f
C7734 avdd.n4932 avss -2.44e-19
C7735 avdd.n4933 avss -8.47e-19
C7736 avdd.n4934 avss -8.15e-19
C7737 avdd.n4935 avss -0.0014f
C7738 avdd.n4936 avss -8.47e-19
C7739 avdd.n4937 avss 0.00466f
C7740 avdd.n4938 avss -3.39e-19
C7741 avdd.n4939 avss -6.67e-19
C7742 avdd.n4940 avss -3.49e-19
C7743 avdd.n4941 avss 0.0184f
C7744 avdd.n4942 avss 0.00873f
C7745 avdd.n4943 avss 0.0148f
C7746 avdd.n4944 avss 0.00873f
C7747 avdd.n4945 avss 0.0111f
C7748 avdd.n4946 avss -2.44e-19
C7749 avdd.n4947 avss -2.33e-19
C7750 avdd.n4948 avss -1.8e-19
C7751 avdd.n4949 avss -1.48e-19
C7752 avdd.n4950 avss -8.47e-19
C7753 avdd.n4951 avss 0.00357f
C7754 avdd.n4952 avss 0.0348f
C7755 avdd.n4953 avss -0.00137f
C7756 avdd.n4954 avss -6.46e-19
C7757 avdd.n4955 avss 0.0189f
C7758 avdd.n4956 avss -3.07e-19
C7759 avdd.n4957 avss -2.01e-19
C7760 avdd.n4958 avss -3.28e-19
C7761 avdd.n4959 avss -3.28e-19
C7762 avdd.n4960 avss -8.47e-19
C7763 avdd.n4961 avss 0.0398f
C7764 avdd.n4962 avss -3.07e-19
C7765 avdd.n4963 avss 0.0181f
C7766 avdd.n4964 avss 0.0167f
C7767 avdd.n4965 avss 0.00875f
C7768 avdd.n4966 avss -2.54e-19
C7769 avdd.n4967 avss -2.54e-19
C7770 avdd.n4968 avss -2.22e-19
C7771 avdd.n4969 avss 0.0192f
C7772 avdd.n4970 avss -4.76e-19
C7773 avdd.n4971 avss -0.00128f
C7774 avdd.n4972 avss 0.0346f
C7775 avdd.n4973 avss -8.47e-19
C7776 avdd.n4974 avss 0.0388f
C7777 avdd.n4975 avss -8.47e-19
C7778 avdd.n4976 avss 0.0049f
C7779 avdd.n4977 avss 3e-19
C7780 avdd.n4978 avss -8.47e-19
C7781 avdd.n4979 avss -3.39e-19
C7782 avdd.n4980 avss -2.33e-19
C7783 avdd.n4981 avss -1.16e-19
C7784 avdd.n4982 avss 0.0182f
C7785 avdd.n4983 avss 0.0148f
C7786 avdd.n4984 avss 0.00875f
C7787 avdd.n4985 avss -2.22e-19
C7788 avdd.n4986 avss -2.22e-19
C7789 avdd.n4987 avss -1.8e-19
C7790 avdd.n4988 avss -1.8e-19
C7791 avdd.n4989 avss -1.59e-19
C7792 avdd.n4990 avss 0.0192f
C7793 avdd.n4991 avss -3.07e-19
C7794 avdd.n4992 avss -6.46e-19
C7795 avdd.n4993 avss -5.82e-19
C7796 avdd.n4994 avss -8.47e-19
C7797 avdd.n4995 avss -3.39e-19
C7798 avdd.n4996 avss -3.18e-19
C7799 avdd.n4997 avss -2.01e-19
C7800 avdd.n4998 avss 0.0183f
C7801 avdd.n4999 avss 0.0154f
C7802 avdd.n5000 avss 0.0154f
C7803 avdd.n5001 avss -1.8e-19
C7804 avdd.n5002 avss 0.0191f
C7805 avdd.n5003 avss -1.8e-19
C7806 avdd.n5004 avss -2.44e-19
C7807 avdd.n5005 avss -1.8e-19
C7808 avdd.n5006 avss -1.8e-19
C7809 avdd.n5007 avss -1.38e-19
C7810 avdd.n5008 avss -3.49e-19
C7811 avdd.n5009 avss 0.0184f
C7812 avdd.n5010 avss 0.00873f
C7813 avdd.n5011 avss 0.0422f
C7814 avdd.n5012 avss 0.00203f
C7815 avdd.n5013 avss 0.019f
C7816 avdd.n5014 avss -1.8e-19
C7817 avdd.n5015 avss -1.48e-19
C7818 avdd.n5016 avss -2.33e-19
C7819 avdd.n5017 avss -2.33e-19
C7820 avdd.n5018 avss -2.44e-19
C7821 avdd.n5019 avss 0.0197f
C7822 avdd.n5020 avss 0.0384f
C7823 avdd.n5021 avss -0.00512f
C7824 avdd.n5023 avss 0.0382f
C7825 avdd.n5024 avss -0.168f
C7826 avdd.n5025 avss -0.203f
C7827 avdd.n5026 avss 0.0269f
C7828 avdd.n5027 avss -1.27e-19
C7829 avdd.n5028 avss -2.96e-19
C7830 avdd.n5029 avss -0.00113f
C7831 avdd.n5031 avss -1.8e-19
C7832 avdd.n5032 avss -8.47e-19
C7833 avdd.n5033 avss 0.00869f
C7834 avdd.n5035 avss -0.00173f
C7835 avdd.n5036 avss -2.44e-19
C7836 avdd.n5037 avss 0.0111f
C7837 avdd.n5038 avss -1.38e-19
C7838 avdd.n5039 avss -2.44e-19
C7839 avdd.n5040 avss 0.0111f
C7840 avdd.n5041 avss -1.8e-19
C7841 avdd.n5042 avss -1.8e-19
C7842 avdd.n5043 avss 0.00908f
C7843 avdd.n5044 avss 0.03f
C7844 avdd.n5045 avss -3.39e-19
C7845 avdd.n5046 avss -3.39e-19
C7846 avdd.n5047 avss -1.59e-19
C7847 avdd.n5048 avss 0.0111f
C7848 avdd.n5049 avss -1.8e-19
C7849 avdd.n5050 avss -1.8e-19
C7850 avdd.n5051 avss 0.0342f
C7851 avdd.n5052 avss 0.00378f
C7852 avdd.n5053 avss -5.77e-19
C7853 avdd.n5054 avss -2.22e-19
C7854 avdd.n5055 avss 0.0168f
C7855 avdd.n5056 avss -3.6e-19
C7856 avdd.n5057 avss -1.8e-19
C7857 avdd.n5058 avss -8.26e-19
C7858 avdd.n5059 avss -0.0013f
C7859 avdd.n5060 avss -3.39e-19
C7860 avdd.n5061 avss -1.27e-19
C7861 avdd.n5062 avss 0.0022f
C7862 avdd.n5063 avss 0.019f
C7863 avdd.n5064 avss 0.0184f
C7864 avdd.n5065 avss -5.19e-19
C7865 avdd.n5066 avss 0.0386f
C7866 avdd.n5067 avss 0.0111f
C7867 avdd.n5068 avss -1.38e-19
C7868 avdd.n5069 avss -1.38e-19
C7869 avdd.n5070 avss -3.39e-19
C7870 avdd.n5071 avss -3.39e-19
C7871 avdd.n5072 avss -1.8e-19
C7872 avdd.n5073 avss 0.0411f
C7873 avdd.n5074 avss 0.0111f
C7874 avdd.n5075 avss -1.8e-19
C7875 avdd.n5076 avss -1.8e-19
C7876 avdd.n5077 avss -0.00173f
C7877 avdd.n5078 avss -0.00122f
C7878 avdd.n5079 avss -2.96e-19
C7879 avdd.n5080 avss -0.00121f
C7880 avdd.n5081 avss -6.35e-19
C7881 avdd.n5082 avss -0.00357f
C7882 avdd.n5083 avss -0.00109f
C7883 avdd.n5084 avss 0.0374f
C7884 avdd.n5085 avss 0.0112f
C7885 avdd.n5086 avss -1.8e-19
C7886 avdd.n5087 avss -1.8e-19
C7887 avdd.n5088 avss -0.00126f
C7888 avdd.n5089 avss 0.0318f
C7889 avdd.n5090 avss -0.00139f
C7890 avdd.n5091 avss -2.22e-19
C7891 avdd.n5092 avss 0.0188f
C7892 avdd.n5093 avss -2.75e-19
C7893 avdd.n5094 avss -3.6e-19
C7894 avdd.n5095 avss -3.07e-19
C7895 avdd.n5096 avss -6.88e-19
C7896 avdd.n5097 avss 0.00725f
C7897 avdd.n5098 avss -0.00336f
C7898 avdd.n5099 avss -1.8e-19
C7899 avdd.n5100 avss -2.01e-19
C7900 avdd.n5101 avss -0.0866f
C7901 avdd.n5102 avss 0.0179f
C7902 avdd.n5103 avss 0.0442f
C7903 avdd.n5104 avss -3.39e-19
C7904 avdd.n5105 avss -2.75e-19
C7905 avdd.n5106 avss 0.0181f
C7906 avdd.n5107 avss 0.00821f
C7907 avdd.n5108 avss 0.00821f
C7908 avdd.n5109 avss -2.75e-19
C7909 avdd.n5110 avss -2.33e-19
C7910 avdd.n5111 avss -2.54e-19
C7911 avdd.n5112 avss -2.54e-19
C7912 avdd.n5113 avss -2.22e-19
C7913 avdd.n5114 avss -1.59e-19
C7914 avdd.n5115 avss 0.0298f
C7915 avdd.n5116 avss 0.0098f
C7916 avdd.n5117 avss -0.00158f
C7917 avdd.n5118 avss -8.47e-19
C7918 avdd.n5119 avss -4.23e-19
C7919 avdd.n5120 avss -3.39e-19
C7920 avdd.n5121 avss -2.33e-19
C7921 avdd.n5122 avss -1.16e-19
C7922 avdd.n5123 avss 0.0182f
C7923 avdd.n5124 avss 0.0148f
C7924 avdd.n5125 avss 0.00875f
C7925 avdd.n5126 avss -2.22e-19
C7926 avdd.n5127 avss -2.22e-19
C7927 avdd.n5128 avss 0.00358f
C7928 avdd.n5129 avss -1.8e-19
C7929 avdd.n5130 avss -1.59e-19
C7930 avdd.n5131 avss 0.0192f
C7931 avdd.n5132 avss -3.07e-19
C7932 avdd.n5133 avss -0.00108f
C7933 avdd.n5134 avss 0.0382f
C7934 avdd.n5135 avss -9.76e-19
C7935 avdd.n5136 avss -2.01e-19
C7936 avdd.n5137 avss 0.0183f
C7937 avdd.n5138 avss 0.0154f
C7938 avdd.n5139 avss 0.0154f
C7939 avdd.n5140 avss 0.0191f
C7940 avdd.n5141 avss -1.8e-19
C7941 avdd.n5142 avss -1.8e-19
C7942 avdd.n5143 avss -2.44e-19
C7943 avdd.n5144 avss -1.8e-19
C7944 avdd.n5145 avss -1.8e-19
C7945 avdd.n5146 avss -5.61e-19
C7946 avdd.n5147 avss 0.0344f
C7947 avdd.n5148 avss -2.44e-19
C7948 avdd.n5149 avss -8.47e-19
C7949 avdd.n5150 avss -8.15e-19
C7950 avdd.n5151 avss -0.0014f
C7951 avdd.n5152 avss -8.47e-19
C7952 avdd.n5153 avss 0.00466f
C7953 avdd.n5154 avss -3.39e-19
C7954 avdd.n5155 avss -6.67e-19
C7955 avdd.n5156 avss -3.49e-19
C7956 avdd.n5157 avss 0.0184f
C7957 avdd.n5158 avss 0.00873f
C7958 avdd.n5159 avss 0.0148f
C7959 avdd.n5160 avss 0.00873f
C7960 avdd.n5161 avss 0.0111f
C7961 avdd.n5162 avss -2.44e-19
C7962 avdd.n5163 avss -2.33e-19
C7963 avdd.n5164 avss -1.8e-19
C7964 avdd.n5165 avss -1.48e-19
C7965 avdd.n5166 avss -8.47e-19
C7966 avdd.n5167 avss 0.00357f
C7967 avdd.n5168 avss 0.0348f
C7968 avdd.n5169 avss -0.00137f
C7969 avdd.n5170 avss -6.46e-19
C7970 avdd.n5171 avss 0.0189f
C7971 avdd.n5172 avss -3.07e-19
C7972 avdd.n5173 avss -2.01e-19
C7973 avdd.n5174 avss -3.28e-19
C7974 avdd.n5175 avss -3.28e-19
C7975 avdd.n5176 avss -8.47e-19
C7976 avdd.n5177 avss 0.0398f
C7977 avdd.n5178 avss -3.07e-19
C7978 avdd.n5179 avss 0.0181f
C7979 avdd.n5180 avss 0.0167f
C7980 avdd.n5181 avss 0.00875f
C7981 avdd.n5182 avss -2.54e-19
C7982 avdd.n5183 avss -2.54e-19
C7983 avdd.n5184 avss -2.22e-19
C7984 avdd.n5185 avss 0.0192f
C7985 avdd.n5186 avss -4.76e-19
C7986 avdd.n5187 avss -0.00128f
C7987 avdd.n5188 avss 0.0346f
C7988 avdd.n5189 avss -8.47e-19
C7989 avdd.n5190 avss 0.0388f
C7990 avdd.n5191 avss -8.47e-19
C7991 avdd.n5192 avss 0.0049f
C7992 avdd.n5193 avss 3e-19
C7993 avdd.n5194 avss -8.47e-19
C7994 avdd.n5195 avss -3.39e-19
C7995 avdd.n5196 avss -2.33e-19
C7996 avdd.n5197 avss -1.16e-19
C7997 avdd.n5198 avss 0.0182f
C7998 avdd.n5199 avss 0.0148f
C7999 avdd.n5200 avss 0.00875f
C8000 avdd.n5201 avss -2.22e-19
C8001 avdd.n5202 avss -2.22e-19
C8002 avdd.n5203 avss -1.8e-19
C8003 avdd.n5204 avss -1.8e-19
C8004 avdd.n5205 avss -1.59e-19
C8005 avdd.n5206 avss 0.0192f
C8006 avdd.n5207 avss -3.07e-19
C8007 avdd.n5208 avss -6.46e-19
C8008 avdd.n5209 avss -5.82e-19
C8009 avdd.n5210 avss -8.47e-19
C8010 avdd.n5211 avss -3.39e-19
C8011 avdd.n5212 avss -3.18e-19
C8012 avdd.n5213 avss -2.01e-19
C8013 avdd.n5214 avss 0.0183f
C8014 avdd.n5215 avss 0.0154f
C8015 avdd.n5216 avss 0.0154f
C8016 avdd.n5217 avss -1.8e-19
C8017 avdd.n5218 avss 0.0191f
C8018 avdd.n5219 avss -1.8e-19
C8019 avdd.n5220 avss -2.44e-19
C8020 avdd.n5221 avss -1.8e-19
C8021 avdd.n5222 avss -1.8e-19
C8022 avdd.n5223 avss -1.38e-19
C8023 avdd.n5224 avss -3.49e-19
C8024 avdd.n5225 avss 0.0184f
C8025 avdd.n5226 avss 0.00873f
C8026 avdd.n5227 avss 0.0422f
C8027 avdd.n5228 avss 0.00203f
C8028 avdd.n5229 avss 0.019f
C8029 avdd.n5230 avss -1.8e-19
C8030 avdd.n5231 avss -1.48e-19
C8031 avdd.n5232 avss -2.33e-19
C8032 avdd.n5233 avss -2.33e-19
C8033 avdd.n5234 avss -2.44e-19
C8034 avdd.n5235 avss 0.0197f
C8035 avdd.n5236 avss 0.0384f
C8036 avdd.n5237 avss -0.00512f
C8037 avdd.n5239 avss 0.0382f
C8038 avdd.n5240 avss -0.168f
C8039 avdd.n5241 avss -0.202f
C8040 avdd.n5242 avss 0.0269f
C8041 avdd.n5243 avss -1.27e-19
C8042 avdd.n5244 avss -2.96e-19
C8043 avdd.n5245 avss -0.00113f
C8044 avdd.n5247 avss -1.8e-19
C8045 avdd.n5248 avss -8.47e-19
C8046 avdd.n5249 avss 0.00869f
C8047 avdd.n5251 avss -0.00173f
C8048 avdd.n5252 avss -2.44e-19
C8049 avdd.n5253 avss 0.0111f
C8050 avdd.n5254 avss -1.38e-19
C8051 avdd.n5255 avss -2.44e-19
C8052 avdd.n5256 avss 0.0111f
C8053 avdd.n5257 avss -1.8e-19
C8054 avdd.n5258 avss -1.8e-19
C8055 avdd.n5259 avss 0.00908f
C8056 avdd.n5260 avss 0.03f
C8057 avdd.n5261 avss -3.39e-19
C8058 avdd.n5262 avss -3.39e-19
C8059 avdd.n5263 avss -1.59e-19
C8060 avdd.n5264 avss 0.0111f
C8061 avdd.n5265 avss -1.8e-19
C8062 avdd.n5266 avss -1.8e-19
C8063 avdd.n5267 avss 0.0342f
C8064 avdd.n5268 avss 0.00378f
C8065 avdd.n5269 avss -5.77e-19
C8066 avdd.n5270 avss -2.22e-19
C8067 avdd.n5271 avss 0.0168f
C8068 avdd.n5272 avss -3.6e-19
C8069 avdd.n5273 avss -1.8e-19
C8070 avdd.n5274 avss -8.26e-19
C8071 avdd.n5275 avss -0.0013f
C8072 avdd.n5276 avss -3.39e-19
C8073 avdd.n5277 avss -1.27e-19
C8074 avdd.n5278 avss 0.0022f
C8075 avdd.n5279 avss 0.019f
C8076 avdd.n5280 avss 0.0184f
C8077 avdd.n5281 avss -5.19e-19
C8078 avdd.n5282 avss 0.0386f
C8079 avdd.n5283 avss 0.0111f
C8080 avdd.n5284 avss -1.38e-19
C8081 avdd.n5285 avss -1.38e-19
C8082 avdd.n5286 avss -3.39e-19
C8083 avdd.n5287 avss -3.39e-19
C8084 avdd.n5288 avss -1.8e-19
C8085 avdd.n5289 avss 0.0411f
C8086 avdd.n5290 avss 0.0111f
C8087 avdd.n5291 avss -1.8e-19
C8088 avdd.n5292 avss -1.8e-19
C8089 avdd.n5293 avss -0.00173f
C8090 avdd.n5294 avss -0.00122f
C8091 avdd.n5295 avss -2.96e-19
C8092 avdd.n5296 avss -0.00121f
C8093 avdd.n5297 avss -6.35e-19
C8094 avdd.n5298 avss -0.00357f
C8095 avdd.n5299 avss -0.00109f
C8096 avdd.n5300 avss 0.0374f
C8097 avdd.n5301 avss 0.0112f
C8098 avdd.n5302 avss -1.8e-19
C8099 avdd.n5303 avss -1.8e-19
C8100 avdd.n5304 avss -0.00126f
C8101 avdd.n5305 avss 0.0318f
C8102 avdd.n5306 avss -0.00139f
C8103 avdd.n5307 avss -2.22e-19
C8104 avdd.n5308 avss 0.0188f
C8105 avdd.n5309 avss -2.75e-19
C8106 avdd.n5310 avss -3.6e-19
C8107 avdd.n5311 avss -3.07e-19
C8108 avdd.n5312 avss -6.88e-19
C8109 avdd.n5313 avss 0.00725f
C8110 avdd.n5314 avss -0.00336f
C8111 avdd.n5315 avss -1.8e-19
C8112 avdd.n5316 avss -2.01e-19
C8113 avdd.n5317 avss -0.0866f
C8114 avdd.n5318 avss 0.0179f
C8115 avdd.n5319 avss 0.0442f
C8116 avdd.n5320 avss -3.39e-19
C8117 avdd.n5321 avss -2.75e-19
C8118 avdd.n5322 avss 0.0181f
C8119 avdd.n5323 avss 0.00821f
C8120 avdd.n5324 avss 0.00821f
C8121 avdd.n5325 avss -2.75e-19
C8122 avdd.n5326 avss -2.33e-19
C8123 avdd.n5327 avss -2.54e-19
C8124 avdd.n5328 avss -2.54e-19
C8125 avdd.n5329 avss -2.22e-19
C8126 avdd.n5330 avss -1.59e-19
C8127 avdd.n5331 avss 0.0298f
C8128 avdd.n5332 avss 0.0098f
C8129 avdd.n5333 avss -0.00158f
C8130 avdd.n5334 avss -8.47e-19
C8131 avdd.n5335 avss -4.23e-19
C8132 avdd.n5336 avss -3.39e-19
C8133 avdd.n5337 avss -2.33e-19
C8134 avdd.n5338 avss -1.16e-19
C8135 avdd.n5339 avss 0.0182f
C8136 avdd.n5340 avss 0.0148f
C8137 avdd.n5341 avss 0.00875f
C8138 avdd.n5342 avss -2.22e-19
C8139 avdd.n5343 avss -2.22e-19
C8140 avdd.n5344 avss 0.00358f
C8141 avdd.n5345 avss -1.8e-19
C8142 avdd.n5346 avss -1.59e-19
C8143 avdd.n5347 avss 0.0192f
C8144 avdd.n5348 avss -3.07e-19
C8145 avdd.n5349 avss -0.00108f
C8146 avdd.n5350 avss 0.0382f
C8147 avdd.n5351 avss -9.76e-19
C8148 avdd.n5352 avss -2.01e-19
C8149 avdd.n5353 avss 0.0183f
C8150 avdd.n5354 avss 0.0154f
C8151 avdd.n5355 avss 0.0154f
C8152 avdd.n5356 avss 0.0191f
C8153 avdd.n5357 avss -1.8e-19
C8154 avdd.n5358 avss -1.8e-19
C8155 avdd.n5359 avss -2.44e-19
C8156 avdd.n5360 avss -1.8e-19
C8157 avdd.n5361 avss -1.8e-19
C8158 avdd.n5362 avss -5.61e-19
C8159 avdd.n5363 avss 0.0344f
C8160 avdd.n5364 avss -2.44e-19
C8161 avdd.n5365 avss -8.47e-19
C8162 avdd.n5366 avss -8.15e-19
C8163 avdd.n5367 avss -0.0014f
C8164 avdd.n5368 avss -8.47e-19
C8165 avdd.n5369 avss 0.00466f
C8166 avdd.n5370 avss -3.39e-19
C8167 avdd.n5371 avss -6.67e-19
C8168 avdd.n5372 avss -3.49e-19
C8169 avdd.n5373 avss 0.0184f
C8170 avdd.n5374 avss 0.00873f
C8171 avdd.n5375 avss 0.0148f
C8172 avdd.n5376 avss 0.00873f
C8173 avdd.n5377 avss 0.0111f
C8174 avdd.n5378 avss -2.44e-19
C8175 avdd.n5379 avss -2.33e-19
C8176 avdd.n5380 avss -1.8e-19
C8177 avdd.n5381 avss -1.48e-19
C8178 avdd.n5382 avss -8.47e-19
C8179 avdd.n5383 avss 0.00357f
C8180 avdd.n5384 avss 0.0348f
C8181 avdd.n5385 avss -0.00137f
C8182 avdd.n5386 avss -6.46e-19
C8183 avdd.n5387 avss 0.0189f
C8184 avdd.n5388 avss -3.07e-19
C8185 avdd.n5389 avss -2.01e-19
C8186 avdd.n5390 avss -3.28e-19
C8187 avdd.n5391 avss -3.28e-19
C8188 avdd.n5392 avss -8.47e-19
C8189 avdd.n5393 avss 0.0398f
C8190 avdd.n5394 avss -3.07e-19
C8191 avdd.n5395 avss 0.0181f
C8192 avdd.n5396 avss 0.0167f
C8193 avdd.n5397 avss 0.00875f
C8194 avdd.n5398 avss -2.54e-19
C8195 avdd.n5399 avss -2.54e-19
C8196 avdd.n5400 avss -2.22e-19
C8197 avdd.n5401 avss 0.0192f
C8198 avdd.n5402 avss -4.76e-19
C8199 avdd.n5403 avss -0.00128f
C8200 avdd.n5404 avss 0.0346f
C8201 avdd.n5405 avss -8.47e-19
C8202 avdd.n5406 avss 0.0388f
C8203 avdd.n5407 avss -8.47e-19
C8204 avdd.n5408 avss 0.0049f
C8205 avdd.n5409 avss 3e-19
C8206 avdd.n5410 avss -8.47e-19
C8207 avdd.n5411 avss -3.39e-19
C8208 avdd.n5412 avss -2.33e-19
C8209 avdd.n5413 avss -1.16e-19
C8210 avdd.n5414 avss 0.0182f
C8211 avdd.n5415 avss 0.0148f
C8212 avdd.n5416 avss 0.00875f
C8213 avdd.n5417 avss -2.22e-19
C8214 avdd.n5418 avss -2.22e-19
C8215 avdd.n5419 avss -1.8e-19
C8216 avdd.n5420 avss -1.8e-19
C8217 avdd.n5421 avss -1.59e-19
C8218 avdd.n5422 avss 0.0192f
C8219 avdd.n5423 avss -3.07e-19
C8220 avdd.n5424 avss -6.46e-19
C8221 avdd.n5425 avss -5.82e-19
C8222 avdd.n5426 avss -8.47e-19
C8223 avdd.n5427 avss -3.39e-19
C8224 avdd.n5428 avss -3.18e-19
C8225 avdd.n5429 avss -2.01e-19
C8226 avdd.n5430 avss 0.0183f
C8227 avdd.n5431 avss 0.0154f
C8228 avdd.n5432 avss 0.0154f
C8229 avdd.n5433 avss -1.8e-19
C8230 avdd.n5434 avss 0.0191f
C8231 avdd.n5435 avss -1.8e-19
C8232 avdd.n5436 avss -2.44e-19
C8233 avdd.n5437 avss -1.8e-19
C8234 avdd.n5438 avss -1.8e-19
C8235 avdd.n5439 avss -1.38e-19
C8236 avdd.n5440 avss -3.49e-19
C8237 avdd.n5441 avss 0.0184f
C8238 avdd.n5442 avss 0.00873f
C8239 avdd.n5443 avss 0.0422f
C8240 avdd.n5444 avss 0.00203f
C8241 avdd.n5445 avss 0.019f
C8242 avdd.n5446 avss -1.8e-19
C8243 avdd.n5447 avss -1.48e-19
C8244 avdd.n5448 avss -2.33e-19
C8245 avdd.n5449 avss -2.33e-19
C8246 avdd.n5450 avss -2.44e-19
C8247 avdd.n5451 avss 0.0197f
C8248 avdd.n5452 avss 0.0384f
C8249 avdd.n5453 avss -0.00512f
C8250 avdd.n5455 avss 0.0382f
C8251 avdd.n5456 avss -0.166f
C8252 avdd.n5457 avss -0.202f
C8253 avdd.n5458 avss 0.0269f
C8254 avdd.n5459 avss -1.27e-19
C8255 avdd.n5460 avss -2.96e-19
C8256 avdd.n5461 avss -0.00113f
C8257 avdd.n5463 avss -1.8e-19
C8258 avdd.n5464 avss -8.47e-19
C8259 avdd.n5465 avss 0.00869f
C8260 avdd.n5467 avss -0.00173f
C8261 avdd.n5468 avss -2.44e-19
C8262 avdd.n5469 avss 0.0111f
C8263 avdd.n5470 avss -1.38e-19
C8264 avdd.n5471 avss -2.44e-19
C8265 avdd.n5472 avss 0.0111f
C8266 avdd.n5473 avss -1.8e-19
C8267 avdd.n5474 avss -1.8e-19
C8268 avdd.n5475 avss 0.00908f
C8269 avdd.n5476 avss 0.03f
C8270 avdd.n5477 avss -3.39e-19
C8271 avdd.n5478 avss -3.39e-19
C8272 avdd.n5479 avss -1.59e-19
C8273 avdd.n5480 avss 0.0111f
C8274 avdd.n5481 avss -1.8e-19
C8275 avdd.n5482 avss -1.8e-19
C8276 avdd.n5483 avss 0.0342f
C8277 avdd.n5484 avss 0.00378f
C8278 avdd.n5485 avss -5.77e-19
C8279 avdd.n5486 avss -2.22e-19
C8280 avdd.n5487 avss 0.0168f
C8281 avdd.n5488 avss -3.6e-19
C8282 avdd.n5489 avss -1.8e-19
C8283 avdd.n5490 avss -8.26e-19
C8284 avdd.n5491 avss -0.0013f
C8285 avdd.n5492 avss -3.39e-19
C8286 avdd.n5493 avss -1.27e-19
C8287 avdd.n5494 avss 0.0022f
C8288 avdd.n5495 avss 0.019f
C8289 avdd.n5496 avss 0.0184f
C8290 avdd.n5497 avss -5.19e-19
C8291 avdd.n5498 avss 0.0386f
C8292 avdd.n5499 avss 0.0111f
C8293 avdd.n5500 avss -1.38e-19
C8294 avdd.n5501 avss -1.38e-19
C8295 avdd.n5502 avss -3.39e-19
C8296 avdd.n5503 avss -3.39e-19
C8297 avdd.n5504 avss -1.8e-19
C8298 avdd.n5505 avss 0.0411f
C8299 avdd.n5506 avss 0.0111f
C8300 avdd.n5507 avss -1.8e-19
C8301 avdd.n5508 avss -1.8e-19
C8302 avdd.n5509 avss -0.00173f
C8303 avdd.n5510 avss -0.00122f
C8304 avdd.n5511 avss -2.96e-19
C8305 avdd.n5512 avss -0.00121f
C8306 avdd.n5513 avss -6.35e-19
C8307 avdd.n5514 avss -0.00357f
C8308 avdd.n5515 avss -0.00109f
C8309 avdd.n5516 avss 0.0374f
C8310 avdd.n5517 avss 0.0112f
C8311 avdd.n5518 avss -1.8e-19
C8312 avdd.n5519 avss -1.8e-19
C8313 avdd.n5520 avss -0.00126f
C8314 avdd.n5521 avss 0.0318f
C8315 avdd.n5522 avss -0.00139f
C8316 avdd.n5523 avss -2.22e-19
C8317 avdd.n5524 avss 0.0188f
C8318 avdd.n5525 avss -2.75e-19
C8319 avdd.n5526 avss -3.6e-19
C8320 avdd.n5527 avss -3.07e-19
C8321 avdd.n5528 avss -6.88e-19
C8322 avdd.n5529 avss 0.00725f
C8323 avdd.n5530 avss -0.00336f
C8324 avdd.n5531 avss -1.8e-19
C8325 avdd.n5532 avss -2.01e-19
C8326 avdd.n5533 avss -0.0866f
C8327 avdd.n5534 avss 0.0179f
C8328 avdd.n5535 avss 0.0442f
C8329 avdd.n5536 avss -3.39e-19
C8330 avdd.n5537 avss -2.75e-19
C8331 avdd.n5538 avss 0.0181f
C8332 avdd.n5539 avss 0.00821f
C8333 avdd.n5540 avss 0.00821f
C8334 avdd.n5541 avss -2.75e-19
C8335 avdd.n5542 avss -2.33e-19
C8336 avdd.n5543 avss -2.54e-19
C8337 avdd.n5544 avss -2.54e-19
C8338 avdd.n5545 avss -2.22e-19
C8339 avdd.n5546 avss -1.59e-19
C8340 avdd.n5547 avss 0.0298f
C8341 avdd.n5548 avss 0.0098f
C8342 avdd.n5549 avss -0.00158f
C8343 avdd.n5550 avss -8.47e-19
C8344 avdd.n5551 avss -4.23e-19
C8345 avdd.n5552 avss -3.39e-19
C8346 avdd.n5553 avss -2.33e-19
C8347 avdd.n5554 avss -1.16e-19
C8348 avdd.n5555 avss 0.0182f
C8349 avdd.n5556 avss 0.0148f
C8350 avdd.n5557 avss 0.00875f
C8351 avdd.n5558 avss -2.22e-19
C8352 avdd.n5559 avss -2.22e-19
C8353 avdd.n5560 avss 0.00358f
C8354 avdd.n5561 avss -1.8e-19
C8355 avdd.n5562 avss -1.59e-19
C8356 avdd.n5563 avss 0.0192f
C8357 avdd.n5564 avss -3.07e-19
C8358 avdd.n5565 avss -0.00108f
C8359 avdd.n5566 avss 0.0382f
C8360 avdd.n5567 avss -9.76e-19
C8361 avdd.n5568 avss -2.01e-19
C8362 avdd.n5569 avss 0.0183f
C8363 avdd.n5570 avss 0.0154f
C8364 avdd.n5571 avss 0.0154f
C8365 avdd.n5572 avss 0.0191f
C8366 avdd.n5573 avss -1.8e-19
C8367 avdd.n5574 avss -1.8e-19
C8368 avdd.n5575 avss -2.44e-19
C8369 avdd.n5576 avss -1.8e-19
C8370 avdd.n5577 avss -1.8e-19
C8371 avdd.n5578 avss -5.61e-19
C8372 avdd.n5579 avss 0.0344f
C8373 avdd.n5580 avss -2.44e-19
C8374 avdd.n5581 avss -8.47e-19
C8375 avdd.n5582 avss -8.15e-19
C8376 avdd.n5583 avss -0.0014f
C8377 avdd.n5584 avss -8.47e-19
C8378 avdd.n5585 avss 0.00466f
C8379 avdd.n5586 avss -3.39e-19
C8380 avdd.n5587 avss -6.67e-19
C8381 avdd.n5588 avss -3.49e-19
C8382 avdd.n5589 avss 0.0184f
C8383 avdd.n5590 avss 0.00873f
C8384 avdd.n5591 avss 0.0148f
C8385 avdd.n5592 avss 0.00873f
C8386 avdd.n5593 avss 0.0111f
C8387 avdd.n5594 avss -2.44e-19
C8388 avdd.n5595 avss -2.33e-19
C8389 avdd.n5596 avss -1.8e-19
C8390 avdd.n5597 avss -1.48e-19
C8391 avdd.n5598 avss -8.47e-19
C8392 avdd.n5599 avss 0.00357f
C8393 avdd.n5600 avss 0.0348f
C8394 avdd.n5601 avss -0.00137f
C8395 avdd.n5602 avss -6.46e-19
C8396 avdd.n5603 avss 0.0189f
C8397 avdd.n5604 avss -3.07e-19
C8398 avdd.n5605 avss -2.01e-19
C8399 avdd.n5606 avss -3.28e-19
C8400 avdd.n5607 avss -3.28e-19
C8401 avdd.n5608 avss -8.47e-19
C8402 avdd.n5609 avss 0.0398f
C8403 avdd.n5610 avss -3.07e-19
C8404 avdd.n5611 avss 0.0181f
C8405 avdd.n5612 avss 0.0167f
C8406 avdd.n5613 avss 0.00875f
C8407 avdd.n5614 avss -2.54e-19
C8408 avdd.n5615 avss -2.54e-19
C8409 avdd.n5616 avss -2.22e-19
C8410 avdd.n5617 avss 0.0192f
C8411 avdd.n5618 avss -4.76e-19
C8412 avdd.n5619 avss -0.00128f
C8413 avdd.n5620 avss 0.0346f
C8414 avdd.n5621 avss -8.47e-19
C8415 avdd.n5622 avss 0.0388f
C8416 avdd.n5623 avss -8.47e-19
C8417 avdd.n5624 avss 0.0049f
C8418 avdd.n5625 avss 3e-19
C8419 avdd.n5626 avss -8.47e-19
C8420 avdd.n5627 avss -3.39e-19
C8421 avdd.n5628 avss -2.33e-19
C8422 avdd.n5629 avss -1.16e-19
C8423 avdd.n5630 avss 0.0182f
C8424 avdd.n5631 avss 0.0148f
C8425 avdd.n5632 avss 0.00875f
C8426 avdd.n5633 avss -2.22e-19
C8427 avdd.n5634 avss -2.22e-19
C8428 avdd.n5635 avss -1.8e-19
C8429 avdd.n5636 avss -1.8e-19
C8430 avdd.n5637 avss -1.59e-19
C8431 avdd.n5638 avss 0.0192f
C8432 avdd.n5639 avss -3.07e-19
C8433 avdd.n5640 avss -6.46e-19
C8434 avdd.n5641 avss -5.82e-19
C8435 avdd.n5642 avss -8.47e-19
C8436 avdd.n5643 avss -3.39e-19
C8437 avdd.n5644 avss -3.18e-19
C8438 avdd.n5645 avss -2.01e-19
C8439 avdd.n5646 avss 0.0183f
C8440 avdd.n5647 avss 0.0154f
C8441 avdd.n5648 avss 0.0154f
C8442 avdd.n5649 avss -1.8e-19
C8443 avdd.n5650 avss 0.0191f
C8444 avdd.n5651 avss -1.8e-19
C8445 avdd.n5652 avss -2.44e-19
C8446 avdd.n5653 avss -1.8e-19
C8447 avdd.n5654 avss -1.8e-19
C8448 avdd.n5655 avss -1.38e-19
C8449 avdd.n5656 avss -3.49e-19
C8450 avdd.n5657 avss 0.0184f
C8451 avdd.n5658 avss 0.00873f
C8452 avdd.n5659 avss 0.0422f
C8453 avdd.n5660 avss 0.00203f
C8454 avdd.n5661 avss 0.019f
C8455 avdd.n5662 avss -1.8e-19
C8456 avdd.n5663 avss -1.48e-19
C8457 avdd.n5664 avss -2.33e-19
C8458 avdd.n5665 avss -2.33e-19
C8459 avdd.n5666 avss -2.44e-19
C8460 avdd.n5667 avss 0.0197f
C8461 avdd.n5668 avss 0.0384f
C8462 avdd.n5669 avss -0.00512f
C8463 avdd.n5671 avss 0.0382f
C8464 avdd.n5672 avss -0.166f
C8465 avdd.n5673 avss -0.202f
C8466 avdd.n5674 avss 0.0269f
C8467 avdd.n5675 avss -1.27e-19
C8468 avdd.n5676 avss -2.96e-19
C8469 avdd.n5677 avss -0.00113f
C8470 avdd.n5679 avss -1.8e-19
C8471 avdd.n5680 avss -8.47e-19
C8472 avdd.n5681 avss 0.00869f
C8473 avdd.n5683 avss -0.00173f
C8474 avdd.n5684 avss -2.44e-19
C8475 avdd.n5685 avss 0.0111f
C8476 avdd.n5686 avss -1.38e-19
C8477 avdd.n5687 avss -2.44e-19
C8478 avdd.n5688 avss 0.0111f
C8479 avdd.n5689 avss -1.8e-19
C8480 avdd.n5690 avss -1.8e-19
C8481 avdd.n5691 avss 0.00908f
C8482 avdd.n5692 avss 0.03f
C8483 avdd.n5693 avss -3.39e-19
C8484 avdd.n5694 avss -3.39e-19
C8485 avdd.n5695 avss -1.59e-19
C8486 avdd.n5696 avss 0.0111f
C8487 avdd.n5697 avss -1.8e-19
C8488 avdd.n5698 avss -1.8e-19
C8489 avdd.n5699 avss 0.0342f
C8490 avdd.n5700 avss 0.00378f
C8491 avdd.n5701 avss -5.77e-19
C8492 avdd.n5702 avss -2.22e-19
C8493 avdd.n5703 avss 0.0168f
C8494 avdd.n5704 avss -3.6e-19
C8495 avdd.n5705 avss -1.8e-19
C8496 avdd.n5706 avss -8.26e-19
C8497 avdd.n5707 avss -0.0013f
C8498 avdd.n5708 avss -3.39e-19
C8499 avdd.n5709 avss -1.27e-19
C8500 avdd.n5710 avss 0.0022f
C8501 avdd.n5711 avss 0.019f
C8502 avdd.n5712 avss 0.0184f
C8503 avdd.n5713 avss -5.19e-19
C8504 avdd.n5714 avss 0.0386f
C8505 avdd.n5715 avss 0.0111f
C8506 avdd.n5716 avss -1.38e-19
C8507 avdd.n5717 avss -1.38e-19
C8508 avdd.n5718 avss -3.39e-19
C8509 avdd.n5719 avss -3.39e-19
C8510 avdd.n5720 avss -1.8e-19
C8511 avdd.n5721 avss 0.0411f
C8512 avdd.n5722 avss 0.0111f
C8513 avdd.n5723 avss -1.8e-19
C8514 avdd.n5724 avss -1.8e-19
C8515 avdd.n5725 avss -0.00173f
C8516 avdd.n5726 avss -0.00122f
C8517 avdd.n5727 avss -2.96e-19
C8518 avdd.n5728 avss -0.00121f
C8519 avdd.n5729 avss -6.35e-19
C8520 avdd.n5730 avss -0.00357f
C8521 avdd.n5731 avss -0.00109f
C8522 avdd.n5732 avss 0.0374f
C8523 avdd.n5733 avss 0.0112f
C8524 avdd.n5734 avss -1.8e-19
C8525 avdd.n5735 avss -1.8e-19
C8526 avdd.n5736 avss -0.00126f
C8527 avdd.n5737 avss 0.0318f
C8528 avdd.n5738 avss -0.00139f
C8529 avdd.n5739 avss -2.22e-19
C8530 avdd.n5740 avss 0.0188f
C8531 avdd.n5741 avss -2.75e-19
C8532 avdd.n5742 avss -3.6e-19
C8533 avdd.n5743 avss -3.07e-19
C8534 avdd.n5744 avss -6.88e-19
C8535 avdd.n5745 avss 0.00725f
C8536 avdd.n5746 avss -0.00336f
C8537 avdd.n5747 avss -1.8e-19
C8538 avdd.n5748 avss -2.01e-19
C8539 avdd.n5749 avss -0.0866f
C8540 avdd.n5750 avss 0.0179f
C8541 avdd.n5751 avss 0.0442f
C8542 avdd.n5752 avss -3.39e-19
C8543 avdd.n5753 avss -2.75e-19
C8544 avdd.n5754 avss 0.0181f
C8545 avdd.n5755 avss 0.00821f
C8546 avdd.n5756 avss 0.00821f
C8547 avdd.n5757 avss -2.75e-19
C8548 avdd.n5758 avss -2.33e-19
C8549 avdd.n5759 avss -2.54e-19
C8550 avdd.n5760 avss -2.54e-19
C8551 avdd.n5761 avss -2.22e-19
C8552 avdd.n5762 avss -1.59e-19
C8553 avdd.n5763 avss 0.0298f
C8554 avdd.n5764 avss 0.0098f
C8555 avdd.n5765 avss -0.00158f
C8556 avdd.n5766 avss -8.47e-19
C8557 avdd.n5767 avss -4.23e-19
C8558 avdd.n5768 avss -3.39e-19
C8559 avdd.n5769 avss -2.33e-19
C8560 avdd.n5770 avss -1.16e-19
C8561 avdd.n5771 avss 0.0182f
C8562 avdd.n5772 avss 0.0148f
C8563 avdd.n5773 avss 0.00875f
C8564 avdd.n5774 avss -2.22e-19
C8565 avdd.n5775 avss -2.22e-19
C8566 avdd.n5776 avss 0.00358f
C8567 avdd.n5777 avss -1.8e-19
C8568 avdd.n5778 avss -1.59e-19
C8569 avdd.n5779 avss 0.0192f
C8570 avdd.n5780 avss -3.07e-19
C8571 avdd.n5781 avss -0.00108f
C8572 avdd.n5782 avss 0.0382f
C8573 avdd.n5783 avss -9.76e-19
C8574 avdd.n5784 avss -2.01e-19
C8575 avdd.n5785 avss 0.0183f
C8576 avdd.n5786 avss 0.0154f
C8577 avdd.n5787 avss 0.0154f
C8578 avdd.n5788 avss 0.0191f
C8579 avdd.n5789 avss -1.8e-19
C8580 avdd.n5790 avss -1.8e-19
C8581 avdd.n5791 avss -2.44e-19
C8582 avdd.n5792 avss -1.8e-19
C8583 avdd.n5793 avss -1.8e-19
C8584 avdd.n5794 avss -5.61e-19
C8585 avdd.n5795 avss 0.0344f
C8586 avdd.n5796 avss -2.44e-19
C8587 avdd.n5797 avss -8.47e-19
C8588 avdd.n5798 avss -8.15e-19
C8589 avdd.n5799 avss -0.0014f
C8590 avdd.n5800 avss -8.47e-19
C8591 avdd.n5801 avss 0.00466f
C8592 avdd.n5802 avss -3.39e-19
C8593 avdd.n5803 avss -6.67e-19
C8594 avdd.n5804 avss -3.49e-19
C8595 avdd.n5805 avss 0.0184f
C8596 avdd.n5806 avss 0.00873f
C8597 avdd.n5807 avss 0.0148f
C8598 avdd.n5808 avss 0.00873f
C8599 avdd.n5809 avss 0.0111f
C8600 avdd.n5810 avss -2.44e-19
C8601 avdd.n5811 avss -2.33e-19
C8602 avdd.n5812 avss -1.8e-19
C8603 avdd.n5813 avss -1.48e-19
C8604 avdd.n5814 avss -8.47e-19
C8605 avdd.n5815 avss 0.00357f
C8606 avdd.n5816 avss 0.0348f
C8607 avdd.n5817 avss -0.00137f
C8608 avdd.n5818 avss -6.46e-19
C8609 avdd.n5819 avss 0.0189f
C8610 avdd.n5820 avss -3.07e-19
C8611 avdd.n5821 avss -2.01e-19
C8612 avdd.n5822 avss -3.28e-19
C8613 avdd.n5823 avss -3.28e-19
C8614 avdd.n5824 avss -8.47e-19
C8615 avdd.n5825 avss 0.0398f
C8616 avdd.n5826 avss -3.07e-19
C8617 avdd.n5827 avss 0.0181f
C8618 avdd.n5828 avss 0.0167f
C8619 avdd.n5829 avss 0.00875f
C8620 avdd.n5830 avss -2.54e-19
C8621 avdd.n5831 avss -2.54e-19
C8622 avdd.n5832 avss -2.22e-19
C8623 avdd.n5833 avss 0.0192f
C8624 avdd.n5834 avss -4.76e-19
C8625 avdd.n5835 avss -0.00128f
C8626 avdd.n5836 avss 0.0346f
C8627 avdd.n5837 avss -8.47e-19
C8628 avdd.n5838 avss 0.0388f
C8629 avdd.n5839 avss -8.47e-19
C8630 avdd.n5840 avss 0.0049f
C8631 avdd.n5841 avss 3e-19
C8632 avdd.n5842 avss -8.47e-19
C8633 avdd.n5843 avss -3.39e-19
C8634 avdd.n5844 avss -2.33e-19
C8635 avdd.n5845 avss -1.16e-19
C8636 avdd.n5846 avss 0.0182f
C8637 avdd.n5847 avss 0.0148f
C8638 avdd.n5848 avss 0.00875f
C8639 avdd.n5849 avss -2.22e-19
C8640 avdd.n5850 avss -2.22e-19
C8641 avdd.n5851 avss -1.8e-19
C8642 avdd.n5852 avss -1.8e-19
C8643 avdd.n5853 avss -1.59e-19
C8644 avdd.n5854 avss 0.0192f
C8645 avdd.n5855 avss -3.07e-19
C8646 avdd.n5856 avss -6.46e-19
C8647 avdd.n5857 avss -5.82e-19
C8648 avdd.n5858 avss -8.47e-19
C8649 avdd.n5859 avss -3.39e-19
C8650 avdd.n5860 avss -3.18e-19
C8651 avdd.n5861 avss -2.01e-19
C8652 avdd.n5862 avss 0.0183f
C8653 avdd.n5863 avss 0.0154f
C8654 avdd.n5864 avss 0.0154f
C8655 avdd.n5865 avss -1.8e-19
C8656 avdd.n5866 avss 0.0191f
C8657 avdd.n5867 avss -1.8e-19
C8658 avdd.n5868 avss -2.44e-19
C8659 avdd.n5869 avss -1.8e-19
C8660 avdd.n5870 avss -1.8e-19
C8661 avdd.n5871 avss -1.38e-19
C8662 avdd.n5872 avss -3.49e-19
C8663 avdd.n5873 avss 0.0184f
C8664 avdd.n5874 avss 0.00873f
C8665 avdd.n5875 avss 0.0422f
C8666 avdd.n5876 avss 0.00203f
C8667 avdd.n5877 avss 0.019f
C8668 avdd.n5878 avss -1.8e-19
C8669 avdd.n5879 avss -1.48e-19
C8670 avdd.n5880 avss -2.33e-19
C8671 avdd.n5881 avss -2.33e-19
C8672 avdd.n5882 avss -2.44e-19
C8673 avdd.n5883 avss 0.0197f
C8674 avdd.n5884 avss 0.0384f
C8675 avdd.n5885 avss -0.00512f
C8676 avdd.n5887 avss 0.0382f
C8677 avdd.n5888 avss -0.166f
C8678 avdd.n5889 avss -0.202f
C8679 avdd.n5890 avss 0.0269f
C8680 avdd.n5891 avss -1.27e-19
C8681 avdd.n5892 avss -2.96e-19
C8682 avdd.n5893 avss -0.00113f
C8683 avdd.n5895 avss -1.8e-19
C8684 avdd.n5896 avss -8.47e-19
C8685 avdd.n5897 avss 0.00869f
C8686 avdd.n5899 avss -0.00173f
C8687 avdd.n5900 avss -2.44e-19
C8688 avdd.n5901 avss 0.0111f
C8689 avdd.n5902 avss -1.38e-19
C8690 avdd.n5903 avss -2.44e-19
C8691 avdd.n5904 avss 0.0111f
C8692 avdd.n5905 avss -1.8e-19
C8693 avdd.n5906 avss -1.8e-19
C8694 avdd.n5907 avss 0.00908f
C8695 avdd.n5908 avss 0.03f
C8696 avdd.n5909 avss -3.39e-19
C8697 avdd.n5910 avss -3.39e-19
C8698 avdd.n5911 avss -1.59e-19
C8699 avdd.n5912 avss 0.0111f
C8700 avdd.n5913 avss -1.8e-19
C8701 avdd.n5914 avss -1.8e-19
C8702 avdd.n5915 avss 0.0342f
C8703 avdd.n5916 avss 0.00378f
C8704 avdd.n5917 avss -5.77e-19
C8705 avdd.n5918 avss -2.22e-19
C8706 avdd.n5919 avss 0.0168f
C8707 avdd.n5920 avss -3.6e-19
C8708 avdd.n5921 avss -1.8e-19
C8709 avdd.n5922 avss -8.26e-19
C8710 avdd.n5923 avss -0.0013f
C8711 avdd.n5924 avss -3.39e-19
C8712 avdd.n5925 avss -1.27e-19
C8713 avdd.n5926 avss 0.0022f
C8714 avdd.n5927 avss 0.019f
C8715 avdd.n5928 avss 0.0184f
C8716 avdd.n5929 avss -5.19e-19
C8717 avdd.n5930 avss 0.0386f
C8718 avdd.n5931 avss 0.0111f
C8719 avdd.n5932 avss -1.38e-19
C8720 avdd.n5933 avss -1.38e-19
C8721 avdd.n5934 avss -3.39e-19
C8722 avdd.n5935 avss -3.39e-19
C8723 avdd.n5936 avss -1.8e-19
C8724 avdd.n5937 avss 0.0411f
C8725 avdd.n5938 avss 0.0111f
C8726 avdd.n5939 avss -1.8e-19
C8727 avdd.n5940 avss -1.8e-19
C8728 avdd.n5941 avss -0.00173f
C8729 avdd.n5942 avss -0.00122f
C8730 avdd.n5943 avss -2.96e-19
C8731 avdd.n5944 avss -0.00121f
C8732 avdd.n5945 avss -6.35e-19
C8733 avdd.n5946 avss -0.00357f
C8734 avdd.n5947 avss -0.00109f
C8735 avdd.n5948 avss 0.0374f
C8736 avdd.n5949 avss 0.0112f
C8737 avdd.n5950 avss -1.8e-19
C8738 avdd.n5951 avss -1.8e-19
C8739 avdd.n5952 avss -0.00126f
C8740 avdd.n5953 avss 0.0318f
C8741 avdd.n5954 avss -0.00139f
C8742 avdd.n5955 avss -2.22e-19
C8743 avdd.n5956 avss 0.0188f
C8744 avdd.n5957 avss -2.75e-19
C8745 avdd.n5958 avss -3.6e-19
C8746 avdd.n5959 avss -3.07e-19
C8747 avdd.n5960 avss -6.88e-19
C8748 avdd.n5961 avss 0.00725f
C8749 avdd.n5962 avss -0.00336f
C8750 avdd.n5963 avss -1.8e-19
C8751 avdd.n5964 avss -2.01e-19
C8752 avdd.n5965 avss -0.0866f
C8753 avdd.n5966 avss 0.0179f
C8754 avdd.n5967 avss 0.0442f
C8755 avdd.n5968 avss -3.39e-19
C8756 avdd.n5969 avss -2.75e-19
C8757 avdd.n5970 avss 0.0181f
C8758 avdd.n5971 avss 0.00821f
C8759 avdd.n5972 avss 0.00821f
C8760 avdd.n5973 avss -2.75e-19
C8761 avdd.n5974 avss -2.33e-19
C8762 avdd.n5975 avss -2.54e-19
C8763 avdd.n5976 avss -2.54e-19
C8764 avdd.n5977 avss -2.22e-19
C8765 avdd.n5978 avss -1.59e-19
C8766 avdd.n5979 avss 0.0298f
C8767 avdd.n5980 avss 0.0098f
C8768 avdd.n5981 avss -0.00158f
C8769 avdd.n5982 avss -8.47e-19
C8770 avdd.n5983 avss -4.23e-19
C8771 avdd.n5984 avss -3.39e-19
C8772 avdd.n5985 avss -2.33e-19
C8773 avdd.n5986 avss -1.16e-19
C8774 avdd.n5987 avss 0.0182f
C8775 avdd.n5988 avss 0.0148f
C8776 avdd.n5989 avss 0.00875f
C8777 avdd.n5990 avss -2.22e-19
C8778 avdd.n5991 avss -2.22e-19
C8779 avdd.n5992 avss 0.00358f
C8780 avdd.n5993 avss -1.8e-19
C8781 avdd.n5994 avss -1.59e-19
C8782 avdd.n5995 avss 0.0192f
C8783 avdd.n5996 avss -3.07e-19
C8784 avdd.n5997 avss -0.00108f
C8785 avdd.n5998 avss 0.0382f
C8786 avdd.n5999 avss -9.76e-19
C8787 avdd.n6000 avss -2.01e-19
C8788 avdd.n6001 avss 0.0183f
C8789 avdd.n6002 avss 0.0154f
C8790 avdd.n6003 avss 0.0154f
C8791 avdd.n6004 avss 0.0191f
C8792 avdd.n6005 avss -1.8e-19
C8793 avdd.n6006 avss -1.8e-19
C8794 avdd.n6007 avss -2.44e-19
C8795 avdd.n6008 avss -1.8e-19
C8796 avdd.n6009 avss -1.8e-19
C8797 avdd.n6010 avss -5.61e-19
C8798 avdd.n6011 avss 0.0344f
C8799 avdd.n6012 avss -2.44e-19
C8800 avdd.n6013 avss -8.47e-19
C8801 avdd.n6014 avss -8.15e-19
C8802 avdd.n6015 avss -0.0014f
C8803 avdd.n6016 avss -8.47e-19
C8804 avdd.n6017 avss 0.00466f
C8805 avdd.n6018 avss -3.39e-19
C8806 avdd.n6019 avss -6.67e-19
C8807 avdd.n6020 avss -3.49e-19
C8808 avdd.n6021 avss 0.0184f
C8809 avdd.n6022 avss 0.00873f
C8810 avdd.n6023 avss 0.0148f
C8811 avdd.n6024 avss 0.00873f
C8812 avdd.n6025 avss 0.0111f
C8813 avdd.n6026 avss -2.44e-19
C8814 avdd.n6027 avss -2.33e-19
C8815 avdd.n6028 avss -1.8e-19
C8816 avdd.n6029 avss -1.48e-19
C8817 avdd.n6030 avss -8.47e-19
C8818 avdd.n6031 avss 0.00357f
C8819 avdd.n6032 avss 0.0348f
C8820 avdd.n6033 avss -0.00137f
C8821 avdd.n6034 avss -6.46e-19
C8822 avdd.n6035 avss 0.0189f
C8823 avdd.n6036 avss -3.07e-19
C8824 avdd.n6037 avss -2.01e-19
C8825 avdd.n6038 avss -3.28e-19
C8826 avdd.n6039 avss -3.28e-19
C8827 avdd.n6040 avss -8.47e-19
C8828 avdd.n6041 avss 0.0398f
C8829 avdd.n6042 avss -3.07e-19
C8830 avdd.n6043 avss 0.0181f
C8831 avdd.n6044 avss 0.0167f
C8832 avdd.n6045 avss 0.00875f
C8833 avdd.n6046 avss -2.54e-19
C8834 avdd.n6047 avss -2.54e-19
C8835 avdd.n6048 avss -2.22e-19
C8836 avdd.n6049 avss 0.0192f
C8837 avdd.n6050 avss -4.76e-19
C8838 avdd.n6051 avss -0.00128f
C8839 avdd.n6052 avss 0.0346f
C8840 avdd.n6053 avss -8.47e-19
C8841 avdd.n6054 avss 0.0388f
C8842 avdd.n6055 avss -8.47e-19
C8843 avdd.n6056 avss 0.0049f
C8844 avdd.n6057 avss 3e-19
C8845 avdd.n6058 avss -8.47e-19
C8846 avdd.n6059 avss -3.39e-19
C8847 avdd.n6060 avss -2.33e-19
C8848 avdd.n6061 avss -1.16e-19
C8849 avdd.n6062 avss 0.0182f
C8850 avdd.n6063 avss 0.0148f
C8851 avdd.n6064 avss 0.00875f
C8852 avdd.n6065 avss -2.22e-19
C8853 avdd.n6066 avss -2.22e-19
C8854 avdd.n6067 avss -1.8e-19
C8855 avdd.n6068 avss -1.8e-19
C8856 avdd.n6069 avss -1.59e-19
C8857 avdd.n6070 avss 0.0192f
C8858 avdd.n6071 avss -3.07e-19
C8859 avdd.n6072 avss -6.46e-19
C8860 avdd.n6073 avss -5.82e-19
C8861 avdd.n6074 avss -8.47e-19
C8862 avdd.n6075 avss -3.39e-19
C8863 avdd.n6076 avss -3.18e-19
C8864 avdd.n6077 avss -2.01e-19
C8865 avdd.n6078 avss 0.0183f
C8866 avdd.n6079 avss 0.0154f
C8867 avdd.n6080 avss 0.0154f
C8868 avdd.n6081 avss -1.8e-19
C8869 avdd.n6082 avss 0.0191f
C8870 avdd.n6083 avss -1.8e-19
C8871 avdd.n6084 avss -2.44e-19
C8872 avdd.n6085 avss -1.8e-19
C8873 avdd.n6086 avss -1.8e-19
C8874 avdd.n6087 avss -1.38e-19
C8875 avdd.n6088 avss -3.49e-19
C8876 avdd.n6089 avss 0.0184f
C8877 avdd.n6090 avss 0.00873f
C8878 avdd.n6091 avss 0.0422f
C8879 avdd.n6092 avss 0.00203f
C8880 avdd.n6093 avss 0.019f
C8881 avdd.n6094 avss -1.8e-19
C8882 avdd.n6095 avss -1.48e-19
C8883 avdd.n6096 avss -2.33e-19
C8884 avdd.n6097 avss -2.33e-19
C8885 avdd.n6098 avss -2.44e-19
C8886 avdd.n6099 avss 0.0197f
C8887 avdd.n6100 avss 0.0384f
C8888 avdd.n6101 avss -0.00512f
C8889 avdd.n6103 avss 0.0382f
C8890 avdd.n6104 avss -0.166f
C8891 avdd.n6105 avss -0.2f
C8892 avdd.n6106 avss 0.0269f
C8893 avdd.n6107 avss -1.27e-19
C8894 avdd.n6108 avss -2.96e-19
C8895 avdd.n6109 avss -0.00113f
C8896 avdd.n6111 avss -1.8e-19
C8897 avdd.n6112 avss -8.47e-19
C8898 avdd.n6113 avss 0.00869f
C8899 avdd.n6115 avss -0.00173f
C8900 avdd.n6116 avss -2.44e-19
C8901 avdd.n6117 avss 0.0111f
C8902 avdd.n6118 avss -1.38e-19
C8903 avdd.n6119 avss -2.44e-19
C8904 avdd.n6120 avss 0.0111f
C8905 avdd.n6121 avss -1.8e-19
C8906 avdd.n6122 avss -1.8e-19
C8907 avdd.n6123 avss 0.00908f
C8908 avdd.n6124 avss 0.03f
C8909 avdd.n6125 avss -3.39e-19
C8910 avdd.n6126 avss -3.39e-19
C8911 avdd.n6127 avss -1.59e-19
C8912 avdd.n6128 avss 0.0111f
C8913 avdd.n6129 avss -1.8e-19
C8914 avdd.n6130 avss -1.8e-19
C8915 avdd.n6131 avss 0.0342f
C8916 avdd.n6132 avss 0.00378f
C8917 avdd.n6133 avss -5.77e-19
C8918 avdd.n6134 avss -2.22e-19
C8919 avdd.n6135 avss 0.0168f
C8920 avdd.n6136 avss -3.6e-19
C8921 avdd.n6137 avss -1.8e-19
C8922 avdd.n6138 avss -8.26e-19
C8923 avdd.n6139 avss -0.0013f
C8924 avdd.n6140 avss -3.39e-19
C8925 avdd.n6141 avss -1.27e-19
C8926 avdd.n6142 avss 0.0022f
C8927 avdd.n6143 avss 0.019f
C8928 avdd.n6144 avss 0.0184f
C8929 avdd.n6145 avss -5.19e-19
C8930 avdd.n6146 avss 0.0386f
C8931 avdd.n6147 avss 0.0111f
C8932 avdd.n6148 avss -1.38e-19
C8933 avdd.n6149 avss -1.38e-19
C8934 avdd.n6150 avss -3.39e-19
C8935 avdd.n6151 avss -3.39e-19
C8936 avdd.n6152 avss -1.8e-19
C8937 avdd.n6153 avss 0.0411f
C8938 avdd.n6154 avss 0.0111f
C8939 avdd.n6155 avss -1.8e-19
C8940 avdd.n6156 avss -1.8e-19
C8941 avdd.n6157 avss -0.00173f
C8942 avdd.n6158 avss -0.00122f
C8943 avdd.n6159 avss -2.96e-19
C8944 avdd.n6160 avss -0.00121f
C8945 avdd.n6161 avss -6.35e-19
C8946 avdd.n6162 avss -0.00357f
C8947 avdd.n6163 avss -0.00109f
C8948 avdd.n6164 avss 0.0374f
C8949 avdd.n6165 avss 0.0112f
C8950 avdd.n6166 avss -1.8e-19
C8951 avdd.n6167 avss -1.8e-19
C8952 avdd.n6168 avss -0.00126f
C8953 avdd.n6169 avss 0.0318f
C8954 avdd.n6170 avss -0.00139f
C8955 avdd.n6171 avss -2.22e-19
C8956 avdd.n6172 avss 0.0188f
C8957 avdd.n6173 avss -2.75e-19
C8958 avdd.n6174 avss -3.6e-19
C8959 avdd.n6175 avss -3.07e-19
C8960 avdd.n6176 avss -6.88e-19
C8961 avdd.n6177 avss 0.00725f
C8962 avdd.n6178 avss -0.00336f
C8963 avdd.n6179 avss -1.8e-19
C8964 avdd.n6180 avss -2.01e-19
C8965 avdd.n6181 avss -0.0866f
C8966 avdd.n6182 avss 0.0179f
C8967 avdd.n6183 avss 0.0442f
C8968 avdd.n6184 avss -3.39e-19
C8969 avdd.n6185 avss -2.75e-19
C8970 avdd.n6186 avss 0.0181f
C8971 avdd.n6187 avss 0.00821f
C8972 avdd.n6188 avss 0.00821f
C8973 avdd.n6189 avss -2.75e-19
C8974 avdd.n6190 avss -2.33e-19
C8975 avdd.n6191 avss -2.54e-19
C8976 avdd.n6192 avss -2.54e-19
C8977 avdd.n6193 avss -2.22e-19
C8978 avdd.n6194 avss -1.59e-19
C8979 avdd.n6195 avss 0.0298f
C8980 avdd.n6196 avss 0.0098f
C8981 avdd.n6197 avss -0.00158f
C8982 avdd.n6198 avss -8.47e-19
C8983 avdd.n6199 avss -4.23e-19
C8984 avdd.n6200 avss -3.39e-19
C8985 avdd.n6201 avss -2.33e-19
C8986 avdd.n6202 avss -1.16e-19
C8987 avdd.n6203 avss 0.0182f
C8988 avdd.n6204 avss 0.0148f
C8989 avdd.n6205 avss 0.00875f
C8990 avdd.n6206 avss -2.22e-19
C8991 avdd.n6207 avss -2.22e-19
C8992 avdd.n6208 avss 0.00358f
C8993 avdd.n6209 avss -1.8e-19
C8994 avdd.n6210 avss -1.59e-19
C8995 avdd.n6211 avss 0.0192f
C8996 avdd.n6212 avss -3.07e-19
C8997 avdd.n6213 avss -0.00108f
C8998 avdd.n6214 avss 0.0382f
C8999 avdd.n6215 avss -9.76e-19
C9000 avdd.n6216 avss -2.01e-19
C9001 avdd.n6217 avss 0.0183f
C9002 avdd.n6218 avss 0.0154f
C9003 avdd.n6219 avss 0.0154f
C9004 avdd.n6220 avss 0.0191f
C9005 avdd.n6221 avss -1.8e-19
C9006 avdd.n6222 avss -1.8e-19
C9007 avdd.n6223 avss -2.44e-19
C9008 avdd.n6224 avss -1.8e-19
C9009 avdd.n6225 avss -1.8e-19
C9010 avdd.n6226 avss -5.61e-19
C9011 avdd.n6227 avss 0.0344f
C9012 avdd.n6228 avss -2.44e-19
C9013 avdd.n6229 avss -8.47e-19
C9014 avdd.n6230 avss -8.15e-19
C9015 avdd.n6231 avss -0.0014f
C9016 avdd.n6232 avss -8.47e-19
C9017 avdd.n6233 avss 0.00466f
C9018 avdd.n6234 avss -3.39e-19
C9019 avdd.n6235 avss -6.67e-19
C9020 avdd.n6236 avss -3.49e-19
C9021 avdd.n6237 avss 0.0184f
C9022 avdd.n6238 avss 0.00873f
C9023 avdd.n6239 avss 0.0148f
C9024 avdd.n6240 avss 0.00873f
C9025 avdd.n6241 avss 0.0111f
C9026 avdd.n6242 avss -2.44e-19
C9027 avdd.n6243 avss -2.33e-19
C9028 avdd.n6244 avss -1.8e-19
C9029 avdd.n6245 avss -1.48e-19
C9030 avdd.n6246 avss -8.47e-19
C9031 avdd.n6247 avss 0.00357f
C9032 avdd.n6248 avss 0.0348f
C9033 avdd.n6249 avss -0.00137f
C9034 avdd.n6250 avss -6.46e-19
C9035 avdd.n6251 avss 0.0189f
C9036 avdd.n6252 avss -3.07e-19
C9037 avdd.n6253 avss -2.01e-19
C9038 avdd.n6254 avss -3.28e-19
C9039 avdd.n6255 avss -3.28e-19
C9040 avdd.n6256 avss -8.47e-19
C9041 avdd.n6257 avss 0.0398f
C9042 avdd.n6258 avss -3.07e-19
C9043 avdd.n6259 avss 0.0181f
C9044 avdd.n6260 avss 0.0167f
C9045 avdd.n6261 avss 0.00875f
C9046 avdd.n6262 avss -2.54e-19
C9047 avdd.n6263 avss -2.54e-19
C9048 avdd.n6264 avss -2.22e-19
C9049 avdd.n6265 avss 0.0192f
C9050 avdd.n6266 avss -4.76e-19
C9051 avdd.n6267 avss -0.00128f
C9052 avdd.n6268 avss 0.0346f
C9053 avdd.n6269 avss -8.47e-19
C9054 avdd.n6270 avss 0.0388f
C9055 avdd.n6271 avss -8.47e-19
C9056 avdd.n6272 avss 0.0049f
C9057 avdd.n6273 avss 3e-19
C9058 avdd.n6274 avss -8.47e-19
C9059 avdd.n6275 avss -3.39e-19
C9060 avdd.n6276 avss -2.33e-19
C9061 avdd.n6277 avss -1.16e-19
C9062 avdd.n6278 avss 0.0182f
C9063 avdd.n6279 avss 0.0148f
C9064 avdd.n6280 avss 0.00875f
C9065 avdd.n6281 avss -2.22e-19
C9066 avdd.n6282 avss -2.22e-19
C9067 avdd.n6283 avss -1.8e-19
C9068 avdd.n6284 avss -1.8e-19
C9069 avdd.n6285 avss -1.59e-19
C9070 avdd.n6286 avss 0.0192f
C9071 avdd.n6287 avss -3.07e-19
C9072 avdd.n6288 avss -6.46e-19
C9073 avdd.n6289 avss -5.82e-19
C9074 avdd.n6290 avss -8.47e-19
C9075 avdd.n6291 avss -3.39e-19
C9076 avdd.n6292 avss -3.18e-19
C9077 avdd.n6293 avss -2.01e-19
C9078 avdd.n6294 avss 0.0183f
C9079 avdd.n6295 avss 0.0154f
C9080 avdd.n6296 avss 0.0154f
C9081 avdd.n6297 avss -1.8e-19
C9082 avdd.n6298 avss 0.0191f
C9083 avdd.n6299 avss -1.8e-19
C9084 avdd.n6300 avss -2.44e-19
C9085 avdd.n6301 avss -1.8e-19
C9086 avdd.n6302 avss -1.8e-19
C9087 avdd.n6303 avss -1.38e-19
C9088 avdd.n6304 avss -3.49e-19
C9089 avdd.n6305 avss 0.0184f
C9090 avdd.n6306 avss 0.00873f
C9091 avdd.n6307 avss 0.0422f
C9092 avdd.n6308 avss 0.00203f
C9093 avdd.n6309 avss 0.019f
C9094 avdd.n6310 avss -1.8e-19
C9095 avdd.n6311 avss -1.48e-19
C9096 avdd.n6312 avss -2.33e-19
C9097 avdd.n6313 avss -2.33e-19
C9098 avdd.n6314 avss -2.44e-19
C9099 avdd.n6315 avss 0.0197f
C9100 avdd.n6316 avss 0.0384f
C9101 avdd.n6317 avss -0.00512f
C9102 avdd.n6319 avss 0.0382f
C9103 avdd.n6320 avss -0.165f
C9104 avdd.n6321 avss -0.2f
C9105 avdd.n6322 avss 0.0269f
C9106 avdd.n6323 avss -1.27e-19
C9107 avdd.n6324 avss -2.96e-19
C9108 avdd.n6325 avss -0.00113f
C9109 avdd.n6327 avss -1.8e-19
C9110 avdd.n6328 avss -8.47e-19
C9111 avdd.n6329 avss 0.00869f
C9112 avdd.n6331 avss -0.00173f
C9113 avdd.n6332 avss -2.44e-19
C9114 avdd.n6333 avss 0.0111f
C9115 avdd.n6334 avss -1.38e-19
C9116 avdd.n6335 avss -2.44e-19
C9117 avdd.n6336 avss 0.0111f
C9118 avdd.n6337 avss -1.8e-19
C9119 avdd.n6338 avss -1.8e-19
C9120 avdd.n6339 avss 0.00908f
C9121 avdd.n6340 avss 0.03f
C9122 avdd.n6341 avss -3.39e-19
C9123 avdd.n6342 avss -3.39e-19
C9124 avdd.n6343 avss -1.59e-19
C9125 avdd.n6344 avss 0.0111f
C9126 avdd.n6345 avss -1.8e-19
C9127 avdd.n6346 avss -1.8e-19
C9128 avdd.n6347 avss 0.0342f
C9129 avdd.n6348 avss 0.00378f
C9130 avdd.n6349 avss -5.77e-19
C9131 avdd.n6350 avss -2.22e-19
C9132 avdd.n6351 avss 0.0168f
C9133 avdd.n6352 avss -3.6e-19
C9134 avdd.n6353 avss -1.8e-19
C9135 avdd.n6354 avss -8.26e-19
C9136 avdd.n6355 avss -0.0013f
C9137 avdd.n6356 avss -3.39e-19
C9138 avdd.n6357 avss -1.27e-19
C9139 avdd.n6358 avss 0.0022f
C9140 avdd.n6359 avss 0.019f
C9141 avdd.n6360 avss 0.0184f
C9142 avdd.n6361 avss -5.19e-19
C9143 avdd.n6362 avss 0.0386f
C9144 avdd.n6363 avss 0.0111f
C9145 avdd.n6364 avss -1.38e-19
C9146 avdd.n6365 avss -1.38e-19
C9147 avdd.n6366 avss -3.39e-19
C9148 avdd.n6367 avss -3.39e-19
C9149 avdd.n6368 avss -1.8e-19
C9150 avdd.n6369 avss 0.0411f
C9151 avdd.n6370 avss 0.0111f
C9152 avdd.n6371 avss -1.8e-19
C9153 avdd.n6372 avss -1.8e-19
C9154 avdd.n6373 avss -0.00173f
C9155 avdd.n6374 avss -0.00122f
C9156 avdd.n6375 avss -2.96e-19
C9157 avdd.n6376 avss -0.00121f
C9158 avdd.n6377 avss -6.35e-19
C9159 avdd.n6378 avss -0.00357f
C9160 avdd.n6379 avss -0.00109f
C9161 avdd.n6380 avss 0.0374f
C9162 avdd.n6381 avss 0.0112f
C9163 avdd.n6382 avss -1.8e-19
C9164 avdd.n6383 avss -1.8e-19
C9165 avdd.n6384 avss -0.00126f
C9166 avdd.n6385 avss 0.0318f
C9167 avdd.n6386 avss -0.00139f
C9168 avdd.n6387 avss -2.22e-19
C9169 avdd.n6388 avss 0.0188f
C9170 avdd.n6389 avss -2.75e-19
C9171 avdd.n6390 avss -3.6e-19
C9172 avdd.n6391 avss -3.07e-19
C9173 avdd.n6392 avss -6.88e-19
C9174 avdd.n6393 avss 0.00725f
C9175 avdd.n6394 avss -0.00336f
C9176 avdd.n6395 avss -1.8e-19
C9177 avdd.n6396 avss -2.01e-19
C9178 avdd.n6397 avss -0.0866f
C9179 avdd.n6398 avss 0.0179f
C9180 avdd.n6399 avss 0.0442f
C9181 avdd.n6400 avss -3.39e-19
C9182 avdd.n6401 avss -2.75e-19
C9183 avdd.n6402 avss 0.0181f
C9184 avdd.n6403 avss 0.00821f
C9185 avdd.n6404 avss 0.00821f
C9186 avdd.n6405 avss -2.75e-19
C9187 avdd.n6406 avss -2.33e-19
C9188 avdd.n6407 avss -2.54e-19
C9189 avdd.n6408 avss -2.54e-19
C9190 avdd.n6409 avss -2.22e-19
C9191 avdd.n6410 avss -1.59e-19
C9192 avdd.n6411 avss 0.0298f
C9193 avdd.n6412 avss 0.0098f
C9194 avdd.n6413 avss -0.00158f
C9195 avdd.n6414 avss -8.47e-19
C9196 avdd.n6415 avss -4.23e-19
C9197 avdd.n6416 avss -3.39e-19
C9198 avdd.n6417 avss -2.33e-19
C9199 avdd.n6418 avss -1.16e-19
C9200 avdd.n6419 avss 0.0182f
C9201 avdd.n6420 avss 0.0148f
C9202 avdd.n6421 avss 0.00875f
C9203 avdd.n6422 avss -2.22e-19
C9204 avdd.n6423 avss -2.22e-19
C9205 avdd.n6424 avss 0.00358f
C9206 avdd.n6425 avss -1.8e-19
C9207 avdd.n6426 avss -1.59e-19
C9208 avdd.n6427 avss 0.0192f
C9209 avdd.n6428 avss -3.07e-19
C9210 avdd.n6429 avss -0.00108f
C9211 avdd.n6430 avss 0.0382f
C9212 avdd.n6431 avss -9.76e-19
C9213 avdd.n6432 avss -2.01e-19
C9214 avdd.n6433 avss 0.0183f
C9215 avdd.n6434 avss 0.0154f
C9216 avdd.n6435 avss 0.0154f
C9217 avdd.n6436 avss 0.0191f
C9218 avdd.n6437 avss -1.8e-19
C9219 avdd.n6438 avss -1.8e-19
C9220 avdd.n6439 avss -2.44e-19
C9221 avdd.n6440 avss -1.8e-19
C9222 avdd.n6441 avss -1.8e-19
C9223 avdd.n6442 avss -5.61e-19
C9224 avdd.n6443 avss 0.0344f
C9225 avdd.n6444 avss -2.44e-19
C9226 avdd.n6445 avss -8.47e-19
C9227 avdd.n6446 avss -8.15e-19
C9228 avdd.n6447 avss -0.0014f
C9229 avdd.n6448 avss -8.47e-19
C9230 avdd.n6449 avss 0.00466f
C9231 avdd.n6450 avss -3.39e-19
C9232 avdd.n6451 avss -6.67e-19
C9233 avdd.n6452 avss -3.49e-19
C9234 avdd.n6453 avss 0.0184f
C9235 avdd.n6454 avss 0.00873f
C9236 avdd.n6455 avss 0.0148f
C9237 avdd.n6456 avss 0.00873f
C9238 avdd.n6457 avss 0.0111f
C9239 avdd.n6458 avss -2.44e-19
C9240 avdd.n6459 avss -2.33e-19
C9241 avdd.n6460 avss -1.8e-19
C9242 avdd.n6461 avss -1.48e-19
C9243 avdd.n6462 avss -8.47e-19
C9244 avdd.n6463 avss 0.00357f
C9245 avdd.n6464 avss 0.0348f
C9246 avdd.n6465 avss -0.00137f
C9247 avdd.n6466 avss -6.46e-19
C9248 avdd.n6467 avss 0.0189f
C9249 avdd.n6468 avss -3.07e-19
C9250 avdd.n6469 avss -2.01e-19
C9251 avdd.n6470 avss -3.28e-19
C9252 avdd.n6471 avss -3.28e-19
C9253 avdd.n6472 avss -8.47e-19
C9254 avdd.n6473 avss 0.0398f
C9255 avdd.n6474 avss -3.07e-19
C9256 avdd.n6475 avss 0.0181f
C9257 avdd.n6476 avss 0.0167f
C9258 avdd.n6477 avss 0.00875f
C9259 avdd.n6478 avss -2.54e-19
C9260 avdd.n6479 avss -2.54e-19
C9261 avdd.n6480 avss -2.22e-19
C9262 avdd.n6481 avss 0.0192f
C9263 avdd.n6482 avss -4.76e-19
C9264 avdd.n6483 avss -0.00128f
C9265 avdd.n6484 avss 0.0346f
C9266 avdd.n6485 avss -8.47e-19
C9267 avdd.n6486 avss 0.0388f
C9268 avdd.n6487 avss -8.47e-19
C9269 avdd.n6488 avss 0.0049f
C9270 avdd.n6489 avss 3e-19
C9271 avdd.n6490 avss -8.47e-19
C9272 avdd.n6491 avss -3.39e-19
C9273 avdd.n6492 avss -2.33e-19
C9274 avdd.n6493 avss -1.16e-19
C9275 avdd.n6494 avss 0.0182f
C9276 avdd.n6495 avss 0.0148f
C9277 avdd.n6496 avss 0.00875f
C9278 avdd.n6497 avss -2.22e-19
C9279 avdd.n6498 avss -2.22e-19
C9280 avdd.n6499 avss -1.8e-19
C9281 avdd.n6500 avss -1.8e-19
C9282 avdd.n6501 avss -1.59e-19
C9283 avdd.n6502 avss 0.0192f
C9284 avdd.n6503 avss -3.07e-19
C9285 avdd.n6504 avss -6.46e-19
C9286 avdd.n6505 avss -5.82e-19
C9287 avdd.n6506 avss -8.47e-19
C9288 avdd.n6507 avss -3.39e-19
C9289 avdd.n6508 avss -3.18e-19
C9290 avdd.n6509 avss -2.01e-19
C9291 avdd.n6510 avss 0.0183f
C9292 avdd.n6511 avss 0.0154f
C9293 avdd.n6512 avss 0.0154f
C9294 avdd.n6513 avss -1.8e-19
C9295 avdd.n6514 avss 0.0191f
C9296 avdd.n6515 avss -1.8e-19
C9297 avdd.n6516 avss -2.44e-19
C9298 avdd.n6517 avss -1.8e-19
C9299 avdd.n6518 avss -1.8e-19
C9300 avdd.n6519 avss -1.38e-19
C9301 avdd.n6520 avss -3.49e-19
C9302 avdd.n6521 avss 0.0184f
C9303 avdd.n6522 avss 0.00873f
C9304 avdd.n6523 avss 0.0422f
C9305 avdd.n6524 avss 0.00203f
C9306 avdd.n6525 avss 0.019f
C9307 avdd.n6526 avss -1.8e-19
C9308 avdd.n6527 avss -1.48e-19
C9309 avdd.n6528 avss -2.33e-19
C9310 avdd.n6529 avss -2.33e-19
C9311 avdd.n6530 avss -2.44e-19
C9312 avdd.n6531 avss 0.0197f
C9313 avdd.n6532 avss 0.0384f
C9314 avdd.n6533 avss -0.00512f
C9315 avdd.n6535 avss 0.0382f
C9316 avdd.n6536 avss -0.164f
C9317 avdd.n6537 avss -0.199f
C9318 avdd.n6538 avss 0.0269f
C9319 avdd.n6539 avss -1.27e-19
C9320 avdd.n6540 avss -2.96e-19
C9321 avdd.n6541 avss -0.00113f
C9322 avdd.n6543 avss -1.8e-19
C9323 avdd.n6544 avss -8.47e-19
C9324 avdd.n6545 avss 0.00869f
C9325 avdd.n6547 avss -0.00173f
C9326 avdd.n6548 avss -2.44e-19
C9327 avdd.n6549 avss 0.0111f
C9328 avdd.n6550 avss -1.38e-19
C9329 avdd.n6551 avss -2.44e-19
C9330 avdd.n6552 avss 0.0111f
C9331 avdd.n6553 avss -1.8e-19
C9332 avdd.n6554 avss -1.8e-19
C9333 avdd.n6555 avss 0.00908f
C9334 avdd.n6556 avss 0.03f
C9335 avdd.n6557 avss -3.39e-19
C9336 avdd.n6558 avss -3.39e-19
C9337 avdd.n6559 avss -1.59e-19
C9338 avdd.n6560 avss 0.0111f
C9339 avdd.n6561 avss -1.8e-19
C9340 avdd.n6562 avss -1.8e-19
C9341 avdd.n6563 avss 0.0342f
C9342 avdd.n6564 avss 0.00378f
C9343 avdd.n6565 avss -5.77e-19
C9344 avdd.n6566 avss -2.22e-19
C9345 avdd.n6567 avss 0.0168f
C9346 avdd.n6568 avss -3.6e-19
C9347 avdd.n6569 avss -1.8e-19
C9348 avdd.n6570 avss -8.26e-19
C9349 avdd.n6571 avss -0.0013f
C9350 avdd.n6572 avss -3.39e-19
C9351 avdd.n6573 avss -1.27e-19
C9352 avdd.n6574 avss 0.0022f
C9353 avdd.n6575 avss 0.019f
C9354 avdd.n6576 avss 0.0184f
C9355 avdd.n6577 avss -5.19e-19
C9356 avdd.n6578 avss 0.0386f
C9357 avdd.n6579 avss 0.0111f
C9358 avdd.n6580 avss -1.38e-19
C9359 avdd.n6581 avss -1.38e-19
C9360 avdd.n6582 avss -3.39e-19
C9361 avdd.n6583 avss -3.39e-19
C9362 avdd.n6584 avss -1.8e-19
C9363 avdd.n6585 avss 0.0411f
C9364 avdd.n6586 avss 0.0111f
C9365 avdd.n6587 avss -1.8e-19
C9366 avdd.n6588 avss -1.8e-19
C9367 avdd.n6589 avss -0.00173f
C9368 avdd.n6590 avss -0.00122f
C9369 avdd.n6591 avss -2.96e-19
C9370 avdd.n6592 avss -0.00121f
C9371 avdd.n6593 avss -6.35e-19
C9372 avdd.n6594 avss -0.00357f
C9373 avdd.n6595 avss -0.00109f
C9374 avdd.n6596 avss 0.0374f
C9375 avdd.n6597 avss 0.0112f
C9376 avdd.n6598 avss -1.8e-19
C9377 avdd.n6599 avss -1.8e-19
C9378 avdd.n6600 avss -0.00126f
C9379 avdd.n6601 avss 0.0318f
C9380 avdd.n6602 avss -0.00139f
C9381 avdd.n6603 avss -2.22e-19
C9382 avdd.n6604 avss 0.0188f
C9383 avdd.n6605 avss -2.75e-19
C9384 avdd.n6606 avss -3.6e-19
C9385 avdd.n6607 avss -3.07e-19
C9386 avdd.n6608 avss -6.88e-19
C9387 avdd.n6609 avss 0.00725f
C9388 avdd.n6610 avss -0.00336f
C9389 avdd.n6611 avss -1.8e-19
C9390 avdd.n6612 avss -2.01e-19
C9391 avdd.n6613 avss -0.0866f
C9392 avdd.n6614 avss 0.0179f
C9393 avdd.n6615 avss 0.0442f
C9394 avdd.n6616 avss -3.39e-19
C9395 avdd.n6617 avss -2.75e-19
C9396 avdd.n6618 avss 0.0181f
C9397 avdd.n6619 avss 0.00821f
C9398 avdd.n6620 avss 0.00821f
C9399 avdd.n6621 avss -2.75e-19
C9400 avdd.n6622 avss -2.33e-19
C9401 avdd.n6623 avss -2.54e-19
C9402 avdd.n6624 avss -2.54e-19
C9403 avdd.n6625 avss -2.22e-19
C9404 avdd.n6626 avss -1.59e-19
C9405 avdd.n6627 avss 0.0298f
C9406 avdd.n6628 avss 0.0098f
C9407 avdd.n6629 avss -0.00158f
C9408 avdd.n6630 avss -8.47e-19
C9409 avdd.n6631 avss -4.23e-19
C9410 avdd.n6632 avss -3.39e-19
C9411 avdd.n6633 avss -2.33e-19
C9412 avdd.n6634 avss -1.16e-19
C9413 avdd.n6635 avss 0.0182f
C9414 avdd.n6636 avss 0.0148f
C9415 avdd.n6637 avss 0.00875f
C9416 avdd.n6638 avss -2.22e-19
C9417 avdd.n6639 avss -2.22e-19
C9418 avdd.n6640 avss 0.00358f
C9419 avdd.n6641 avss -1.8e-19
C9420 avdd.n6642 avss -1.59e-19
C9421 avdd.n6643 avss 0.0192f
C9422 avdd.n6644 avss -3.07e-19
C9423 avdd.n6645 avss -0.00108f
C9424 avdd.n6646 avss 0.0382f
C9425 avdd.n6647 avss -9.76e-19
C9426 avdd.n6648 avss -2.01e-19
C9427 avdd.n6649 avss 0.0183f
C9428 avdd.n6650 avss 0.0154f
C9429 avdd.n6651 avss 0.0154f
C9430 avdd.n6652 avss 0.0191f
C9431 avdd.n6653 avss -1.8e-19
C9432 avdd.n6654 avss -1.8e-19
C9433 avdd.n6655 avss -2.44e-19
C9434 avdd.n6656 avss -1.8e-19
C9435 avdd.n6657 avss -1.8e-19
C9436 avdd.n6658 avss -5.61e-19
C9437 avdd.n6659 avss 0.0344f
C9438 avdd.n6660 avss -2.44e-19
C9439 avdd.n6661 avss -8.47e-19
C9440 avdd.n6662 avss -8.15e-19
C9441 avdd.n6663 avss -0.0014f
C9442 avdd.n6664 avss -8.47e-19
C9443 avdd.n6665 avss 0.00466f
C9444 avdd.n6666 avss -3.39e-19
C9445 avdd.n6667 avss -6.67e-19
C9446 avdd.n6668 avss -3.49e-19
C9447 avdd.n6669 avss 0.0184f
C9448 avdd.n6670 avss 0.00873f
C9449 avdd.n6671 avss 0.0148f
C9450 avdd.n6672 avss 0.00873f
C9451 avdd.n6673 avss 0.0111f
C9452 avdd.n6674 avss -2.44e-19
C9453 avdd.n6675 avss -2.33e-19
C9454 avdd.n6676 avss -1.8e-19
C9455 avdd.n6677 avss -1.48e-19
C9456 avdd.n6678 avss -8.47e-19
C9457 avdd.n6679 avss 0.00357f
C9458 avdd.n6680 avss 0.0348f
C9459 avdd.n6681 avss -0.00137f
C9460 avdd.n6682 avss -6.46e-19
C9461 avdd.n6683 avss 0.0189f
C9462 avdd.n6684 avss -3.07e-19
C9463 avdd.n6685 avss -2.01e-19
C9464 avdd.n6686 avss -3.28e-19
C9465 avdd.n6687 avss -3.28e-19
C9466 avdd.n6688 avss -8.47e-19
C9467 avdd.n6689 avss 0.0398f
C9468 avdd.n6690 avss -3.07e-19
C9469 avdd.n6691 avss 0.0181f
C9470 avdd.n6692 avss 0.0167f
C9471 avdd.n6693 avss 0.00875f
C9472 avdd.n6694 avss -2.54e-19
C9473 avdd.n6695 avss -2.54e-19
C9474 avdd.n6696 avss -2.22e-19
C9475 avdd.n6697 avss 0.0192f
C9476 avdd.n6698 avss -4.76e-19
C9477 avdd.n6699 avss -0.00128f
C9478 avdd.n6700 avss 0.0346f
C9479 avdd.n6701 avss -8.47e-19
C9480 avdd.n6702 avss 0.0388f
C9481 avdd.n6703 avss -8.47e-19
C9482 avdd.n6704 avss 0.0049f
C9483 avdd.n6705 avss 3e-19
C9484 avdd.n6706 avss -8.47e-19
C9485 avdd.n6707 avss -3.39e-19
C9486 avdd.n6708 avss -2.33e-19
C9487 avdd.n6709 avss -1.16e-19
C9488 avdd.n6710 avss 0.0182f
C9489 avdd.n6711 avss 0.0148f
C9490 avdd.n6712 avss 0.00875f
C9491 avdd.n6713 avss -2.22e-19
C9492 avdd.n6714 avss -2.22e-19
C9493 avdd.n6715 avss -1.8e-19
C9494 avdd.n6716 avss -1.8e-19
C9495 avdd.n6717 avss -1.59e-19
C9496 avdd.n6718 avss 0.0192f
C9497 avdd.n6719 avss -3.07e-19
C9498 avdd.n6720 avss -6.46e-19
C9499 avdd.n6721 avss -5.82e-19
C9500 avdd.n6722 avss -8.47e-19
C9501 avdd.n6723 avss -3.39e-19
C9502 avdd.n6724 avss -3.18e-19
C9503 avdd.n6725 avss -2.01e-19
C9504 avdd.n6726 avss 0.0183f
C9505 avdd.n6727 avss 0.0154f
C9506 avdd.n6728 avss 0.0154f
C9507 avdd.n6729 avss -1.8e-19
C9508 avdd.n6730 avss 0.0191f
C9509 avdd.n6731 avss -1.8e-19
C9510 avdd.n6732 avss -2.44e-19
C9511 avdd.n6733 avss -1.8e-19
C9512 avdd.n6734 avss -1.8e-19
C9513 avdd.n6735 avss -1.38e-19
C9514 avdd.n6736 avss -3.49e-19
C9515 avdd.n6737 avss 0.0184f
C9516 avdd.n6738 avss 0.00873f
C9517 avdd.n6739 avss 0.0422f
C9518 avdd.n6740 avss 0.00203f
C9519 avdd.n6741 avss 0.019f
C9520 avdd.n6742 avss -1.8e-19
C9521 avdd.n6743 avss -1.48e-19
C9522 avdd.n6744 avss -2.33e-19
C9523 avdd.n6745 avss -2.33e-19
C9524 avdd.n6746 avss -2.44e-19
C9525 avdd.n6747 avss 0.0197f
C9526 avdd.n6748 avss 0.0384f
C9527 avdd.n6749 avss -0.00512f
C9528 avdd.n6751 avss 0.0382f
C9529 avdd.n6752 avss -0.165f
C9530 avdd.n6753 avss -0.2f
C9531 avdd.n6754 avss 0.0269f
C9532 avdd.n6755 avss -1.27e-19
C9533 avdd.n6756 avss -2.96e-19
C9534 avdd.n6757 avss -0.00113f
C9535 avdd.n6759 avss -1.8e-19
C9536 avdd.n6760 avss -8.47e-19
C9537 avdd.n6761 avss 0.00869f
C9538 avdd.n6763 avss -0.00173f
C9539 avdd.n6764 avss -2.44e-19
C9540 avdd.n6765 avss 0.0111f
C9541 avdd.n6766 avss -1.38e-19
C9542 avdd.n6767 avss -2.44e-19
C9543 avdd.n6768 avss 0.0111f
C9544 avdd.n6769 avss -1.8e-19
C9545 avdd.n6770 avss -1.8e-19
C9546 avdd.n6771 avss 0.00908f
C9547 avdd.n6772 avss 0.03f
C9548 avdd.n6773 avss -3.39e-19
C9549 avdd.n6774 avss -3.39e-19
C9550 avdd.n6775 avss -1.59e-19
C9551 avdd.n6776 avss 0.0111f
C9552 avdd.n6777 avss -1.8e-19
C9553 avdd.n6778 avss -1.8e-19
C9554 avdd.n6779 avss 0.0342f
C9555 avdd.n6780 avss 0.00378f
C9556 avdd.n6781 avss -5.77e-19
C9557 avdd.n6782 avss -2.22e-19
C9558 avdd.n6783 avss 0.0168f
C9559 avdd.n6784 avss -3.6e-19
C9560 avdd.n6785 avss -1.8e-19
C9561 avdd.n6786 avss -8.26e-19
C9562 avdd.n6787 avss -0.0013f
C9563 avdd.n6788 avss -3.39e-19
C9564 avdd.n6789 avss -1.27e-19
C9565 avdd.n6790 avss 0.0022f
C9566 avdd.n6791 avss 0.019f
C9567 avdd.n6792 avss 0.0184f
C9568 avdd.n6793 avss -5.19e-19
C9569 avdd.n6794 avss 0.0386f
C9570 avdd.n6795 avss 0.0111f
C9571 avdd.n6796 avss -1.38e-19
C9572 avdd.n6797 avss -1.38e-19
C9573 avdd.n6798 avss -3.39e-19
C9574 avdd.n6799 avss -3.39e-19
C9575 avdd.n6800 avss -1.8e-19
C9576 avdd.n6801 avss 0.0411f
C9577 avdd.n6802 avss 0.0111f
C9578 avdd.n6803 avss -1.8e-19
C9579 avdd.n6804 avss -1.8e-19
C9580 avdd.n6805 avss -0.00173f
C9581 avdd.n6806 avss -0.00122f
C9582 avdd.n6807 avss -2.96e-19
C9583 avdd.n6808 avss -0.00121f
C9584 avdd.n6809 avss -6.35e-19
C9585 avdd.n6810 avss -0.00357f
C9586 avdd.n6811 avss -0.00109f
C9587 avdd.n6812 avss 0.0374f
C9588 avdd.n6813 avss 0.0112f
C9589 avdd.n6814 avss -1.8e-19
C9590 avdd.n6815 avss -1.8e-19
C9591 avdd.n6816 avss -0.00126f
C9592 avdd.n6817 avss 0.0318f
C9593 avdd.n6818 avss -0.00139f
C9594 avdd.n6819 avss -2.22e-19
C9595 avdd.n6820 avss 0.0188f
C9596 avdd.n6821 avss -2.75e-19
C9597 avdd.n6822 avss -3.6e-19
C9598 avdd.n6823 avss -3.07e-19
C9599 avdd.n6824 avss -6.88e-19
C9600 avdd.n6825 avss 0.00725f
C9601 avdd.n6826 avss -0.00336f
C9602 avdd.n6827 avss -1.8e-19
C9603 avdd.n6828 avss -2.01e-19
C9604 avdd.n6829 avss -0.0866f
C9605 avdd.n6830 avss 0.0179f
C9606 avdd.n6831 avss 0.0442f
C9607 avdd.n6832 avss -3.39e-19
C9608 avdd.n6833 avss -2.75e-19
C9609 avdd.n6834 avss 0.0181f
C9610 avdd.n6835 avss 0.00821f
C9611 avdd.n6836 avss 0.00821f
C9612 avdd.n6837 avss -2.75e-19
C9613 avdd.n6838 avss -2.33e-19
C9614 avdd.n6839 avss -2.54e-19
C9615 avdd.n6840 avss -2.54e-19
C9616 avdd.n6841 avss -2.22e-19
C9617 avdd.n6842 avss -1.59e-19
C9618 avdd.n6843 avss 0.0298f
C9619 avdd.n6844 avss 0.0098f
C9620 avdd.n6845 avss -0.00158f
C9621 avdd.n6846 avss -8.47e-19
C9622 avdd.n6847 avss -4.23e-19
C9623 avdd.n6848 avss -3.39e-19
C9624 avdd.n6849 avss -2.33e-19
C9625 avdd.n6850 avss -1.16e-19
C9626 avdd.n6851 avss 0.0182f
C9627 avdd.n6852 avss 0.0148f
C9628 avdd.n6853 avss 0.00875f
C9629 avdd.n6854 avss -2.22e-19
C9630 avdd.n6855 avss -2.22e-19
C9631 avdd.n6856 avss 0.00358f
C9632 avdd.n6857 avss -1.8e-19
C9633 avdd.n6858 avss -1.59e-19
C9634 avdd.n6859 avss 0.0192f
C9635 avdd.n6860 avss -3.07e-19
C9636 avdd.n6861 avss -0.00108f
C9637 avdd.n6862 avss 0.0382f
C9638 avdd.n6863 avss -9.76e-19
C9639 avdd.n6864 avss -2.01e-19
C9640 avdd.n6865 avss 0.0183f
C9641 avdd.n6866 avss 0.0154f
C9642 avdd.n6867 avss 0.0154f
C9643 avdd.n6868 avss 0.0191f
C9644 avdd.n6869 avss -1.8e-19
C9645 avdd.n6870 avss -1.8e-19
C9646 avdd.n6871 avss -2.44e-19
C9647 avdd.n6872 avss -1.8e-19
C9648 avdd.n6873 avss -1.8e-19
C9649 avdd.n6874 avss -5.61e-19
C9650 avdd.n6875 avss 0.0344f
C9651 avdd.n6876 avss -2.44e-19
C9652 avdd.n6877 avss -8.47e-19
C9653 avdd.n6878 avss -8.15e-19
C9654 avdd.n6879 avss -0.0014f
C9655 avdd.n6880 avss -8.47e-19
C9656 avdd.n6881 avss 0.00466f
C9657 avdd.n6882 avss -3.39e-19
C9658 avdd.n6883 avss -6.67e-19
C9659 avdd.n6884 avss -3.49e-19
C9660 avdd.n6885 avss 0.0184f
C9661 avdd.n6886 avss 0.00873f
C9662 avdd.n6887 avss 0.0148f
C9663 avdd.n6888 avss 0.00873f
C9664 avdd.n6889 avss 0.0111f
C9665 avdd.n6890 avss -2.44e-19
C9666 avdd.n6891 avss -2.33e-19
C9667 avdd.n6892 avss -1.8e-19
C9668 avdd.n6893 avss -1.48e-19
C9669 avdd.n6894 avss -8.47e-19
C9670 avdd.n6895 avss 0.00357f
C9671 avdd.n6896 avss 0.0348f
C9672 avdd.n6897 avss -0.00137f
C9673 avdd.n6898 avss -6.46e-19
C9674 avdd.n6899 avss 0.0189f
C9675 avdd.n6900 avss -3.07e-19
C9676 avdd.n6901 avss -2.01e-19
C9677 avdd.n6902 avss -3.28e-19
C9678 avdd.n6903 avss -3.28e-19
C9679 avdd.n6904 avss -8.47e-19
C9680 avdd.n6905 avss 0.0398f
C9681 avdd.n6906 avss -3.07e-19
C9682 avdd.n6907 avss 0.0181f
C9683 avdd.n6908 avss 0.0167f
C9684 avdd.n6909 avss 0.00875f
C9685 avdd.n6910 avss -2.54e-19
C9686 avdd.n6911 avss -2.54e-19
C9687 avdd.n6912 avss -2.22e-19
C9688 avdd.n6913 avss 0.0192f
C9689 avdd.n6914 avss -4.76e-19
C9690 avdd.n6915 avss -0.00128f
C9691 avdd.n6916 avss 0.0346f
C9692 avdd.n6917 avss -8.47e-19
C9693 avdd.n6918 avss 0.0388f
C9694 avdd.n6919 avss -8.47e-19
C9695 avdd.n6920 avss 0.0049f
C9696 avdd.n6921 avss 3e-19
C9697 avdd.n6922 avss -8.47e-19
C9698 avdd.n6923 avss -3.39e-19
C9699 avdd.n6924 avss -2.33e-19
C9700 avdd.n6925 avss -1.16e-19
C9701 avdd.n6926 avss 0.0182f
C9702 avdd.n6927 avss 0.0148f
C9703 avdd.n6928 avss 0.00875f
C9704 avdd.n6929 avss -2.22e-19
C9705 avdd.n6930 avss -2.22e-19
C9706 avdd.n6931 avss -1.8e-19
C9707 avdd.n6932 avss -1.8e-19
C9708 avdd.n6933 avss -1.59e-19
C9709 avdd.n6934 avss 0.0192f
C9710 avdd.n6935 avss -3.07e-19
C9711 avdd.n6936 avss -6.46e-19
C9712 avdd.n6937 avss -5.82e-19
C9713 avdd.n6938 avss -8.47e-19
C9714 avdd.n6939 avss -3.39e-19
C9715 avdd.n6940 avss -3.18e-19
C9716 avdd.n6941 avss -2.01e-19
C9717 avdd.n6942 avss 0.0183f
C9718 avdd.n6943 avss 0.0154f
C9719 avdd.n6944 avss 0.0154f
C9720 avdd.n6945 avss -1.8e-19
C9721 avdd.n6946 avss 0.0191f
C9722 avdd.n6947 avss -1.8e-19
C9723 avdd.n6948 avss -2.44e-19
C9724 avdd.n6949 avss -1.8e-19
C9725 avdd.n6950 avss -1.8e-19
C9726 avdd.n6951 avss -1.38e-19
C9727 avdd.n6952 avss -3.49e-19
C9728 avdd.n6953 avss 0.0184f
C9729 avdd.n6954 avss 0.00873f
C9730 avdd.n6955 avss 0.0422f
C9731 avdd.n6956 avss 0.00203f
C9732 avdd.n6957 avss 0.019f
C9733 avdd.n6958 avss -1.8e-19
C9734 avdd.n6959 avss -1.48e-19
C9735 avdd.n6960 avss -2.33e-19
C9736 avdd.n6961 avss -2.33e-19
C9737 avdd.n6962 avss -2.44e-19
C9738 avdd.n6963 avss 0.0197f
C9739 avdd.n6964 avss 0.0384f
C9740 avdd.n6965 avss -0.00512f
C9741 avdd.n6967 avss 0.0382f
C9742 avdd.n6968 avss -0.165f
C9743 avdd.n6969 avss -0.199f
C9744 avdd.n6970 avss 0.0269f
C9745 avdd.n6971 avss -1.27e-19
C9746 avdd.n6972 avss -2.96e-19
C9747 avdd.n6973 avss -0.00113f
C9748 avdd.n6975 avss -1.8e-19
C9749 avdd.n6976 avss -8.47e-19
C9750 avdd.n6977 avss 0.00869f
C9751 avdd.n6979 avss -0.00173f
C9752 avdd.n6980 avss -2.44e-19
C9753 avdd.n6981 avss 0.0111f
C9754 avdd.n6982 avss -1.38e-19
C9755 avdd.n6983 avss -2.44e-19
C9756 avdd.n6984 avss 0.0111f
C9757 avdd.n6985 avss -1.8e-19
C9758 avdd.n6986 avss -1.8e-19
C9759 avdd.n6987 avss 0.00908f
C9760 avdd.n6988 avss 0.03f
C9761 avdd.n6989 avss -3.39e-19
C9762 avdd.n6990 avss -3.39e-19
C9763 avdd.n6991 avss -1.59e-19
C9764 avdd.n6992 avss 0.0111f
C9765 avdd.n6993 avss -1.8e-19
C9766 avdd.n6994 avss -1.8e-19
C9767 avdd.n6995 avss 0.0342f
C9768 avdd.n6996 avss 0.00378f
C9769 avdd.n6997 avss -5.77e-19
C9770 avdd.n6998 avss -2.22e-19
C9771 avdd.n6999 avss 0.0168f
C9772 avdd.n7000 avss -3.6e-19
C9773 avdd.n7001 avss -1.8e-19
C9774 avdd.n7002 avss -8.26e-19
C9775 avdd.n7003 avss -0.0013f
C9776 avdd.n7004 avss -3.39e-19
C9777 avdd.n7005 avss -1.27e-19
C9778 avdd.n7006 avss 0.0022f
C9779 avdd.n7007 avss 0.019f
C9780 avdd.n7008 avss 0.0184f
C9781 avdd.n7009 avss -5.19e-19
C9782 avdd.n7010 avss 0.0386f
C9783 avdd.n7011 avss 0.0111f
C9784 avdd.n7012 avss -1.38e-19
C9785 avdd.n7013 avss -1.38e-19
C9786 avdd.n7014 avss -3.39e-19
C9787 avdd.n7015 avss -3.39e-19
C9788 avdd.n7016 avss -1.8e-19
C9789 avdd.n7017 avss 0.0411f
C9790 avdd.n7018 avss 0.0111f
C9791 avdd.n7019 avss -1.8e-19
C9792 avdd.n7020 avss -1.8e-19
C9793 avdd.n7021 avss -0.00173f
C9794 avdd.n7022 avss -0.00122f
C9795 avdd.n7023 avss -2.96e-19
C9796 avdd.n7024 avss -0.00121f
C9797 avdd.n7025 avss -6.35e-19
C9798 avdd.n7026 avss -0.00357f
C9799 avdd.n7027 avss -0.00109f
C9800 avdd.n7028 avss 0.0374f
C9801 avdd.n7029 avss 0.0112f
C9802 avdd.n7030 avss -1.8e-19
C9803 avdd.n7031 avss -1.8e-19
C9804 avdd.n7032 avss -0.00126f
C9805 avdd.n7033 avss 0.0318f
C9806 avdd.n7034 avss -0.00139f
C9807 avdd.n7035 avss -2.22e-19
C9808 avdd.n7036 avss 0.0188f
C9809 avdd.n7037 avss -2.75e-19
C9810 avdd.n7038 avss -3.6e-19
C9811 avdd.n7039 avss -3.07e-19
C9812 avdd.n7040 avss -6.88e-19
C9813 avdd.n7041 avss 0.00725f
C9814 avdd.n7042 avss -0.00336f
C9815 avdd.n7043 avss -1.8e-19
C9816 avdd.n7044 avss -2.01e-19
C9817 avdd.n7045 avss -0.0866f
C9818 avdd.n7046 avss 0.0179f
C9819 avdd.n7047 avss 0.0442f
C9820 avdd.n7048 avss -3.39e-19
C9821 avdd.n7049 avss -2.75e-19
C9822 avdd.n7050 avss 0.0181f
C9823 avdd.n7051 avss 0.00821f
C9824 avdd.n7052 avss 0.00821f
C9825 avdd.n7053 avss -2.75e-19
C9826 avdd.n7054 avss -2.33e-19
C9827 avdd.n7055 avss -2.54e-19
C9828 avdd.n7056 avss -2.54e-19
C9829 avdd.n7057 avss -2.22e-19
C9830 avdd.n7058 avss -1.59e-19
C9831 avdd.n7059 avss 0.0298f
C9832 avdd.n7060 avss 0.0098f
C9833 avdd.n7061 avss -0.00158f
C9834 avdd.n7062 avss -8.47e-19
C9835 avdd.n7063 avss -4.23e-19
C9836 avdd.n7064 avss -3.39e-19
C9837 avdd.n7065 avss -2.33e-19
C9838 avdd.n7066 avss -1.16e-19
C9839 avdd.n7067 avss 0.0182f
C9840 avdd.n7068 avss 0.0148f
C9841 avdd.n7069 avss 0.00875f
C9842 avdd.n7070 avss -2.22e-19
C9843 avdd.n7071 avss -2.22e-19
C9844 avdd.n7072 avss 0.00358f
C9845 avdd.n7073 avss -1.8e-19
C9846 avdd.n7074 avss -1.59e-19
C9847 avdd.n7075 avss 0.0192f
C9848 avdd.n7076 avss -3.07e-19
C9849 avdd.n7077 avss -0.00108f
C9850 avdd.n7078 avss 0.0382f
C9851 avdd.n7079 avss -9.76e-19
C9852 avdd.n7080 avss -2.01e-19
C9853 avdd.n7081 avss 0.0183f
C9854 avdd.n7082 avss 0.0154f
C9855 avdd.n7083 avss 0.0154f
C9856 avdd.n7084 avss 0.0191f
C9857 avdd.n7085 avss -1.8e-19
C9858 avdd.n7086 avss -1.8e-19
C9859 avdd.n7087 avss -2.44e-19
C9860 avdd.n7088 avss -1.8e-19
C9861 avdd.n7089 avss -1.8e-19
C9862 avdd.n7090 avss -5.61e-19
C9863 avdd.n7091 avss 0.0344f
C9864 avdd.n7092 avss -2.44e-19
C9865 avdd.n7093 avss -8.47e-19
C9866 avdd.n7094 avss -8.15e-19
C9867 avdd.n7095 avss -0.0014f
C9868 avdd.n7096 avss -8.47e-19
C9869 avdd.n7097 avss 0.00466f
C9870 avdd.n7098 avss -3.39e-19
C9871 avdd.n7099 avss -6.67e-19
C9872 avdd.n7100 avss -3.49e-19
C9873 avdd.n7101 avss 0.0184f
C9874 avdd.n7102 avss 0.00873f
C9875 avdd.n7103 avss 0.0148f
C9876 avdd.n7104 avss 0.00873f
C9877 avdd.n7105 avss 0.0111f
C9878 avdd.n7106 avss -2.44e-19
C9879 avdd.n7107 avss -2.33e-19
C9880 avdd.n7108 avss -1.8e-19
C9881 avdd.n7109 avss -1.48e-19
C9882 avdd.n7110 avss -8.47e-19
C9883 avdd.n7111 avss 0.00357f
C9884 avdd.n7112 avss 0.0348f
C9885 avdd.n7113 avss -0.00137f
C9886 avdd.n7114 avss -6.46e-19
C9887 avdd.n7115 avss 0.0189f
C9888 avdd.n7116 avss -3.07e-19
C9889 avdd.n7117 avss -2.01e-19
C9890 avdd.n7118 avss -3.28e-19
C9891 avdd.n7119 avss -3.28e-19
C9892 avdd.n7120 avss -8.47e-19
C9893 avdd.n7121 avss 0.0398f
C9894 avdd.n7122 avss -3.07e-19
C9895 avdd.n7123 avss 0.0181f
C9896 avdd.n7124 avss 0.0167f
C9897 avdd.n7125 avss 0.00875f
C9898 avdd.n7126 avss -2.54e-19
C9899 avdd.n7127 avss -2.54e-19
C9900 avdd.n7128 avss -2.22e-19
C9901 avdd.n7129 avss 0.0192f
C9902 avdd.n7130 avss -4.76e-19
C9903 avdd.n7131 avss -0.00128f
C9904 avdd.n7132 avss 0.0346f
C9905 avdd.n7133 avss -8.47e-19
C9906 avdd.n7134 avss 0.0388f
C9907 avdd.n7135 avss -8.47e-19
C9908 avdd.n7136 avss 0.0049f
C9909 avdd.n7137 avss 3e-19
C9910 avdd.n7138 avss -8.47e-19
C9911 avdd.n7139 avss -3.39e-19
C9912 avdd.n7140 avss -2.33e-19
C9913 avdd.n7141 avss -1.16e-19
C9914 avdd.n7142 avss 0.0182f
C9915 avdd.n7143 avss 0.0148f
C9916 avdd.n7144 avss 0.00875f
C9917 avdd.n7145 avss -2.22e-19
C9918 avdd.n7146 avss -2.22e-19
C9919 avdd.n7147 avss -1.8e-19
C9920 avdd.n7148 avss -1.8e-19
C9921 avdd.n7149 avss -1.59e-19
C9922 avdd.n7150 avss 0.0192f
C9923 avdd.n7151 avss -3.07e-19
C9924 avdd.n7152 avss -6.46e-19
C9925 avdd.n7153 avss -5.82e-19
C9926 avdd.n7154 avss -8.47e-19
C9927 avdd.n7155 avss -3.39e-19
C9928 avdd.n7156 avss -3.18e-19
C9929 avdd.n7157 avss -2.01e-19
C9930 avdd.n7158 avss 0.0183f
C9931 avdd.n7159 avss 0.0154f
C9932 avdd.n7160 avss 0.0154f
C9933 avdd.n7161 avss -1.8e-19
C9934 avdd.n7162 avss 0.0191f
C9935 avdd.n7163 avss -1.8e-19
C9936 avdd.n7164 avss -2.44e-19
C9937 avdd.n7165 avss -1.8e-19
C9938 avdd.n7166 avss -1.8e-19
C9939 avdd.n7167 avss -1.38e-19
C9940 avdd.n7168 avss -3.49e-19
C9941 avdd.n7169 avss 0.0184f
C9942 avdd.n7170 avss 0.00873f
C9943 avdd.n7171 avss 0.0422f
C9944 avdd.n7172 avss 0.00203f
C9945 avdd.n7173 avss 0.019f
C9946 avdd.n7174 avss -1.8e-19
C9947 avdd.n7175 avss -1.48e-19
C9948 avdd.n7176 avss -2.33e-19
C9949 avdd.n7177 avss -2.33e-19
C9950 avdd.n7178 avss -2.44e-19
C9951 avdd.n7179 avss 0.0197f
C9952 avdd.n7180 avss 0.0384f
C9953 avdd.n7181 avss -0.00512f
C9954 avdd.n7183 avss 0.0382f
C9955 avdd.n7184 avss -0.164f
C9956 avdd.n7185 avss -0.199f
C9957 avdd.n7186 avss 0.0269f
C9958 avdd.n7187 avss -1.27e-19
C9959 avdd.n7188 avss -2.96e-19
C9960 avdd.n7189 avss -0.00113f
C9961 avdd.n7191 avss -1.8e-19
C9962 avdd.n7192 avss -8.47e-19
C9963 avdd.n7193 avss 0.00869f
C9964 avdd.n7195 avss -0.00173f
C9965 avdd.n7196 avss -2.44e-19
C9966 avdd.n7197 avss 0.0111f
C9967 avdd.n7198 avss -1.38e-19
C9968 avdd.n7199 avss -2.44e-19
C9969 avdd.n7200 avss 0.0111f
C9970 avdd.n7201 avss -1.8e-19
C9971 avdd.n7202 avss -1.8e-19
C9972 avdd.n7203 avss 0.00908f
C9973 avdd.n7204 avss 0.03f
C9974 avdd.n7205 avss -3.39e-19
C9975 avdd.n7206 avss -3.39e-19
C9976 avdd.n7207 avss -1.59e-19
C9977 avdd.n7208 avss 0.0111f
C9978 avdd.n7209 avss -1.8e-19
C9979 avdd.n7210 avss -1.8e-19
C9980 avdd.n7211 avss 0.0342f
C9981 avdd.n7212 avss 0.00378f
C9982 avdd.n7213 avss -5.77e-19
C9983 avdd.n7214 avss -2.22e-19
C9984 avdd.n7215 avss 0.0168f
C9985 avdd.n7216 avss -3.6e-19
C9986 avdd.n7217 avss -1.8e-19
C9987 avdd.n7218 avss -8.26e-19
C9988 avdd.n7219 avss -0.0013f
C9989 avdd.n7220 avss -3.39e-19
C9990 avdd.n7221 avss -1.27e-19
C9991 avdd.n7222 avss 0.0022f
C9992 avdd.n7223 avss 0.019f
C9993 avdd.n7224 avss 0.0184f
C9994 avdd.n7225 avss -5.19e-19
C9995 avdd.n7226 avss 0.0386f
C9996 avdd.n7227 avss 0.0111f
C9997 avdd.n7228 avss -1.38e-19
C9998 avdd.n7229 avss -1.38e-19
C9999 avdd.n7230 avss -3.39e-19
C10000 avdd.n7231 avss -3.39e-19
C10001 avdd.n7232 avss -1.8e-19
C10002 avdd.n7233 avss 0.0411f
C10003 avdd.n7234 avss 0.0111f
C10004 avdd.n7235 avss -1.8e-19
C10005 avdd.n7236 avss -1.8e-19
C10006 avdd.n7237 avss -0.00173f
C10007 avdd.n7238 avss -0.00122f
C10008 avdd.n7239 avss -2.96e-19
C10009 avdd.n7240 avss -0.00121f
C10010 avdd.n7241 avss -6.35e-19
C10011 avdd.n7242 avss -0.00357f
C10012 avdd.n7243 avss -0.00109f
C10013 avdd.n7244 avss 0.0374f
C10014 avdd.n7245 avss 0.0112f
C10015 avdd.n7246 avss -1.8e-19
C10016 avdd.n7247 avss -1.8e-19
C10017 avdd.n7248 avss -0.00126f
C10018 avdd.n7249 avss 0.0318f
C10019 avdd.n7250 avss -0.00139f
C10020 avdd.n7251 avss -2.22e-19
C10021 avdd.n7252 avss 0.0188f
C10022 avdd.n7253 avss -2.75e-19
C10023 avdd.n7254 avss -3.6e-19
C10024 avdd.n7255 avss -3.07e-19
C10025 avdd.n7256 avss -6.88e-19
C10026 avdd.n7257 avss 0.00725f
C10027 avdd.n7258 avss -0.00336f
C10028 avdd.n7259 avss -1.8e-19
C10029 avdd.n7260 avss -2.01e-19
C10030 avdd.n7261 avss -0.0866f
C10031 avdd.n7262 avss 0.0179f
C10032 avdd.n7263 avss 0.0442f
C10033 avdd.n7264 avss -3.39e-19
C10034 avdd.n7265 avss -2.75e-19
C10035 avdd.n7266 avss 0.0181f
C10036 avdd.n7267 avss 0.00821f
C10037 avdd.n7268 avss 0.00821f
C10038 avdd.n7269 avss -2.75e-19
C10039 avdd.n7270 avss -2.33e-19
C10040 avdd.n7271 avss -2.54e-19
C10041 avdd.n7272 avss -2.54e-19
C10042 avdd.n7273 avss -2.22e-19
C10043 avdd.n7274 avss -1.59e-19
C10044 avdd.n7275 avss 0.0298f
C10045 avdd.n7276 avss 0.0098f
C10046 avdd.n7277 avss -0.00158f
C10047 avdd.n7278 avss -8.47e-19
C10048 avdd.n7279 avss -4.23e-19
C10049 avdd.n7280 avss -3.39e-19
C10050 avdd.n7281 avss -2.33e-19
C10051 avdd.n7282 avss -1.16e-19
C10052 avdd.n7283 avss 0.0182f
C10053 avdd.n7284 avss 0.0148f
C10054 avdd.n7285 avss 0.00875f
C10055 avdd.n7286 avss -2.22e-19
C10056 avdd.n7287 avss -2.22e-19
C10057 avdd.n7288 avss 0.00358f
C10058 avdd.n7289 avss -1.8e-19
C10059 avdd.n7290 avss -1.59e-19
C10060 avdd.n7291 avss 0.0192f
C10061 avdd.n7292 avss -3.07e-19
C10062 avdd.n7293 avss -0.00108f
C10063 avdd.n7294 avss 0.0382f
C10064 avdd.n7295 avss -9.76e-19
C10065 avdd.n7296 avss -2.01e-19
C10066 avdd.n7297 avss 0.0183f
C10067 avdd.n7298 avss 0.0154f
C10068 avdd.n7299 avss 0.0154f
C10069 avdd.n7300 avss 0.0191f
C10070 avdd.n7301 avss -1.8e-19
C10071 avdd.n7302 avss -1.8e-19
C10072 avdd.n7303 avss -2.44e-19
C10073 avdd.n7304 avss -1.8e-19
C10074 avdd.n7305 avss -1.8e-19
C10075 avdd.n7306 avss -5.61e-19
C10076 avdd.n7307 avss 0.0344f
C10077 avdd.n7308 avss -2.44e-19
C10078 avdd.n7309 avss -8.47e-19
C10079 avdd.n7310 avss -8.15e-19
C10080 avdd.n7311 avss -0.0014f
C10081 avdd.n7312 avss -8.47e-19
C10082 avdd.n7313 avss 0.00466f
C10083 avdd.n7314 avss -3.39e-19
C10084 avdd.n7315 avss -6.67e-19
C10085 avdd.n7316 avss -3.49e-19
C10086 avdd.n7317 avss 0.0184f
C10087 avdd.n7318 avss 0.00873f
C10088 avdd.n7319 avss 0.0148f
C10089 avdd.n7320 avss 0.00873f
C10090 avdd.n7321 avss 0.0111f
C10091 avdd.n7322 avss -2.44e-19
C10092 avdd.n7323 avss -2.33e-19
C10093 avdd.n7324 avss -1.8e-19
C10094 avdd.n7325 avss -1.48e-19
C10095 avdd.n7326 avss -8.47e-19
C10096 avdd.n7327 avss 0.00357f
C10097 avdd.n7328 avss 0.0348f
C10098 avdd.n7329 avss -0.00137f
C10099 avdd.n7330 avss -6.46e-19
C10100 avdd.n7331 avss 0.0189f
C10101 avdd.n7332 avss -3.07e-19
C10102 avdd.n7333 avss -2.01e-19
C10103 avdd.n7334 avss -3.28e-19
C10104 avdd.n7335 avss -3.28e-19
C10105 avdd.n7336 avss -8.47e-19
C10106 avdd.n7337 avss 0.0398f
C10107 avdd.n7338 avss -3.07e-19
C10108 avdd.n7339 avss 0.0181f
C10109 avdd.n7340 avss 0.0167f
C10110 avdd.n7341 avss 0.00875f
C10111 avdd.n7342 avss -2.54e-19
C10112 avdd.n7343 avss -2.54e-19
C10113 avdd.n7344 avss -2.22e-19
C10114 avdd.n7345 avss 0.0192f
C10115 avdd.n7346 avss -4.76e-19
C10116 avdd.n7347 avss -0.00128f
C10117 avdd.n7348 avss 0.0346f
C10118 avdd.n7349 avss -8.47e-19
C10119 avdd.n7350 avss 0.0388f
C10120 avdd.n7351 avss -8.47e-19
C10121 avdd.n7352 avss 0.0049f
C10122 avdd.n7353 avss 3e-19
C10123 avdd.n7354 avss -8.47e-19
C10124 avdd.n7355 avss -3.39e-19
C10125 avdd.n7356 avss -2.33e-19
C10126 avdd.n7357 avss -1.16e-19
C10127 avdd.n7358 avss 0.0182f
C10128 avdd.n7359 avss 0.0148f
C10129 avdd.n7360 avss 0.00875f
C10130 avdd.n7361 avss -2.22e-19
C10131 avdd.n7362 avss -2.22e-19
C10132 avdd.n7363 avss -1.8e-19
C10133 avdd.n7364 avss -1.8e-19
C10134 avdd.n7365 avss -1.59e-19
C10135 avdd.n7366 avss 0.0192f
C10136 avdd.n7367 avss -3.07e-19
C10137 avdd.n7368 avss -6.46e-19
C10138 avdd.n7369 avss -5.82e-19
C10139 avdd.n7370 avss -8.47e-19
C10140 avdd.n7371 avss -3.39e-19
C10141 avdd.n7372 avss -3.18e-19
C10142 avdd.n7373 avss -2.01e-19
C10143 avdd.n7374 avss 0.0183f
C10144 avdd.n7375 avss 0.0154f
C10145 avdd.n7376 avss 0.0154f
C10146 avdd.n7377 avss -1.8e-19
C10147 avdd.n7378 avss 0.0191f
C10148 avdd.n7379 avss -1.8e-19
C10149 avdd.n7380 avss -2.44e-19
C10150 avdd.n7381 avss -1.8e-19
C10151 avdd.n7382 avss -1.8e-19
C10152 avdd.n7383 avss -1.38e-19
C10153 avdd.n7384 avss -3.49e-19
C10154 avdd.n7385 avss 0.0184f
C10155 avdd.n7386 avss 0.00873f
C10156 avdd.n7387 avss 0.0422f
C10157 avdd.n7388 avss 0.00203f
C10158 avdd.n7389 avss 0.019f
C10159 avdd.n7390 avss -1.8e-19
C10160 avdd.n7391 avss -1.48e-19
C10161 avdd.n7392 avss -2.33e-19
C10162 avdd.n7393 avss -2.33e-19
C10163 avdd.n7394 avss -2.44e-19
C10164 avdd.n7395 avss 0.0197f
C10165 avdd.n7396 avss 0.0384f
C10166 avdd.n7397 avss -0.00512f
C10167 avdd.n7399 avss 0.0382f
C10168 avdd.n7400 avss -0.152f
C10169 avdd.n7401 avss -0.429f
C10170 avdd.n7402 avss -0.503f
C10171 avdd.t189 avss -0.00215f
C10172 avdd.n7403 avss -0.00826f
C10173 avdd.n7404 avss -0.00562f
C10174 avdd.n7405 avss -0.00797f
C10175 avdd.t202 avss -0.0366f
C10176 avdd.n7406 avss -0.00549f
C10177 avdd.n7407 avss -0.00263f
C10178 avdd.n7408 avss -0.00482f
C10179 avdd.n7409 avss -0.00168f
C10180 avdd.t122 avss -0.00353f
C10181 avdd.t265 avss -8.66e-19
C10182 avdd.t116 avss -8.66e-19
C10183 avdd.n7410 avss -0.00196f
C10184 avdd.n7411 avss -0.00252f
C10185 avdd.n7412 avss -0.00202f
C10186 avdd.t148 avss -0.00288f
C10187 avdd.n7413 avss -0.00168f
C10188 avdd.t39 avss -0.00353f
C10189 avdd.t44 avss -8.66e-19
C10190 avdd.t49 avss -8.66e-19
C10191 avdd.n7414 avss -0.00196f
C10192 avdd.n7415 avss -0.00252f
C10193 avdd.n7416 avss -0.00213f
C10194 avdd.t51 avss -0.00288f
C10195 avdd.t195 avss -0.00212f
C10196 avdd.n7417 avss -0.0045f
C10197 avdd.n7418 avss -0.00213f
C10198 avdd.t321 avss -0.00479f
C10199 avdd.t226 avss -0.00215f
C10200 avdd.n7419 avss -0.00826f
C10201 avdd.n7420 avss -0.00562f
C10202 avdd.n7421 avss -0.00797f
C10203 avdd.n7422 avss -0.0269f
C10204 avdd.t211 avss -0.0231f
C10205 avdd.t97 avss -0.0146f
C10206 avdd.t86 avss -0.0113f
C10207 avdd.t94 avss -0.0113f
C10208 avdd.t91 avss -0.0107f
C10209 avdd.t13 avss -0.0141f
C10210 avdd.t113 avss -0.0113f
C10211 avdd.t119 avss -0.0113f
C10212 avdd.t103 avss -0.0107f
C10213 avdd.t221 avss -0.0366f
C10214 avdd.n7423 avss -0.00549f
C10215 avdd.n7424 avss -0.00263f
C10216 avdd.n7425 avss -0.00484f
C10217 avdd.t312 avss -0.0156f
C10218 avdd.n7426 avss -0.0327f
C10219 avdd.t222 avss -0.0021f
C10220 avdd.n7427 avss -0.00168f
C10221 avdd.t104 avss -0.00353f
C10222 avdd.t114 avss -8.66e-19
C10223 avdd.t120 avss -8.66e-19
C10224 avdd.n7428 avss -0.00196f
C10225 avdd.n7429 avss -0.00252f
C10226 avdd.n7430 avss -0.00202f
C10227 avdd.t14 avss -0.00288f
C10228 avdd.n7431 avss -0.00168f
C10229 avdd.t92 avss -0.00353f
C10230 avdd.t87 avss -8.66e-19
C10231 avdd.t95 avss -8.66e-19
C10232 avdd.n7432 avss -0.00196f
C10233 avdd.n7433 avss -0.00252f
C10234 avdd.n7434 avss -0.00213f
C10235 avdd.t98 avss -0.00288f
C10236 avdd.t213 avss -0.00212f
C10237 avdd.n7435 avss -0.0045f
C10238 avdd.n7436 avss -0.00213f
C10239 avdd.t328 avss -0.00479f
C10240 avdd.n7437 avss -0.003f
C10241 avdd.t212 avss -0.00212f
C10242 avdd.n7438 avss -0.00172f
C10243 avdd.n7439 avss -0.00788f
C10244 avdd.n7440 avss -0.00627f
C10245 avdd.n7441 avss -0.00283f
C10246 avdd.n7442 avss -6.18e-19
C10247 avdd.n7443 avss -0.0109f
C10248 avdd.n7444 avss -3.33e-19
C10249 avdd.n7445 avss -0.00871f
C10250 avdd.t99 avss -0.0161f
C10251 avdd.n7446 avss -0.00514f
C10252 avdd.t85 avss -0.0215f
C10253 avdd.t100 avss -0.0215f
C10254 avdd.t90 avss -0.0215f
C10255 avdd.t88 avss -0.0265f
C10256 avdd.n7447 avss -0.0433f
C10257 avdd.n7448 avss -0.0211f
C10258 avdd.n7449 avss -0.0108f
C10259 avdd.t102 avss -0.0161f
C10260 avdd.t96 avss -0.0215f
C10261 avdd.t101 avss -0.0215f
C10262 avdd.t89 avss -0.0215f
C10263 avdd.t93 avss -0.0264f
C10264 avdd.n7450 avss -0.0158f
C10265 avdd.n7451 avss -0.00151f
C10266 avdd.n7453 avss -5.62e-19
C10267 avdd.n7454 avss -0.00501f
C10268 avdd.n7455 avss -0.00145f
C10269 avdd.n7456 avss -0.00278f
C10270 avdd.n7457 avss -0.00287f
C10271 avdd.n7458 avss -8.24e-19
C10272 avdd.n7459 avss -0.00283f
C10273 avdd.n7460 avss -0.00283f
C10274 avdd.n7461 avss -0.00283f
C10275 avdd.n7462 avss -8.24e-19
C10276 avdd.n7463 avss -0.00489f
C10277 avdd.n7464 avss -0.00278f
C10278 avdd.n7465 avss -8.24e-19
C10279 avdd.n7466 avss -0.00283f
C10280 avdd.n7467 avss -0.00283f
C10281 avdd.n7468 avss -0.00283f
C10282 avdd.n7469 avss -8.24e-19
C10283 avdd.n7470 avss -0.00481f
C10284 avdd.n7471 avss -0.00651f
C10285 avdd.n7472 avss -0.00632f
C10286 avdd.n7473 avss -0.0101f
C10287 avdd.n7474 avss -0.00797f
C10288 avdd.n7475 avss -0.00561f
C10289 avdd.n7476 avss -0.00378f
C10290 avdd.n7477 avss -0.00145f
C10291 avdd.t314 avss -0.00479f
C10292 avdd.t228 avss -0.00212f
C10293 avdd.n7478 avss -0.00172f
C10294 avdd.n7479 avss -0.00788f
C10295 avdd.t229 avss -0.00212f
C10296 avdd.n7480 avss -8.24e-19
C10297 avdd.n7481 avss -6.18e-19
C10298 avdd.n7482 avss -0.0109f
C10299 avdd.n7483 avss -3.33e-19
C10300 avdd.n7484 avss -0.00871f
C10301 avdd.t133 avss -0.0161f
C10302 avdd.n7485 avss -0.00514f
C10303 avdd.t127 avss -0.0215f
C10304 avdd.t134 avss -0.0215f
C10305 avdd.t143 avss -0.0215f
C10306 avdd.t135 avss -0.0265f
C10307 avdd.n7486 avss -0.0433f
C10308 avdd.n7487 avss -0.0211f
C10309 avdd.n7488 avss -0.0108f
C10310 avdd.t139 avss -0.0161f
C10311 avdd.t144 avss -0.0215f
C10312 avdd.t136 avss -0.0215f
C10313 avdd.t142 avss -0.0215f
C10314 avdd.t128 avss -0.0264f
C10315 avdd.n7489 avss -0.0158f
C10316 avdd.n7490 avss -0.00151f
C10317 avdd.n7492 avss -5.62e-19
C10318 avdd.n7493 avss -0.00501f
C10319 avdd.n7494 avss -0.00283f
C10320 avdd.t138 avss -8.66e-19
C10321 avdd.t130 avss -8.66e-19
C10322 avdd.n7495 avss -0.00196f
C10323 avdd.t82 avss -0.00288f
C10324 avdd.n7496 avss -0.00278f
C10325 avdd.n7497 avss -0.00283f
C10326 avdd.t118 avss -8.66e-19
C10327 avdd.t76 avss -8.66e-19
C10328 avdd.n7498 avss -0.00196f
C10329 avdd.t267 avss -0.00353f
C10330 avdd.n7499 avss -0.00481f
C10331 avdd.t225 avss -0.0021f
C10332 avdd.t313 avss -0.0156f
C10333 avdd.n7500 avss -0.0327f
C10334 avdd.n7501 avss -0.0101f
C10335 avdd.n7502 avss -0.00632f
C10336 avdd.n7503 avss -0.00651f
C10337 avdd.n7504 avss -0.00482f
C10338 avdd.n7505 avss -0.00168f
C10339 avdd.n7506 avss -0.00283f
C10340 avdd.n7507 avss -8.24e-19
C10341 avdd.n7508 avss -0.00252f
C10342 avdd.n7509 avss -8.24e-19
C10343 avdd.n7510 avss -0.00283f
C10344 avdd.n7511 avss -0.00202f
C10345 avdd.n7512 avss -0.00168f
C10346 avdd.t141 avss -0.00353f
C10347 avdd.n7513 avss -0.00489f
C10348 avdd.n7514 avss -8.24e-19
C10349 avdd.n7515 avss -0.00252f
C10350 avdd.n7516 avss -0.00283f
C10351 avdd.n7517 avss -0.00283f
C10352 avdd.n7518 avss -0.00213f
C10353 avdd.t132 avss -0.00288f
C10354 avdd.n7519 avss -0.00287f
C10355 avdd.n7520 avss -0.00278f
C10356 avdd.n7521 avss -0.0045f
C10357 avdd.n7522 avss -0.00627f
C10358 avdd.n7523 avss -0.00283f
C10359 avdd.n7524 avss -0.00213f
C10360 avdd.n7525 avss -0.00234f
C10361 avdd.n7526 avss -0.00364f
C10362 avdd.t223 avss -0.00215f
C10363 avdd.n7527 avss -0.00826f
C10364 avdd.n7528 avss -0.00924f
C10365 avdd.n7529 avss -0.0248f
C10366 avdd.t227 avss -0.0186f
C10367 avdd.t131 avss -0.0146f
C10368 avdd.t137 avss -0.0113f
C10369 avdd.t129 avss -0.0113f
C10370 avdd.t140 avss -0.0107f
C10371 avdd.t81 avss -0.0141f
C10372 avdd.t117 avss -0.0113f
C10373 avdd.t75 avss -0.0113f
C10374 avdd.t266 avss -0.0107f
C10375 avdd.t224 avss -0.0366f
C10376 avdd.t121 avss -0.0107f
C10377 avdd.t115 avss -0.0113f
C10378 avdd.t264 avss -0.0113f
C10379 avdd.t147 avss -0.0141f
C10380 avdd.t38 avss -0.0107f
C10381 avdd.t48 avss -0.0113f
C10382 avdd.t43 avss -0.0113f
C10383 avdd.t50 avss -0.0146f
C10384 avdd.t193 avss -0.0186f
C10385 avdd.n7530 avss -0.0248f
C10386 avdd.n7531 avss -0.00924f
C10387 avdd.n7532 avss -0.00549f
C10388 avdd.n7533 avss -0.00378f
C10389 avdd.n7534 avss -0.00234f
C10390 avdd.n7535 avss -0.00364f
C10391 avdd.n7536 avss -0.00263f
C10392 avdd.t194 avss -0.00212f
C10393 avdd.n7537 avss -0.00172f
C10394 avdd.n7538 avss -0.00788f
C10395 avdd.n7539 avss -0.00627f
C10396 avdd.n7540 avss -0.00283f
C10397 avdd.n7541 avss -6.18e-19
C10398 avdd.n7542 avss -0.0109f
C10399 avdd.n7543 avss -3.33e-19
C10400 avdd.n7544 avss -0.00871f
C10401 avdd.t35 avss -0.0161f
C10402 avdd.n7545 avss -0.00514f
C10403 avdd.t45 avss -0.0215f
C10404 avdd.t36 avss -0.0215f
C10405 avdd.t46 avss -0.0215f
C10406 avdd.t37 avss -0.0265f
C10407 avdd.n7546 avss -0.0433f
C10408 avdd.n7547 avss -0.0211f
C10409 avdd.n7548 avss -0.0108f
C10410 avdd.t42 avss -0.0161f
C10411 avdd.t52 avss -0.0215f
C10412 avdd.t41 avss -0.0215f
C10413 avdd.t40 avss -0.0215f
C10414 avdd.t47 avss -0.0264f
C10415 avdd.n7549 avss -0.0158f
C10416 avdd.n7550 avss -0.00151f
C10417 avdd.n7552 avss -5.62e-19
C10418 avdd.n7553 avss -0.00501f
C10419 avdd.n7554 avss -0.00145f
C10420 avdd.n7555 avss -0.00278f
C10421 avdd.n7556 avss -0.00287f
C10422 avdd.n7557 avss -8.24e-19
C10423 avdd.n7558 avss -0.00283f
C10424 avdd.n7559 avss -0.00283f
C10425 avdd.n7560 avss -0.00283f
C10426 avdd.n7561 avss -8.24e-19
C10427 avdd.n7562 avss -0.00489f
C10428 avdd.n7563 avss -0.00278f
C10429 avdd.n7564 avss -8.24e-19
C10430 avdd.n7565 avss -0.00283f
C10431 avdd.n7566 avss -0.00283f
C10432 avdd.n7567 avss -0.00283f
C10433 avdd.n7568 avss -8.24e-19
C10434 avdd.n7569 avss -0.00481f
C10435 avdd.n7570 avss -0.00651f
C10436 avdd.n7571 avss -0.00632f
C10437 avdd.t327 avss -0.0156f
C10438 avdd.t203 avss -0.0021f
C10439 avdd.n7572 avss -0.0327f
C10440 avdd.n7573 avss -0.0101f
C10441 avdd.n7574 avss -0.00797f
C10442 avdd.n7575 avss -0.00562f
C10443 avdd.n7576 avss -0.00378f
C10444 avdd.n7577 avss -0.00145f
C10445 avdd.t322 avss -0.00479f
C10446 avdd.t197 avss -0.00212f
C10447 avdd.n7578 avss -0.00172f
C10448 avdd.n7579 avss -0.00788f
C10449 avdd.t198 avss -0.00212f
C10450 avdd.n7580 avss -8.24e-19
C10451 avdd.n7581 avss -6.18e-19
C10452 avdd.n7582 avss -0.0109f
C10453 avdd.n7583 avss -3.33e-19
C10454 avdd.n7584 avss -0.00871f
C10455 avdd.t306 avss -0.0161f
C10456 avdd.n7585 avss -0.00514f
C10457 avdd.t291 avss -0.0215f
C10458 avdd.t307 avss -0.0215f
C10459 avdd.t299 avss -0.0215f
C10460 avdd.t292 avss -0.0265f
C10461 avdd.n7586 avss -0.0433f
C10462 avdd.n7587 avss -0.0211f
C10463 avdd.n7588 avss -0.0108f
C10464 avdd.t298 avss -0.0161f
C10465 avdd.t305 avss -0.0215f
C10466 avdd.t302 avss -0.0215f
C10467 avdd.t308 avss -0.0215f
C10468 avdd.t297 avss -0.0264f
C10469 avdd.n7589 avss -0.0158f
C10470 avdd.n7590 avss -0.00151f
C10471 avdd.n7592 avss -5.62e-19
C10472 avdd.n7593 avss -0.00501f
C10473 avdd.n7594 avss -0.00283f
C10474 avdd.t296 avss -8.66e-19
C10475 avdd.t301 avss -8.66e-19
C10476 avdd.n7595 avss -0.00196f
C10477 avdd.t150 avss -0.00288f
C10478 avdd.n7596 avss -0.00278f
C10479 avdd.n7597 avss -0.00283f
C10480 avdd.t184 avss -8.66e-19
C10481 avdd.t12 avss -8.66e-19
C10482 avdd.n7598 avss -0.00196f
C10483 avdd.t261 avss -0.00353f
C10484 avdd.n7599 avss -0.00481f
C10485 avdd.t188 avss -0.0021f
C10486 avdd.t320 avss -0.0156f
C10487 avdd.n7600 avss -0.0327f
C10488 avdd.n7601 avss -0.0101f
C10489 avdd.n7602 avss -0.00632f
C10490 avdd.n7603 avss -0.00651f
C10491 avdd.n7604 avss -0.00482f
C10492 avdd.n7605 avss -0.00168f
C10493 avdd.n7606 avss -0.00283f
C10494 avdd.n7607 avss -8.24e-19
C10495 avdd.n7608 avss -0.00252f
C10496 avdd.n7609 avss -8.24e-19
C10497 avdd.n7610 avss -0.00283f
C10498 avdd.n7611 avss -0.00202f
C10499 avdd.n7612 avss -0.00168f
C10500 avdd.t294 avss -0.00353f
C10501 avdd.n7613 avss -0.00489f
C10502 avdd.n7614 avss -8.24e-19
C10503 avdd.n7615 avss -0.00252f
C10504 avdd.n7616 avss -0.00283f
C10505 avdd.n7617 avss -0.00283f
C10506 avdd.n7618 avss -0.00213f
C10507 avdd.t304 avss -0.00288f
C10508 avdd.n7619 avss -0.00287f
C10509 avdd.n7620 avss -0.00278f
C10510 avdd.n7621 avss -0.0045f
C10511 avdd.n7622 avss -0.00627f
C10512 avdd.n7623 avss -0.00283f
C10513 avdd.n7624 avss -0.00213f
C10514 avdd.n7625 avss -0.00234f
C10515 avdd.n7626 avss -0.00364f
C10516 avdd.t204 avss -0.00215f
C10517 avdd.n7627 avss -0.00826f
C10518 avdd.n7628 avss -0.00924f
C10519 avdd.n7629 avss -0.0248f
C10520 avdd.t196 avss -0.0186f
C10521 avdd.t303 avss -0.0146f
C10522 avdd.t295 avss -0.0113f
C10523 avdd.t300 avss -0.0113f
C10524 avdd.t293 avss -0.0107f
C10525 avdd.t149 avss -0.0141f
C10526 avdd.t183 avss -0.0113f
C10527 avdd.t11 avss -0.0113f
C10528 avdd.t260 avss -0.0107f
C10529 avdd.t187 avss -0.0366f
C10530 avdd.n7630 avss -0.0192f
C10531 avdd.n7631 avss -0.0248f
C10532 avdd.n7632 avss -0.00924f
C10533 avdd.n7633 avss -0.00549f
C10534 avdd.n7634 avss -0.00378f
C10535 avdd.n7635 avss -6.67e-19
C10536 avdd.n7636 avss -0.00234f
C10537 avdd.n7637 avss -0.0038f
C10538 avdd.n7638 avss -0.00323f
C10539 avdd.n7639 avss -0.0886f
C10540 avdd.n7640 avss -8.26e-19
C10541 avdd.n7641 avss 0.0348f
C10542 avdd.n7642 avss 0.00357f
C10543 avdd.n7643 avss -8.47e-19
C10544 avdd.n7644 avss -3.39e-19
C10545 avdd.n7645 avss -8.47e-19
C10546 avdd.n7646 avss 0.0344f
C10547 avdd.n7647 avss 0.00466f
C10548 avdd.n7648 avss -3.39e-19
C10549 avdd.n7649 avss -6.67e-19
C10550 avdd.n7650 avss -5.61e-19
C10551 avdd.n7651 avss -3.39e-19
C10552 avdd.n7652 avss -6.35e-19
C10553 avdd.n7653 avss 0.0398f
C10554 avdd.n7654 avss -3.07e-19
C10555 avdd.n7655 avss -1.8e-19
C10556 avdd.n7656 avss 0.0168f
C10557 avdd.n7657 avss 0.0189f
C10558 avdd.n7658 avss 0.00875f
C10559 avdd.n7659 avss 0.0167f
C10560 avdd.n7660 avss 0.0181f
C10561 avdd.n7661 avss -3.6e-19
C10562 avdd.n7662 avss -2.01e-19
C10563 avdd.n7663 avss -3.07e-19
C10564 avdd.n7664 avss -6.46e-19
C10565 avdd.n7665 avss -0.00137f
C10566 avdd.n7666 avss -0.0013f
C10567 avdd.n7667 avss -5.19e-19
C10568 avdd.n7668 avss 0.0386f
C10569 avdd.n7669 avss 0.00873f
C10570 avdd.n7670 avss 0.0111f
C10571 avdd.n7671 avss 0.0148f
C10572 avdd.n7672 avss 0.019f
C10573 avdd.n7673 avss -1.8e-19
C10574 avdd.n7674 avss 0.0184f
C10575 avdd.n7675 avss -2.44e-19
C10576 avdd.n7676 avss -2.33e-19
C10577 avdd.n7677 avss 0.0022f
C10578 avdd.n7678 avss -1.48e-19
C10579 avdd.n7679 avss -1.27e-19
C10580 avdd.n7680 avss -2.44e-19
C10581 avdd.n7681 avss -8.15e-19
C10582 avdd.n7682 avss -0.0014f
C10583 avdd.n7683 avss -8.47e-19
C10584 avdd.n7684 avss -3.39e-19
C10585 avdd.n7685 avss -3.49e-19
C10586 avdd.n7686 avss -1.38e-19
C10587 avdd.n7687 avss -1.8e-19
C10588 avdd.n7688 avss 0.00873f
C10589 avdd.n7689 avss 0.0111f
C10590 avdd.n7690 avss 0.0154f
C10591 avdd.n7691 avss 0.0191f
C10592 avdd.n7692 avss -1.8e-19
C10593 avdd.n7693 avss 0.0184f
C10594 avdd.n7694 avss -1.38e-19
C10595 avdd.n7695 avss -1.8e-19
C10596 avdd.n7696 avss -2.44e-19
C10597 avdd.n7697 avss 0.0411f
C10598 avdd.n7698 avss -1.8e-19
C10599 avdd.n7699 avss -1.8e-19
C10600 avdd.n7700 avss -2.96e-19
C10601 avdd.n7701 avss -0.00139f
C10602 avdd.n7702 avss 0.0098f
C10603 avdd.n7703 avss 0.0298f
C10604 avdd.n7704 avss -2.22e-19
C10605 avdd.n7705 avss 0.0188f
C10606 avdd.n7706 avss -2.33e-19
C10607 avdd.n7707 avss -1.59e-19
C10608 avdd.n7708 avss -2.22e-19
C10609 avdd.n7709 avss 0.00821f
C10610 avdd.n7710 avss -2.75e-19
C10611 avdd.n7711 avss 0.0112f
C10612 avdd.n7712 avss 0.0148f
C10613 avdd.n7713 avss 0.0182f
C10614 avdd.n7714 avss -1.8e-19
C10615 avdd.n7715 avss -2.54e-19
C10616 avdd.n7716 avss -2.54e-19
C10617 avdd.n7717 avss -1.8e-19
C10618 avdd.n7718 avss -1.16e-19
C10619 avdd.n7719 avss -2.33e-19
C10620 avdd.n7720 avss -0.00126f
C10621 avdd.n7721 avss -0.00109f
C10622 avdd.n7722 avss -0.00108f
C10623 avdd.n7723 avss -3.07e-19
C10624 avdd.n7724 avss 0.0374f
C10625 avdd.n7725 avss 0.00358f
C10626 avdd.n7726 avss 0.0192f
C10627 avdd.n7727 avss -1.59e-19
C10628 avdd.n7728 avss -1.8e-19
C10629 avdd.n7729 avss 0.00875f
C10630 avdd.n7730 avss 0.0111f
C10631 avdd.n7731 avss 0.0154f
C10632 avdd.n7732 avss 0.0183f
C10633 avdd.n7733 avss -1.8e-19
C10634 avdd.n7734 avss -2.22e-19
C10635 avdd.n7735 avss -2.22e-19
C10636 avdd.n7736 avss -1.8e-19
C10637 avdd.n7737 avss -2.01e-19
C10638 avdd.n7738 avss -9.59e-19
C10639 avdd.n7739 avss -0.00106f
C10640 avdd.n7740 avss -0.00173f
C10641 avdd.n7741 avss -0.00139f
C10642 avdd.n7742 avss -6.88e-19
C10643 avdd.n7743 avss -3.07e-19
C10644 avdd.n7744 avss -1.8e-19
C10645 avdd.n7745 avss 0.00821f
C10646 avdd.n7746 avss -2.75e-19
C10647 avdd.n7747 avss 0.0442f
C10648 avdd.n7748 avss 0.0179f
C10649 avdd.n7749 avss 0.0181f
C10650 avdd.n7750 avss -2.75e-19
C10651 avdd.n7751 avss -3.39e-19
C10652 avdd.n7752 avss -3.6e-19
C10653 avdd.n7753 avss -2.01e-19
C10654 avdd.n7754 avss -0.0866f
C10655 avdd.n7755 avss -0.00336f
C10656 avdd.n7756 avss 0.00725f
C10657 avdd.n7757 avss 0.0318f
C10658 avdd.n7758 avss -0.00158f
C10659 avdd.n7759 avss -8.47e-19
C10660 avdd.n7760 avss -3.39e-19
C10661 avdd.n7761 avss -4.23e-19
C10662 avdd.n7762 avss -0.00357f
C10663 avdd.n7764 avss 0.0382f
C10664 avdd.n7765 avss -0.167f
C10665 avdd.n7766 avss -3.28e-19
C10666 avdd.n7767 avss -3.28e-19
C10667 avdd.n7768 avss -8.47e-19
C10668 avdd.n7769 avss 0.00378f
C10669 avdd.n7770 avss 0.0346f
C10670 avdd.n7771 avss -8.47e-19
C10671 avdd.n7772 avss -3.39e-19
C10672 avdd.n7773 avss -8.47e-19
C10673 avdd.n7774 avss 3e-19
C10674 avdd.n7775 avss 0.0388f
C10675 avdd.n7776 avss -3.39e-19
C10676 avdd.n7777 avss -6.46e-19
C10677 avdd.n7778 avss -5.82e-19
C10678 avdd.n7779 avss -3.39e-19
C10679 avdd.n7780 avss -8.47e-19
C10680 avdd.n7781 avss -0.00113f
C10681 avdd.n7782 avss 0.0384f
C10682 avdd.n7783 avss -2.44e-19
C10683 avdd.n7784 avss 0.0422f
C10684 avdd.n7785 avss 0.019f
C10685 avdd.n7786 avss -1.8e-19
C10686 avdd.n7787 avss 0.0197f
C10687 avdd.n7788 avss -2.44e-19
C10688 avdd.n7789 avss -2.33e-19
C10689 avdd.n7790 avss -2.33e-19
C10690 avdd.n7791 avss -1.48e-19
C10691 avdd.n7792 avss -1.27e-19
C10692 avdd.n7793 avss 0.00203f
C10693 avdd.n7794 avss -5.77e-19
C10694 avdd.n7795 avss -0.00128f
C10695 avdd.n7796 avss -4.76e-19
C10696 avdd.n7797 avss -2.22e-19
C10697 avdd.n7798 avss 0.0192f
C10698 avdd.n7799 avss -2.22e-19
C10699 avdd.n7800 avss 0.0111f
C10700 avdd.n7801 avss 0.0148f
C10701 avdd.n7802 avss 0.0182f
C10702 avdd.n7803 avss -1.8e-19
C10703 avdd.n7804 avss -2.54e-19
C10704 avdd.n7805 avss -2.54e-19
C10705 avdd.n7806 avss -1.8e-19
C10706 avdd.n7807 avss -1.16e-19
C10707 avdd.n7808 avss -2.33e-19
C10708 avdd.n7809 avss 0.0342f
C10709 avdd.n7810 avss 0.0049f
C10710 avdd.n7811 avss -8.47e-19
C10711 avdd.n7812 avss -3.39e-19
C10712 avdd.n7813 avss -3.07e-19
C10713 avdd.n7814 avss -1.59e-19
C10714 avdd.n7815 avss -1.8e-19
C10715 avdd.n7816 avss 0.0192f
C10716 avdd.n7817 avss -1.59e-19
C10717 avdd.n7818 avss -1.8e-19
C10718 avdd.n7819 avss 0.00875f
C10719 avdd.n7820 avss 0.0111f
C10720 avdd.n7821 avss 0.0154f
C10721 avdd.n7822 avss 0.0183f
C10722 avdd.n7823 avss -1.8e-19
C10723 avdd.n7824 avss -2.22e-19
C10724 avdd.n7825 avss -2.22e-19
C10725 avdd.n7826 avss -1.8e-19
C10726 avdd.n7827 avss -2.01e-19
C10727 avdd.n7828 avss -3.18e-19
C10728 avdd.n7829 avss 0.03f
C10729 avdd.n7830 avss 0.00899f
C10730 avdd.n7831 avss -7.52e-19
C10731 avdd.n7832 avss -2.96e-19
C10732 avdd.n7833 avss -1.8e-19
C10733 avdd.n7834 avss -1.8e-19
C10734 avdd.n7835 avss 0.00873f
C10735 avdd.n7836 avss 0.0111f
C10736 avdd.n7837 avss 0.0154f
C10737 avdd.n7838 avss 0.0191f
C10738 avdd.n7839 avss -1.8e-19
C10739 avdd.n7840 avss 0.0184f
C10740 avdd.n7841 avss -1.38e-19
C10741 avdd.n7842 avss -1.8e-19
C10742 avdd.n7843 avss -2.44e-19
C10743 avdd.n7844 avss -2.44e-19
C10744 avdd.n7845 avss -1.8e-19
C10745 avdd.n7846 avss -1.38e-19
C10746 avdd.n7847 avss -3.49e-19
C10747 avdd.n7848 avss 0.0269f
C10748 avdd.n7849 avss 0.00869f
C10749 avdd.n7850 avss -0.00173f
C10750 avdd.n7852 avss -0.00512f
C10751 avdd.n7854 avss 0.0382f
C10752 avdd.n7855 avss -0.564f
C10753 avdd.n7856 avss -0.511f
C10754 avdd.n7857 avss -0.00173f
C10755 avdd.n7859 avss 0.0384f
C10756 avdd.n7860 avss -2.44e-19
C10757 avdd.n7861 avss 0.0422f
C10758 avdd.n7862 avss 0.019f
C10759 avdd.n7863 avss -1.8e-19
C10760 avdd.n7864 avss 0.0197f
C10761 avdd.n7865 avss -2.44e-19
C10762 avdd.n7866 avss -2.33e-19
C10763 avdd.n7867 avss -2.33e-19
C10764 avdd.n7868 avss -1.48e-19
C10765 avdd.n7869 avss -1.27e-19
C10766 avdd.n7870 avss 0.00203f
C10767 avdd.n7871 avss -0.00128f
C10768 avdd.n7872 avss -4.76e-19
C10769 avdd.n7873 avss -2.22e-19
C10770 avdd.n7874 avss 0.0192f
C10771 avdd.n7875 avss -2.22e-19
C10772 avdd.n7876 avss 0.0148f
C10773 avdd.n7877 avss 0.0182f
C10774 avdd.n7878 avss -1.8e-19
C10775 avdd.n7879 avss -2.54e-19
C10776 avdd.n7880 avss -2.54e-19
C10777 avdd.n7881 avss -1.8e-19
C10778 avdd.n7882 avss -1.16e-19
C10779 avdd.n7883 avss -2.33e-19
C10780 avdd.n7884 avss 0.0342f
C10781 avdd.n7885 avss 0.0049f
C10782 avdd.n7886 avss -8.47e-19
C10783 avdd.n7887 avss -3.39e-19
C10784 avdd.n7888 avss -3.07e-19
C10785 avdd.n7889 avss -1.59e-19
C10786 avdd.n7890 avss -1.8e-19
C10787 avdd.n7891 avss 0.0192f
C10788 avdd.n7892 avss -1.59e-19
C10789 avdd.n7893 avss -1.8e-19
C10790 avdd.n7894 avss 0.00875f
C10791 avdd.n7895 avss 0.0111f
C10792 avdd.n7896 avss 0.0154f
C10793 avdd.n7897 avss 0.0183f
C10794 avdd.n7898 avss -1.8e-19
C10795 avdd.n7899 avss -2.22e-19
C10796 avdd.n7900 avss -2.22e-19
C10797 avdd.n7901 avss -1.8e-19
C10798 avdd.n7902 avss -2.01e-19
C10799 avdd.n7903 avss -3.18e-19
C10800 avdd.n7904 avss 0.03f
C10801 avdd.n7905 avss 0.00899f
C10802 avdd.n7906 avss -7.52e-19
C10803 avdd.n7907 avss -2.96e-19
C10804 avdd.n7908 avss -1.8e-19
C10805 avdd.n7909 avss -1.8e-19
C10806 avdd.n7910 avss 0.00873f
C10807 avdd.n7911 avss 0.0111f
C10808 avdd.n7912 avss 0.0154f
C10809 avdd.n7913 avss 0.0191f
C10810 avdd.n7914 avss -1.8e-19
C10811 avdd.n7915 avss 0.0184f
C10812 avdd.n7916 avss -1.38e-19
C10813 avdd.n7917 avss -1.8e-19
C10814 avdd.n7918 avss -2.44e-19
C10815 avdd.n7919 avss -2.44e-19
C10816 avdd.n7920 avss -1.8e-19
C10817 avdd.n7921 avss -1.38e-19
C10818 avdd.n7922 avss -3.49e-19
C10819 avdd.n7924 avss 0.0269f
C10820 avdd.n7925 avss 0.00869f
C10821 avdd.n7926 avss 0.00378f
C10822 avdd.n7927 avss 0.0346f
C10823 avdd.n7928 avss -8.47e-19
C10824 avdd.n7929 avss -3.39e-19
C10825 avdd.n7930 avss -8.47e-19
C10826 avdd.n7931 avss 3e-19
C10827 avdd.n7932 avss 0.0388f
C10828 avdd.n7933 avss -3.39e-19
C10829 avdd.n7934 avss -6.46e-19
C10830 avdd.n7935 avss -5.82e-19
C10831 avdd.n7936 avss -3.39e-19
C10832 avdd.n7937 avss -8.47e-19
C10833 avdd.n7938 avss -0.00113f
C10834 avdd.n7939 avss -0.00512f
C10835 avdd.n7940 avss 0.0382f
C10836 avdd.n7941 avss -0.144f
C10837 avdd.n7942 avss -0.179f
C10838 avdd.n7943 avss -0.00173f
C10839 avdd.n7945 avss 0.0384f
C10840 avdd.n7946 avss -2.44e-19
C10841 avdd.n7947 avss 0.0422f
C10842 avdd.n7948 avss 0.019f
C10843 avdd.n7949 avss -1.8e-19
C10844 avdd.n7950 avss 0.0197f
C10845 avdd.n7951 avss -2.44e-19
C10846 avdd.n7952 avss -2.33e-19
C10847 avdd.n7953 avss -2.33e-19
C10848 avdd.n7954 avss -1.48e-19
C10849 avdd.n7955 avss -1.27e-19
C10850 avdd.n7956 avss 0.00203f
C10851 avdd.n7957 avss -0.00128f
C10852 avdd.n7958 avss -4.76e-19
C10853 avdd.n7959 avss -2.22e-19
C10854 avdd.n7960 avss 0.0192f
C10855 avdd.n7961 avss -2.22e-19
C10856 avdd.n7962 avss 0.0148f
C10857 avdd.n7963 avss 0.0182f
C10858 avdd.n7964 avss -1.8e-19
C10859 avdd.n7965 avss -2.54e-19
C10860 avdd.n7966 avss -2.54e-19
C10861 avdd.n7967 avss -1.8e-19
C10862 avdd.n7968 avss -1.16e-19
C10863 avdd.n7969 avss -2.33e-19
C10864 avdd.n7970 avss 0.0342f
C10865 avdd.n7971 avss 0.0049f
C10866 avdd.n7972 avss -8.47e-19
C10867 avdd.n7973 avss -3.39e-19
C10868 avdd.n7974 avss -3.07e-19
C10869 avdd.n7975 avss -1.59e-19
C10870 avdd.n7976 avss -1.8e-19
C10871 avdd.n7977 avss 0.0192f
C10872 avdd.n7978 avss -1.59e-19
C10873 avdd.n7979 avss -1.8e-19
C10874 avdd.n7980 avss 0.00875f
C10875 avdd.n7981 avss 0.0111f
C10876 avdd.n7982 avss 0.0154f
C10877 avdd.n7983 avss 0.0183f
C10878 avdd.n7984 avss -1.8e-19
C10879 avdd.n7985 avss -2.22e-19
C10880 avdd.n7986 avss -2.22e-19
C10881 avdd.n7987 avss -1.8e-19
C10882 avdd.n7988 avss -2.01e-19
C10883 avdd.n7989 avss -3.18e-19
C10884 avdd.n7990 avss 0.03f
C10885 avdd.n7991 avss 0.00899f
C10886 avdd.n7992 avss -7.52e-19
C10887 avdd.n7993 avss -2.96e-19
C10888 avdd.n7994 avss -1.8e-19
C10889 avdd.n7995 avss -1.8e-19
C10890 avdd.n7996 avss 0.00873f
C10891 avdd.n7997 avss 0.0111f
C10892 avdd.n7998 avss 0.0154f
C10893 avdd.n7999 avss 0.0191f
C10894 avdd.n8000 avss -1.8e-19
C10895 avdd.n8001 avss 0.0184f
C10896 avdd.n8002 avss -1.38e-19
C10897 avdd.n8003 avss -1.8e-19
C10898 avdd.n8004 avss -2.44e-19
C10899 avdd.n8005 avss -2.44e-19
C10900 avdd.n8006 avss -1.8e-19
C10901 avdd.n8007 avss -1.38e-19
C10902 avdd.n8008 avss -3.49e-19
C10903 avdd.n8010 avss 0.0269f
C10904 avdd.n8011 avss 0.00869f
C10905 avdd.n8012 avss 0.00378f
C10906 avdd.n8013 avss 0.0346f
C10907 avdd.n8014 avss -8.47e-19
C10908 avdd.n8015 avss -3.39e-19
C10909 avdd.n8016 avss -8.47e-19
C10910 avdd.n8017 avss 3e-19
C10911 avdd.n8018 avss 0.0388f
C10912 avdd.n8019 avss -3.39e-19
C10913 avdd.n8020 avss -6.46e-19
C10914 avdd.n8021 avss -5.82e-19
C10915 avdd.n8022 avss -3.39e-19
C10916 avdd.n8023 avss -8.47e-19
C10917 avdd.n8024 avss -0.00113f
C10918 avdd.n8025 avss -0.00512f
C10919 avdd.n8026 avss 0.0382f
C10920 avdd.n8027 avss -0.148f
C10921 avdd.n8028 avss -0.179f
C10922 avdd.n8029 avss -0.00173f
C10923 avdd.n8031 avss 0.0384f
C10924 avdd.n8032 avss -2.44e-19
C10925 avdd.n8033 avss 0.0422f
C10926 avdd.n8034 avss 0.019f
C10927 avdd.n8035 avss -1.8e-19
C10928 avdd.n8036 avss 0.0197f
C10929 avdd.n8037 avss -2.44e-19
C10930 avdd.n8038 avss -2.33e-19
C10931 avdd.n8039 avss -2.33e-19
C10932 avdd.n8040 avss -1.48e-19
C10933 avdd.n8041 avss -1.27e-19
C10934 avdd.n8042 avss 0.00203f
C10935 avdd.n8043 avss -0.00128f
C10936 avdd.n8044 avss -4.76e-19
C10937 avdd.n8045 avss -2.22e-19
C10938 avdd.n8046 avss 0.0192f
C10939 avdd.n8047 avss -2.22e-19
C10940 avdd.n8048 avss 0.0148f
C10941 avdd.n8049 avss 0.0182f
C10942 avdd.n8050 avss -1.8e-19
C10943 avdd.n8051 avss -2.54e-19
C10944 avdd.n8052 avss -2.54e-19
C10945 avdd.n8053 avss -1.8e-19
C10946 avdd.n8054 avss -1.16e-19
C10947 avdd.n8055 avss -2.33e-19
C10948 avdd.n8056 avss 0.0342f
C10949 avdd.n8057 avss 0.0049f
C10950 avdd.n8058 avss -8.47e-19
C10951 avdd.n8059 avss -3.39e-19
C10952 avdd.n8060 avss -3.07e-19
C10953 avdd.n8061 avss -1.59e-19
C10954 avdd.n8062 avss -1.8e-19
C10955 avdd.n8063 avss 0.0192f
C10956 avdd.n8064 avss -1.59e-19
C10957 avdd.n8065 avss -1.8e-19
C10958 avdd.n8066 avss 0.00875f
C10959 avdd.n8067 avss 0.0111f
C10960 avdd.n8068 avss 0.0154f
C10961 avdd.n8069 avss 0.0183f
C10962 avdd.n8070 avss -1.8e-19
C10963 avdd.n8071 avss -2.22e-19
C10964 avdd.n8072 avss -2.22e-19
C10965 avdd.n8073 avss -1.8e-19
C10966 avdd.n8074 avss -2.01e-19
C10967 avdd.n8075 avss -3.18e-19
C10968 avdd.n8076 avss 0.03f
C10969 avdd.n8077 avss 0.00899f
C10970 avdd.n8078 avss -7.52e-19
C10971 avdd.n8079 avss -2.96e-19
C10972 avdd.n8080 avss -1.8e-19
C10973 avdd.n8081 avss -1.8e-19
C10974 avdd.n8082 avss 0.00873f
C10975 avdd.n8083 avss 0.0111f
C10976 avdd.n8084 avss 0.0154f
C10977 avdd.n8085 avss 0.0191f
C10978 avdd.n8086 avss -1.8e-19
C10979 avdd.n8087 avss 0.0184f
C10980 avdd.n8088 avss -1.38e-19
C10981 avdd.n8089 avss -1.8e-19
C10982 avdd.n8090 avss -2.44e-19
C10983 avdd.n8091 avss -2.44e-19
C10984 avdd.n8092 avss -1.8e-19
C10985 avdd.n8093 avss -1.38e-19
C10986 avdd.n8094 avss -3.49e-19
C10987 avdd.n8096 avss 0.0269f
C10988 avdd.n8097 avss 0.00869f
C10989 avdd.n8098 avss 0.00378f
C10990 avdd.n8099 avss 0.0346f
C10991 avdd.n8100 avss -8.47e-19
C10992 avdd.n8101 avss -3.39e-19
C10993 avdd.n8102 avss -8.47e-19
C10994 avdd.n8103 avss 3e-19
C10995 avdd.n8104 avss 0.0388f
C10996 avdd.n8105 avss -3.39e-19
C10997 avdd.n8106 avss -6.46e-19
C10998 avdd.n8107 avss -5.82e-19
C10999 avdd.n8108 avss -3.39e-19
C11000 avdd.n8109 avss -8.47e-19
C11001 avdd.n8110 avss -0.00113f
C11002 avdd.n8111 avss -0.00512f
C11003 avdd.n8112 avss 0.0382f
C11004 avdd.n8113 avss -0.149f
C11005 avdd.n8114 avss -0.181f
C11006 avdd.n8115 avss -0.00173f
C11007 avdd.n8117 avss 0.0384f
C11008 avdd.n8118 avss -2.44e-19
C11009 avdd.n8119 avss 0.0422f
C11010 avdd.n8120 avss 0.019f
C11011 avdd.n8121 avss -1.8e-19
C11012 avdd.n8122 avss 0.0197f
C11013 avdd.n8123 avss -2.44e-19
C11014 avdd.n8124 avss -2.33e-19
C11015 avdd.n8125 avss -2.33e-19
C11016 avdd.n8126 avss -1.48e-19
C11017 avdd.n8127 avss -1.27e-19
C11018 avdd.n8128 avss 0.00203f
C11019 avdd.n8129 avss -0.00128f
C11020 avdd.n8130 avss -4.76e-19
C11021 avdd.n8131 avss -2.22e-19
C11022 avdd.n8132 avss 0.0192f
C11023 avdd.n8133 avss -2.22e-19
C11024 avdd.n8134 avss 0.0148f
C11025 avdd.n8135 avss 0.0182f
C11026 avdd.n8136 avss -1.8e-19
C11027 avdd.n8137 avss -2.54e-19
C11028 avdd.n8138 avss -2.54e-19
C11029 avdd.n8139 avss -1.8e-19
C11030 avdd.n8140 avss -1.16e-19
C11031 avdd.n8141 avss -2.33e-19
C11032 avdd.n8142 avss 0.0342f
C11033 avdd.n8143 avss 0.0049f
C11034 avdd.n8144 avss -8.47e-19
C11035 avdd.n8145 avss -3.39e-19
C11036 avdd.n8146 avss -3.07e-19
C11037 avdd.n8147 avss -1.59e-19
C11038 avdd.n8148 avss -1.8e-19
C11039 avdd.n8149 avss 0.0192f
C11040 avdd.n8150 avss -1.59e-19
C11041 avdd.n8151 avss -1.8e-19
C11042 avdd.n8152 avss 0.00875f
C11043 avdd.n8153 avss 0.0111f
C11044 avdd.n8154 avss 0.0154f
C11045 avdd.n8155 avss 0.0183f
C11046 avdd.n8156 avss -1.8e-19
C11047 avdd.n8157 avss -2.22e-19
C11048 avdd.n8158 avss -2.22e-19
C11049 avdd.n8159 avss -1.8e-19
C11050 avdd.n8160 avss -2.01e-19
C11051 avdd.n8161 avss -3.18e-19
C11052 avdd.n8162 avss 0.03f
C11053 avdd.n8163 avss 0.00899f
C11054 avdd.n8164 avss -7.52e-19
C11055 avdd.n8165 avss -2.96e-19
C11056 avdd.n8166 avss -1.8e-19
C11057 avdd.n8167 avss -1.8e-19
C11058 avdd.n8168 avss 0.00873f
C11059 avdd.n8169 avss 0.0111f
C11060 avdd.n8170 avss 0.0154f
C11061 avdd.n8171 avss 0.0191f
C11062 avdd.n8172 avss -1.8e-19
C11063 avdd.n8173 avss 0.0184f
C11064 avdd.n8174 avss -1.38e-19
C11065 avdd.n8175 avss -1.8e-19
C11066 avdd.n8176 avss -2.44e-19
C11067 avdd.n8177 avss -2.44e-19
C11068 avdd.n8178 avss -1.8e-19
C11069 avdd.n8179 avss -1.38e-19
C11070 avdd.n8180 avss -3.49e-19
C11071 avdd.n8182 avss 0.0269f
C11072 avdd.n8183 avss 0.00869f
C11073 avdd.n8184 avss 0.00378f
C11074 avdd.n8185 avss 0.0346f
C11075 avdd.n8186 avss -8.47e-19
C11076 avdd.n8187 avss -3.39e-19
C11077 avdd.n8188 avss -8.47e-19
C11078 avdd.n8189 avss 3e-19
C11079 avdd.n8190 avss 0.0388f
C11080 avdd.n8191 avss -3.39e-19
C11081 avdd.n8192 avss -6.46e-19
C11082 avdd.n8193 avss -5.82e-19
C11083 avdd.n8194 avss -3.39e-19
C11084 avdd.n8195 avss -8.47e-19
C11085 avdd.n8196 avss -0.00113f
C11086 avdd.n8197 avss -0.00512f
C11087 avdd.n8198 avss 0.0382f
C11088 avdd.n8199 avss -0.149f
C11089 avdd.n8200 avss -0.18f
C11090 avdd.n8201 avss -0.00173f
C11091 avdd.n8203 avss 0.0384f
C11092 avdd.n8204 avss -2.44e-19
C11093 avdd.n8205 avss 0.0422f
C11094 avdd.n8206 avss 0.019f
C11095 avdd.n8207 avss -1.8e-19
C11096 avdd.n8208 avss 0.0197f
C11097 avdd.n8209 avss -2.44e-19
C11098 avdd.n8210 avss -2.33e-19
C11099 avdd.n8211 avss -2.33e-19
C11100 avdd.n8212 avss -1.48e-19
C11101 avdd.n8213 avss -1.27e-19
C11102 avdd.n8214 avss 0.00203f
C11103 avdd.n8215 avss -0.00128f
C11104 avdd.n8216 avss -4.76e-19
C11105 avdd.n8217 avss -2.22e-19
C11106 avdd.n8218 avss 0.0192f
C11107 avdd.n8219 avss -2.22e-19
C11108 avdd.n8220 avss 0.0148f
C11109 avdd.n8221 avss 0.0182f
C11110 avdd.n8222 avss -1.8e-19
C11111 avdd.n8223 avss -2.54e-19
C11112 avdd.n8224 avss -2.54e-19
C11113 avdd.n8225 avss -1.8e-19
C11114 avdd.n8226 avss -1.16e-19
C11115 avdd.n8227 avss -2.33e-19
C11116 avdd.n8228 avss 0.0342f
C11117 avdd.n8229 avss 0.0049f
C11118 avdd.n8230 avss -8.47e-19
C11119 avdd.n8231 avss -3.39e-19
C11120 avdd.n8232 avss -3.07e-19
C11121 avdd.n8233 avss -1.59e-19
C11122 avdd.n8234 avss -1.8e-19
C11123 avdd.n8235 avss 0.0192f
C11124 avdd.n8236 avss -1.59e-19
C11125 avdd.n8237 avss -1.8e-19
C11126 avdd.n8238 avss 0.00875f
C11127 avdd.n8239 avss 0.0111f
C11128 avdd.n8240 avss 0.0154f
C11129 avdd.n8241 avss 0.0183f
C11130 avdd.n8242 avss -1.8e-19
C11131 avdd.n8243 avss -2.22e-19
C11132 avdd.n8244 avss -2.22e-19
C11133 avdd.n8245 avss -1.8e-19
C11134 avdd.n8246 avss -2.01e-19
C11135 avdd.n8247 avss -3.18e-19
C11136 avdd.n8248 avss 0.03f
C11137 avdd.n8249 avss 0.00899f
C11138 avdd.n8250 avss -7.52e-19
C11139 avdd.n8251 avss -2.96e-19
C11140 avdd.n8252 avss -1.8e-19
C11141 avdd.n8253 avss -1.8e-19
C11142 avdd.n8254 avss 0.00873f
C11143 avdd.n8255 avss 0.0111f
C11144 avdd.n8256 avss 0.0154f
C11145 avdd.n8257 avss 0.0191f
C11146 avdd.n8258 avss -1.8e-19
C11147 avdd.n8259 avss 0.0184f
C11148 avdd.n8260 avss -1.38e-19
C11149 avdd.n8261 avss -1.8e-19
C11150 avdd.n8262 avss -2.44e-19
C11151 avdd.n8263 avss -2.44e-19
C11152 avdd.n8264 avss -1.8e-19
C11153 avdd.n8265 avss -1.38e-19
C11154 avdd.n8266 avss -3.49e-19
C11155 avdd.n8268 avss 0.0269f
C11156 avdd.n8269 avss 0.00869f
C11157 avdd.n8270 avss 0.00378f
C11158 avdd.n8271 avss 0.0346f
C11159 avdd.n8272 avss -8.47e-19
C11160 avdd.n8273 avss -3.39e-19
C11161 avdd.n8274 avss -8.47e-19
C11162 avdd.n8275 avss 3e-19
C11163 avdd.n8276 avss 0.0388f
C11164 avdd.n8277 avss -3.39e-19
C11165 avdd.n8278 avss -6.46e-19
C11166 avdd.n8279 avss -5.82e-19
C11167 avdd.n8280 avss -3.39e-19
C11168 avdd.n8281 avss -8.47e-19
C11169 avdd.n8282 avss -0.00113f
C11170 avdd.n8283 avss -0.00512f
C11171 avdd.n8284 avss 0.0382f
C11172 avdd.n8285 avss -0.149f
C11173 avdd.n8286 avss -0.181f
C11174 avdd.n8287 avss -0.00173f
C11175 avdd.n8289 avss 0.0384f
C11176 avdd.n8290 avss -2.44e-19
C11177 avdd.n8291 avss 0.0422f
C11178 avdd.n8292 avss 0.019f
C11179 avdd.n8293 avss -1.8e-19
C11180 avdd.n8294 avss 0.0197f
C11181 avdd.n8295 avss -2.44e-19
C11182 avdd.n8296 avss -2.33e-19
C11183 avdd.n8297 avss -2.33e-19
C11184 avdd.n8298 avss -1.48e-19
C11185 avdd.n8299 avss -1.27e-19
C11186 avdd.n8300 avss 0.00203f
C11187 avdd.n8301 avss -0.00128f
C11188 avdd.n8302 avss -4.76e-19
C11189 avdd.n8303 avss -2.22e-19
C11190 avdd.n8304 avss 0.0192f
C11191 avdd.n8305 avss -2.22e-19
C11192 avdd.n8306 avss 0.0148f
C11193 avdd.n8307 avss 0.0182f
C11194 avdd.n8308 avss -1.8e-19
C11195 avdd.n8309 avss -2.54e-19
C11196 avdd.n8310 avss -2.54e-19
C11197 avdd.n8311 avss -1.8e-19
C11198 avdd.n8312 avss -1.16e-19
C11199 avdd.n8313 avss -2.33e-19
C11200 avdd.n8314 avss 0.0342f
C11201 avdd.n8315 avss 0.0049f
C11202 avdd.n8316 avss -8.47e-19
C11203 avdd.n8317 avss -3.39e-19
C11204 avdd.n8318 avss -3.07e-19
C11205 avdd.n8319 avss -1.59e-19
C11206 avdd.n8320 avss -1.8e-19
C11207 avdd.n8321 avss 0.0192f
C11208 avdd.n8322 avss -1.59e-19
C11209 avdd.n8323 avss -1.8e-19
C11210 avdd.n8324 avss 0.00875f
C11211 avdd.n8325 avss 0.0111f
C11212 avdd.n8326 avss 0.0154f
C11213 avdd.n8327 avss 0.0183f
C11214 avdd.n8328 avss -1.8e-19
C11215 avdd.n8329 avss -2.22e-19
C11216 avdd.n8330 avss -2.22e-19
C11217 avdd.n8331 avss -1.8e-19
C11218 avdd.n8332 avss -2.01e-19
C11219 avdd.n8333 avss -3.18e-19
C11220 avdd.n8334 avss 0.03f
C11221 avdd.n8335 avss 0.00899f
C11222 avdd.n8336 avss -7.52e-19
C11223 avdd.n8337 avss -2.96e-19
C11224 avdd.n8338 avss -1.8e-19
C11225 avdd.n8339 avss -1.8e-19
C11226 avdd.n8340 avss 0.00873f
C11227 avdd.n8341 avss 0.0111f
C11228 avdd.n8342 avss 0.0154f
C11229 avdd.n8343 avss 0.0191f
C11230 avdd.n8344 avss -1.8e-19
C11231 avdd.n8345 avss 0.0184f
C11232 avdd.n8346 avss -1.38e-19
C11233 avdd.n8347 avss -1.8e-19
C11234 avdd.n8348 avss -2.44e-19
C11235 avdd.n8349 avss -2.44e-19
C11236 avdd.n8350 avss -1.8e-19
C11237 avdd.n8351 avss -1.38e-19
C11238 avdd.n8352 avss -3.49e-19
C11239 avdd.n8354 avss 0.0269f
C11240 avdd.n8355 avss 0.00869f
C11241 avdd.n8356 avss 0.00378f
C11242 avdd.n8357 avss 0.0346f
C11243 avdd.n8358 avss -8.47e-19
C11244 avdd.n8359 avss -3.39e-19
C11245 avdd.n8360 avss -8.47e-19
C11246 avdd.n8361 avss 3e-19
C11247 avdd.n8362 avss 0.0388f
C11248 avdd.n8363 avss -3.39e-19
C11249 avdd.n8364 avss -6.46e-19
C11250 avdd.n8365 avss -5.82e-19
C11251 avdd.n8366 avss -3.39e-19
C11252 avdd.n8367 avss -8.47e-19
C11253 avdd.n8368 avss -0.00113f
C11254 avdd.n8369 avss -0.00512f
C11255 avdd.n8370 avss 0.0382f
C11256 avdd.n8371 avss -0.149f
C11257 avdd.n8372 avss -0.181f
C11258 avdd.n8373 avss -0.00173f
C11259 avdd.n8375 avss 0.0384f
C11260 avdd.n8376 avss -2.44e-19
C11261 avdd.n8377 avss 0.0422f
C11262 avdd.n8378 avss 0.019f
C11263 avdd.n8379 avss -1.8e-19
C11264 avdd.n8380 avss 0.0197f
C11265 avdd.n8381 avss -2.44e-19
C11266 avdd.n8382 avss -2.33e-19
C11267 avdd.n8383 avss -2.33e-19
C11268 avdd.n8384 avss -1.48e-19
C11269 avdd.n8385 avss -1.27e-19
C11270 avdd.n8386 avss 0.00203f
C11271 avdd.n8387 avss -0.00128f
C11272 avdd.n8388 avss -4.76e-19
C11273 avdd.n8389 avss -2.22e-19
C11274 avdd.n8390 avss 0.0192f
C11275 avdd.n8391 avss -2.22e-19
C11276 avdd.n8392 avss 0.0148f
C11277 avdd.n8393 avss 0.0182f
C11278 avdd.n8394 avss -1.8e-19
C11279 avdd.n8395 avss -2.54e-19
C11280 avdd.n8396 avss -2.54e-19
C11281 avdd.n8397 avss -1.8e-19
C11282 avdd.n8398 avss -1.16e-19
C11283 avdd.n8399 avss -2.33e-19
C11284 avdd.n8400 avss 0.0342f
C11285 avdd.n8401 avss 0.0049f
C11286 avdd.n8402 avss -8.47e-19
C11287 avdd.n8403 avss -3.39e-19
C11288 avdd.n8404 avss -3.07e-19
C11289 avdd.n8405 avss -1.59e-19
C11290 avdd.n8406 avss -1.8e-19
C11291 avdd.n8407 avss 0.0192f
C11292 avdd.n8408 avss -1.59e-19
C11293 avdd.n8409 avss -1.8e-19
C11294 avdd.n8410 avss 0.00875f
C11295 avdd.n8411 avss 0.0111f
C11296 avdd.n8412 avss 0.0154f
C11297 avdd.n8413 avss 0.0183f
C11298 avdd.n8414 avss -1.8e-19
C11299 avdd.n8415 avss -2.22e-19
C11300 avdd.n8416 avss -2.22e-19
C11301 avdd.n8417 avss -1.8e-19
C11302 avdd.n8418 avss -2.01e-19
C11303 avdd.n8419 avss -3.18e-19
C11304 avdd.n8420 avss 0.03f
C11305 avdd.n8421 avss 0.00899f
C11306 avdd.n8422 avss -7.52e-19
C11307 avdd.n8423 avss -2.96e-19
C11308 avdd.n8424 avss -1.8e-19
C11309 avdd.n8425 avss -1.8e-19
C11310 avdd.n8426 avss 0.00873f
C11311 avdd.n8427 avss 0.0111f
C11312 avdd.n8428 avss 0.0154f
C11313 avdd.n8429 avss 0.0191f
C11314 avdd.n8430 avss -1.8e-19
C11315 avdd.n8431 avss 0.0184f
C11316 avdd.n8432 avss -1.38e-19
C11317 avdd.n8433 avss -1.8e-19
C11318 avdd.n8434 avss -2.44e-19
C11319 avdd.n8435 avss -2.44e-19
C11320 avdd.n8436 avss -1.8e-19
C11321 avdd.n8437 avss -1.38e-19
C11322 avdd.n8438 avss -3.49e-19
C11323 avdd.n8440 avss 0.0269f
C11324 avdd.n8441 avss 0.00869f
C11325 avdd.n8442 avss 0.00378f
C11326 avdd.n8443 avss 0.0346f
C11327 avdd.n8444 avss -8.47e-19
C11328 avdd.n8445 avss -3.39e-19
C11329 avdd.n8446 avss -8.47e-19
C11330 avdd.n8447 avss 3e-19
C11331 avdd.n8448 avss 0.0388f
C11332 avdd.n8449 avss -3.39e-19
C11333 avdd.n8450 avss -6.46e-19
C11334 avdd.n8451 avss -5.82e-19
C11335 avdd.n8452 avss -3.39e-19
C11336 avdd.n8453 avss -8.47e-19
C11337 avdd.n8454 avss -0.00113f
C11338 avdd.n8455 avss -0.00512f
C11339 avdd.n8456 avss 0.0382f
C11340 avdd.n8457 avss -0.151f
C11341 avdd.n8458 avss -0.183f
C11342 avdd.n8459 avss -0.00173f
C11343 avdd.n8461 avss 0.0384f
C11344 avdd.n8462 avss -2.44e-19
C11345 avdd.n8463 avss 0.0422f
C11346 avdd.n8464 avss 0.019f
C11347 avdd.n8465 avss -1.8e-19
C11348 avdd.n8466 avss 0.0197f
C11349 avdd.n8467 avss -2.44e-19
C11350 avdd.n8468 avss -2.33e-19
C11351 avdd.n8469 avss -2.33e-19
C11352 avdd.n8470 avss -1.48e-19
C11353 avdd.n8471 avss -1.27e-19
C11354 avdd.n8472 avss 0.00203f
C11355 avdd.n8473 avss -0.00128f
C11356 avdd.n8474 avss -4.76e-19
C11357 avdd.n8475 avss -2.22e-19
C11358 avdd.n8476 avss 0.0192f
C11359 avdd.n8477 avss -2.22e-19
C11360 avdd.n8478 avss 0.0148f
C11361 avdd.n8479 avss 0.0182f
C11362 avdd.n8480 avss -1.8e-19
C11363 avdd.n8481 avss -2.54e-19
C11364 avdd.n8482 avss -2.54e-19
C11365 avdd.n8483 avss -1.8e-19
C11366 avdd.n8484 avss -1.16e-19
C11367 avdd.n8485 avss -2.33e-19
C11368 avdd.n8486 avss 0.0342f
C11369 avdd.n8487 avss 0.0049f
C11370 avdd.n8488 avss -8.47e-19
C11371 avdd.n8489 avss -3.39e-19
C11372 avdd.n8490 avss -3.07e-19
C11373 avdd.n8491 avss -1.59e-19
C11374 avdd.n8492 avss -1.8e-19
C11375 avdd.n8493 avss 0.0192f
C11376 avdd.n8494 avss -1.59e-19
C11377 avdd.n8495 avss -1.8e-19
C11378 avdd.n8496 avss 0.00875f
C11379 avdd.n8497 avss 0.0111f
C11380 avdd.n8498 avss 0.0154f
C11381 avdd.n8499 avss 0.0183f
C11382 avdd.n8500 avss -1.8e-19
C11383 avdd.n8501 avss -2.22e-19
C11384 avdd.n8502 avss -2.22e-19
C11385 avdd.n8503 avss -1.8e-19
C11386 avdd.n8504 avss -2.01e-19
C11387 avdd.n8505 avss -3.18e-19
C11388 avdd.n8506 avss 0.03f
C11389 avdd.n8507 avss 0.00899f
C11390 avdd.n8508 avss -7.52e-19
C11391 avdd.n8509 avss -2.96e-19
C11392 avdd.n8510 avss -1.8e-19
C11393 avdd.n8511 avss -1.8e-19
C11394 avdd.n8512 avss 0.00873f
C11395 avdd.n8513 avss 0.0111f
C11396 avdd.n8514 avss 0.0154f
C11397 avdd.n8515 avss 0.0191f
C11398 avdd.n8516 avss -1.8e-19
C11399 avdd.n8517 avss 0.0184f
C11400 avdd.n8518 avss -1.38e-19
C11401 avdd.n8519 avss -1.8e-19
C11402 avdd.n8520 avss -2.44e-19
C11403 avdd.n8521 avss -2.44e-19
C11404 avdd.n8522 avss -1.8e-19
C11405 avdd.n8523 avss -1.38e-19
C11406 avdd.n8524 avss -3.49e-19
C11407 avdd.n8526 avss 0.0269f
C11408 avdd.n8527 avss 0.00869f
C11409 avdd.n8528 avss 0.00378f
C11410 avdd.n8529 avss 0.0346f
C11411 avdd.n8530 avss -8.47e-19
C11412 avdd.n8531 avss -3.39e-19
C11413 avdd.n8532 avss -8.47e-19
C11414 avdd.n8533 avss 3e-19
C11415 avdd.n8534 avss 0.0388f
C11416 avdd.n8535 avss -3.39e-19
C11417 avdd.n8536 avss -6.46e-19
C11418 avdd.n8537 avss -5.82e-19
C11419 avdd.n8538 avss -3.39e-19
C11420 avdd.n8539 avss -8.47e-19
C11421 avdd.n8540 avss -0.00113f
C11422 avdd.n8541 avss -0.00512f
C11423 avdd.n8542 avss 0.0382f
C11424 avdd.n8543 avss -0.151f
C11425 avdd.n8544 avss -0.183f
C11426 avdd.n8545 avss -0.00173f
C11427 avdd.n8547 avss 0.0384f
C11428 avdd.n8548 avss -2.44e-19
C11429 avdd.n8549 avss 0.0422f
C11430 avdd.n8550 avss 0.019f
C11431 avdd.n8551 avss -1.8e-19
C11432 avdd.n8552 avss 0.0197f
C11433 avdd.n8553 avss -2.44e-19
C11434 avdd.n8554 avss -2.33e-19
C11435 avdd.n8555 avss -2.33e-19
C11436 avdd.n8556 avss -1.48e-19
C11437 avdd.n8557 avss -1.27e-19
C11438 avdd.n8558 avss 0.00203f
C11439 avdd.n8559 avss -0.00128f
C11440 avdd.n8560 avss -4.76e-19
C11441 avdd.n8561 avss -2.22e-19
C11442 avdd.n8562 avss 0.0192f
C11443 avdd.n8563 avss -2.22e-19
C11444 avdd.n8564 avss 0.0148f
C11445 avdd.n8565 avss 0.0182f
C11446 avdd.n8566 avss -1.8e-19
C11447 avdd.n8567 avss -2.54e-19
C11448 avdd.n8568 avss -2.54e-19
C11449 avdd.n8569 avss -1.8e-19
C11450 avdd.n8570 avss -1.16e-19
C11451 avdd.n8571 avss -2.33e-19
C11452 avdd.n8572 avss 0.0342f
C11453 avdd.n8573 avss 0.0049f
C11454 avdd.n8574 avss -8.47e-19
C11455 avdd.n8575 avss -3.39e-19
C11456 avdd.n8576 avss -3.07e-19
C11457 avdd.n8577 avss -1.59e-19
C11458 avdd.n8578 avss -1.8e-19
C11459 avdd.n8579 avss 0.0192f
C11460 avdd.n8580 avss -1.59e-19
C11461 avdd.n8581 avss -1.8e-19
C11462 avdd.n8582 avss 0.00875f
C11463 avdd.n8583 avss 0.0111f
C11464 avdd.n8584 avss 0.0154f
C11465 avdd.n8585 avss 0.0183f
C11466 avdd.n8586 avss -1.8e-19
C11467 avdd.n8587 avss -2.22e-19
C11468 avdd.n8588 avss -2.22e-19
C11469 avdd.n8589 avss -1.8e-19
C11470 avdd.n8590 avss -2.01e-19
C11471 avdd.n8591 avss -3.18e-19
C11472 avdd.n8592 avss 0.03f
C11473 avdd.n8593 avss 0.00899f
C11474 avdd.n8594 avss -7.52e-19
C11475 avdd.n8595 avss -2.96e-19
C11476 avdd.n8596 avss -1.8e-19
C11477 avdd.n8597 avss -1.8e-19
C11478 avdd.n8598 avss 0.00873f
C11479 avdd.n8599 avss 0.0111f
C11480 avdd.n8600 avss 0.0154f
C11481 avdd.n8601 avss 0.0191f
C11482 avdd.n8602 avss -1.8e-19
C11483 avdd.n8603 avss 0.0184f
C11484 avdd.n8604 avss -1.38e-19
C11485 avdd.n8605 avss -1.8e-19
C11486 avdd.n8606 avss -2.44e-19
C11487 avdd.n8607 avss -2.44e-19
C11488 avdd.n8608 avss -1.8e-19
C11489 avdd.n8609 avss -1.38e-19
C11490 avdd.n8610 avss -3.49e-19
C11491 avdd.n8612 avss 0.0269f
C11492 avdd.n8613 avss 0.00869f
C11493 avdd.n8614 avss 0.00378f
C11494 avdd.n8615 avss 0.0346f
C11495 avdd.n8616 avss -8.47e-19
C11496 avdd.n8617 avss -3.39e-19
C11497 avdd.n8618 avss -8.47e-19
C11498 avdd.n8619 avss 3e-19
C11499 avdd.n8620 avss 0.0388f
C11500 avdd.n8621 avss -3.39e-19
C11501 avdd.n8622 avss -6.46e-19
C11502 avdd.n8623 avss -5.82e-19
C11503 avdd.n8624 avss -3.39e-19
C11504 avdd.n8625 avss -8.47e-19
C11505 avdd.n8626 avss -0.00113f
C11506 avdd.n8627 avss -0.00512f
C11507 avdd.n8628 avss 0.0382f
C11508 avdd.n8629 avss -0.151f
C11509 avdd.n8630 avss -0.183f
C11510 avdd.n8631 avss -0.00173f
C11511 avdd.n8633 avss 0.0384f
C11512 avdd.n8634 avss -2.44e-19
C11513 avdd.n8635 avss 0.0422f
C11514 avdd.n8636 avss 0.019f
C11515 avdd.n8637 avss -1.8e-19
C11516 avdd.n8638 avss 0.0197f
C11517 avdd.n8639 avss -2.44e-19
C11518 avdd.n8640 avss -2.33e-19
C11519 avdd.n8641 avss -2.33e-19
C11520 avdd.n8642 avss -1.48e-19
C11521 avdd.n8643 avss -1.27e-19
C11522 avdd.n8644 avss 0.00203f
C11523 avdd.n8645 avss -0.00128f
C11524 avdd.n8646 avss -4.76e-19
C11525 avdd.n8647 avss -2.22e-19
C11526 avdd.n8648 avss 0.0192f
C11527 avdd.n8649 avss -2.22e-19
C11528 avdd.n8650 avss 0.0148f
C11529 avdd.n8651 avss 0.0182f
C11530 avdd.n8652 avss -1.8e-19
C11531 avdd.n8653 avss -2.54e-19
C11532 avdd.n8654 avss -2.54e-19
C11533 avdd.n8655 avss -1.8e-19
C11534 avdd.n8656 avss -1.16e-19
C11535 avdd.n8657 avss -2.33e-19
C11536 avdd.n8658 avss 0.0342f
C11537 avdd.n8659 avss 0.0049f
C11538 avdd.n8660 avss -8.47e-19
C11539 avdd.n8661 avss -3.39e-19
C11540 avdd.n8662 avss -3.07e-19
C11541 avdd.n8663 avss -1.59e-19
C11542 avdd.n8664 avss -1.8e-19
C11543 avdd.n8665 avss 0.0192f
C11544 avdd.n8666 avss -1.59e-19
C11545 avdd.n8667 avss -1.8e-19
C11546 avdd.n8668 avss 0.00875f
C11547 avdd.n8669 avss 0.0111f
C11548 avdd.n8670 avss 0.0154f
C11549 avdd.n8671 avss 0.0183f
C11550 avdd.n8672 avss -1.8e-19
C11551 avdd.n8673 avss -2.22e-19
C11552 avdd.n8674 avss -2.22e-19
C11553 avdd.n8675 avss -1.8e-19
C11554 avdd.n8676 avss -2.01e-19
C11555 avdd.n8677 avss -3.18e-19
C11556 avdd.n8678 avss 0.03f
C11557 avdd.n8679 avss 0.00899f
C11558 avdd.n8680 avss -7.52e-19
C11559 avdd.n8681 avss -2.96e-19
C11560 avdd.n8682 avss -1.8e-19
C11561 avdd.n8683 avss -1.8e-19
C11562 avdd.n8684 avss 0.00873f
C11563 avdd.n8685 avss 0.0111f
C11564 avdd.n8686 avss 0.0154f
C11565 avdd.n8687 avss 0.0191f
C11566 avdd.n8688 avss -1.8e-19
C11567 avdd.n8689 avss 0.0184f
C11568 avdd.n8690 avss -1.38e-19
C11569 avdd.n8691 avss -1.8e-19
C11570 avdd.n8692 avss -2.44e-19
C11571 avdd.n8693 avss -2.44e-19
C11572 avdd.n8694 avss -1.8e-19
C11573 avdd.n8695 avss -1.38e-19
C11574 avdd.n8696 avss -3.49e-19
C11575 avdd.n8698 avss 0.0269f
C11576 avdd.n8699 avss 0.00869f
C11577 avdd.n8700 avss 0.00378f
C11578 avdd.n8701 avss 0.0346f
C11579 avdd.n8702 avss -8.47e-19
C11580 avdd.n8703 avss -3.39e-19
C11581 avdd.n8704 avss -8.47e-19
C11582 avdd.n8705 avss 3e-19
C11583 avdd.n8706 avss 0.0388f
C11584 avdd.n8707 avss -3.39e-19
C11585 avdd.n8708 avss -6.46e-19
C11586 avdd.n8709 avss -5.82e-19
C11587 avdd.n8710 avss -3.39e-19
C11588 avdd.n8711 avss -8.47e-19
C11589 avdd.n8712 avss -0.00113f
C11590 avdd.n8713 avss -0.00512f
C11591 avdd.n8714 avss 0.0382f
C11592 avdd.n8715 avss -0.151f
C11593 avdd.n8716 avss -0.182f
C11594 avdd.n8717 avss -0.00173f
C11595 avdd.n8719 avss 0.0384f
C11596 avdd.n8720 avss -2.44e-19
C11597 avdd.n8721 avss 0.0422f
C11598 avdd.n8722 avss 0.019f
C11599 avdd.n8723 avss -1.8e-19
C11600 avdd.n8724 avss 0.0197f
C11601 avdd.n8725 avss -2.44e-19
C11602 avdd.n8726 avss -2.33e-19
C11603 avdd.n8727 avss -2.33e-19
C11604 avdd.n8728 avss -1.48e-19
C11605 avdd.n8729 avss -1.27e-19
C11606 avdd.n8730 avss 0.00203f
C11607 avdd.n8731 avss -0.00128f
C11608 avdd.n8732 avss -4.76e-19
C11609 avdd.n8733 avss -2.22e-19
C11610 avdd.n8734 avss 0.0192f
C11611 avdd.n8735 avss -2.22e-19
C11612 avdd.n8736 avss 0.0148f
C11613 avdd.n8737 avss 0.0182f
C11614 avdd.n8738 avss -1.8e-19
C11615 avdd.n8739 avss -2.54e-19
C11616 avdd.n8740 avss -2.54e-19
C11617 avdd.n8741 avss -1.8e-19
C11618 avdd.n8742 avss -1.16e-19
C11619 avdd.n8743 avss -2.33e-19
C11620 avdd.n8744 avss 0.0342f
C11621 avdd.n8745 avss 0.0049f
C11622 avdd.n8746 avss -8.47e-19
C11623 avdd.n8747 avss -3.39e-19
C11624 avdd.n8748 avss -3.07e-19
C11625 avdd.n8749 avss -1.59e-19
C11626 avdd.n8750 avss -1.8e-19
C11627 avdd.n8751 avss 0.0192f
C11628 avdd.n8752 avss -1.59e-19
C11629 avdd.n8753 avss -1.8e-19
C11630 avdd.n8754 avss 0.00875f
C11631 avdd.n8755 avss 0.0111f
C11632 avdd.n8756 avss 0.0154f
C11633 avdd.n8757 avss 0.0183f
C11634 avdd.n8758 avss -1.8e-19
C11635 avdd.n8759 avss -2.22e-19
C11636 avdd.n8760 avss -2.22e-19
C11637 avdd.n8761 avss -1.8e-19
C11638 avdd.n8762 avss -2.01e-19
C11639 avdd.n8763 avss -3.18e-19
C11640 avdd.n8764 avss 0.03f
C11641 avdd.n8765 avss 0.00899f
C11642 avdd.n8766 avss -7.52e-19
C11643 avdd.n8767 avss -2.96e-19
C11644 avdd.n8768 avss -1.8e-19
C11645 avdd.n8769 avss -1.8e-19
C11646 avdd.n8770 avss 0.00873f
C11647 avdd.n8771 avss 0.0111f
C11648 avdd.n8772 avss 0.0154f
C11649 avdd.n8773 avss 0.0191f
C11650 avdd.n8774 avss -1.8e-19
C11651 avdd.n8775 avss 0.0184f
C11652 avdd.n8776 avss -1.38e-19
C11653 avdd.n8777 avss -1.8e-19
C11654 avdd.n8778 avss -2.44e-19
C11655 avdd.n8779 avss -2.44e-19
C11656 avdd.n8780 avss -1.8e-19
C11657 avdd.n8781 avss -1.38e-19
C11658 avdd.n8782 avss -3.49e-19
C11659 avdd.n8784 avss 0.0269f
C11660 avdd.n8785 avss 0.00869f
C11661 avdd.n8786 avss 0.00378f
C11662 avdd.n8787 avss 0.0346f
C11663 avdd.n8788 avss -8.47e-19
C11664 avdd.n8789 avss -3.39e-19
C11665 avdd.n8790 avss -8.47e-19
C11666 avdd.n8791 avss 3e-19
C11667 avdd.n8792 avss 0.0388f
C11668 avdd.n8793 avss -3.39e-19
C11669 avdd.n8794 avss -6.46e-19
C11670 avdd.n8795 avss -5.82e-19
C11671 avdd.n8796 avss -3.39e-19
C11672 avdd.n8797 avss -8.47e-19
C11673 avdd.n8798 avss -0.00113f
C11674 avdd.n8799 avss -0.00512f
C11675 avdd.n8800 avss 0.0382f
C11676 avdd.n8801 avss -0.152f
C11677 avdd.n8802 avss -0.184f
C11678 avdd.n8803 avss -0.00173f
C11679 avdd.n8805 avss 0.0384f
C11680 avdd.n8806 avss -2.44e-19
C11681 avdd.n8807 avss 0.0422f
C11682 avdd.n8808 avss 0.019f
C11683 avdd.n8809 avss -1.8e-19
C11684 avdd.n8810 avss 0.0197f
C11685 avdd.n8811 avss -2.44e-19
C11686 avdd.n8812 avss -2.33e-19
C11687 avdd.n8813 avss -2.33e-19
C11688 avdd.n8814 avss -1.48e-19
C11689 avdd.n8815 avss -1.27e-19
C11690 avdd.n8816 avss 0.00203f
C11691 avdd.n8817 avss -0.00128f
C11692 avdd.n8818 avss -4.76e-19
C11693 avdd.n8819 avss -2.22e-19
C11694 avdd.n8820 avss 0.0192f
C11695 avdd.n8821 avss -2.22e-19
C11696 avdd.n8822 avss 0.0148f
C11697 avdd.n8823 avss 0.0182f
C11698 avdd.n8824 avss -1.8e-19
C11699 avdd.n8825 avss -2.54e-19
C11700 avdd.n8826 avss -2.54e-19
C11701 avdd.n8827 avss -1.8e-19
C11702 avdd.n8828 avss -1.16e-19
C11703 avdd.n8829 avss -2.33e-19
C11704 avdd.n8830 avss 0.0342f
C11705 avdd.n8831 avss 0.0049f
C11706 avdd.n8832 avss -8.47e-19
C11707 avdd.n8833 avss -3.39e-19
C11708 avdd.n8834 avss -3.07e-19
C11709 avdd.n8835 avss -1.59e-19
C11710 avdd.n8836 avss -1.8e-19
C11711 avdd.n8837 avss 0.0192f
C11712 avdd.n8838 avss -1.59e-19
C11713 avdd.n8839 avss -1.8e-19
C11714 avdd.n8840 avss 0.00875f
C11715 avdd.n8841 avss 0.0111f
C11716 avdd.n8842 avss 0.0154f
C11717 avdd.n8843 avss 0.0183f
C11718 avdd.n8844 avss -1.8e-19
C11719 avdd.n8845 avss -2.22e-19
C11720 avdd.n8846 avss -2.22e-19
C11721 avdd.n8847 avss -1.8e-19
C11722 avdd.n8848 avss -2.01e-19
C11723 avdd.n8849 avss -3.18e-19
C11724 avdd.n8850 avss 0.03f
C11725 avdd.n8851 avss 0.00899f
C11726 avdd.n8852 avss -7.52e-19
C11727 avdd.n8853 avss -2.96e-19
C11728 avdd.n8854 avss -1.8e-19
C11729 avdd.n8855 avss -1.8e-19
C11730 avdd.n8856 avss 0.00873f
C11731 avdd.n8857 avss 0.0111f
C11732 avdd.n8858 avss 0.0154f
C11733 avdd.n8859 avss 0.0191f
C11734 avdd.n8860 avss -1.8e-19
C11735 avdd.n8861 avss 0.0184f
C11736 avdd.n8862 avss -1.38e-19
C11737 avdd.n8863 avss -1.8e-19
C11738 avdd.n8864 avss -2.44e-19
C11739 avdd.n8865 avss -2.44e-19
C11740 avdd.n8866 avss -1.8e-19
C11741 avdd.n8867 avss -1.38e-19
C11742 avdd.n8868 avss -3.49e-19
C11743 avdd.n8870 avss 0.0269f
C11744 avdd.n8871 avss 0.00869f
C11745 avdd.n8872 avss 0.00378f
C11746 avdd.n8873 avss 0.0346f
C11747 avdd.n8874 avss -8.47e-19
C11748 avdd.n8875 avss -3.39e-19
C11749 avdd.n8876 avss -8.47e-19
C11750 avdd.n8877 avss 3e-19
C11751 avdd.n8878 avss 0.0388f
C11752 avdd.n8879 avss -3.39e-19
C11753 avdd.n8880 avss -6.46e-19
C11754 avdd.n8881 avss -5.82e-19
C11755 avdd.n8882 avss -3.39e-19
C11756 avdd.n8883 avss -8.47e-19
C11757 avdd.n8884 avss -0.00113f
C11758 avdd.n8885 avss -0.00512f
C11759 avdd.n8886 avss 0.0382f
C11760 avdd.n8887 avss -0.152f
C11761 avdd.n8888 avss -0.229f
C11762 avdd.n8889 avss -8.47e-19
C11763 avdd.n8890 avss -3.28e-19
C11764 avdd.n8891 avss -3.28e-19
C11765 avdd.n8892 avss -8.26e-19
C11766 avdd.n8893 avss 0.0348f
C11767 avdd.n8894 avss 0.00357f
C11768 avdd.n8895 avss -8.47e-19
C11769 avdd.n8896 avss -3.39e-19
C11770 avdd.n8897 avss -8.47e-19
C11771 avdd.n8898 avss 0.0344f
C11772 avdd.n8899 avss 0.00466f
C11773 avdd.n8900 avss -3.39e-19
C11774 avdd.n8901 avss -6.67e-19
C11775 avdd.n8902 avss -5.61e-19
C11776 avdd.n8903 avss -0.00137f
C11777 avdd.n8904 avss -0.0013f
C11778 avdd.n8905 avss -5.19e-19
C11779 avdd.n8906 avss 0.0386f
C11780 avdd.n8907 avss 0.0111f
C11781 avdd.n8908 avss 0.0148f
C11782 avdd.n8909 avss 0.019f
C11783 avdd.n8910 avss -1.8e-19
C11784 avdd.n8911 avss 0.0184f
C11785 avdd.n8912 avss -2.44e-19
C11786 avdd.n8913 avss -2.33e-19
C11787 avdd.n8914 avss 0.0022f
C11788 avdd.n8915 avss -1.48e-19
C11789 avdd.n8916 avss -1.27e-19
C11790 avdd.n8917 avss -2.44e-19
C11791 avdd.n8918 avss -8.15e-19
C11792 avdd.n8919 avss -0.0014f
C11793 avdd.n8920 avss -8.47e-19
C11794 avdd.n8921 avss -3.39e-19
C11795 avdd.n8922 avss -3.49e-19
C11796 avdd.n8923 avss -1.38e-19
C11797 avdd.n8924 avss -1.8e-19
C11798 avdd.n8925 avss 0.00873f
C11799 avdd.n8926 avss 0.0111f
C11800 avdd.n8927 avss 0.0154f
C11801 avdd.n8928 avss 0.0191f
C11802 avdd.n8929 avss -1.8e-19
C11803 avdd.n8930 avss 0.0184f
C11804 avdd.n8931 avss -1.38e-19
C11805 avdd.n8932 avss -1.8e-19
C11806 avdd.n8933 avss -2.44e-19
C11807 avdd.n8934 avss 0.0411f
C11808 avdd.n8935 avss -1.8e-19
C11809 avdd.n8936 avss -1.8e-19
C11810 avdd.n8937 avss -2.96e-19
C11811 avdd.n8938 avss -3.39e-19
C11812 avdd.n8939 avss -6.35e-19
C11813 avdd.n8940 avss 0.0098f
C11814 avdd.n8941 avss -0.00139f
C11815 avdd.n8942 avss -6.88e-19
C11816 avdd.n8943 avss -3.07e-19
C11817 avdd.n8944 avss -1.8e-19
C11818 avdd.n8945 avss 0.0112f
C11819 avdd.n8946 avss -2.75e-19
C11820 avdd.n8947 avss 0.00821f
C11821 avdd.n8948 avss 0.00821f
C11822 avdd.n8949 avss -2.75e-19
C11823 avdd.n8950 avss 0.0442f
C11824 avdd.n8951 avss 0.0179f
C11825 avdd.n8952 avss -2.22e-19
C11826 avdd.n8953 avss -1.59e-19
C11827 avdd.n8954 avss -2.33e-19
C11828 avdd.n8955 avss 0.0188f
C11829 avdd.n8956 avss 0.0181f
C11830 avdd.n8957 avss -2.75e-19
C11831 avdd.n8958 avss -3.39e-19
C11832 avdd.n8959 avss -3.6e-19
C11833 avdd.n8960 avss -2.01e-19
C11834 avdd.n8961 avss -0.0866f
C11835 avdd.n8962 avss -0.00336f
C11836 avdd.n8963 avss 0.00725f
C11837 avdd.n8964 avss 0.0318f
C11838 avdd.n8965 avss -0.00158f
C11839 avdd.n8966 avss -8.47e-19
C11840 avdd.n8967 avss 0.0298f
C11841 avdd.n8968 avss -2.22e-19
C11842 avdd.n8969 avss 0.0148f
C11843 avdd.n8970 avss 0.0182f
C11844 avdd.n8971 avss -1.8e-19
C11845 avdd.n8972 avss -2.54e-19
C11846 avdd.n8973 avss -2.54e-19
C11847 avdd.n8974 avss -1.8e-19
C11848 avdd.n8975 avss -1.16e-19
C11849 avdd.n8976 avss -0.00126f
C11850 avdd.n8977 avss -2.33e-19
C11851 avdd.n8978 avss -3.39e-19
C11852 avdd.n8979 avss -4.23e-19
C11853 avdd.n8980 avss 0.00358f
C11854 avdd.n8981 avss 0.0374f
C11855 avdd.n8982 avss -3.07e-19
C11856 avdd.n8983 avss -0.00108f
C11857 avdd.n8984 avss -0.00109f
C11858 avdd.n8985 avss 0.0192f
C11859 avdd.n8986 avss -1.59e-19
C11860 avdd.n8987 avss -1.8e-19
C11861 avdd.n8988 avss 0.00875f
C11862 avdd.n8989 avss 0.0111f
C11863 avdd.n8990 avss 0.0154f
C11864 avdd.n8991 avss 0.0183f
C11865 avdd.n8992 avss -1.8e-19
C11866 avdd.n8993 avss -2.22e-19
C11867 avdd.n8994 avss -2.22e-19
C11868 avdd.n8995 avss -1.8e-19
C11869 avdd.n8996 avss -2.01e-19
C11870 avdd.n8997 avss -9.76e-19
C11871 avdd.n8998 avss -0.00121f
C11872 avdd.n8999 avss -0.00122f
C11873 avdd.n9000 avss -0.00173f
C11874 avdd.n9001 avss -0.00357f
C11875 avdd.n9002 avss 0.0382f
C11876 avdd.n9003 avss -8.47e-19
C11877 avdd.n9004 avss -3.28e-19
C11878 avdd.n9005 avss -3.28e-19
C11879 avdd.n9006 avss -8.26e-19
C11880 avdd.n9007 avss 0.0348f
C11881 avdd.n9008 avss 0.00357f
C11882 avdd.n9009 avss -8.47e-19
C11883 avdd.n9010 avss -3.39e-19
C11884 avdd.n9011 avss -8.47e-19
C11885 avdd.n9012 avss 0.0344f
C11886 avdd.n9013 avss 0.00466f
C11887 avdd.n9014 avss -3.39e-19
C11888 avdd.n9015 avss -6.67e-19
C11889 avdd.n9016 avss -5.61e-19
C11890 avdd.n9017 avss -0.00137f
C11891 avdd.n9018 avss -0.0013f
C11892 avdd.n9019 avss -5.19e-19
C11893 avdd.n9020 avss 0.0386f
C11894 avdd.n9021 avss 0.0111f
C11895 avdd.n9022 avss 0.0148f
C11896 avdd.n9023 avss 0.019f
C11897 avdd.n9024 avss -1.8e-19
C11898 avdd.n9025 avss 0.0184f
C11899 avdd.n9026 avss -2.44e-19
C11900 avdd.n9027 avss -2.33e-19
C11901 avdd.n9028 avss 0.0022f
C11902 avdd.n9029 avss -1.48e-19
C11903 avdd.n9030 avss -1.27e-19
C11904 avdd.n9031 avss -2.44e-19
C11905 avdd.n9032 avss -8.15e-19
C11906 avdd.n9033 avss -0.0014f
C11907 avdd.n9034 avss -8.47e-19
C11908 avdd.n9035 avss -3.39e-19
C11909 avdd.n9036 avss -3.49e-19
C11910 avdd.n9037 avss -1.38e-19
C11911 avdd.n9038 avss -1.8e-19
C11912 avdd.n9039 avss 0.00873f
C11913 avdd.n9040 avss 0.0111f
C11914 avdd.n9041 avss 0.0154f
C11915 avdd.n9042 avss 0.0191f
C11916 avdd.n9043 avss -1.8e-19
C11917 avdd.n9044 avss 0.0184f
C11918 avdd.n9045 avss -1.38e-19
C11919 avdd.n9046 avss -1.8e-19
C11920 avdd.n9047 avss -2.44e-19
C11921 avdd.n9048 avss 0.0411f
C11922 avdd.n9049 avss -1.8e-19
C11923 avdd.n9050 avss -1.8e-19
C11924 avdd.n9051 avss -2.96e-19
C11925 avdd.n9052 avss -3.39e-19
C11926 avdd.n9053 avss -6.35e-19
C11927 avdd.n9054 avss 0.0098f
C11928 avdd.n9055 avss -0.00139f
C11929 avdd.n9056 avss -6.88e-19
C11930 avdd.n9057 avss -3.07e-19
C11931 avdd.n9058 avss -1.8e-19
C11932 avdd.n9059 avss 0.0112f
C11933 avdd.n9060 avss -2.75e-19
C11934 avdd.n9061 avss 0.00821f
C11935 avdd.n9062 avss 0.00821f
C11936 avdd.n9063 avss -2.75e-19
C11937 avdd.n9064 avss 0.0442f
C11938 avdd.n9065 avss 0.0179f
C11939 avdd.n9066 avss -2.22e-19
C11940 avdd.n9067 avss -1.59e-19
C11941 avdd.n9068 avss -2.33e-19
C11942 avdd.n9069 avss 0.0188f
C11943 avdd.n9070 avss 0.0181f
C11944 avdd.n9071 avss -2.75e-19
C11945 avdd.n9072 avss -3.39e-19
C11946 avdd.n9073 avss -3.6e-19
C11947 avdd.n9074 avss -2.01e-19
C11948 avdd.n9075 avss -0.0866f
C11949 avdd.n9076 avss -0.00336f
C11950 avdd.n9077 avss 0.00725f
C11951 avdd.n9078 avss 0.0318f
C11952 avdd.n9079 avss -0.00158f
C11953 avdd.n9080 avss -8.47e-19
C11954 avdd.n9081 avss 0.0298f
C11955 avdd.n9082 avss -2.22e-19
C11956 avdd.n9083 avss 0.0148f
C11957 avdd.n9084 avss 0.0182f
C11958 avdd.n9085 avss -1.8e-19
C11959 avdd.n9086 avss -2.54e-19
C11960 avdd.n9087 avss -2.54e-19
C11961 avdd.n9088 avss -1.8e-19
C11962 avdd.n9089 avss -1.16e-19
C11963 avdd.n9090 avss -0.00126f
C11964 avdd.n9091 avss -2.33e-19
C11965 avdd.n9092 avss -3.39e-19
C11966 avdd.n9093 avss -4.23e-19
C11967 avdd.n9094 avss 0.00358f
C11968 avdd.n9095 avss 0.0374f
C11969 avdd.n9096 avss -3.07e-19
C11970 avdd.n9097 avss -0.00108f
C11971 avdd.n9098 avss -0.00109f
C11972 avdd.n9099 avss 0.0192f
C11973 avdd.n9100 avss -1.59e-19
C11974 avdd.n9101 avss -1.8e-19
C11975 avdd.n9102 avss 0.00875f
C11976 avdd.n9103 avss 0.0111f
C11977 avdd.n9104 avss 0.0154f
C11978 avdd.n9105 avss 0.0183f
C11979 avdd.n9106 avss -1.8e-19
C11980 avdd.n9107 avss -2.22e-19
C11981 avdd.n9108 avss -2.22e-19
C11982 avdd.n9109 avss -1.8e-19
C11983 avdd.n9110 avss -2.01e-19
C11984 avdd.n9111 avss -9.76e-19
C11985 avdd.n9112 avss -0.00121f
C11986 avdd.n9113 avss -0.00122f
C11987 avdd.n9114 avss -0.00173f
C11988 avdd.n9115 avss -0.00357f
C11989 avdd.n9116 avss 0.0382f
C11990 avdd.n9117 avss -8.47e-19
C11991 avdd.n9118 avss -3.28e-19
C11992 avdd.n9119 avss -3.28e-19
C11993 avdd.n9120 avss -8.26e-19
C11994 avdd.n9121 avss 0.0348f
C11995 avdd.n9122 avss 0.00357f
C11996 avdd.n9123 avss -8.47e-19
C11997 avdd.n9124 avss -3.39e-19
C11998 avdd.n9125 avss -8.47e-19
C11999 avdd.n9126 avss 0.0344f
C12000 avdd.n9127 avss 0.00466f
C12001 avdd.n9128 avss -3.39e-19
C12002 avdd.n9129 avss -6.67e-19
C12003 avdd.n9130 avss -5.61e-19
C12004 avdd.n9131 avss -0.00137f
C12005 avdd.n9132 avss -0.0013f
C12006 avdd.n9133 avss -5.19e-19
C12007 avdd.n9134 avss 0.0386f
C12008 avdd.n9135 avss 0.0111f
C12009 avdd.n9136 avss 0.0148f
C12010 avdd.n9137 avss 0.019f
C12011 avdd.n9138 avss -1.8e-19
C12012 avdd.n9139 avss 0.0184f
C12013 avdd.n9140 avss -2.44e-19
C12014 avdd.n9141 avss -2.33e-19
C12015 avdd.n9142 avss 0.0022f
C12016 avdd.n9143 avss -1.48e-19
C12017 avdd.n9144 avss -1.27e-19
C12018 avdd.n9145 avss -2.44e-19
C12019 avdd.n9146 avss -8.15e-19
C12020 avdd.n9147 avss -0.0014f
C12021 avdd.n9148 avss -8.47e-19
C12022 avdd.n9149 avss -3.39e-19
C12023 avdd.n9150 avss -3.49e-19
C12024 avdd.n9151 avss -1.38e-19
C12025 avdd.n9152 avss -1.8e-19
C12026 avdd.n9153 avss 0.00873f
C12027 avdd.n9154 avss 0.0111f
C12028 avdd.n9155 avss 0.0154f
C12029 avdd.n9156 avss 0.0191f
C12030 avdd.n9157 avss -1.8e-19
C12031 avdd.n9158 avss 0.0184f
C12032 avdd.n9159 avss -1.38e-19
C12033 avdd.n9160 avss -1.8e-19
C12034 avdd.n9161 avss -2.44e-19
C12035 avdd.n9162 avss 0.0411f
C12036 avdd.n9163 avss -1.8e-19
C12037 avdd.n9164 avss -1.8e-19
C12038 avdd.n9165 avss -2.96e-19
C12039 avdd.n9166 avss -3.39e-19
C12040 avdd.n9167 avss -6.35e-19
C12041 avdd.n9168 avss 0.0098f
C12042 avdd.n9169 avss -0.00139f
C12043 avdd.n9170 avss -6.88e-19
C12044 avdd.n9171 avss -3.07e-19
C12045 avdd.n9172 avss -1.8e-19
C12046 avdd.n9173 avss 0.0112f
C12047 avdd.n9174 avss -2.75e-19
C12048 avdd.n9175 avss 0.00821f
C12049 avdd.n9176 avss 0.00821f
C12050 avdd.n9177 avss -2.75e-19
C12051 avdd.n9178 avss 0.0442f
C12052 avdd.n9179 avss 0.0179f
C12053 avdd.n9180 avss -2.22e-19
C12054 avdd.n9181 avss -1.59e-19
C12055 avdd.n9182 avss -2.33e-19
C12056 avdd.n9183 avss 0.0188f
C12057 avdd.n9184 avss 0.0181f
C12058 avdd.n9185 avss -2.75e-19
C12059 avdd.n9186 avss -3.39e-19
C12060 avdd.n9187 avss -3.6e-19
C12061 avdd.n9188 avss -2.01e-19
C12062 avdd.n9189 avss -0.0866f
C12063 avdd.n9190 avss -0.00336f
C12064 avdd.n9191 avss 0.00725f
C12065 avdd.n9192 avss 0.0318f
C12066 avdd.n9193 avss -0.00158f
C12067 avdd.n9194 avss -8.47e-19
C12068 avdd.n9195 avss 0.0298f
C12069 avdd.n9196 avss -2.22e-19
C12070 avdd.n9197 avss 0.0148f
C12071 avdd.n9198 avss 0.0182f
C12072 avdd.n9199 avss -1.8e-19
C12073 avdd.n9200 avss -2.54e-19
C12074 avdd.n9201 avss -2.54e-19
C12075 avdd.n9202 avss -1.8e-19
C12076 avdd.n9203 avss -1.16e-19
C12077 avdd.n9204 avss -0.00126f
C12078 avdd.n9205 avss -2.33e-19
C12079 avdd.n9206 avss -3.39e-19
C12080 avdd.n9207 avss -4.23e-19
C12081 avdd.n9208 avss 0.00358f
C12082 avdd.n9209 avss 0.0374f
C12083 avdd.n9210 avss -3.07e-19
C12084 avdd.n9211 avss -0.00108f
C12085 avdd.n9212 avss -0.00109f
C12086 avdd.n9213 avss 0.0192f
C12087 avdd.n9214 avss -1.59e-19
C12088 avdd.n9215 avss -1.8e-19
C12089 avdd.n9216 avss 0.00875f
C12090 avdd.n9217 avss 0.0111f
C12091 avdd.n9218 avss 0.0154f
C12092 avdd.n9219 avss 0.0183f
C12093 avdd.n9220 avss -1.8e-19
C12094 avdd.n9221 avss -2.22e-19
C12095 avdd.n9222 avss -2.22e-19
C12096 avdd.n9223 avss -1.8e-19
C12097 avdd.n9224 avss -2.01e-19
C12098 avdd.n9225 avss -9.76e-19
C12099 avdd.n9226 avss -0.00121f
C12100 avdd.n9227 avss -0.00122f
C12101 avdd.n9228 avss -0.00173f
C12102 avdd.n9229 avss -0.00357f
C12103 avdd.n9230 avss 0.0382f
C12104 avdd.n9231 avss -8.47e-19
C12105 avdd.n9232 avss -3.28e-19
C12106 avdd.n9233 avss -3.28e-19
C12107 avdd.n9234 avss -8.26e-19
C12108 avdd.n9235 avss 0.0348f
C12109 avdd.n9236 avss 0.00357f
C12110 avdd.n9237 avss -8.47e-19
C12111 avdd.n9238 avss -3.39e-19
C12112 avdd.n9239 avss -8.47e-19
C12113 avdd.n9240 avss 0.0344f
C12114 avdd.n9241 avss 0.00466f
C12115 avdd.n9242 avss -3.39e-19
C12116 avdd.n9243 avss -6.67e-19
C12117 avdd.n9244 avss -5.61e-19
C12118 avdd.n9245 avss -0.00137f
C12119 avdd.n9246 avss -0.0013f
C12120 avdd.n9247 avss -5.19e-19
C12121 avdd.n9248 avss 0.0386f
C12122 avdd.n9249 avss 0.0111f
C12123 avdd.n9250 avss 0.0148f
C12124 avdd.n9251 avss 0.019f
C12125 avdd.n9252 avss -1.8e-19
C12126 avdd.n9253 avss 0.0184f
C12127 avdd.n9254 avss -2.44e-19
C12128 avdd.n9255 avss -2.33e-19
C12129 avdd.n9256 avss 0.0022f
C12130 avdd.n9257 avss -1.48e-19
C12131 avdd.n9258 avss -1.27e-19
C12132 avdd.n9259 avss -2.44e-19
C12133 avdd.n9260 avss -8.15e-19
C12134 avdd.n9261 avss -0.0014f
C12135 avdd.n9262 avss -8.47e-19
C12136 avdd.n9263 avss -3.39e-19
C12137 avdd.n9264 avss -3.49e-19
C12138 avdd.n9265 avss -1.38e-19
C12139 avdd.n9266 avss -1.8e-19
C12140 avdd.n9267 avss 0.00873f
C12141 avdd.n9268 avss 0.0111f
C12142 avdd.n9269 avss 0.0154f
C12143 avdd.n9270 avss 0.0191f
C12144 avdd.n9271 avss -1.8e-19
C12145 avdd.n9272 avss 0.0184f
C12146 avdd.n9273 avss -1.38e-19
C12147 avdd.n9274 avss -1.8e-19
C12148 avdd.n9275 avss -2.44e-19
C12149 avdd.n9276 avss 0.0411f
C12150 avdd.n9277 avss -1.8e-19
C12151 avdd.n9278 avss -1.8e-19
C12152 avdd.n9279 avss -2.96e-19
C12153 avdd.n9280 avss -3.39e-19
C12154 avdd.n9281 avss -6.35e-19
C12155 avdd.n9282 avss 0.0098f
C12156 avdd.n9283 avss -0.00139f
C12157 avdd.n9284 avss -6.88e-19
C12158 avdd.n9285 avss -3.07e-19
C12159 avdd.n9286 avss -1.8e-19
C12160 avdd.n9287 avss 0.0112f
C12161 avdd.n9288 avss -2.75e-19
C12162 avdd.n9289 avss 0.00821f
C12163 avdd.n9290 avss 0.00821f
C12164 avdd.n9291 avss -2.75e-19
C12165 avdd.n9292 avss 0.0442f
C12166 avdd.n9293 avss 0.0179f
C12167 avdd.n9294 avss -2.22e-19
C12168 avdd.n9295 avss -1.59e-19
C12169 avdd.n9296 avss -2.33e-19
C12170 avdd.n9297 avss 0.0188f
C12171 avdd.n9298 avss 0.0181f
C12172 avdd.n9299 avss -2.75e-19
C12173 avdd.n9300 avss -3.39e-19
C12174 avdd.n9301 avss -3.6e-19
C12175 avdd.n9302 avss -2.01e-19
C12176 avdd.n9303 avss -0.0866f
C12177 avdd.n9304 avss -0.00336f
C12178 avdd.n9305 avss 0.00725f
C12179 avdd.n9306 avss 0.0318f
C12180 avdd.n9307 avss -0.00158f
C12181 avdd.n9308 avss -8.47e-19
C12182 avdd.n9309 avss 0.0298f
C12183 avdd.n9310 avss -2.22e-19
C12184 avdd.n9311 avss 0.0148f
C12185 avdd.n9312 avss 0.0182f
C12186 avdd.n9313 avss -1.8e-19
C12187 avdd.n9314 avss -2.54e-19
C12188 avdd.n9315 avss -2.54e-19
C12189 avdd.n9316 avss -1.8e-19
C12190 avdd.n9317 avss -1.16e-19
C12191 avdd.n9318 avss -0.00126f
C12192 avdd.n9319 avss -2.33e-19
C12193 avdd.n9320 avss -3.39e-19
C12194 avdd.n9321 avss -4.23e-19
C12195 avdd.n9322 avss 0.00358f
C12196 avdd.n9323 avss 0.0374f
C12197 avdd.n9324 avss -3.07e-19
C12198 avdd.n9325 avss -0.00108f
C12199 avdd.n9326 avss -0.00109f
C12200 avdd.n9327 avss 0.0192f
C12201 avdd.n9328 avss -1.59e-19
C12202 avdd.n9329 avss -1.8e-19
C12203 avdd.n9330 avss 0.00875f
C12204 avdd.n9331 avss 0.0111f
C12205 avdd.n9332 avss 0.0154f
C12206 avdd.n9333 avss 0.0183f
C12207 avdd.n9334 avss -1.8e-19
C12208 avdd.n9335 avss -2.22e-19
C12209 avdd.n9336 avss -2.22e-19
C12210 avdd.n9337 avss -1.8e-19
C12211 avdd.n9338 avss -2.01e-19
C12212 avdd.n9339 avss -9.76e-19
C12213 avdd.n9340 avss -0.00121f
C12214 avdd.n9341 avss -0.00122f
C12215 avdd.n9342 avss -0.00173f
C12216 avdd.n9343 avss -0.00357f
C12217 avdd.n9344 avss 0.0382f
C12218 avdd.n9345 avss -8.47e-19
C12219 avdd.n9346 avss -3.28e-19
C12220 avdd.n9347 avss -3.28e-19
C12221 avdd.n9348 avss -8.26e-19
C12222 avdd.n9349 avss 0.0348f
C12223 avdd.n9350 avss 0.00357f
C12224 avdd.n9351 avss -8.47e-19
C12225 avdd.n9352 avss -3.39e-19
C12226 avdd.n9353 avss -8.47e-19
C12227 avdd.n9354 avss 0.0344f
C12228 avdd.n9355 avss 0.00466f
C12229 avdd.n9356 avss -3.39e-19
C12230 avdd.n9357 avss -6.67e-19
C12231 avdd.n9358 avss -5.61e-19
C12232 avdd.n9359 avss -0.00137f
C12233 avdd.n9360 avss -0.0013f
C12234 avdd.n9361 avss -5.19e-19
C12235 avdd.n9362 avss 0.0386f
C12236 avdd.n9363 avss 0.0111f
C12237 avdd.n9364 avss 0.0148f
C12238 avdd.n9365 avss 0.019f
C12239 avdd.n9366 avss -1.8e-19
C12240 avdd.n9367 avss 0.0184f
C12241 avdd.n9368 avss -2.44e-19
C12242 avdd.n9369 avss -2.33e-19
C12243 avdd.n9370 avss 0.0022f
C12244 avdd.n9371 avss -1.48e-19
C12245 avdd.n9372 avss -1.27e-19
C12246 avdd.n9373 avss -2.44e-19
C12247 avdd.n9374 avss -8.15e-19
C12248 avdd.n9375 avss -0.0014f
C12249 avdd.n9376 avss -8.47e-19
C12250 avdd.n9377 avss -3.39e-19
C12251 avdd.n9378 avss -3.49e-19
C12252 avdd.n9379 avss -1.38e-19
C12253 avdd.n9380 avss -1.8e-19
C12254 avdd.n9381 avss 0.00873f
C12255 avdd.n9382 avss 0.0111f
C12256 avdd.n9383 avss 0.0154f
C12257 avdd.n9384 avss 0.0191f
C12258 avdd.n9385 avss -1.8e-19
C12259 avdd.n9386 avss 0.0184f
C12260 avdd.n9387 avss -1.38e-19
C12261 avdd.n9388 avss -1.8e-19
C12262 avdd.n9389 avss -2.44e-19
C12263 avdd.n9390 avss 0.0411f
C12264 avdd.n9391 avss -1.8e-19
C12265 avdd.n9392 avss -1.8e-19
C12266 avdd.n9393 avss -2.96e-19
C12267 avdd.n9394 avss -3.39e-19
C12268 avdd.n9395 avss -6.35e-19
C12269 avdd.n9396 avss 0.0098f
C12270 avdd.n9397 avss -0.00139f
C12271 avdd.n9398 avss -6.88e-19
C12272 avdd.n9399 avss -3.07e-19
C12273 avdd.n9400 avss -1.8e-19
C12274 avdd.n9401 avss 0.0112f
C12275 avdd.n9402 avss -2.75e-19
C12276 avdd.n9403 avss 0.00821f
C12277 avdd.n9404 avss 0.00821f
C12278 avdd.n9405 avss -2.75e-19
C12279 avdd.n9406 avss 0.0442f
C12280 avdd.n9407 avss 0.0179f
C12281 avdd.n9408 avss -2.22e-19
C12282 avdd.n9409 avss -1.59e-19
C12283 avdd.n9410 avss -2.33e-19
C12284 avdd.n9411 avss 0.0188f
C12285 avdd.n9412 avss 0.0181f
C12286 avdd.n9413 avss -2.75e-19
C12287 avdd.n9414 avss -3.39e-19
C12288 avdd.n9415 avss -3.6e-19
C12289 avdd.n9416 avss -2.01e-19
C12290 avdd.n9417 avss -0.0866f
C12291 avdd.n9418 avss -0.00336f
C12292 avdd.n9419 avss 0.00725f
C12293 avdd.n9420 avss 0.0318f
C12294 avdd.n9421 avss -0.00158f
C12295 avdd.n9422 avss -8.47e-19
C12296 avdd.n9423 avss 0.0298f
C12297 avdd.n9424 avss -2.22e-19
C12298 avdd.n9425 avss 0.0148f
C12299 avdd.n9426 avss 0.0182f
C12300 avdd.n9427 avss -1.8e-19
C12301 avdd.n9428 avss -2.54e-19
C12302 avdd.n9429 avss -2.54e-19
C12303 avdd.n9430 avss -1.8e-19
C12304 avdd.n9431 avss -1.16e-19
C12305 avdd.n9432 avss -0.00126f
C12306 avdd.n9433 avss -2.33e-19
C12307 avdd.n9434 avss -3.39e-19
C12308 avdd.n9435 avss -4.23e-19
C12309 avdd.n9436 avss 0.00358f
C12310 avdd.n9437 avss 0.0374f
C12311 avdd.n9438 avss -3.07e-19
C12312 avdd.n9439 avss -0.00108f
C12313 avdd.n9440 avss -0.00109f
C12314 avdd.n9441 avss 0.0192f
C12315 avdd.n9442 avss -1.59e-19
C12316 avdd.n9443 avss -1.8e-19
C12317 avdd.n9444 avss 0.00875f
C12318 avdd.n9445 avss 0.0111f
C12319 avdd.n9446 avss 0.0154f
C12320 avdd.n9447 avss 0.0183f
C12321 avdd.n9448 avss -1.8e-19
C12322 avdd.n9449 avss -2.22e-19
C12323 avdd.n9450 avss -2.22e-19
C12324 avdd.n9451 avss -1.8e-19
C12325 avdd.n9452 avss -2.01e-19
C12326 avdd.n9453 avss -9.76e-19
C12327 avdd.n9454 avss -0.00121f
C12328 avdd.n9455 avss -0.00122f
C12329 avdd.n9456 avss -0.00173f
C12330 avdd.n9457 avss -0.00357f
C12331 avdd.n9458 avss 0.0382f
C12332 avdd.n9459 avss -8.47e-19
C12333 avdd.n9460 avss -3.28e-19
C12334 avdd.n9461 avss -3.28e-19
C12335 avdd.n9462 avss -8.26e-19
C12336 avdd.n9463 avss 0.0348f
C12337 avdd.n9464 avss 0.00357f
C12338 avdd.n9465 avss -8.47e-19
C12339 avdd.n9466 avss -3.39e-19
C12340 avdd.n9467 avss -8.47e-19
C12341 avdd.n9468 avss 0.0344f
C12342 avdd.n9469 avss 0.00466f
C12343 avdd.n9470 avss -3.39e-19
C12344 avdd.n9471 avss -6.67e-19
C12345 avdd.n9472 avss -5.61e-19
C12346 avdd.n9473 avss -0.00137f
C12347 avdd.n9474 avss -0.0013f
C12348 avdd.n9475 avss -5.19e-19
C12349 avdd.n9476 avss 0.0386f
C12350 avdd.n9477 avss 0.0111f
C12351 avdd.n9478 avss 0.0148f
C12352 avdd.n9479 avss 0.019f
C12353 avdd.n9480 avss -1.8e-19
C12354 avdd.n9481 avss 0.0184f
C12355 avdd.n9482 avss -2.44e-19
C12356 avdd.n9483 avss -2.33e-19
C12357 avdd.n9484 avss 0.0022f
C12358 avdd.n9485 avss -1.48e-19
C12359 avdd.n9486 avss -1.27e-19
C12360 avdd.n9487 avss -2.44e-19
C12361 avdd.n9488 avss -8.15e-19
C12362 avdd.n9489 avss -0.0014f
C12363 avdd.n9490 avss -8.47e-19
C12364 avdd.n9491 avss -3.39e-19
C12365 avdd.n9492 avss -3.49e-19
C12366 avdd.n9493 avss -1.38e-19
C12367 avdd.n9494 avss -1.8e-19
C12368 avdd.n9495 avss 0.00873f
C12369 avdd.n9496 avss 0.0111f
C12370 avdd.n9497 avss 0.0154f
C12371 avdd.n9498 avss 0.0191f
C12372 avdd.n9499 avss -1.8e-19
C12373 avdd.n9500 avss 0.0184f
C12374 avdd.n9501 avss -1.38e-19
C12375 avdd.n9502 avss -1.8e-19
C12376 avdd.n9503 avss -2.44e-19
C12377 avdd.n9504 avss 0.0411f
C12378 avdd.n9505 avss -1.8e-19
C12379 avdd.n9506 avss -1.8e-19
C12380 avdd.n9507 avss -2.96e-19
C12381 avdd.n9508 avss -3.39e-19
C12382 avdd.n9509 avss -6.35e-19
C12383 avdd.n9510 avss 0.0098f
C12384 avdd.n9511 avss -0.00139f
C12385 avdd.n9512 avss -6.88e-19
C12386 avdd.n9513 avss -3.07e-19
C12387 avdd.n9514 avss -1.8e-19
C12388 avdd.n9515 avss 0.0112f
C12389 avdd.n9516 avss -2.75e-19
C12390 avdd.n9517 avss 0.00821f
C12391 avdd.n9518 avss 0.00821f
C12392 avdd.n9519 avss -2.75e-19
C12393 avdd.n9520 avss 0.0442f
C12394 avdd.n9521 avss 0.0179f
C12395 avdd.n9522 avss -2.22e-19
C12396 avdd.n9523 avss -1.59e-19
C12397 avdd.n9524 avss -2.33e-19
C12398 avdd.n9525 avss 0.0188f
C12399 avdd.n9526 avss 0.0181f
C12400 avdd.n9527 avss -2.75e-19
C12401 avdd.n9528 avss -3.39e-19
C12402 avdd.n9529 avss -3.6e-19
C12403 avdd.n9530 avss -2.01e-19
C12404 avdd.n9531 avss -0.0866f
C12405 avdd.n9532 avss -0.00336f
C12406 avdd.n9533 avss 0.00725f
C12407 avdd.n9534 avss 0.0318f
C12408 avdd.n9535 avss -0.00158f
C12409 avdd.n9536 avss -8.47e-19
C12410 avdd.n9537 avss 0.0298f
C12411 avdd.n9538 avss -2.22e-19
C12412 avdd.n9539 avss 0.0148f
C12413 avdd.n9540 avss 0.0182f
C12414 avdd.n9541 avss -1.8e-19
C12415 avdd.n9542 avss -2.54e-19
C12416 avdd.n9543 avss -2.54e-19
C12417 avdd.n9544 avss -1.8e-19
C12418 avdd.n9545 avss -1.16e-19
C12419 avdd.n9546 avss -0.00126f
C12420 avdd.n9547 avss -2.33e-19
C12421 avdd.n9548 avss -3.39e-19
C12422 avdd.n9549 avss -4.23e-19
C12423 avdd.n9550 avss 0.00358f
C12424 avdd.n9551 avss 0.0374f
C12425 avdd.n9552 avss -3.07e-19
C12426 avdd.n9553 avss -0.00108f
C12427 avdd.n9554 avss -0.00109f
C12428 avdd.n9555 avss 0.0192f
C12429 avdd.n9556 avss -1.59e-19
C12430 avdd.n9557 avss -1.8e-19
C12431 avdd.n9558 avss 0.00875f
C12432 avdd.n9559 avss 0.0111f
C12433 avdd.n9560 avss 0.0154f
C12434 avdd.n9561 avss 0.0183f
C12435 avdd.n9562 avss -1.8e-19
C12436 avdd.n9563 avss -2.22e-19
C12437 avdd.n9564 avss -2.22e-19
C12438 avdd.n9565 avss -1.8e-19
C12439 avdd.n9566 avss -2.01e-19
C12440 avdd.n9567 avss -9.76e-19
C12441 avdd.n9568 avss -0.00121f
C12442 avdd.n9569 avss -0.00122f
C12443 avdd.n9570 avss -0.00173f
C12444 avdd.n9571 avss -0.00357f
C12445 avdd.n9572 avss 0.0382f
C12446 avdd.n9573 avss -8.47e-19
C12447 avdd.n9574 avss -3.28e-19
C12448 avdd.n9575 avss -3.28e-19
C12449 avdd.n9576 avss -8.26e-19
C12450 avdd.n9577 avss 0.0348f
C12451 avdd.n9578 avss 0.00357f
C12452 avdd.n9579 avss -8.47e-19
C12453 avdd.n9580 avss -3.39e-19
C12454 avdd.n9581 avss -8.47e-19
C12455 avdd.n9582 avss 0.0344f
C12456 avdd.n9583 avss 0.00466f
C12457 avdd.n9584 avss -3.39e-19
C12458 avdd.n9585 avss -6.67e-19
C12459 avdd.n9586 avss -5.61e-19
C12460 avdd.n9587 avss -0.00121f
C12461 avdd.n9588 avss -0.00137f
C12462 avdd.n9589 avss -0.0013f
C12463 avdd.n9590 avss -5.19e-19
C12464 avdd.n9591 avss 0.0386f
C12465 avdd.n9592 avss 0.0111f
C12466 avdd.n9593 avss 0.0148f
C12467 avdd.n9594 avss 0.019f
C12468 avdd.n9595 avss -1.8e-19
C12469 avdd.n9596 avss 0.0184f
C12470 avdd.n9597 avss -2.44e-19
C12471 avdd.n9598 avss -2.33e-19
C12472 avdd.n9599 avss 0.0022f
C12473 avdd.n9600 avss -1.48e-19
C12474 avdd.n9601 avss -1.27e-19
C12475 avdd.n9602 avss -2.44e-19
C12476 avdd.n9603 avss -8.15e-19
C12477 avdd.n9604 avss -0.0014f
C12478 avdd.n9605 avss -8.47e-19
C12479 avdd.n9606 avss -3.39e-19
C12480 avdd.n9607 avss -3.49e-19
C12481 avdd.n9608 avss -1.38e-19
C12482 avdd.n9609 avss -1.8e-19
C12483 avdd.n9610 avss 0.00873f
C12484 avdd.n9611 avss 0.0111f
C12485 avdd.n9612 avss 0.0154f
C12486 avdd.n9613 avss 0.0191f
C12487 avdd.n9614 avss -1.8e-19
C12488 avdd.n9615 avss 0.0184f
C12489 avdd.n9616 avss -1.38e-19
C12490 avdd.n9617 avss -1.8e-19
C12491 avdd.n9618 avss -2.44e-19
C12492 avdd.n9619 avss 0.0411f
C12493 avdd.n9620 avss -1.8e-19
C12494 avdd.n9621 avss -1.8e-19
C12495 avdd.n9622 avss -2.96e-19
C12496 avdd.n9623 avss -3.39e-19
C12497 avdd.n9624 avss -6.35e-19
C12498 avdd.n9625 avss 0.0098f
C12499 avdd.n9626 avss -0.00139f
C12500 avdd.n9627 avss -6.88e-19
C12501 avdd.n9628 avss -3.07e-19
C12502 avdd.n9629 avss -1.8e-19
C12503 avdd.n9630 avss 0.0112f
C12504 avdd.n9631 avss -2.75e-19
C12505 avdd.n9632 avss 0.00821f
C12506 avdd.n9633 avss 0.00821f
C12507 avdd.n9634 avss -2.75e-19
C12508 avdd.n9635 avss 0.0442f
C12509 avdd.n9636 avss 0.0179f
C12510 avdd.n9637 avss -2.22e-19
C12511 avdd.n9638 avss -1.59e-19
C12512 avdd.n9639 avss -2.33e-19
C12513 avdd.n9640 avss 0.0188f
C12514 avdd.n9641 avss 0.0181f
C12515 avdd.n9642 avss -2.75e-19
C12516 avdd.n9643 avss -3.39e-19
C12517 avdd.n9644 avss -3.6e-19
C12518 avdd.n9645 avss -2.01e-19
C12519 avdd.n9646 avss -0.0866f
C12520 avdd.n9647 avss -0.00336f
C12521 avdd.n9648 avss 0.00725f
C12522 avdd.n9649 avss 0.0318f
C12523 avdd.n9650 avss -0.00158f
C12524 avdd.n9651 avss -8.47e-19
C12525 avdd.n9652 avss 0.0298f
C12526 avdd.n9653 avss -2.22e-19
C12527 avdd.n9654 avss 0.0148f
C12528 avdd.n9655 avss 0.0182f
C12529 avdd.n9656 avss -1.8e-19
C12530 avdd.n9657 avss -2.54e-19
C12531 avdd.n9658 avss -2.54e-19
C12532 avdd.n9659 avss -1.8e-19
C12533 avdd.n9660 avss -1.16e-19
C12534 avdd.n9661 avss -0.00126f
C12535 avdd.n9662 avss -2.33e-19
C12536 avdd.n9663 avss -3.39e-19
C12537 avdd.n9664 avss -4.23e-19
C12538 avdd.n9665 avss 0.00358f
C12539 avdd.n9666 avss 0.0374f
C12540 avdd.n9667 avss -3.07e-19
C12541 avdd.n9668 avss -0.00108f
C12542 avdd.n9669 avss -0.00109f
C12543 avdd.n9670 avss 0.0192f
C12544 avdd.n9671 avss -1.59e-19
C12545 avdd.n9672 avss -1.8e-19
C12546 avdd.n9673 avss 0.00875f
C12547 avdd.n9674 avss 0.0111f
C12548 avdd.n9675 avss 0.0154f
C12549 avdd.n9676 avss 0.0183f
C12550 avdd.n9677 avss -1.8e-19
C12551 avdd.n9678 avss -2.22e-19
C12552 avdd.n9679 avss -2.22e-19
C12553 avdd.n9680 avss -1.8e-19
C12554 avdd.n9681 avss -2.01e-19
C12555 avdd.n9682 avss -9.76e-19
C12556 avdd.n9683 avss -0.00122f
C12557 avdd.n9684 avss -0.00173f
C12558 avdd.n9685 avss -0.00357f
C12559 avdd.n9686 avss 0.0382f
C12560 avdd.n9687 avss -8.47e-19
C12561 avdd.n9688 avss -3.28e-19
C12562 avdd.n9689 avss -3.28e-19
C12563 avdd.n9690 avss -8.26e-19
C12564 avdd.n9691 avss 0.0348f
C12565 avdd.n9692 avss 0.00357f
C12566 avdd.n9693 avss -8.47e-19
C12567 avdd.n9694 avss -3.39e-19
C12568 avdd.n9695 avss -8.47e-19
C12569 avdd.n9696 avss 0.0344f
C12570 avdd.n9697 avss 0.00466f
C12571 avdd.n9698 avss -3.39e-19
C12572 avdd.n9699 avss -6.67e-19
C12573 avdd.n9700 avss -5.61e-19
C12574 avdd.n9701 avss -0.00137f
C12575 avdd.n9702 avss -0.0013f
C12576 avdd.n9703 avss -5.19e-19
C12577 avdd.n9704 avss 0.0386f
C12578 avdd.n9705 avss 0.0111f
C12579 avdd.n9706 avss 0.0148f
C12580 avdd.n9707 avss 0.019f
C12581 avdd.n9708 avss -1.8e-19
C12582 avdd.n9709 avss 0.0184f
C12583 avdd.n9710 avss -2.44e-19
C12584 avdd.n9711 avss -2.33e-19
C12585 avdd.n9712 avss 0.0022f
C12586 avdd.n9713 avss -1.48e-19
C12587 avdd.n9714 avss -1.27e-19
C12588 avdd.n9715 avss -2.44e-19
C12589 avdd.n9716 avss -8.15e-19
C12590 avdd.n9717 avss -0.0014f
C12591 avdd.n9718 avss -8.47e-19
C12592 avdd.n9719 avss -3.39e-19
C12593 avdd.n9720 avss -3.49e-19
C12594 avdd.n9721 avss -1.38e-19
C12595 avdd.n9722 avss -1.8e-19
C12596 avdd.n9723 avss 0.00873f
C12597 avdd.n9724 avss 0.0111f
C12598 avdd.n9725 avss 0.0154f
C12599 avdd.n9726 avss 0.0191f
C12600 avdd.n9727 avss -1.8e-19
C12601 avdd.n9728 avss 0.0184f
C12602 avdd.n9729 avss -1.38e-19
C12603 avdd.n9730 avss -1.8e-19
C12604 avdd.n9731 avss -2.44e-19
C12605 avdd.n9732 avss 0.0411f
C12606 avdd.n9733 avss -1.8e-19
C12607 avdd.n9734 avss -1.8e-19
C12608 avdd.n9735 avss -2.96e-19
C12609 avdd.n9736 avss -3.39e-19
C12610 avdd.n9737 avss -6.35e-19
C12611 avdd.n9738 avss 0.0098f
C12612 avdd.n9739 avss -0.00139f
C12613 avdd.n9740 avss -6.88e-19
C12614 avdd.n9741 avss -3.07e-19
C12615 avdd.n9742 avss -1.8e-19
C12616 avdd.n9743 avss 0.0112f
C12617 avdd.n9744 avss -2.75e-19
C12618 avdd.n9745 avss 0.00821f
C12619 avdd.n9746 avss 0.00821f
C12620 avdd.n9747 avss -2.75e-19
C12621 avdd.n9748 avss 0.0442f
C12622 avdd.n9749 avss 0.0179f
C12623 avdd.n9750 avss -2.22e-19
C12624 avdd.n9751 avss -1.59e-19
C12625 avdd.n9752 avss -2.33e-19
C12626 avdd.n9753 avss 0.0188f
C12627 avdd.n9754 avss 0.0181f
C12628 avdd.n9755 avss -2.75e-19
C12629 avdd.n9756 avss -3.39e-19
C12630 avdd.n9757 avss -3.6e-19
C12631 avdd.n9758 avss -2.01e-19
C12632 avdd.n9759 avss -0.0866f
C12633 avdd.n9760 avss -0.00336f
C12634 avdd.n9761 avss 0.00725f
C12635 avdd.n9762 avss 0.0318f
C12636 avdd.n9763 avss -0.00158f
C12637 avdd.n9764 avss -8.47e-19
C12638 avdd.n9765 avss 0.0298f
C12639 avdd.n9766 avss -2.22e-19
C12640 avdd.n9767 avss 0.0148f
C12641 avdd.n9768 avss 0.0182f
C12642 avdd.n9769 avss -1.8e-19
C12643 avdd.n9770 avss -2.54e-19
C12644 avdd.n9771 avss -2.54e-19
C12645 avdd.n9772 avss -1.8e-19
C12646 avdd.n9773 avss -1.16e-19
C12647 avdd.n9774 avss -0.00126f
C12648 avdd.n9775 avss -2.33e-19
C12649 avdd.n9776 avss -3.39e-19
C12650 avdd.n9777 avss -4.23e-19
C12651 avdd.n9778 avss 0.00358f
C12652 avdd.n9779 avss 0.0374f
C12653 avdd.n9780 avss -3.07e-19
C12654 avdd.n9781 avss -0.00108f
C12655 avdd.n9782 avss -0.00109f
C12656 avdd.n9783 avss 0.0192f
C12657 avdd.n9784 avss -1.59e-19
C12658 avdd.n9785 avss -1.8e-19
C12659 avdd.n9786 avss 0.00875f
C12660 avdd.n9787 avss 0.0111f
C12661 avdd.n9788 avss 0.0154f
C12662 avdd.n9789 avss 0.0183f
C12663 avdd.n9790 avss -1.8e-19
C12664 avdd.n9791 avss -2.22e-19
C12665 avdd.n9792 avss -2.22e-19
C12666 avdd.n9793 avss -1.8e-19
C12667 avdd.n9794 avss -2.01e-19
C12668 avdd.n9795 avss -9.76e-19
C12669 avdd.n9796 avss -0.00121f
C12670 avdd.n9797 avss -0.00122f
C12671 avdd.n9798 avss -0.00173f
C12672 avdd.n9799 avss -0.00357f
C12673 avdd.n9800 avss 0.0382f
C12674 avdd.n9801 avss -8.47e-19
C12675 avdd.n9802 avss -3.28e-19
C12676 avdd.n9803 avss -3.28e-19
C12677 avdd.n9804 avss -8.26e-19
C12678 avdd.n9805 avss 0.0348f
C12679 avdd.n9806 avss 0.00357f
C12680 avdd.n9807 avss -8.47e-19
C12681 avdd.n9808 avss -3.39e-19
C12682 avdd.n9809 avss -8.47e-19
C12683 avdd.n9810 avss 0.0344f
C12684 avdd.n9811 avss 0.00466f
C12685 avdd.n9812 avss -3.39e-19
C12686 avdd.n9813 avss -6.67e-19
C12687 avdd.n9814 avss -5.61e-19
C12688 avdd.n9815 avss -0.00137f
C12689 avdd.n9816 avss -0.0013f
C12690 avdd.n9817 avss -5.19e-19
C12691 avdd.n9818 avss 0.0386f
C12692 avdd.n9819 avss 0.0111f
C12693 avdd.n9820 avss 0.0148f
C12694 avdd.n9821 avss 0.019f
C12695 avdd.n9822 avss -1.8e-19
C12696 avdd.n9823 avss 0.0184f
C12697 avdd.n9824 avss -2.44e-19
C12698 avdd.n9825 avss -2.33e-19
C12699 avdd.n9826 avss 0.0022f
C12700 avdd.n9827 avss -1.48e-19
C12701 avdd.n9828 avss -1.27e-19
C12702 avdd.n9829 avss -2.44e-19
C12703 avdd.n9830 avss -8.15e-19
C12704 avdd.n9831 avss -0.0014f
C12705 avdd.n9832 avss -8.47e-19
C12706 avdd.n9833 avss -3.39e-19
C12707 avdd.n9834 avss -3.49e-19
C12708 avdd.n9835 avss -1.38e-19
C12709 avdd.n9836 avss -1.8e-19
C12710 avdd.n9837 avss 0.00873f
C12711 avdd.n9838 avss 0.0111f
C12712 avdd.n9839 avss 0.0154f
C12713 avdd.n9840 avss 0.0191f
C12714 avdd.n9841 avss -1.8e-19
C12715 avdd.n9842 avss 0.0184f
C12716 avdd.n9843 avss -1.38e-19
C12717 avdd.n9844 avss -1.8e-19
C12718 avdd.n9845 avss -2.44e-19
C12719 avdd.n9846 avss 0.0411f
C12720 avdd.n9847 avss -1.8e-19
C12721 avdd.n9848 avss -1.8e-19
C12722 avdd.n9849 avss -2.96e-19
C12723 avdd.n9850 avss -3.39e-19
C12724 avdd.n9851 avss -6.35e-19
C12725 avdd.n9852 avss 0.0098f
C12726 avdd.n9853 avss -0.00139f
C12727 avdd.n9854 avss -6.88e-19
C12728 avdd.n9855 avss -3.07e-19
C12729 avdd.n9856 avss -1.8e-19
C12730 avdd.n9857 avss 0.0112f
C12731 avdd.n9858 avss -2.75e-19
C12732 avdd.n9859 avss 0.00821f
C12733 avdd.n9860 avss 0.00821f
C12734 avdd.n9861 avss -2.75e-19
C12735 avdd.n9862 avss 0.0442f
C12736 avdd.n9863 avss 0.0179f
C12737 avdd.n9864 avss -2.22e-19
C12738 avdd.n9865 avss -1.59e-19
C12739 avdd.n9866 avss -2.33e-19
C12740 avdd.n9867 avss 0.0188f
C12741 avdd.n9868 avss 0.0181f
C12742 avdd.n9869 avss -2.75e-19
C12743 avdd.n9870 avss -3.39e-19
C12744 avdd.n9871 avss -3.6e-19
C12745 avdd.n9872 avss -2.01e-19
C12746 avdd.n9873 avss -0.0866f
C12747 avdd.n9874 avss -0.00336f
C12748 avdd.n9875 avss 0.00725f
C12749 avdd.n9876 avss 0.0318f
C12750 avdd.n9877 avss -0.00158f
C12751 avdd.n9878 avss -8.47e-19
C12752 avdd.n9879 avss 0.0298f
C12753 avdd.n9880 avss -2.22e-19
C12754 avdd.n9881 avss 0.0148f
C12755 avdd.n9882 avss 0.0182f
C12756 avdd.n9883 avss -1.8e-19
C12757 avdd.n9884 avss -2.54e-19
C12758 avdd.n9885 avss -2.54e-19
C12759 avdd.n9886 avss -1.8e-19
C12760 avdd.n9887 avss -1.16e-19
C12761 avdd.n9888 avss -0.00126f
C12762 avdd.n9889 avss -2.33e-19
C12763 avdd.n9890 avss -3.39e-19
C12764 avdd.n9891 avss -4.23e-19
C12765 avdd.n9892 avss 0.00358f
C12766 avdd.n9893 avss 0.0374f
C12767 avdd.n9894 avss -3.07e-19
C12768 avdd.n9895 avss -0.00108f
C12769 avdd.n9896 avss -0.00109f
C12770 avdd.n9897 avss 0.0192f
C12771 avdd.n9898 avss -1.59e-19
C12772 avdd.n9899 avss -1.8e-19
C12773 avdd.n9900 avss 0.00875f
C12774 avdd.n9901 avss 0.0111f
C12775 avdd.n9902 avss 0.0154f
C12776 avdd.n9903 avss 0.0183f
C12777 avdd.n9904 avss -1.8e-19
C12778 avdd.n9905 avss -2.22e-19
C12779 avdd.n9906 avss -2.22e-19
C12780 avdd.n9907 avss -1.8e-19
C12781 avdd.n9908 avss -2.01e-19
C12782 avdd.n9909 avss -9.76e-19
C12783 avdd.n9910 avss -0.00121f
C12784 avdd.n9911 avss -0.00122f
C12785 avdd.n9912 avss -0.00173f
C12786 avdd.n9913 avss -0.00357f
C12787 avdd.n9914 avss 0.0382f
C12788 avdd.n9915 avss -8.47e-19
C12789 avdd.n9916 avss -3.28e-19
C12790 avdd.n9917 avss -3.28e-19
C12791 avdd.n9918 avss -8.26e-19
C12792 avdd.n9919 avss 0.0348f
C12793 avdd.n9920 avss 0.00357f
C12794 avdd.n9921 avss -8.47e-19
C12795 avdd.n9922 avss -3.39e-19
C12796 avdd.n9923 avss -8.47e-19
C12797 avdd.n9924 avss 0.0344f
C12798 avdd.n9925 avss 0.00466f
C12799 avdd.n9926 avss -3.39e-19
C12800 avdd.n9927 avss -6.67e-19
C12801 avdd.n9928 avss -5.61e-19
C12802 avdd.n9929 avss -0.00137f
C12803 avdd.n9930 avss -0.0013f
C12804 avdd.n9931 avss -5.19e-19
C12805 avdd.n9932 avss 0.0386f
C12806 avdd.n9933 avss 0.0111f
C12807 avdd.n9934 avss 0.0148f
C12808 avdd.n9935 avss 0.019f
C12809 avdd.n9936 avss -1.8e-19
C12810 avdd.n9937 avss 0.0184f
C12811 avdd.n9938 avss -2.44e-19
C12812 avdd.n9939 avss -2.33e-19
C12813 avdd.n9940 avss 0.0022f
C12814 avdd.n9941 avss -1.48e-19
C12815 avdd.n9942 avss -1.27e-19
C12816 avdd.n9943 avss -2.44e-19
C12817 avdd.n9944 avss -8.15e-19
C12818 avdd.n9945 avss -0.0014f
C12819 avdd.n9946 avss -8.47e-19
C12820 avdd.n9947 avss -3.39e-19
C12821 avdd.n9948 avss -3.49e-19
C12822 avdd.n9949 avss -1.38e-19
C12823 avdd.n9950 avss -1.8e-19
C12824 avdd.n9951 avss 0.00873f
C12825 avdd.n9952 avss 0.0111f
C12826 avdd.n9953 avss 0.0154f
C12827 avdd.n9954 avss 0.0191f
C12828 avdd.n9955 avss -1.8e-19
C12829 avdd.n9956 avss 0.0184f
C12830 avdd.n9957 avss -1.38e-19
C12831 avdd.n9958 avss -1.8e-19
C12832 avdd.n9959 avss -2.44e-19
C12833 avdd.n9960 avss 0.0411f
C12834 avdd.n9961 avss -1.8e-19
C12835 avdd.n9962 avss -1.8e-19
C12836 avdd.n9963 avss -2.96e-19
C12837 avdd.n9964 avss -3.39e-19
C12838 avdd.n9965 avss -6.35e-19
C12839 avdd.n9966 avss 0.0098f
C12840 avdd.n9967 avss -0.00139f
C12841 avdd.n9968 avss -6.88e-19
C12842 avdd.n9969 avss -3.07e-19
C12843 avdd.n9970 avss -1.8e-19
C12844 avdd.n9971 avss 0.0112f
C12845 avdd.n9972 avss -2.75e-19
C12846 avdd.n9973 avss 0.00821f
C12847 avdd.n9974 avss 0.00821f
C12848 avdd.n9975 avss -2.75e-19
C12849 avdd.n9976 avss 0.0442f
C12850 avdd.n9977 avss 0.0179f
C12851 avdd.n9978 avss -2.22e-19
C12852 avdd.n9979 avss -1.59e-19
C12853 avdd.n9980 avss -2.33e-19
C12854 avdd.n9981 avss 0.0188f
C12855 avdd.n9982 avss 0.0181f
C12856 avdd.n9983 avss -2.75e-19
C12857 avdd.n9984 avss -3.39e-19
C12858 avdd.n9985 avss -3.6e-19
C12859 avdd.n9986 avss -2.01e-19
C12860 avdd.n9987 avss -0.0866f
C12861 avdd.n9988 avss -0.00336f
C12862 avdd.n9989 avss 0.00725f
C12863 avdd.n9990 avss 0.0318f
C12864 avdd.n9991 avss -0.00158f
C12865 avdd.n9992 avss -8.47e-19
C12866 avdd.n9993 avss 0.0298f
C12867 avdd.n9994 avss -2.22e-19
C12868 avdd.n9995 avss 0.0148f
C12869 avdd.n9996 avss 0.0182f
C12870 avdd.n9997 avss -1.8e-19
C12871 avdd.n9998 avss -2.54e-19
C12872 avdd.n9999 avss -2.54e-19
C12873 avdd.n10000 avss -1.8e-19
C12874 avdd.n10001 avss -1.16e-19
C12875 avdd.n10002 avss -0.00126f
C12876 avdd.n10003 avss -2.33e-19
C12877 avdd.n10004 avss -3.39e-19
C12878 avdd.n10005 avss -4.23e-19
C12879 avdd.n10006 avss 0.00358f
C12880 avdd.n10007 avss 0.0374f
C12881 avdd.n10008 avss -3.07e-19
C12882 avdd.n10009 avss -0.00108f
C12883 avdd.n10010 avss -0.00109f
C12884 avdd.n10011 avss 0.0192f
C12885 avdd.n10012 avss -1.59e-19
C12886 avdd.n10013 avss -1.8e-19
C12887 avdd.n10014 avss 0.00875f
C12888 avdd.n10015 avss 0.0111f
C12889 avdd.n10016 avss 0.0154f
C12890 avdd.n10017 avss 0.0183f
C12891 avdd.n10018 avss -1.8e-19
C12892 avdd.n10019 avss -2.22e-19
C12893 avdd.n10020 avss -2.22e-19
C12894 avdd.n10021 avss -1.8e-19
C12895 avdd.n10022 avss -2.01e-19
C12896 avdd.n10023 avss -9.76e-19
C12897 avdd.n10024 avss -0.00121f
C12898 avdd.n10025 avss -0.00122f
C12899 avdd.n10026 avss -0.00173f
C12900 avdd.n10027 avss -0.00357f
C12901 avdd.n10028 avss 0.0382f
C12902 avdd.n10029 avss 0.00378f
C12903 avdd.n10030 avss 0.0346f
C12904 avdd.n10031 avss -8.47e-19
C12905 avdd.n10032 avss -3.39e-19
C12906 avdd.n10033 avss -8.47e-19
C12907 avdd.n10034 avss 3e-19
C12908 avdd.n10035 avss 0.0388f
C12909 avdd.n10036 avss -3.39e-19
C12910 avdd.n10037 avss -6.46e-19
C12911 avdd.n10038 avss -5.82e-19
C12912 avdd.n10039 avss -3.39e-19
C12913 avdd.n10040 avss -8.47e-19
C12914 avdd.n10041 avss -0.00113f
C12915 avdd.n10042 avss 0.0384f
C12916 avdd.n10043 avss -2.44e-19
C12917 avdd.n10044 avss 0.0422f
C12918 avdd.n10045 avss 0.019f
C12919 avdd.n10046 avss -1.8e-19
C12920 avdd.n10047 avss 0.0197f
C12921 avdd.n10048 avss -2.44e-19
C12922 avdd.n10049 avss -2.33e-19
C12923 avdd.n10050 avss -2.33e-19
C12924 avdd.n10051 avss -1.48e-19
C12925 avdd.n10052 avss -1.27e-19
C12926 avdd.n10053 avss 0.00203f
C12927 avdd.n10054 avss -0.00128f
C12928 avdd.n10055 avss -4.76e-19
C12929 avdd.n10056 avss -2.22e-19
C12930 avdd.n10057 avss 0.0192f
C12931 avdd.n10058 avss -2.22e-19
C12932 avdd.n10059 avss 0.0148f
C12933 avdd.n10060 avss 0.0182f
C12934 avdd.n10061 avss -1.8e-19
C12935 avdd.n10062 avss -2.54e-19
C12936 avdd.n10063 avss -2.54e-19
C12937 avdd.n10064 avss -1.8e-19
C12938 avdd.n10065 avss -1.16e-19
C12939 avdd.n10066 avss -2.33e-19
C12940 avdd.n10067 avss 0.0342f
C12941 avdd.n10068 avss 0.0049f
C12942 avdd.n10069 avss -8.47e-19
C12943 avdd.n10070 avss -3.39e-19
C12944 avdd.n10071 avss -3.07e-19
C12945 avdd.n10072 avss -1.59e-19
C12946 avdd.n10073 avss -1.8e-19
C12947 avdd.n10074 avss 0.0192f
C12948 avdd.n10075 avss -1.59e-19
C12949 avdd.n10076 avss -1.8e-19
C12950 avdd.n10077 avss 0.00875f
C12951 avdd.n10078 avss 0.0111f
C12952 avdd.n10079 avss 0.0154f
C12953 avdd.n10080 avss 0.0183f
C12954 avdd.n10081 avss -1.8e-19
C12955 avdd.n10082 avss -2.22e-19
C12956 avdd.n10083 avss -2.22e-19
C12957 avdd.n10084 avss -1.8e-19
C12958 avdd.n10085 avss -2.01e-19
C12959 avdd.n10086 avss -3.18e-19
C12960 avdd.n10087 avss 0.03f
C12961 avdd.n10088 avss 0.00899f
C12962 avdd.n10089 avss -7.52e-19
C12963 avdd.n10090 avss -2.96e-19
C12964 avdd.n10091 avss -1.8e-19
C12965 avdd.n10092 avss -1.8e-19
C12966 avdd.n10093 avss 0.00873f
C12967 avdd.n10094 avss 0.0111f
C12968 avdd.n10095 avss 0.0154f
C12969 avdd.n10096 avss 0.0191f
C12970 avdd.n10097 avss -1.8e-19
C12971 avdd.n10098 avss 0.0184f
C12972 avdd.n10099 avss -1.38e-19
C12973 avdd.n10100 avss -1.8e-19
C12974 avdd.n10101 avss -2.44e-19
C12975 avdd.n10102 avss -2.44e-19
C12976 avdd.n10103 avss -1.8e-19
C12977 avdd.n10104 avss -1.38e-19
C12978 avdd.n10105 avss -3.49e-19
C12979 avdd.n10106 avss 0.0269f
C12980 avdd.n10107 avss 0.00869f
C12981 avdd.n10108 avss -0.00173f
C12982 avdd.n10110 avss -0.00512f
C12983 avdd.n10112 avss 0.0382f
C12984 avdd.n10113 avss -0.137f
C12985 avdd.n10114 avss -8.47e-19
C12986 avdd.n10115 avss -3.28e-19
C12987 avdd.n10116 avss -3.28e-19
C12988 avdd.n10117 avss -8.26e-19
C12989 avdd.n10118 avss 0.0348f
C12990 avdd.n10119 avss 0.00357f
C12991 avdd.n10120 avss -8.47e-19
C12992 avdd.n10121 avss -3.39e-19
C12993 avdd.n10122 avss -8.47e-19
C12994 avdd.n10123 avss 0.0344f
C12995 avdd.n10124 avss 0.00466f
C12996 avdd.n10125 avss -3.39e-19
C12997 avdd.n10126 avss -6.67e-19
C12998 avdd.n10127 avss -5.61e-19
C12999 avdd.n10128 avss -3.39e-19
C13000 avdd.n10129 avss -6.35e-19
C13001 avdd.n10130 avss -5.77e-19
C13002 avdd.n10131 avss 0.0398f
C13003 avdd.n10132 avss -3.07e-19
C13004 avdd.n10133 avss -1.8e-19
C13005 avdd.n10134 avss 0.0168f
C13006 avdd.n10135 avss 0.0189f
C13007 avdd.n10136 avss 0.0111f
C13008 avdd.n10137 avss 0.00875f
C13009 avdd.n10138 avss 0.0167f
C13010 avdd.n10139 avss 0.0181f
C13011 avdd.n10140 avss -3.6e-19
C13012 avdd.n10141 avss -2.01e-19
C13013 avdd.n10142 avss -3.07e-19
C13014 avdd.n10143 avss -6.46e-19
C13015 avdd.n10144 avss -0.00137f
C13016 avdd.n10145 avss -0.0013f
C13017 avdd.n10146 avss -5.19e-19
C13018 avdd.n10147 avss 0.0386f
C13019 avdd.n10148 avss 0.00873f
C13020 avdd.n10149 avss 0.0111f
C13021 avdd.n10150 avss 0.0148f
C13022 avdd.n10151 avss 0.019f
C13023 avdd.n10152 avss -1.8e-19
C13024 avdd.n10153 avss 0.0184f
C13025 avdd.n10154 avss -2.44e-19
C13026 avdd.n10155 avss -2.33e-19
C13027 avdd.n10156 avss 0.0022f
C13028 avdd.n10157 avss -1.48e-19
C13029 avdd.n10158 avss -1.27e-19
C13030 avdd.n10159 avss -2.44e-19
C13031 avdd.n10160 avss -8.15e-19
C13032 avdd.n10161 avss -0.0014f
C13033 avdd.n10162 avss -8.47e-19
C13034 avdd.n10163 avss -3.39e-19
C13035 avdd.n10164 avss -3.49e-19
C13036 avdd.n10165 avss -1.38e-19
C13037 avdd.n10166 avss -1.8e-19
C13038 avdd.n10167 avss 0.00873f
C13039 avdd.n10168 avss 0.0111f
C13040 avdd.n10169 avss 0.0154f
C13041 avdd.n10170 avss 0.0191f
C13042 avdd.n10171 avss -1.8e-19
C13043 avdd.n10172 avss 0.0184f
C13044 avdd.n10173 avss -1.38e-19
C13045 avdd.n10174 avss -1.8e-19
C13046 avdd.n10175 avss -2.44e-19
C13047 avdd.n10176 avss 0.0411f
C13048 avdd.n10177 avss -1.8e-19
C13049 avdd.n10178 avss -1.8e-19
C13050 avdd.n10179 avss -2.96e-19
C13051 avdd.n10180 avss -0.00139f
C13052 avdd.n10181 avss 0.0098f
C13053 avdd.n10182 avss 0.0298f
C13054 avdd.n10183 avss -2.22e-19
C13055 avdd.n10184 avss 0.0188f
C13056 avdd.n10185 avss -2.33e-19
C13057 avdd.n10186 avss -1.59e-19
C13058 avdd.n10187 avss -2.22e-19
C13059 avdd.n10188 avss 0.00821f
C13060 avdd.n10189 avss -2.75e-19
C13061 avdd.n10190 avss 0.0112f
C13062 avdd.n10191 avss 0.0148f
C13063 avdd.n10192 avss 0.0182f
C13064 avdd.n10193 avss -1.8e-19
C13065 avdd.n10194 avss -2.54e-19
C13066 avdd.n10195 avss -2.54e-19
C13067 avdd.n10196 avss -1.8e-19
C13068 avdd.n10197 avss -1.16e-19
C13069 avdd.n10198 avss -2.33e-19
C13070 avdd.n10199 avss -0.00126f
C13071 avdd.n10200 avss -0.00109f
C13072 avdd.n10201 avss -0.00108f
C13073 avdd.n10202 avss -3.07e-19
C13074 avdd.n10203 avss 0.0374f
C13075 avdd.n10204 avss 0.00358f
C13076 avdd.n10205 avss 0.0192f
C13077 avdd.n10206 avss -1.59e-19
C13078 avdd.n10207 avss -1.8e-19
C13079 avdd.n10208 avss 0.00875f
C13080 avdd.n10209 avss 0.0111f
C13081 avdd.n10210 avss 0.0154f
C13082 avdd.n10211 avss 0.0183f
C13083 avdd.n10212 avss -1.8e-19
C13084 avdd.n10213 avss -2.22e-19
C13085 avdd.n10214 avss -2.22e-19
C13086 avdd.n10215 avss -1.8e-19
C13087 avdd.n10216 avss -2.01e-19
C13088 avdd.n10217 avss -9.59e-19
C13089 avdd.n10218 avss -0.00106f
C13090 avdd.n10219 avss -0.00173f
C13091 avdd.n10220 avss -0.00139f
C13092 avdd.n10221 avss -6.88e-19
C13093 avdd.n10222 avss -3.07e-19
C13094 avdd.n10223 avss -1.8e-19
C13095 avdd.n10224 avss 0.00821f
C13096 avdd.n10225 avss -2.75e-19
C13097 avdd.n10226 avss 0.0442f
C13098 avdd.n10227 avss 0.0179f
C13099 avdd.n10228 avss 0.0181f
C13100 avdd.n10229 avss -2.75e-19
C13101 avdd.n10230 avss -3.39e-19
C13102 avdd.n10231 avss -3.6e-19
C13103 avdd.n10232 avss -2.01e-19
C13104 avdd.n10233 avss -0.0866f
C13105 avdd.n10234 avss -0.00336f
C13106 avdd.n10235 avss 0.00725f
C13107 avdd.n10236 avss 0.0318f
C13108 avdd.n10237 avss -0.00158f
C13109 avdd.n10238 avss -8.47e-19
C13110 avdd.n10239 avss -3.39e-19
C13111 avdd.n10240 avss -4.23e-19
C13112 avdd.n10241 avss -0.00357f
C13113 avdd.n10243 avss 0.0382f
C13114 avdd.n10244 avss -0.166f
C13115 avdd.n10245 avss 0.00378f
C13116 avdd.n10246 avss 0.0346f
C13117 avdd.n10247 avss -8.47e-19
C13118 avdd.n10248 avss -3.39e-19
C13119 avdd.n10249 avss -8.47e-19
C13120 avdd.n10250 avss 3e-19
C13121 avdd.n10251 avss 0.0388f
C13122 avdd.n10252 avss -3.39e-19
C13123 avdd.n10253 avss -6.46e-19
C13124 avdd.n10254 avss -5.82e-19
C13125 avdd.n10255 avss -3.39e-19
C13126 avdd.n10256 avss -8.47e-19
C13127 avdd.n10257 avss -0.00113f
C13128 avdd.n10258 avss 0.0384f
C13129 avdd.n10259 avss -2.44e-19
C13130 avdd.n10260 avss 0.0422f
C13131 avdd.n10261 avss 0.019f
C13132 avdd.n10262 avss -1.8e-19
C13133 avdd.n10263 avss 0.0197f
C13134 avdd.n10264 avss -2.44e-19
C13135 avdd.n10265 avss -2.33e-19
C13136 avdd.n10266 avss -2.33e-19
C13137 avdd.n10267 avss -1.48e-19
C13138 avdd.n10269 avss -1.27e-19
C13139 avdd.n10270 avss 0.00203f
C13140 avdd.n10271 avss -6.46e-19
C13141 avdd.n10272 avss -3.07e-19
C13142 avdd.n10273 avss 0.00873f
C13143 avdd.n10274 avss 0.0168f
C13144 avdd.n10275 avss 0.0189f
C13145 avdd.n10276 avss 0.0167f
C13146 avdd.n10277 avss 0.0181f
C13147 avdd.n10278 avss -3.6e-19
C13148 avdd.n10279 avss -2.01e-19
C13149 avdd.n10280 avss -1.8e-19
C13150 avdd.n10281 avss -3.07e-19
C13151 avdd.n10282 avss 0.0398f
C13152 avdd.n10283 avss -5.77e-19
C13153 avdd.n10284 avss -0.00128f
C13154 avdd.n10285 avss -4.76e-19
C13155 avdd.n10286 avss -2.22e-19
C13156 avdd.n10287 avss 0.0192f
C13157 avdd.n10288 avss -2.22e-19
C13158 avdd.n10289 avss 0.00875f
C13159 avdd.n10290 avss 0.0111f
C13160 avdd.n10291 avss 0.0148f
C13161 avdd.n10292 avss 0.0182f
C13162 avdd.n10293 avss -1.8e-19
C13163 avdd.n10294 avss -2.54e-19
C13164 avdd.n10295 avss -2.54e-19
C13165 avdd.n10296 avss -1.8e-19
C13166 avdd.n10297 avss -1.16e-19
C13167 avdd.n10298 avss -2.33e-19
C13168 avdd.n10299 avss 0.0342f
C13169 avdd.n10300 avss 0.0049f
C13170 avdd.n10301 avss -8.47e-19
C13171 avdd.n10302 avss -3.39e-19
C13172 avdd.n10303 avss -3.07e-19
C13173 avdd.n10304 avss -1.59e-19
C13174 avdd.n10305 avss -1.8e-19
C13175 avdd.n10306 avss 0.0192f
C13176 avdd.n10307 avss -1.59e-19
C13177 avdd.n10308 avss -1.8e-19
C13178 avdd.n10309 avss 0.00875f
C13179 avdd.n10310 avss 0.0111f
C13180 avdd.n10311 avss 0.0154f
C13181 avdd.n10312 avss 0.0183f
C13182 avdd.n10313 avss -1.8e-19
C13183 avdd.n10314 avss -2.22e-19
C13184 avdd.n10315 avss -2.22e-19
C13185 avdd.n10316 avss -1.8e-19
C13186 avdd.n10317 avss -2.01e-19
C13187 avdd.n10318 avss -3.18e-19
C13188 avdd.n10319 avss 0.03f
C13189 avdd.n10320 avss 0.00908f
C13190 avdd.n10321 avss -8.47e-19
C13191 avdd.n10322 avss -2.96e-19
C13192 avdd.n10323 avss -1.8e-19
C13193 avdd.n10324 avss -1.8e-19
C13194 avdd.n10325 avss 0.00873f
C13195 avdd.n10326 avss 0.0111f
C13196 avdd.n10327 avss 0.0154f
C13197 avdd.n10328 avss 0.0191f
C13198 avdd.n10329 avss -1.8e-19
C13199 avdd.n10330 avss 0.0184f
C13200 avdd.n10331 avss -1.38e-19
C13201 avdd.n10332 avss -1.8e-19
C13202 avdd.n10333 avss -2.44e-19
C13203 avdd.n10334 avss -2.44e-19
C13204 avdd.n10335 avss -1.8e-19
C13205 avdd.n10336 avss -1.38e-19
C13206 avdd.n10337 avss -3.49e-19
C13207 avdd.n10339 avss 0.0269f
C13208 avdd.n10340 avss 0.00869f
C13209 avdd.n10341 avss -0.00173f
C13210 avdd.n10342 avss -0.00512f
C13211 avdd.n10344 avss 0.0382f
C13212 avdd.n10345 avss -0.139f
C13213 avdd.n10346 avss -0.168f
C13214 avdd.n10347 avss 0.00378f
C13215 avdd.n10348 avss 0.0346f
C13216 avdd.n10349 avss -8.47e-19
C13217 avdd.n10350 avss -3.39e-19
C13218 avdd.n10351 avss -8.47e-19
C13219 avdd.n10352 avss 3e-19
C13220 avdd.n10353 avss 0.0388f
C13221 avdd.n10354 avss -3.39e-19
C13222 avdd.n10355 avss -6.46e-19
C13223 avdd.n10356 avss -5.82e-19
C13224 avdd.n10357 avss -3.39e-19
C13225 avdd.n10358 avss -8.47e-19
C13226 avdd.n10359 avss -0.00113f
C13227 avdd.n10360 avss 0.0384f
C13228 avdd.n10361 avss -2.44e-19
C13229 avdd.n10362 avss 0.0422f
C13230 avdd.n10363 avss 0.019f
C13231 avdd.n10364 avss -1.8e-19
C13232 avdd.n10365 avss 0.0197f
C13233 avdd.n10366 avss -2.44e-19
C13234 avdd.n10367 avss -2.33e-19
C13235 avdd.n10368 avss -2.33e-19
C13236 avdd.n10369 avss -1.48e-19
C13237 avdd.n10371 avss -1.27e-19
C13238 avdd.n10372 avss 0.00203f
C13239 avdd.n10373 avss -6.46e-19
C13240 avdd.n10374 avss -3.07e-19
C13241 avdd.n10375 avss 0.00873f
C13242 avdd.n10376 avss 0.0168f
C13243 avdd.n10377 avss 0.0189f
C13244 avdd.n10378 avss 0.0167f
C13245 avdd.n10379 avss 0.0181f
C13246 avdd.n10380 avss -3.6e-19
C13247 avdd.n10381 avss -2.01e-19
C13248 avdd.n10382 avss -1.8e-19
C13249 avdd.n10383 avss -3.07e-19
C13250 avdd.n10384 avss 0.0398f
C13251 avdd.n10385 avss -5.77e-19
C13252 avdd.n10386 avss -0.00128f
C13253 avdd.n10387 avss -4.76e-19
C13254 avdd.n10388 avss -2.22e-19
C13255 avdd.n10389 avss 0.0192f
C13256 avdd.n10390 avss -2.22e-19
C13257 avdd.n10391 avss 0.00875f
C13258 avdd.n10392 avss 0.0111f
C13259 avdd.n10393 avss 0.0148f
C13260 avdd.n10394 avss 0.0182f
C13261 avdd.n10395 avss -1.8e-19
C13262 avdd.n10396 avss -2.54e-19
C13263 avdd.n10397 avss -2.54e-19
C13264 avdd.n10398 avss -1.8e-19
C13265 avdd.n10399 avss -1.16e-19
C13266 avdd.n10400 avss -2.33e-19
C13267 avdd.n10401 avss 0.0342f
C13268 avdd.n10402 avss 0.0049f
C13269 avdd.n10403 avss -8.47e-19
C13270 avdd.n10404 avss -3.39e-19
C13271 avdd.n10405 avss -3.07e-19
C13272 avdd.n10406 avss -1.59e-19
C13273 avdd.n10407 avss -1.8e-19
C13274 avdd.n10408 avss 0.0192f
C13275 avdd.n10409 avss -1.59e-19
C13276 avdd.n10410 avss -1.8e-19
C13277 avdd.n10411 avss 0.00875f
C13278 avdd.n10412 avss 0.0111f
C13279 avdd.n10413 avss 0.0154f
C13280 avdd.n10414 avss 0.0183f
C13281 avdd.n10415 avss -1.8e-19
C13282 avdd.n10416 avss -2.22e-19
C13283 avdd.n10417 avss -2.22e-19
C13284 avdd.n10418 avss -1.8e-19
C13285 avdd.n10419 avss -2.01e-19
C13286 avdd.n10420 avss -3.18e-19
C13287 avdd.n10421 avss 0.03f
C13288 avdd.n10422 avss 0.00908f
C13289 avdd.n10423 avss -8.47e-19
C13290 avdd.n10424 avss -2.96e-19
C13291 avdd.n10425 avss -1.8e-19
C13292 avdd.n10426 avss -1.8e-19
C13293 avdd.n10427 avss 0.00873f
C13294 avdd.n10428 avss 0.0111f
C13295 avdd.n10429 avss 0.0154f
C13296 avdd.n10430 avss 0.0191f
C13297 avdd.n10431 avss -1.8e-19
C13298 avdd.n10432 avss 0.0184f
C13299 avdd.n10433 avss -1.38e-19
C13300 avdd.n10434 avss -1.8e-19
C13301 avdd.n10435 avss -2.44e-19
C13302 avdd.n10436 avss -2.44e-19
C13303 avdd.n10437 avss -1.8e-19
C13304 avdd.n10438 avss -1.38e-19
C13305 avdd.n10439 avss -3.49e-19
C13306 avdd.n10441 avss 0.0269f
C13307 avdd.n10442 avss 0.00869f
C13308 avdd.n10443 avss -0.00173f
C13309 avdd.n10444 avss -0.00512f
C13310 avdd.n10446 avss 0.0382f
C13311 avdd.n10447 avss -0.139f
C13312 avdd.n10448 avss -0.167f
C13313 avdd.n10449 avss 0.00378f
C13314 avdd.n10450 avss 0.0346f
C13315 avdd.n10451 avss -8.47e-19
C13316 avdd.n10452 avss -3.39e-19
C13317 avdd.n10453 avss -8.47e-19
C13318 avdd.n10454 avss 3e-19
C13319 avdd.n10455 avss 0.0388f
C13320 avdd.n10456 avss -3.39e-19
C13321 avdd.n10457 avss -6.46e-19
C13322 avdd.n10458 avss -5.82e-19
C13323 avdd.n10459 avss -3.39e-19
C13324 avdd.n10460 avss -8.47e-19
C13325 avdd.n10461 avss -0.00113f
C13326 avdd.n10462 avss 0.0384f
C13327 avdd.n10463 avss -2.44e-19
C13328 avdd.n10464 avss 0.0422f
C13329 avdd.n10465 avss 0.019f
C13330 avdd.n10466 avss -1.8e-19
C13331 avdd.n10467 avss 0.0197f
C13332 avdd.n10468 avss -2.44e-19
C13333 avdd.n10469 avss -2.33e-19
C13334 avdd.n10470 avss -2.33e-19
C13335 avdd.n10471 avss -1.48e-19
C13336 avdd.n10473 avss -1.27e-19
C13337 avdd.n10474 avss 0.00203f
C13338 avdd.n10475 avss -6.46e-19
C13339 avdd.n10476 avss -3.07e-19
C13340 avdd.n10477 avss 0.00873f
C13341 avdd.n10478 avss 0.0168f
C13342 avdd.n10479 avss 0.0189f
C13343 avdd.n10480 avss 0.0167f
C13344 avdd.n10481 avss 0.0181f
C13345 avdd.n10482 avss -3.6e-19
C13346 avdd.n10483 avss -2.01e-19
C13347 avdd.n10484 avss -1.8e-19
C13348 avdd.n10485 avss -3.07e-19
C13349 avdd.n10486 avss 0.0398f
C13350 avdd.n10487 avss -5.77e-19
C13351 avdd.n10488 avss -0.00128f
C13352 avdd.n10489 avss -4.76e-19
C13353 avdd.n10490 avss -2.22e-19
C13354 avdd.n10491 avss 0.0192f
C13355 avdd.n10492 avss -2.22e-19
C13356 avdd.n10493 avss 0.00875f
C13357 avdd.n10494 avss 0.0111f
C13358 avdd.n10495 avss 0.0148f
C13359 avdd.n10496 avss 0.0182f
C13360 avdd.n10497 avss -1.8e-19
C13361 avdd.n10498 avss -2.54e-19
C13362 avdd.n10499 avss -2.54e-19
C13363 avdd.n10500 avss -1.8e-19
C13364 avdd.n10501 avss -1.16e-19
C13365 avdd.n10502 avss -2.33e-19
C13366 avdd.n10503 avss 0.0342f
C13367 avdd.n10504 avss 0.0049f
C13368 avdd.n10505 avss -8.47e-19
C13369 avdd.n10506 avss -3.39e-19
C13370 avdd.n10507 avss -3.07e-19
C13371 avdd.n10508 avss -1.59e-19
C13372 avdd.n10509 avss -1.8e-19
C13373 avdd.n10510 avss 0.0192f
C13374 avdd.n10511 avss -1.59e-19
C13375 avdd.n10512 avss -1.8e-19
C13376 avdd.n10513 avss 0.00875f
C13377 avdd.n10514 avss 0.0111f
C13378 avdd.n10515 avss 0.0154f
C13379 avdd.n10516 avss 0.0183f
C13380 avdd.n10517 avss -1.8e-19
C13381 avdd.n10518 avss -2.22e-19
C13382 avdd.n10519 avss -2.22e-19
C13383 avdd.n10520 avss -1.8e-19
C13384 avdd.n10521 avss -2.01e-19
C13385 avdd.n10522 avss -3.18e-19
C13386 avdd.n10523 avss 0.03f
C13387 avdd.n10524 avss 0.00908f
C13388 avdd.n10525 avss -8.47e-19
C13389 avdd.n10526 avss -2.96e-19
C13390 avdd.n10527 avss -1.8e-19
C13391 avdd.n10528 avss -1.8e-19
C13392 avdd.n10529 avss 0.00873f
C13393 avdd.n10530 avss 0.0111f
C13394 avdd.n10531 avss 0.0154f
C13395 avdd.n10532 avss 0.0191f
C13396 avdd.n10533 avss -1.8e-19
C13397 avdd.n10534 avss 0.0184f
C13398 avdd.n10535 avss -1.38e-19
C13399 avdd.n10536 avss -1.8e-19
C13400 avdd.n10537 avss -2.44e-19
C13401 avdd.n10538 avss -2.44e-19
C13402 avdd.n10539 avss -1.8e-19
C13403 avdd.n10540 avss -1.38e-19
C13404 avdd.n10541 avss -3.49e-19
C13405 avdd.n10543 avss 0.0269f
C13406 avdd.n10544 avss 0.00869f
C13407 avdd.n10545 avss -0.00173f
C13408 avdd.n10546 avss -0.00512f
C13409 avdd.n10548 avss 0.0382f
C13410 avdd.n10549 avss -0.138f
C13411 avdd.n10550 avss -0.168f
C13412 avdd.n10551 avss 0.00378f
C13413 avdd.n10552 avss 0.0346f
C13414 avdd.n10553 avss -8.47e-19
C13415 avdd.n10554 avss -3.39e-19
C13416 avdd.n10555 avss -8.47e-19
C13417 avdd.n10556 avss 3e-19
C13418 avdd.n10557 avss 0.0388f
C13419 avdd.n10558 avss -3.39e-19
C13420 avdd.n10559 avss -6.46e-19
C13421 avdd.n10560 avss -5.82e-19
C13422 avdd.n10561 avss -3.39e-19
C13423 avdd.n10562 avss -8.47e-19
C13424 avdd.n10563 avss -0.00113f
C13425 avdd.n10564 avss 0.0384f
C13426 avdd.n10565 avss -2.44e-19
C13427 avdd.n10566 avss 0.0422f
C13428 avdd.n10567 avss 0.019f
C13429 avdd.n10568 avss -1.8e-19
C13430 avdd.n10569 avss 0.0197f
C13431 avdd.n10570 avss -2.44e-19
C13432 avdd.n10571 avss -2.33e-19
C13433 avdd.n10572 avss -2.33e-19
C13434 avdd.n10573 avss -1.48e-19
C13435 avdd.n10575 avss -1.27e-19
C13436 avdd.n10576 avss 0.00203f
C13437 avdd.n10577 avss -6.46e-19
C13438 avdd.n10578 avss -3.07e-19
C13439 avdd.n10579 avss 0.00873f
C13440 avdd.n10580 avss 0.0168f
C13441 avdd.n10581 avss 0.0189f
C13442 avdd.n10582 avss 0.0167f
C13443 avdd.n10583 avss 0.0181f
C13444 avdd.n10584 avss -3.6e-19
C13445 avdd.n10585 avss -2.01e-19
C13446 avdd.n10586 avss -1.8e-19
C13447 avdd.n10587 avss -3.07e-19
C13448 avdd.n10588 avss 0.0398f
C13449 avdd.n10589 avss -5.77e-19
C13450 avdd.n10590 avss -0.00128f
C13451 avdd.n10591 avss -4.76e-19
C13452 avdd.n10592 avss -2.22e-19
C13453 avdd.n10593 avss 0.0192f
C13454 avdd.n10594 avss -2.22e-19
C13455 avdd.n10595 avss 0.00875f
C13456 avdd.n10596 avss 0.0111f
C13457 avdd.n10597 avss 0.0148f
C13458 avdd.n10598 avss 0.0182f
C13459 avdd.n10599 avss -1.8e-19
C13460 avdd.n10600 avss -2.54e-19
C13461 avdd.n10601 avss -2.54e-19
C13462 avdd.n10602 avss -1.8e-19
C13463 avdd.n10603 avss -1.16e-19
C13464 avdd.n10604 avss -2.33e-19
C13465 avdd.n10605 avss 0.0342f
C13466 avdd.n10606 avss 0.0049f
C13467 avdd.n10607 avss -8.47e-19
C13468 avdd.n10608 avss -3.39e-19
C13469 avdd.n10609 avss -3.07e-19
C13470 avdd.n10610 avss -1.59e-19
C13471 avdd.n10611 avss -1.8e-19
C13472 avdd.n10612 avss 0.0192f
C13473 avdd.n10613 avss -1.59e-19
C13474 avdd.n10614 avss -1.8e-19
C13475 avdd.n10615 avss 0.00875f
C13476 avdd.n10616 avss 0.0111f
C13477 avdd.n10617 avss 0.0154f
C13478 avdd.n10618 avss 0.0183f
C13479 avdd.n10619 avss -1.8e-19
C13480 avdd.n10620 avss -2.22e-19
C13481 avdd.n10621 avss -2.22e-19
C13482 avdd.n10622 avss -1.8e-19
C13483 avdd.n10623 avss -2.01e-19
C13484 avdd.n10624 avss -3.18e-19
C13485 avdd.n10625 avss 0.03f
C13486 avdd.n10626 avss 0.00908f
C13487 avdd.n10627 avss -8.47e-19
C13488 avdd.n10628 avss -2.96e-19
C13489 avdd.n10629 avss -1.8e-19
C13490 avdd.n10630 avss -1.8e-19
C13491 avdd.n10631 avss 0.00873f
C13492 avdd.n10632 avss 0.0111f
C13493 avdd.n10633 avss 0.0154f
C13494 avdd.n10634 avss 0.0191f
C13495 avdd.n10635 avss -1.8e-19
C13496 avdd.n10636 avss 0.0184f
C13497 avdd.n10637 avss -1.38e-19
C13498 avdd.n10638 avss -1.8e-19
C13499 avdd.n10639 avss -2.44e-19
C13500 avdd.n10640 avss -2.44e-19
C13501 avdd.n10641 avss -1.8e-19
C13502 avdd.n10642 avss -1.38e-19
C13503 avdd.n10643 avss -3.49e-19
C13504 avdd.n10645 avss 0.0269f
C13505 avdd.n10646 avss 0.00869f
C13506 avdd.n10647 avss -0.00173f
C13507 avdd.n10648 avss -0.00512f
C13508 avdd.n10650 avss 0.0382f
C13509 avdd.n10651 avss -0.139f
C13510 avdd.n10652 avss -0.168f
C13511 avdd.n10653 avss 0.00378f
C13512 avdd.n10654 avss 0.0346f
C13513 avdd.n10655 avss -8.47e-19
C13514 avdd.n10656 avss -3.39e-19
C13515 avdd.n10657 avss -8.47e-19
C13516 avdd.n10658 avss 3e-19
C13517 avdd.n10659 avss 0.0388f
C13518 avdd.n10660 avss -3.39e-19
C13519 avdd.n10661 avss -6.46e-19
C13520 avdd.n10662 avss -5.82e-19
C13521 avdd.n10663 avss -3.39e-19
C13522 avdd.n10664 avss -8.47e-19
C13523 avdd.n10665 avss -0.00113f
C13524 avdd.n10666 avss 0.0384f
C13525 avdd.n10667 avss -2.44e-19
C13526 avdd.n10668 avss 0.0422f
C13527 avdd.n10669 avss 0.019f
C13528 avdd.n10670 avss -1.8e-19
C13529 avdd.n10671 avss 0.0197f
C13530 avdd.n10672 avss -2.44e-19
C13531 avdd.n10673 avss -2.33e-19
C13532 avdd.n10674 avss -2.33e-19
C13533 avdd.n10675 avss -1.48e-19
C13534 avdd.n10677 avss -1.27e-19
C13535 avdd.n10678 avss 0.00203f
C13536 avdd.n10679 avss -6.46e-19
C13537 avdd.n10680 avss -3.07e-19
C13538 avdd.n10681 avss 0.00873f
C13539 avdd.n10682 avss 0.0168f
C13540 avdd.n10683 avss 0.0189f
C13541 avdd.n10684 avss 0.0167f
C13542 avdd.n10685 avss 0.0181f
C13543 avdd.n10686 avss -3.6e-19
C13544 avdd.n10687 avss -2.01e-19
C13545 avdd.n10688 avss -1.8e-19
C13546 avdd.n10689 avss -3.07e-19
C13547 avdd.n10690 avss 0.0398f
C13548 avdd.n10691 avss -5.77e-19
C13549 avdd.n10692 avss -0.00128f
C13550 avdd.n10693 avss -4.76e-19
C13551 avdd.n10694 avss -2.22e-19
C13552 avdd.n10695 avss 0.0192f
C13553 avdd.n10696 avss -2.22e-19
C13554 avdd.n10697 avss 0.00875f
C13555 avdd.n10698 avss 0.0111f
C13556 avdd.n10699 avss 0.0148f
C13557 avdd.n10700 avss 0.0182f
C13558 avdd.n10701 avss -1.8e-19
C13559 avdd.n10702 avss -2.54e-19
C13560 avdd.n10703 avss -2.54e-19
C13561 avdd.n10704 avss -1.8e-19
C13562 avdd.n10705 avss -1.16e-19
C13563 avdd.n10706 avss -2.33e-19
C13564 avdd.n10707 avss 0.0342f
C13565 avdd.n10708 avss 0.0049f
C13566 avdd.n10709 avss -8.47e-19
C13567 avdd.n10710 avss -3.39e-19
C13568 avdd.n10711 avss -3.07e-19
C13569 avdd.n10712 avss -1.59e-19
C13570 avdd.n10713 avss -1.8e-19
C13571 avdd.n10714 avss 0.0192f
C13572 avdd.n10715 avss -1.59e-19
C13573 avdd.n10716 avss -1.8e-19
C13574 avdd.n10717 avss 0.00875f
C13575 avdd.n10718 avss 0.0111f
C13576 avdd.n10719 avss 0.0154f
C13577 avdd.n10720 avss 0.0183f
C13578 avdd.n10721 avss -1.8e-19
C13579 avdd.n10722 avss -2.22e-19
C13580 avdd.n10723 avss -2.22e-19
C13581 avdd.n10724 avss -1.8e-19
C13582 avdd.n10725 avss -2.01e-19
C13583 avdd.n10726 avss -3.18e-19
C13584 avdd.n10727 avss 0.03f
C13585 avdd.n10728 avss 0.00908f
C13586 avdd.n10729 avss -8.47e-19
C13587 avdd.n10730 avss -2.96e-19
C13588 avdd.n10731 avss -1.8e-19
C13589 avdd.n10732 avss -1.8e-19
C13590 avdd.n10733 avss 0.00873f
C13591 avdd.n10734 avss 0.0111f
C13592 avdd.n10735 avss 0.0154f
C13593 avdd.n10736 avss 0.0191f
C13594 avdd.n10737 avss -1.8e-19
C13595 avdd.n10738 avss 0.0184f
C13596 avdd.n10739 avss -1.38e-19
C13597 avdd.n10740 avss -1.8e-19
C13598 avdd.n10741 avss -2.44e-19
C13599 avdd.n10742 avss -2.44e-19
C13600 avdd.n10743 avss -1.8e-19
C13601 avdd.n10744 avss -1.38e-19
C13602 avdd.n10745 avss -3.49e-19
C13603 avdd.n10747 avss 0.0269f
C13604 avdd.n10748 avss 0.00869f
C13605 avdd.n10749 avss -0.00173f
C13606 avdd.n10750 avss -0.00512f
C13607 avdd.n10752 avss 0.0382f
C13608 avdd.n10753 avss -0.14f
C13609 avdd.n10754 avss -0.17f
C13610 avdd.n10755 avss 0.00378f
C13611 avdd.n10756 avss 0.0346f
C13612 avdd.n10757 avss -8.47e-19
C13613 avdd.n10758 avss -3.39e-19
C13614 avdd.n10759 avss -8.47e-19
C13615 avdd.n10760 avss 3e-19
C13616 avdd.n10761 avss 0.0388f
C13617 avdd.n10762 avss -3.39e-19
C13618 avdd.n10763 avss -6.46e-19
C13619 avdd.n10764 avss -5.82e-19
C13620 avdd.n10765 avss -3.39e-19
C13621 avdd.n10766 avss -8.47e-19
C13622 avdd.n10767 avss -0.00113f
C13623 avdd.n10768 avss 0.0384f
C13624 avdd.n10769 avss -2.44e-19
C13625 avdd.n10770 avss 0.0422f
C13626 avdd.n10771 avss 0.019f
C13627 avdd.n10772 avss -1.8e-19
C13628 avdd.n10773 avss 0.0197f
C13629 avdd.n10774 avss -2.44e-19
C13630 avdd.n10775 avss -2.33e-19
C13631 avdd.n10776 avss -2.33e-19
C13632 avdd.n10777 avss -1.48e-19
C13633 avdd.n10779 avss -1.27e-19
C13634 avdd.n10780 avss 0.00203f
C13635 avdd.n10781 avss -6.46e-19
C13636 avdd.n10782 avss -3.07e-19
C13637 avdd.n10783 avss 0.00873f
C13638 avdd.n10784 avss 0.0168f
C13639 avdd.n10785 avss 0.0189f
C13640 avdd.n10786 avss 0.0167f
C13641 avdd.n10787 avss 0.0181f
C13642 avdd.n10788 avss -3.6e-19
C13643 avdd.n10789 avss -2.01e-19
C13644 avdd.n10790 avss -1.8e-19
C13645 avdd.n10791 avss -3.07e-19
C13646 avdd.n10792 avss 0.0398f
C13647 avdd.n10793 avss -5.77e-19
C13648 avdd.n10794 avss -0.00128f
C13649 avdd.n10795 avss -4.76e-19
C13650 avdd.n10796 avss -2.22e-19
C13651 avdd.n10797 avss 0.0192f
C13652 avdd.n10798 avss -2.22e-19
C13653 avdd.n10799 avss 0.00875f
C13654 avdd.n10800 avss 0.0111f
C13655 avdd.n10801 avss 0.0148f
C13656 avdd.n10802 avss 0.0182f
C13657 avdd.n10803 avss -1.8e-19
C13658 avdd.n10804 avss -2.54e-19
C13659 avdd.n10805 avss -2.54e-19
C13660 avdd.n10806 avss -1.8e-19
C13661 avdd.n10807 avss -1.16e-19
C13662 avdd.n10808 avss -2.33e-19
C13663 avdd.n10809 avss 0.0342f
C13664 avdd.n10810 avss 0.0049f
C13665 avdd.n10811 avss -8.47e-19
C13666 avdd.n10812 avss -3.39e-19
C13667 avdd.n10813 avss -3.07e-19
C13668 avdd.n10814 avss -1.59e-19
C13669 avdd.n10815 avss -1.8e-19
C13670 avdd.n10816 avss 0.0192f
C13671 avdd.n10817 avss -1.59e-19
C13672 avdd.n10818 avss -1.8e-19
C13673 avdd.n10819 avss 0.00875f
C13674 avdd.n10820 avss 0.0111f
C13675 avdd.n10821 avss 0.0154f
C13676 avdd.n10822 avss 0.0183f
C13677 avdd.n10823 avss -1.8e-19
C13678 avdd.n10824 avss -2.22e-19
C13679 avdd.n10825 avss -2.22e-19
C13680 avdd.n10826 avss -1.8e-19
C13681 avdd.n10827 avss -2.01e-19
C13682 avdd.n10828 avss -3.18e-19
C13683 avdd.n10829 avss 0.03f
C13684 avdd.n10830 avss 0.00908f
C13685 avdd.n10831 avss -8.47e-19
C13686 avdd.n10832 avss -2.96e-19
C13687 avdd.n10833 avss -1.8e-19
C13688 avdd.n10834 avss -1.8e-19
C13689 avdd.n10835 avss 0.00873f
C13690 avdd.n10836 avss 0.0111f
C13691 avdd.n10837 avss 0.0154f
C13692 avdd.n10838 avss 0.0191f
C13693 avdd.n10839 avss -1.8e-19
C13694 avdd.n10840 avss 0.0184f
C13695 avdd.n10841 avss -1.38e-19
C13696 avdd.n10842 avss -1.8e-19
C13697 avdd.n10843 avss -2.44e-19
C13698 avdd.n10844 avss -2.44e-19
C13699 avdd.n10845 avss -1.8e-19
C13700 avdd.n10846 avss -1.38e-19
C13701 avdd.n10847 avss -3.49e-19
C13702 avdd.n10849 avss 0.0269f
C13703 avdd.n10850 avss 0.00869f
C13704 avdd.n10851 avss -0.00173f
C13705 avdd.n10852 avss -0.00512f
C13706 avdd.n10854 avss 0.0382f
C13707 avdd.n10855 avss -0.14f
C13708 avdd.n10856 avss -0.17f
C13709 avdd.n10857 avss 0.00378f
C13710 avdd.n10858 avss 0.0346f
C13711 avdd.n10859 avss -8.47e-19
C13712 avdd.n10860 avss -3.39e-19
C13713 avdd.n10861 avss -8.47e-19
C13714 avdd.n10862 avss 3e-19
C13715 avdd.n10863 avss 0.0388f
C13716 avdd.n10864 avss -3.39e-19
C13717 avdd.n10865 avss -6.46e-19
C13718 avdd.n10866 avss -5.82e-19
C13719 avdd.n10867 avss -3.39e-19
C13720 avdd.n10868 avss -8.47e-19
C13721 avdd.n10869 avss -0.00113f
C13722 avdd.n10870 avss 0.0384f
C13723 avdd.n10871 avss -2.44e-19
C13724 avdd.n10872 avss 0.0422f
C13725 avdd.n10873 avss 0.019f
C13726 avdd.n10874 avss -1.8e-19
C13727 avdd.n10875 avss 0.0197f
C13728 avdd.n10876 avss -2.44e-19
C13729 avdd.n10877 avss -2.33e-19
C13730 avdd.n10878 avss -2.33e-19
C13731 avdd.n10879 avss -1.48e-19
C13732 avdd.n10881 avss -1.27e-19
C13733 avdd.n10882 avss 0.00203f
C13734 avdd.n10883 avss -6.46e-19
C13735 avdd.n10884 avss -3.07e-19
C13736 avdd.n10885 avss 0.00873f
C13737 avdd.n10886 avss 0.0168f
C13738 avdd.n10887 avss 0.0189f
C13739 avdd.n10888 avss 0.0167f
C13740 avdd.n10889 avss 0.0181f
C13741 avdd.n10890 avss -3.6e-19
C13742 avdd.n10891 avss -2.01e-19
C13743 avdd.n10892 avss -1.8e-19
C13744 avdd.n10893 avss -3.07e-19
C13745 avdd.n10894 avss 0.0398f
C13746 avdd.n10895 avss -5.77e-19
C13747 avdd.n10896 avss -0.00128f
C13748 avdd.n10897 avss -4.76e-19
C13749 avdd.n10898 avss -2.22e-19
C13750 avdd.n10899 avss 0.0192f
C13751 avdd.n10900 avss -2.22e-19
C13752 avdd.n10901 avss 0.00875f
C13753 avdd.n10902 avss 0.0111f
C13754 avdd.n10903 avss 0.0148f
C13755 avdd.n10904 avss 0.0182f
C13756 avdd.n10905 avss -1.8e-19
C13757 avdd.n10906 avss -2.54e-19
C13758 avdd.n10907 avss -2.54e-19
C13759 avdd.n10908 avss -1.8e-19
C13760 avdd.n10909 avss -1.16e-19
C13761 avdd.n10910 avss -2.33e-19
C13762 avdd.n10911 avss 0.0342f
C13763 avdd.n10912 avss 0.0049f
C13764 avdd.n10913 avss -8.47e-19
C13765 avdd.n10914 avss -3.39e-19
C13766 avdd.n10915 avss -3.07e-19
C13767 avdd.n10916 avss -1.59e-19
C13768 avdd.n10917 avss -1.8e-19
C13769 avdd.n10918 avss 0.0192f
C13770 avdd.n10919 avss -1.59e-19
C13771 avdd.n10920 avss -1.8e-19
C13772 avdd.n10921 avss 0.00875f
C13773 avdd.n10922 avss 0.0111f
C13774 avdd.n10923 avss 0.0154f
C13775 avdd.n10924 avss 0.0183f
C13776 avdd.n10925 avss -1.8e-19
C13777 avdd.n10926 avss -2.22e-19
C13778 avdd.n10927 avss -2.22e-19
C13779 avdd.n10928 avss -1.8e-19
C13780 avdd.n10929 avss -2.01e-19
C13781 avdd.n10930 avss -3.18e-19
C13782 avdd.n10931 avss 0.03f
C13783 avdd.n10932 avss 0.00908f
C13784 avdd.n10933 avss -8.47e-19
C13785 avdd.n10934 avss -2.96e-19
C13786 avdd.n10935 avss -1.8e-19
C13787 avdd.n10936 avss -1.8e-19
C13788 avdd.n10937 avss 0.00873f
C13789 avdd.n10938 avss 0.0111f
C13790 avdd.n10939 avss 0.0154f
C13791 avdd.n10940 avss 0.0191f
C13792 avdd.n10941 avss -1.8e-19
C13793 avdd.n10942 avss 0.0184f
C13794 avdd.n10943 avss -1.38e-19
C13795 avdd.n10944 avss -1.8e-19
C13796 avdd.n10945 avss -2.44e-19
C13797 avdd.n10946 avss -2.44e-19
C13798 avdd.n10947 avss -1.8e-19
C13799 avdd.n10948 avss -1.38e-19
C13800 avdd.n10949 avss -3.49e-19
C13801 avdd.n10951 avss 0.0269f
C13802 avdd.n10952 avss 0.00869f
C13803 avdd.n10953 avss -0.00173f
C13804 avdd.n10954 avss -0.00512f
C13805 avdd.n10956 avss 0.0382f
C13806 avdd.n10957 avss -0.14f
C13807 avdd.n10958 avss -0.17f
C13808 avdd.n10959 avss 0.00378f
C13809 avdd.n10960 avss 0.0346f
C13810 avdd.n10961 avss -8.47e-19
C13811 avdd.n10962 avss -3.39e-19
C13812 avdd.n10963 avss -8.47e-19
C13813 avdd.n10964 avss 3e-19
C13814 avdd.n10965 avss 0.0388f
C13815 avdd.n10966 avss -3.39e-19
C13816 avdd.n10967 avss -6.46e-19
C13817 avdd.n10968 avss -5.82e-19
C13818 avdd.n10969 avss -3.39e-19
C13819 avdd.n10970 avss -8.47e-19
C13820 avdd.n10971 avss -0.00113f
C13821 avdd.n10972 avss 0.0384f
C13822 avdd.n10973 avss -2.44e-19
C13823 avdd.n10974 avss 0.0422f
C13824 avdd.n10975 avss 0.019f
C13825 avdd.n10976 avss -1.8e-19
C13826 avdd.n10977 avss 0.0197f
C13827 avdd.n10978 avss -2.44e-19
C13828 avdd.n10979 avss -2.33e-19
C13829 avdd.n10980 avss -2.33e-19
C13830 avdd.n10981 avss -1.48e-19
C13831 avdd.n10983 avss -1.27e-19
C13832 avdd.n10984 avss 0.00203f
C13833 avdd.n10985 avss -6.46e-19
C13834 avdd.n10986 avss -3.07e-19
C13835 avdd.n10987 avss 0.00873f
C13836 avdd.n10988 avss 0.0168f
C13837 avdd.n10989 avss 0.0189f
C13838 avdd.n10990 avss 0.0167f
C13839 avdd.n10991 avss 0.0181f
C13840 avdd.n10992 avss -3.6e-19
C13841 avdd.n10993 avss -2.01e-19
C13842 avdd.n10994 avss -1.8e-19
C13843 avdd.n10995 avss -3.07e-19
C13844 avdd.n10996 avss 0.0398f
C13845 avdd.n10997 avss -5.77e-19
C13846 avdd.n10998 avss -0.00128f
C13847 avdd.n10999 avss -4.76e-19
C13848 avdd.n11000 avss -2.22e-19
C13849 avdd.n11001 avss 0.0192f
C13850 avdd.n11002 avss -2.22e-19
C13851 avdd.n11003 avss 0.00875f
C13852 avdd.n11004 avss 0.0111f
C13853 avdd.n11005 avss 0.0148f
C13854 avdd.n11006 avss 0.0182f
C13855 avdd.n11007 avss -1.8e-19
C13856 avdd.n11008 avss -2.54e-19
C13857 avdd.n11009 avss -2.54e-19
C13858 avdd.n11010 avss -1.8e-19
C13859 avdd.n11011 avss -1.16e-19
C13860 avdd.n11012 avss -2.33e-19
C13861 avdd.n11013 avss 0.0342f
C13862 avdd.n11014 avss 0.0049f
C13863 avdd.n11015 avss -8.47e-19
C13864 avdd.n11016 avss -3.39e-19
C13865 avdd.n11017 avss -3.07e-19
C13866 avdd.n11018 avss -1.59e-19
C13867 avdd.n11019 avss -1.8e-19
C13868 avdd.n11020 avss 0.0192f
C13869 avdd.n11021 avss -1.59e-19
C13870 avdd.n11022 avss -1.8e-19
C13871 avdd.n11023 avss 0.00875f
C13872 avdd.n11024 avss 0.0111f
C13873 avdd.n11025 avss 0.0154f
C13874 avdd.n11026 avss 0.0183f
C13875 avdd.n11027 avss -1.8e-19
C13876 avdd.n11028 avss -2.22e-19
C13877 avdd.n11029 avss -2.22e-19
C13878 avdd.n11030 avss -1.8e-19
C13879 avdd.n11031 avss -2.01e-19
C13880 avdd.n11032 avss -3.18e-19
C13881 avdd.n11033 avss 0.03f
C13882 avdd.n11034 avss 0.00908f
C13883 avdd.n11035 avss -8.47e-19
C13884 avdd.n11036 avss -2.96e-19
C13885 avdd.n11037 avss -1.8e-19
C13886 avdd.n11038 avss -1.8e-19
C13887 avdd.n11039 avss 0.00873f
C13888 avdd.n11040 avss 0.0111f
C13889 avdd.n11041 avss 0.0154f
C13890 avdd.n11042 avss 0.0191f
C13891 avdd.n11043 avss -1.8e-19
C13892 avdd.n11044 avss 0.0184f
C13893 avdd.n11045 avss -1.38e-19
C13894 avdd.n11046 avss -1.8e-19
C13895 avdd.n11047 avss -2.44e-19
C13896 avdd.n11048 avss -2.44e-19
C13897 avdd.n11049 avss -1.8e-19
C13898 avdd.n11050 avss -1.38e-19
C13899 avdd.n11051 avss -3.49e-19
C13900 avdd.n11053 avss 0.0269f
C13901 avdd.n11054 avss 0.00869f
C13902 avdd.n11055 avss -0.00173f
C13903 avdd.n11056 avss -0.00512f
C13904 avdd.n11058 avss 0.0382f
C13905 avdd.n11059 avss -0.14f
C13906 avdd.n11060 avss -0.17f
C13907 avdd.n11061 avss 0.00378f
C13908 avdd.n11062 avss 0.0346f
C13909 avdd.n11063 avss -8.47e-19
C13910 avdd.n11064 avss -3.39e-19
C13911 avdd.n11065 avss -8.47e-19
C13912 avdd.n11066 avss 3e-19
C13913 avdd.n11067 avss 0.0388f
C13914 avdd.n11068 avss -3.39e-19
C13915 avdd.n11069 avss -6.46e-19
C13916 avdd.n11070 avss -5.82e-19
C13917 avdd.n11071 avss -3.39e-19
C13918 avdd.n11072 avss -8.47e-19
C13919 avdd.n11073 avss -0.00113f
C13920 avdd.n11074 avss 0.0384f
C13921 avdd.n11075 avss -2.44e-19
C13922 avdd.n11076 avss 0.0422f
C13923 avdd.n11077 avss 0.019f
C13924 avdd.n11078 avss -1.8e-19
C13925 avdd.n11079 avss 0.0197f
C13926 avdd.n11080 avss -2.44e-19
C13927 avdd.n11081 avss -2.33e-19
C13928 avdd.n11082 avss -2.33e-19
C13929 avdd.n11083 avss -1.48e-19
C13930 avdd.n11085 avss -1.27e-19
C13931 avdd.n11086 avss 0.00203f
C13932 avdd.n11087 avss -6.46e-19
C13933 avdd.n11088 avss -3.07e-19
C13934 avdd.n11089 avss 0.00873f
C13935 avdd.n11090 avss 0.0168f
C13936 avdd.n11091 avss 0.0189f
C13937 avdd.n11092 avss 0.0167f
C13938 avdd.n11093 avss 0.0181f
C13939 avdd.n11094 avss -3.6e-19
C13940 avdd.n11095 avss -2.01e-19
C13941 avdd.n11096 avss -1.8e-19
C13942 avdd.n11097 avss -3.07e-19
C13943 avdd.n11098 avss 0.0398f
C13944 avdd.n11099 avss -5.77e-19
C13945 avdd.n11100 avss -0.00128f
C13946 avdd.n11101 avss -4.76e-19
C13947 avdd.n11102 avss -2.22e-19
C13948 avdd.n11103 avss 0.0192f
C13949 avdd.n11104 avss -2.22e-19
C13950 avdd.n11105 avss 0.00875f
C13951 avdd.n11106 avss 0.0111f
C13952 avdd.n11107 avss 0.0148f
C13953 avdd.n11108 avss 0.0182f
C13954 avdd.n11109 avss -1.8e-19
C13955 avdd.n11110 avss -2.54e-19
C13956 avdd.n11111 avss -2.54e-19
C13957 avdd.n11112 avss -1.8e-19
C13958 avdd.n11113 avss -1.16e-19
C13959 avdd.n11114 avss -2.33e-19
C13960 avdd.n11115 avss 0.0342f
C13961 avdd.n11116 avss 0.0049f
C13962 avdd.n11117 avss -8.47e-19
C13963 avdd.n11118 avss -3.39e-19
C13964 avdd.n11119 avss -3.07e-19
C13965 avdd.n11120 avss -1.59e-19
C13966 avdd.n11121 avss -1.8e-19
C13967 avdd.n11122 avss 0.0192f
C13968 avdd.n11123 avss -1.59e-19
C13969 avdd.n11124 avss -1.8e-19
C13970 avdd.n11125 avss 0.00875f
C13971 avdd.n11126 avss 0.0111f
C13972 avdd.n11127 avss 0.0154f
C13973 avdd.n11128 avss 0.0183f
C13974 avdd.n11129 avss -1.8e-19
C13975 avdd.n11130 avss -2.22e-19
C13976 avdd.n11131 avss -2.22e-19
C13977 avdd.n11132 avss -1.8e-19
C13978 avdd.n11133 avss -2.01e-19
C13979 avdd.n11134 avss -3.18e-19
C13980 avdd.n11135 avss 0.03f
C13981 avdd.n11136 avss 0.00908f
C13982 avdd.n11137 avss -8.47e-19
C13983 avdd.n11138 avss -2.96e-19
C13984 avdd.n11139 avss -1.8e-19
C13985 avdd.n11140 avss -1.8e-19
C13986 avdd.n11141 avss 0.00873f
C13987 avdd.n11142 avss 0.0111f
C13988 avdd.n11143 avss 0.0154f
C13989 avdd.n11144 avss 0.0191f
C13990 avdd.n11145 avss -1.8e-19
C13991 avdd.n11146 avss 0.0184f
C13992 avdd.n11147 avss -1.38e-19
C13993 avdd.n11148 avss -1.8e-19
C13994 avdd.n11149 avss -2.44e-19
C13995 avdd.n11150 avss -2.44e-19
C13996 avdd.n11151 avss -1.8e-19
C13997 avdd.n11152 avss -1.38e-19
C13998 avdd.n11153 avss -3.49e-19
C13999 avdd.n11155 avss 0.0269f
C14000 avdd.n11156 avss 0.00869f
C14001 avdd.n11157 avss -0.00173f
C14002 avdd.n11158 avss -0.00512f
C14003 avdd.n11160 avss 0.0382f
C14004 avdd.n11161 avss -0.141f
C14005 avdd.n11162 avss -0.171f
C14006 avdd.n11163 avss 0.00378f
C14007 avdd.n11164 avss 0.0346f
C14008 avdd.n11165 avss -8.47e-19
C14009 avdd.n11166 avss -3.39e-19
C14010 avdd.n11167 avss -8.47e-19
C14011 avdd.n11168 avss 3e-19
C14012 avdd.n11169 avss 0.0388f
C14013 avdd.n11170 avss -3.39e-19
C14014 avdd.n11171 avss -6.46e-19
C14015 avdd.n11172 avss -5.82e-19
C14016 avdd.n11173 avss -3.39e-19
C14017 avdd.n11174 avss -8.47e-19
C14018 avdd.n11175 avss -0.00113f
C14019 avdd.n11176 avss 0.0384f
C14020 avdd.n11177 avss -2.44e-19
C14021 avdd.n11178 avss 0.0422f
C14022 avdd.n11179 avss 0.019f
C14023 avdd.n11180 avss -1.8e-19
C14024 avdd.n11181 avss 0.0197f
C14025 avdd.n11182 avss -2.44e-19
C14026 avdd.n11183 avss -2.33e-19
C14027 avdd.n11184 avss -2.33e-19
C14028 avdd.n11185 avss -1.48e-19
C14029 avdd.n11187 avss -1.27e-19
C14030 avdd.n11188 avss 0.00203f
C14031 avdd.n11189 avss -6.46e-19
C14032 avdd.n11190 avss -3.07e-19
C14033 avdd.n11191 avss 0.00873f
C14034 avdd.n11192 avss 0.0168f
C14035 avdd.n11193 avss 0.0189f
C14036 avdd.n11194 avss 0.0167f
C14037 avdd.n11195 avss 0.0181f
C14038 avdd.n11196 avss -3.6e-19
C14039 avdd.n11197 avss -2.01e-19
C14040 avdd.n11198 avss -1.8e-19
C14041 avdd.n11199 avss -3.07e-19
C14042 avdd.n11200 avss 0.0398f
C14043 avdd.n11201 avss -5.77e-19
C14044 avdd.n11202 avss -0.00128f
C14045 avdd.n11203 avss -4.76e-19
C14046 avdd.n11204 avss -2.22e-19
C14047 avdd.n11205 avss 0.0192f
C14048 avdd.n11206 avss -2.22e-19
C14049 avdd.n11207 avss 0.00875f
C14050 avdd.n11208 avss 0.0111f
C14051 avdd.n11209 avss 0.0148f
C14052 avdd.n11210 avss 0.0182f
C14053 avdd.n11211 avss -1.8e-19
C14054 avdd.n11212 avss -2.54e-19
C14055 avdd.n11213 avss -2.54e-19
C14056 avdd.n11214 avss -1.8e-19
C14057 avdd.n11215 avss -1.16e-19
C14058 avdd.n11216 avss -2.33e-19
C14059 avdd.n11217 avss 0.0342f
C14060 avdd.n11218 avss 0.0049f
C14061 avdd.n11219 avss -8.47e-19
C14062 avdd.n11220 avss -3.39e-19
C14063 avdd.n11221 avss -3.07e-19
C14064 avdd.n11222 avss -1.59e-19
C14065 avdd.n11223 avss -1.8e-19
C14066 avdd.n11224 avss 0.0192f
C14067 avdd.n11225 avss -1.59e-19
C14068 avdd.n11226 avss -1.8e-19
C14069 avdd.n11227 avss 0.00875f
C14070 avdd.n11228 avss 0.0111f
C14071 avdd.n11229 avss 0.0154f
C14072 avdd.n11230 avss 0.0183f
C14073 avdd.n11231 avss -1.8e-19
C14074 avdd.n11232 avss -2.22e-19
C14075 avdd.n11233 avss -2.22e-19
C14076 avdd.n11234 avss -1.8e-19
C14077 avdd.n11235 avss -2.01e-19
C14078 avdd.n11236 avss -3.18e-19
C14079 avdd.n11237 avss 0.03f
C14080 avdd.n11238 avss 0.00908f
C14081 avdd.n11239 avss -8.47e-19
C14082 avdd.n11240 avss -2.96e-19
C14083 avdd.n11241 avss -1.8e-19
C14084 avdd.n11242 avss -1.8e-19
C14085 avdd.n11243 avss 0.00873f
C14086 avdd.n11244 avss 0.0111f
C14087 avdd.n11245 avss 0.0154f
C14088 avdd.n11246 avss 0.0191f
C14089 avdd.n11247 avss -1.8e-19
C14090 avdd.n11248 avss 0.0184f
C14091 avdd.n11249 avss -1.38e-19
C14092 avdd.n11250 avss -1.8e-19
C14093 avdd.n11251 avss -2.44e-19
C14094 avdd.n11252 avss -2.44e-19
C14095 avdd.n11253 avss -1.8e-19
C14096 avdd.n11254 avss -1.38e-19
C14097 avdd.n11255 avss -3.49e-19
C14098 avdd.n11257 avss 0.0269f
C14099 avdd.n11258 avss 0.00869f
C14100 avdd.n11259 avss -0.00173f
C14101 avdd.n11260 avss -0.00512f
C14102 avdd.n11262 avss 0.0382f
C14103 avdd.n11263 avss -0.141f
C14104 avdd.n11264 avss -0.625f
C14105 avdd.n11265 avss -0.543f
C14106 avdd.n11266 avss -0.0512f
C14107 vinp.t18 avss 0.0241f
C14108 vinp.t67 avss 0.0219f
C14109 vinp.t15 avss 0.0182f
C14110 vinp.t10 avss 0.0182f
C14111 vinp.n0 avss 0.127f
C14112 vinp.t64 avss 0.0182f
C14113 vinp.t60 avss 0.0182f
C14114 vinp.n1 avss 0.128f
C14115 vinp.t14 avss 0.0182f
C14116 vinp.t17 avss 0.0182f
C14117 vinp.n2 avss 0.127f
C14118 vinp.t63 avss 0.0182f
C14119 vinp.t66 avss 0.0182f
C14120 vinp.n3 avss 0.128f
C14121 vinp.t13 avss 0.0182f
C14122 vinp.t19 avss 0.0182f
C14123 vinp.n4 avss 0.127f
C14124 vinp.t62 avss 0.0182f
C14125 vinp.t69 avss 0.0182f
C14126 vinp.n5 avss 0.128f
C14127 vinp.t16 avss 0.0182f
C14128 vinp.t12 avss 0.0182f
C14129 vinp.n6 avss 0.127f
C14130 vinp.t65 avss 0.0182f
C14131 vinp.t61 avss 0.0182f
C14132 vinp.n7 avss 0.128f
C14133 vinp.t11 avss 0.0241f
C14134 vinp.t68 avss 0.0219f
C14135 vinp.n8 avss 0.365f
C14136 vinp.n9 avss 0.107f
C14137 vinp.n10 avss 0.107f
C14138 vinp.n11 avss 0.107f
C14139 vinp.n12 avss 0.107f
C14140 vinp.n13 avss 0.382f
C14141 vinp.t50 avss 0.0241f
C14142 vinp.t46 avss 0.0219f
C14143 vinp.t57 avss 0.0182f
C14144 vinp.t53 avss 0.0182f
C14145 vinp.n14 avss 0.127f
C14146 vinp.t45 avss 0.0182f
C14147 vinp.t41 avss 0.0182f
C14148 vinp.n15 avss 0.128f
C14149 vinp.t56 avss 0.0182f
C14150 vinp.t52 avss 0.0182f
C14151 vinp.n16 avss 0.127f
C14152 vinp.t44 avss 0.0182f
C14153 vinp.t40 avss 0.0182f
C14154 vinp.n17 avss 0.128f
C14155 vinp.t55 avss 0.0182f
C14156 vinp.t51 avss 0.0182f
C14157 vinp.n18 avss 0.127f
C14158 vinp.t43 avss 0.0182f
C14159 vinp.t49 avss 0.0182f
C14160 vinp.n19 avss 0.128f
C14161 vinp.t58 avss 0.0182f
C14162 vinp.t59 avss 0.0182f
C14163 vinp.n20 avss 0.127f
C14164 vinp.t47 avss 0.0182f
C14165 vinp.t48 avss 0.0182f
C14166 vinp.n21 avss 0.128f
C14167 vinp.t54 avss 0.0241f
C14168 vinp.t42 avss 0.0219f
C14169 vinp.n22 avss 0.365f
C14170 vinp.n23 avss 0.107f
C14171 vinp.n24 avss 0.107f
C14172 vinp.n25 avss 0.107f
C14173 vinp.n26 avss 0.107f
C14174 vinp.n27 avss 0.381f
C14175 vinp.n28 avss 0.0807f
C14176 vinp.t70 avss 0.0241f
C14177 vinp.t30 avss 0.0219f
C14178 vinp.t73 avss 0.0182f
C14179 vinp.t75 avss 0.0182f
C14180 vinp.n29 avss 0.127f
C14181 vinp.t39 avss 0.0182f
C14182 vinp.t34 avss 0.0182f
C14183 vinp.n30 avss 0.128f
C14184 vinp.t79 avss 0.0182f
C14185 vinp.t77 avss 0.0182f
C14186 vinp.n31 avss 0.127f
C14187 vinp.t38 avss 0.0182f
C14188 vinp.t36 avss 0.0182f
C14189 vinp.n32 avss 0.128f
C14190 vinp.t76 avss 0.0182f
C14191 vinp.t72 avss 0.0182f
C14192 vinp.n33 avss 0.127f
C14193 vinp.t35 avss 0.0182f
C14194 vinp.t32 avss 0.0182f
C14195 vinp.n34 avss 0.128f
C14196 vinp.t74 avss 0.0182f
C14197 vinp.t71 avss 0.0182f
C14198 vinp.n35 avss 0.127f
C14199 vinp.t33 avss 0.0182f
C14200 vinp.t31 avss 0.0182f
C14201 vinp.n36 avss 0.128f
C14202 vinp.t78 avss 0.0241f
C14203 vinp.t37 avss 0.0219f
C14204 vinp.n37 avss 0.365f
C14205 vinp.n38 avss 0.107f
C14206 vinp.n39 avss 0.107f
C14207 vinp.n40 avss 0.107f
C14208 vinp.n41 avss 0.107f
C14209 vinp.n42 avss 0.381f
C14210 vinp.n43 avss 0.0817f
C14211 vinp.t28 avss 0.0241f
C14212 vinp.t6 avss 0.0219f
C14213 vinp.t25 avss 0.0182f
C14214 vinp.t20 avss 0.0182f
C14215 vinp.n44 avss 0.127f
C14216 vinp.t2 avss 0.0182f
C14217 vinp.t8 avss 0.0182f
C14218 vinp.n45 avss 0.128f
C14219 vinp.t24 avss 0.0182f
C14220 vinp.t29 avss 0.0182f
C14221 vinp.n46 avss 0.127f
C14222 vinp.t1 avss 0.0182f
C14223 vinp.t5 avss 0.0182f
C14224 vinp.n47 avss 0.128f
C14225 vinp.t23 avss 0.0182f
C14226 vinp.t27 avss 0.0182f
C14227 vinp.n48 avss 0.127f
C14228 vinp.t0 avss 0.0182f
C14229 vinp.t4 avss 0.0182f
C14230 vinp.n49 avss 0.128f
C14231 vinp.t22 avss 0.0182f
C14232 vinp.t26 avss 0.0182f
C14233 vinp.n50 avss 0.127f
C14234 vinp.t7 avss 0.0182f
C14235 vinp.t3 avss 0.0182f
C14236 vinp.n51 avss 0.128f
C14237 vinp.t21 avss 0.0241f
C14238 vinp.t9 avss 0.0219f
C14239 vinp.n52 avss 0.365f
C14240 vinp.n53 avss 0.107f
C14241 vinp.n54 avss 0.107f
C14242 vinp.n55 avss 0.107f
C14243 vinp.n56 avss 0.107f
C14244 vinp.n57 avss 0.38f
C14245 vinp.n58 avss 0.303f
C14246 vinp.n59 avss 0.559f
C14247 vinp.n60 avss 0.506f
C14248 vinp.n61 avss 0.394f
C14249 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t4 avss 0.459f
C14250 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t0 avss 0.00732f
C14251 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t2 avss 0.00732f
C14252 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n0 avss 0.0187f
C14253 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n1 avss 0.0323f
C14254 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t1 avss 0.00476f
C14255 dac_0.sky130_fd_sc_hd__inv_2_2.Y.t3 avss 0.00476f
C14256 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n2 avss 0.0113f
C14257 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n3 avss 0.00676f
C14258 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n4 avss 0.288f
C14259 dac_0.sky130_fd_sc_hd__inv_2_2.Y.n5 avss 0.211f
C14260 comparator_0.vp.t82 avss 0.908f
C14261 comparator_0.vp.t80 avss 3.09f
C14262 comparator_0.vp.t86 avss 3.87f
C14263 comparator_0.vp.t84 avss 0.584f
C14264 comparator_0.vp.n0 avss 0.0368f
C14265 comparator_0.vp.n1 avss 0.0358f
C14266 comparator_0.vp.n2 avss 0.0391f
C14267 comparator_0.vp.n3 avss 0.0368f
C14268 comparator_0.vp.n4 avss 0.0358f
C14269 comparator_0.vp.n5 avss 0.0391f
C14270 comparator_0.vp.n6 avss 0.0372f
C14271 comparator_0.vp.n7 avss 0.0336f
C14272 comparator_0.vp.n8 avss 0.0372f
C14273 comparator_0.vp.n9 avss 0.0336f
C14274 comparator_0.vp.t81 avss 0.955f
C14275 comparator_0.vp.t87 avss 0.955f
C14276 comparator_0.vp.t83 avss 0.955f
C14277 comparator_0.vp.t85 avss 0.0162f
C14278 comparator_0.vp.n10 avss 0.0848f
C14279 comparator_0.vp.t55 avss 0.00494f
C14280 comparator_0.vp.t51 avss 0.00494f
C14281 comparator_0.vp.n11 avss 0.0407f
C14282 comparator_0.vp.t40 avss 0.00494f
C14283 comparator_0.vp.t44 avss 0.00494f
C14284 comparator_0.vp.n12 avss 0.0347f
C14285 comparator_0.vp.t58 avss 0.00494f
C14286 comparator_0.vp.t50 avss 0.00494f
C14287 comparator_0.vp.n13 avss 0.0414f
C14288 comparator_0.vp.t59 avss 0.00494f
C14289 comparator_0.vp.t57 avss 0.00494f
C14290 comparator_0.vp.n14 avss 0.0384f
C14291 comparator_0.vp.t46 avss 0.00494f
C14292 comparator_0.vp.t41 avss 0.00494f
C14293 comparator_0.vp.n15 avss 0.0347f
C14294 comparator_0.vp.n16 avss 0.0299f
C14295 comparator_0.vp.t48 avss 0.00494f
C14296 comparator_0.vp.t47 avss 0.00494f
C14297 comparator_0.vp.n17 avss 0.0345f
C14298 comparator_0.vp.n18 avss 0.0358f
C14299 comparator_0.vp.t52 avss 0.00494f
C14300 comparator_0.vp.t54 avss 0.00494f
C14301 comparator_0.vp.n19 avss 0.0428f
C14302 comparator_0.vp.t42 avss 0.00494f
C14303 comparator_0.vp.t49 avss 0.00494f
C14304 comparator_0.vp.n20 avss 0.035f
C14305 comparator_0.vp.t53 avss 0.00494f
C14306 comparator_0.vp.t56 avss 0.00494f
C14307 comparator_0.vp.n21 avss 0.0426f
C14308 comparator_0.vp.t45 avss 0.00494f
C14309 comparator_0.vp.t43 avss 0.00494f
C14310 comparator_0.vp.n22 avss 0.035f
C14311 comparator_0.vp.t73 avss 0.00494f
C14312 comparator_0.vp.t71 avss 0.00494f
C14313 comparator_0.vp.n23 avss 0.0491f
C14314 comparator_0.vp.t32 avss 0.00494f
C14315 comparator_0.vp.t34 avss 0.00494f
C14316 comparator_0.vp.n24 avss 0.0347f
C14317 comparator_0.vp.t79 avss 0.00494f
C14318 comparator_0.vp.t74 avss 0.00494f
C14319 comparator_0.vp.n25 avss 0.0422f
C14320 comparator_0.vp.t76 avss 0.00494f
C14321 comparator_0.vp.t77 avss 0.00494f
C14322 comparator_0.vp.n26 avss 0.0407f
C14323 comparator_0.vp.t31 avss 0.00494f
C14324 comparator_0.vp.t30 avss 0.00494f
C14325 comparator_0.vp.n27 avss 0.0347f
C14326 comparator_0.vp.t70 avss 0.00494f
C14327 comparator_0.vp.t72 avss 0.00494f
C14328 comparator_0.vp.n28 avss 0.0407f
C14329 comparator_0.vp.t78 avss 0.00494f
C14330 comparator_0.vp.t75 avss 0.00494f
C14331 comparator_0.vp.n29 avss 0.0384f
C14332 comparator_0.vp.t36 avss 0.00494f
C14333 comparator_0.vp.t33 avss 0.00494f
C14334 comparator_0.vp.n30 avss 0.0347f
C14335 comparator_0.vp.n31 avss 0.0299f
C14336 comparator_0.vp.t38 avss 0.00494f
C14337 comparator_0.vp.t37 avss 0.00494f
C14338 comparator_0.vp.n32 avss 0.0341f
C14339 comparator_0.vp.n33 avss 0.037f
C14340 comparator_0.vp.n34 avss 0.0145f
C14341 comparator_0.vp.t39 avss 0.00494f
C14342 comparator_0.vp.t35 avss 0.00494f
C14343 comparator_0.vp.n35 avss 0.0461f
C14344 comparator_0.vp.n36 avss 0.0161f
C14345 comparator_0.vp.t20 avss 0.00494f
C14346 comparator_0.vp.t29 avss 0.00494f
C14347 comparator_0.vp.n37 avss 0.0407f
C14348 comparator_0.vp.t7 avss 0.00494f
C14349 comparator_0.vp.t3 avss 0.00494f
C14350 comparator_0.vp.n38 avss 0.0347f
C14351 comparator_0.vp.t22 avss 0.00494f
C14352 comparator_0.vp.t28 avss 0.00494f
C14353 comparator_0.vp.n39 avss 0.0414f
C14354 comparator_0.vp.t25 avss 0.00494f
C14355 comparator_0.vp.t23 avss 0.00494f
C14356 comparator_0.vp.n40 avss 0.0384f
C14357 comparator_0.vp.t8 avss 0.00494f
C14358 comparator_0.vp.t2 avss 0.00494f
C14359 comparator_0.vp.n41 avss 0.0347f
C14360 comparator_0.vp.n42 avss 0.0299f
C14361 comparator_0.vp.t0 avss 0.00494f
C14362 comparator_0.vp.t5 avss 0.00494f
C14363 comparator_0.vp.n43 avss 0.0345f
C14364 comparator_0.vp.n44 avss 0.0358f
C14365 comparator_0.vp.t26 avss 0.00494f
C14366 comparator_0.vp.t27 avss 0.00494f
C14367 comparator_0.vp.n45 avss 0.0428f
C14368 comparator_0.vp.t4 avss 0.00494f
C14369 comparator_0.vp.t6 avss 0.00494f
C14370 comparator_0.vp.n46 avss 0.035f
C14371 comparator_0.vp.t24 avss 0.00494f
C14372 comparator_0.vp.t21 avss 0.00494f
C14373 comparator_0.vp.n47 avss 0.0426f
C14374 comparator_0.vp.t9 avss 0.00494f
C14375 comparator_0.vp.t1 avss 0.00494f
C14376 comparator_0.vp.n48 avss 0.035f
C14377 comparator_0.vp.n49 avss 0.181f
C14378 comparator_0.vp.n50 avss 0.128f
C14379 comparator_0.vp.n51 avss 0.0731f
C14380 comparator_0.vp.t63 avss 0.00494f
C14381 comparator_0.vp.t61 avss 0.00494f
C14382 comparator_0.vp.n52 avss 0.0463f
C14383 comparator_0.vp.t62 avss 0.00494f
C14384 comparator_0.vp.t69 avss 0.00494f
C14385 comparator_0.vp.n53 avss 0.0347f
C14386 comparator_0.vp.t14 avss 0.00494f
C14387 comparator_0.vp.t19 avss 0.00494f
C14388 comparator_0.vp.n54 avss 0.0422f
C14389 comparator_0.vp.t13 avss 0.00494f
C14390 comparator_0.vp.t12 avss 0.00494f
C14391 comparator_0.vp.n55 avss 0.0407f
C14392 comparator_0.vp.t64 avss 0.00494f
C14393 comparator_0.vp.t65 avss 0.00494f
C14394 comparator_0.vp.n56 avss 0.0347f
C14395 comparator_0.vp.t11 avss 0.00494f
C14396 comparator_0.vp.t16 avss 0.00494f
C14397 comparator_0.vp.n57 avss 0.0407f
C14398 comparator_0.vp.t15 avss 0.00494f
C14399 comparator_0.vp.t18 avss 0.00494f
C14400 comparator_0.vp.n58 avss 0.0384f
C14401 comparator_0.vp.t68 avss 0.00494f
C14402 comparator_0.vp.t66 avss 0.00494f
C14403 comparator_0.vp.n59 avss 0.0347f
C14404 comparator_0.vp.n60 avss 0.0299f
C14405 comparator_0.vp.t60 avss 0.00494f
C14406 comparator_0.vp.t67 avss 0.00494f
C14407 comparator_0.vp.n61 avss 0.0341f
C14408 comparator_0.vp.n62 avss 0.037f
C14409 comparator_0.vp.t17 avss 0.00494f
C14410 comparator_0.vp.t10 avss 0.00494f
C14411 comparator_0.vp.n63 avss 0.0491f
C14412 comparator_0.vp.n64 avss 0.0153f
C14413 comparator_0.vp.n65 avss 0.0159f
.ends

