magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -36 101 36 107
rect -36 67 -17 101
rect -36 61 36 67
<< pwell >>
rect -124 -197 124 55
<< nmoslvt >>
rect -40 -171 40 29
<< ndiff >>
rect -98 14 -40 29
rect -98 -20 -86 14
rect -52 -20 -40 14
rect -98 -54 -40 -20
rect -98 -88 -86 -54
rect -52 -88 -40 -54
rect -98 -122 -40 -88
rect -98 -156 -86 -122
rect -52 -156 -40 -122
rect -98 -171 -40 -156
rect 40 14 98 29
rect 40 -20 52 14
rect 86 -20 98 14
rect 40 -54 98 -20
rect 40 -88 52 -54
rect 86 -88 98 -54
rect 40 -122 98 -88
rect 40 -156 52 -122
rect 86 -156 98 -122
rect 40 -171 98 -156
<< ndiffc >>
rect -86 -20 -52 14
rect -86 -88 -52 -54
rect -86 -156 -52 -122
rect 52 -20 86 14
rect 52 -88 86 -54
rect 52 -156 86 -122
<< poly >>
rect -40 101 40 117
rect -40 67 -17 101
rect 17 67 40 101
rect -40 29 40 67
rect -40 -197 40 -171
<< polycont >>
rect -17 67 17 101
<< locali >>
rect -40 67 -17 101
rect 17 67 40 101
rect -86 14 -52 33
rect -86 -54 -52 -52
rect -86 -90 -52 -88
rect -86 -175 -52 -156
rect 52 14 86 33
rect 52 -54 86 -52
rect 52 -90 86 -88
rect 52 -175 86 -156
<< viali >>
rect -17 67 17 101
rect -86 -20 -52 -18
rect -86 -52 -52 -20
rect -86 -122 -52 -90
rect -86 -124 -52 -122
rect 52 -20 86 -18
rect 52 -52 86 -20
rect 52 -122 86 -90
rect 52 -124 86 -122
<< metal1 >>
rect -36 101 36 107
rect -36 67 -17 101
rect 17 67 36 101
rect -36 61 36 67
rect -92 -18 -46 29
rect -92 -52 -86 -18
rect -52 -52 -46 -18
rect -92 -90 -46 -52
rect -92 -124 -86 -90
rect -52 -124 -46 -90
rect -92 -171 -46 -124
rect 46 -18 92 29
rect 46 -52 52 -18
rect 86 -52 92 -18
rect 46 -90 92 -52
rect 46 -124 52 -90
rect 86 -124 92 -90
rect 46 -171 92 -124
<< end >>
