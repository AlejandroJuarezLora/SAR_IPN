* NGSPICE file created from comp_temp.ext - technology: sky130B

.subckt comparator vn clk trim0 trim1 trim3 trimb0 trimb1 vp outp outn trim2 trimb4
+ trimb3 vdd trim4 trimb2 vss
X0 vdd clk outp sky130_fd_pr__pfet_01v8_2.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D trim3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X2 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X3 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 diff clk vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X6 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D trim0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X7 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 vss trimb3 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X9 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 vss trim4 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X12 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 IP vp diff vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X16 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trimb4 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X17 vss trimb1 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X18 vdd clk IN sky130_fd_pr__pfet_01v8_4.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X19 vdd outp outn sky130_fd_pr__pfet_01v8_1.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X20 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 outn outp IN vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X24 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 vss trimb2 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X28 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X38 vss trimb0 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X39 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 outp outn IP vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X41 diff clk vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X42 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 vdd outn outp sky130_fd_pr__pfet_01v8_0.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X47 IN vn diff vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X48 IN trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 vdd clk outn sky130_fd_pr__pfet_01v8_3.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X50 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 vdd clk IP sky130_fd_pr__pfet_01v8_5.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X53 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D IP sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

