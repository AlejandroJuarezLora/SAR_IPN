magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 1 117 185 163
rect 1 -19 718 117
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 196 7 226 91
rect 280 7 310 91
rect 442 7 472 91
rect 526 7 556 91
rect 610 7 640 91
<< scpmoshvt >>
rect 79 257 109 457
rect 459 373 489 457
rect 543 373 573 457
rect 627 373 657 457
rect 196 257 226 341
rect 268 257 298 341
<< ndiff >>
rect 27 89 79 137
rect 27 55 35 89
rect 69 55 79 89
rect 27 7 79 55
rect 109 91 159 137
rect 109 66 196 91
rect 109 32 119 66
rect 153 32 196 66
rect 109 7 196 32
rect 226 66 280 91
rect 226 32 236 66
rect 270 32 280 66
rect 226 7 280 32
rect 310 57 442 91
rect 310 23 320 57
rect 354 23 398 57
rect 432 23 442 57
rect 310 7 442 23
rect 472 66 526 91
rect 472 32 482 66
rect 516 32 526 66
rect 472 7 526 32
rect 556 7 610 91
rect 640 63 692 91
rect 640 29 650 63
rect 684 29 692 63
rect 640 7 692 29
<< pdiff >>
rect 27 418 79 457
rect 27 384 35 418
rect 69 384 79 418
rect 27 329 79 384
rect 27 295 35 329
rect 69 295 79 329
rect 27 257 79 295
rect 109 441 161 457
rect 109 407 119 441
rect 153 407 161 441
rect 109 341 161 407
rect 407 432 459 457
rect 407 398 415 432
rect 449 398 459 432
rect 407 373 459 398
rect 489 445 543 457
rect 489 411 499 445
rect 533 411 543 445
rect 489 373 543 411
rect 573 445 627 457
rect 573 411 583 445
rect 617 411 627 445
rect 573 373 627 411
rect 657 432 709 457
rect 657 398 667 432
rect 701 398 709 432
rect 657 373 709 398
rect 109 257 196 341
rect 226 257 268 341
rect 298 319 351 341
rect 298 285 308 319
rect 342 285 351 319
rect 298 257 351 285
<< ndiffc >>
rect 35 55 69 89
rect 119 32 153 66
rect 236 32 270 66
rect 320 23 354 57
rect 398 23 432 57
rect 482 32 516 66
rect 650 29 684 63
<< pdiffc >>
rect 35 384 69 418
rect 35 295 69 329
rect 119 407 153 441
rect 415 398 449 432
rect 499 411 533 445
rect 583 411 617 445
rect 667 398 701 432
rect 308 285 342 319
<< poly >>
rect 79 457 109 483
rect 459 457 489 483
rect 543 457 573 483
rect 627 457 657 483
rect 196 341 226 367
rect 268 341 298 367
rect 459 341 489 373
rect 442 311 489 341
rect 79 225 109 257
rect 196 225 226 257
rect 76 209 130 225
rect 76 175 86 209
rect 120 175 130 209
rect 76 159 130 175
rect 172 209 226 225
rect 172 175 182 209
rect 216 175 226 209
rect 268 235 298 257
rect 442 247 472 311
rect 543 287 573 373
rect 268 225 310 235
rect 268 209 326 225
rect 268 202 282 209
rect 172 159 226 175
rect 272 175 282 202
rect 316 175 326 209
rect 272 159 326 175
rect 368 191 472 247
rect 79 137 109 159
rect 196 91 226 159
rect 280 91 310 159
rect 368 157 378 191
rect 412 157 472 191
rect 368 113 472 157
rect 442 91 472 113
rect 526 271 580 287
rect 526 237 536 271
rect 570 237 580 271
rect 526 221 580 237
rect 627 225 657 373
rect 526 91 556 221
rect 627 209 700 225
rect 627 189 656 209
rect 610 175 656 189
rect 690 175 700 209
rect 610 159 700 175
rect 610 91 640 159
rect 79 -19 109 7
rect 196 -19 226 7
rect 280 -19 310 7
rect 442 -19 472 7
rect 526 -19 556 7
rect 610 -19 640 7
<< polycont >>
rect 86 175 120 209
rect 182 175 216 209
rect 282 175 316 209
rect 378 157 412 191
rect 536 237 570 271
rect 656 175 690 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 17 418 69 453
rect 17 384 35 418
rect 103 441 169 487
rect 103 407 119 441
rect 153 407 169 441
rect 398 434 449 453
rect 583 445 633 487
rect 221 432 449 434
rect 17 329 69 384
rect 221 400 415 432
rect 221 355 255 400
rect 17 295 35 329
rect 17 265 69 295
rect 103 321 255 355
rect 398 398 415 400
rect 483 411 499 445
rect 533 411 549 445
rect 398 373 449 398
rect 17 122 52 265
rect 103 225 137 321
rect 308 319 342 341
rect 398 339 480 373
rect 342 285 412 303
rect 86 209 137 225
rect 120 175 137 209
rect 86 159 137 175
rect 182 209 248 283
rect 308 269 412 285
rect 216 175 248 209
rect 182 159 248 175
rect 282 209 340 235
rect 316 175 340 209
rect 282 159 340 175
rect 378 191 412 269
rect 378 125 412 157
rect 17 89 69 122
rect 17 55 35 89
rect 236 91 412 125
rect 446 134 480 339
rect 515 361 549 411
rect 617 411 633 445
rect 583 395 633 411
rect 667 432 703 453
rect 701 398 703 432
rect 667 361 703 398
rect 515 327 703 361
rect 520 271 616 291
rect 520 237 536 271
rect 570 237 616 271
rect 520 231 616 237
rect 446 100 516 134
rect 564 113 616 231
rect 656 209 708 291
rect 690 175 708 209
rect 656 113 708 175
rect 236 66 270 91
rect 17 11 69 55
rect 103 32 119 66
rect 153 32 189 66
rect 103 -23 189 32
rect 482 66 516 100
rect 236 11 270 32
rect 304 23 320 57
rect 354 23 398 57
rect 432 23 448 57
rect 304 -23 448 23
rect 482 11 516 32
rect 631 63 711 79
rect 631 29 650 63
rect 684 29 711 63
rect 631 -23 711 29
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a2bb2o_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel locali s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel locali s 674 181 708 215 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 674 249 708 283 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 674 113 708 147 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A1_N
port 10 nsew
flabel locali s 306 181 340 215 0 FreeSans 200 0 0 0 A2_N
port 9 nsew
flabel locali s 30 45 64 79 0 FreeSans 200 0 0 0 X
port 11 nsew
flabel locali s 582 249 616 283 0 FreeSans 200 0 0 0 B2
port 8 nsew
flabel locali s 214 249 248 283 0 FreeSans 200 0 0 0 A1_N
port 10 nsew
flabel locali s 30 385 64 419 0 FreeSans 200 0 0 0 X
port 11 nsew
flabel locali s 30 317 64 351 0 FreeSans 200 0 0 0 X
port 11 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
