magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 222 542
<< pwell >>
rect 31 -50 63 -28
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 184 521
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 184 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 29 -57 63 -23
rect 121 -57 155 -23
<< metal1 >>
rect 0 521 184 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 184 521
rect 0 456 184 487
rect 0 -23 184 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 184 -23
rect 0 -88 184 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 fill_2
flabel metal1 s 20 -54 73 -22 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 21 490 73 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 28 495 62 513 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 31 -50 63 -28 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 184 504
string path 0.000 -1.000 4.600 -1.000 
<< end >>
