* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt M2_1 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n109# a_n98_n109# 0.104f
C1 a_n40_n197# a_n98_n109# 0.0145f
C2 a_n40_n197# a_40_n109# 0.0145f
C3 a_40_n109# VSUBS 0.122f
C4 a_n98_n109# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt M2_inv a_n40_n201# a_40_n104# w_n236_n324# a_n98_n104# VSUBS
X0 a_40_n104# a_n40_n201# a_n98_n104# w_n236_n324# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_n98_n104# a_40_n104# 0.104f
C1 a_n98_n104# a_n40_n201# 0.0145f
C2 w_n236_n324# a_40_n104# 0.0219f
C3 w_n236_n324# a_n40_n201# 0.12f
C4 a_40_n104# a_n40_n201# 0.0145f
C5 w_n236_n324# a_n98_n104# 0.0219f
C6 a_40_n104# VSUBS 0.1f
C7 a_n98_n104# VSUBS 0.1f
C8 a_n40_n201# VSUBS 0.146f
C9 w_n236_n324# VSUBS 0.804f
.ends

.subckt M1_inv a_40_n171# a_n40_n197# a_n98_n171# VSUBS
X0 a_40_n171# a_n40_n197# a_n98_n171# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n171# a_n98_n171# 0.104f
C1 a_n40_n197# a_n98_n171# 0.0145f
C2 a_n40_n197# a_40_n171# 0.0145f
C3 a_40_n171# VSUBS 0.122f
C4 a_n98_n171# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt inv_lvt M2_inv_0/a_n98_n104# M2_inv_0/w_n236_n324# M1_inv_0/a_n98_n171# m1_170_505#
+ m2_289_257# VSUBS
XM2_inv_0 m1_170_505# m2_289_257# M2_inv_0/w_n236_n324# M2_inv_0/a_n98_n104# VSUBS
+ M2_inv
XM1_inv_0 m2_289_257# m1_170_505# M1_inv_0/a_n98_n171# VSUBS M1_inv
C0 M2_inv_0/a_n98_n104# m2_289_257# 0.00845f
C1 M1_inv_0/a_n98_n171# M2_inv_0/w_n236_n324# 0.00225f
C2 M2_inv_0/a_n98_n104# m1_170_505# 0.0037f
C3 M1_inv_0/a_n98_n171# m2_289_257# 0.00845f
C4 M1_inv_0/a_n98_n171# m1_170_505# 0.00383f
C5 M2_inv_0/w_n236_n324# m2_289_257# 0.055f
C6 M2_inv_0/w_n236_n324# m1_170_505# 0.0237f
C7 M1_inv_0/a_n98_n171# M2_inv_0/a_n98_n104# 0.00387f
C8 m2_289_257# m1_170_505# 0.153f
C9 M2_inv_0/w_n236_n324# M2_inv_0/a_n98_n104# -1.52e-20
C10 M1_inv_0/a_n98_n171# VSUBS 0.122f
C11 m2_289_257# VSUBS 0.582f
C12 M2_inv_0/a_n98_n104# VSUBS 0.1f
C13 m1_170_505# VSUBS 0.453f
C14 M2_inv_0/w_n236_n324# VSUBS 0.804f
.ends

.subckt M1_2 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_n98_n109# a_n40_n197# 0.0145f
C1 a_40_n109# a_n98_n109# 0.104f
C2 a_40_n109# a_n40_n197# 0.0145f
C3 a_40_n109# VSUBS 0.122f
C4 a_n98_n109# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt latch vdd Qn S R Q m1_458_623# m1_1673_493# vss
XM2_1_0 vss m1_1673_493# Q vss M2_1
Xinv_lvt_0 vdd vdd vss R m1_1673_493# vss inv_lvt
Xinv_lvt_1 vdd vdd vss S m1_458_623# vss inv_lvt
Xinv_lvt_2 vdd vdd vss Qn Q vss inv_lvt
Xinv_lvt_3 vdd vdd vss Q Qn vss inv_lvt
XM1_2_0 Qn m1_458_623# vss vss M1_2
C0 S Q 1.46e-19
C1 m1_458_623# Qn 0.104f
C2 m1_1673_493# Qn 0.0703f
C3 m1_458_623# Q 0.0703f
C4 m1_1673_493# Q 0.104f
C5 R Q 0.0155f
C6 vdd Qn 0.221f
C7 m1_458_623# S 0.0354f
C8 vdd Q 0.528f
C9 vdd S 0.161f
C10 R m1_1673_493# 0.0354f
C11 vdd m1_458_623# 0.214f
C12 vdd m1_1673_493# 0.215f
C13 vdd R 0.159f
C14 Q Qn 0.655f
C15 S Qn 0.0154f
C16 Qn vss 0.899f
C17 Q vss 0.835f
C18 m1_458_623# vss 0.689f
C19 S vss 0.48f
C20 m1_1673_493# vss 0.686f
C21 R vss 0.479f
C22 vdd vss 7.03f
.ends

.subckt inv2 w_0_269# a_67_305# a_59_207# a_149_55# a_67_55# VSUBS
X0 a_67_55# a_59_207# a_149_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_149_55# a_59_207# a_67_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_67_305# a_59_207# a_149_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_149_55# a_59_207# a_67_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 a_67_305# a_67_55# 0.0423f
C1 a_67_305# w_0_269# 0.0521f
C2 w_0_269# a_67_55# 0.00649f
C3 a_149_55# a_67_55# 0.155f
C4 a_67_305# a_149_55# 0.209f
C5 a_149_55# w_0_269# 0.0061f
C6 a_67_305# a_59_207# 0.0631f
C7 a_59_207# a_67_55# 0.0638f
C8 a_59_207# w_0_269# 0.0742f
C9 a_59_207# a_149_55# 0.0894f
C10 a_67_55# VSUBS 0.266f
C11 a_149_55# VSUBS 0.0332f
C12 a_67_305# VSUBS 0.246f
C13 a_59_207# VSUBS 0.263f
C14 w_0_269# VSUBS 0.339f
.ends

.subckt decap_8 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=2.89
C0 w_0_269# a_65_331# 0.105f
C1 a_65_331# a_65_55# 1.27f
C2 w_0_269# a_65_55# 0.22f
C3 a_65_331# VSUBS 1.14f
C4 a_65_55# VSUBS 0.992f
C5 w_0_269# VSUBS 0.782f
.ends

.subckt M1_3 a_207_n176# a_n29_n176# a_26_55# a_n328_55# a_89_n176# a_n446_55# a_n564_55#
+ a_n210_55# a_n501_n176# a_561_n176# a_n383_n176# a_498_55# a_144_55# a_443_n176#
+ a_n265_n176# a_262_55# a_380_55# a_n619_n176# a_n92_55# w_n757_n324# a_325_n176#
+ a_n147_n176# VSUBS
X0 a_n383_n176# a_n446_55# a_n501_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n29_n176# a_n92_55# a_n147_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_325_n176# a_262_55# a_207_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_561_n176# a_498_55# a_443_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X4 a_n265_n176# a_n328_55# a_n383_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_89_n176# a_26_55# a_n29_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_207_n176# a_144_55# a_89_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_n501_n176# a_n564_55# a_n619_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X8 a_n147_n176# a_n210_55# a_n265_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_443_n176# a_380_55# a_325_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
C0 a_207_n176# a_325_n176# 0.121f
C1 a_n501_n176# a_n446_55# 0.0116f
C2 a_n265_n176# a_n383_n176# 0.121f
C3 a_26_55# w_n757_n324# 0.105f
C4 a_n92_55# a_n210_55# 0.0657f
C5 a_89_n176# a_207_n176# 0.121f
C6 a_n383_n176# a_n501_n176# 0.121f
C7 a_n92_55# a_n29_n176# 0.0116f
C8 a_n265_n176# w_n757_n324# 0.0274f
C9 a_n210_55# a_n328_55# 0.0657f
C10 a_n501_n176# w_n757_n324# 0.0247f
C11 w_n757_n324# a_262_55# 0.104f
C12 a_443_n176# a_561_n176# 0.121f
C13 a_n619_n176# a_n564_55# 0.0116f
C14 a_207_n176# w_n757_n324# 0.0274f
C15 a_325_n176# a_443_n176# 0.121f
C16 a_498_55# a_561_n176# 0.0116f
C17 a_144_55# a_89_n176# 0.0116f
C18 a_498_55# a_443_n176# 0.0116f
C19 a_n92_55# a_26_55# 0.0657f
C20 a_n265_n176# a_n328_55# 0.0116f
C21 a_380_55# a_262_55# 0.0657f
C22 a_26_55# a_n29_n176# 0.0116f
C23 a_144_55# w_n757_n324# 0.104f
C24 a_n265_n176# a_n210_55# 0.0116f
C25 a_n501_n176# a_n564_55# 0.0116f
C26 w_n757_n324# a_561_n176# 0.0913f
C27 w_n757_n324# a_443_n176# 0.0247f
C28 w_n757_n324# a_325_n176# 0.0258f
C29 a_n383_n176# a_n446_55# 0.0116f
C30 w_n757_n324# a_498_55# 0.13f
C31 a_n147_n176# w_n757_n324# 0.0258f
C32 a_n619_n176# a_n501_n176# 0.121f
C33 a_89_n176# w_n757_n324# 0.0258f
C34 w_n757_n324# a_n446_55# 0.105f
C35 a_n383_n176# w_n757_n324# 0.0258f
C36 a_380_55# a_443_n176# 0.0116f
C37 a_380_55# a_325_n176# 0.0116f
C38 a_n92_55# a_n147_n176# 0.0116f
C39 a_380_55# a_498_55# 0.0657f
C40 a_n210_55# a_n147_n176# 0.0116f
C41 a_207_n176# a_262_55# 0.0116f
C42 a_n147_n176# a_n29_n176# 0.121f
C43 a_n446_55# a_n564_55# 0.0657f
C44 a_n328_55# a_n446_55# 0.0657f
C45 a_89_n176# a_n29_n176# 0.121f
C46 a_144_55# a_26_55# 0.0657f
C47 a_n92_55# w_n757_n324# 0.105f
C48 a_n383_n176# a_n328_55# 0.0116f
C49 a_380_55# w_n757_n324# 0.105f
C50 w_n757_n324# a_n564_55# 0.13f
C51 a_n328_55# w_n757_n324# 0.104f
C52 a_144_55# a_262_55# 0.0657f
C53 a_n210_55# w_n757_n324# 0.104f
C54 w_n757_n324# a_n29_n176# 0.0238f
C55 a_n265_n176# a_n147_n176# 0.121f
C56 a_144_55# a_207_n176# 0.0116f
C57 a_89_n176# a_26_55# 0.0116f
C58 a_n619_n176# w_n757_n324# 0.0913f
C59 a_262_55# a_325_n176# 0.0116f
C60 a_561_n176# VSUBS 0.056f
C61 a_443_n176# VSUBS 0.0249f
C62 a_325_n176# VSUBS 0.0249f
C63 a_207_n176# VSUBS 0.0249f
C64 a_89_n176# VSUBS 0.0249f
C65 a_n29_n176# VSUBS 0.0249f
C66 a_n147_n176# VSUBS 0.0249f
C67 a_n265_n176# VSUBS 0.0249f
C68 a_n383_n176# VSUBS 0.0249f
C69 a_n501_n176# VSUBS 0.0249f
C70 a_n619_n176# VSUBS 0.056f
C71 a_498_55# VSUBS 0.0832f
C72 a_380_55# VSUBS 0.0669f
C73 a_262_55# VSUBS 0.0669f
C74 a_144_55# VSUBS 0.0669f
C75 a_26_55# VSUBS 0.0669f
C76 a_n92_55# VSUBS 0.0669f
C77 a_n210_55# VSUBS 0.0669f
C78 a_n328_55# VSUBS 0.0669f
C79 a_n446_55# VSUBS 0.0669f
C80 a_n564_55# VSUBS 0.0832f
C81 w_n757_n324# VSUBS 3.39f
.ends

.subckt M2_2 a_26_51# a_89_n171# a_n328_51# a_n446_51# a_n564_51# a_n501_n171# a_n210_51#
+ a_561_n171# a_n383_n171# a_498_51# a_443_n171# a_144_51# a_n265_n171# a_262_51#
+ a_n619_n171# a_380_51# a_n92_51# a_n721_n283# a_325_n171# a_n147_n171# a_207_n171#
+ a_n29_n171#
X0 a_89_n171# a_26_51# a_n29_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_207_n171# a_144_51# a_89_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n147_n171# a_n210_51# a_n265_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_n501_n171# a_n564_51# a_n619_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X4 a_443_n171# a_380_51# a_325_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n383_n171# a_n446_51# a_n501_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_n29_n171# a_n92_51# a_n147_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_325_n171# a_262_51# a_207_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_561_n171# a_498_51# a_443_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X9 a_n265_n171# a_n328_51# a_n383_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
C0 a_n29_n171# a_89_n171# 0.121f
C1 a_n328_51# a_n210_51# 0.0633f
C2 a_n265_n171# a_n147_n171# 0.121f
C3 a_n446_51# a_n383_n171# 0.0116f
C4 a_325_n171# a_380_51# 0.0116f
C5 a_498_51# a_443_n171# 0.0116f
C6 a_n446_51# a_n328_51# 0.0633f
C7 a_561_n171# a_498_51# 0.0116f
C8 a_n265_n171# a_n383_n171# 0.121f
C9 a_144_51# a_89_n171# 0.0116f
C10 a_561_n171# a_443_n171# 0.121f
C11 a_n265_n171# a_n328_51# 0.0116f
C12 a_n92_51# a_26_51# 0.0633f
C13 a_n210_51# a_n92_51# 0.0633f
C14 a_n501_n171# a_n564_51# 0.0116f
C15 a_262_51# a_325_n171# 0.0116f
C16 a_144_51# a_207_n171# 0.0116f
C17 a_498_51# a_380_51# 0.0633f
C18 a_n265_n171# a_n210_51# 0.0116f
C19 a_n29_n171# a_n147_n171# 0.121f
C20 a_443_n171# a_380_51# 0.0116f
C21 a_89_n171# a_26_51# 0.0116f
C22 a_n501_n171# a_n383_n171# 0.121f
C23 a_262_51# a_207_n171# 0.0116f
C24 a_n383_n171# a_n328_51# 0.0116f
C25 a_n29_n171# a_26_51# 0.0116f
C26 a_n564_51# a_n619_n171# 0.0116f
C27 a_n29_n171# a_n92_51# 0.0116f
C28 a_325_n171# a_207_n171# 0.121f
C29 a_443_n171# a_325_n171# 0.121f
C30 a_n501_n171# a_n619_n171# 0.121f
C31 a_n446_51# a_n564_51# 0.0633f
C32 a_n501_n171# a_n446_51# 0.0116f
C33 a_262_51# a_144_51# 0.0633f
C34 a_n147_n171# a_n92_51# 0.0116f
C35 a_n147_n171# a_n210_51# 0.0116f
C36 a_144_51# a_26_51# 0.0633f
C37 a_89_n171# a_207_n171# 0.121f
C38 a_262_51# a_380_51# 0.0633f
C39 a_561_n171# a_n721_n283# 0.148f
C40 a_443_n171# a_n721_n283# 0.0499f
C41 a_325_n171# a_n721_n283# 0.051f
C42 a_207_n171# a_n721_n283# 0.0526f
C43 a_89_n171# a_n721_n283# 0.051f
C44 a_n29_n171# a_n721_n283# 0.0489f
C45 a_n147_n171# a_n721_n283# 0.051f
C46 a_n265_n171# a_n721_n283# 0.0526f
C47 a_n383_n171# a_n721_n283# 0.051f
C48 a_n501_n171# a_n721_n283# 0.0499f
C49 a_n619_n171# a_n721_n283# 0.148f
C50 a_498_51# a_n721_n283# 0.208f
C51 a_380_51# a_n721_n283# 0.169f
C52 a_262_51# a_n721_n283# 0.168f
C53 a_144_51# a_n721_n283# 0.168f
C54 a_26_51# a_n721_n283# 0.169f
C55 a_n92_51# a_n721_n283# 0.169f
C56 a_n210_51# a_n721_n283# 0.168f
C57 a_n328_51# a_n721_n283# 0.168f
C58 a_n446_51# a_n721_n283# 0.169f
C59 a_n564_51# a_n721_n283# 0.208f
.ends

.subckt inv_4 w_0_269# a_59_207# a_75_55# a_75_305# a_157_55# VSUBS
X0 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 a_157_55# a_59_207# 0.36f
C1 a_75_55# a_59_207# 0.0819f
C2 a_75_55# a_157_55# 0.263f
C3 w_0_269# a_75_305# 0.0654f
C4 a_75_305# a_59_207# 0.0982f
C5 a_157_55# a_75_305# 0.362f
C6 a_75_55# a_75_305# 0.0501f
C7 w_0_269# a_59_207# 0.142f
C8 a_157_55# w_0_269# 0.0159f
C9 a_75_55# w_0_269# 0.00667f
C10 a_75_55# VSUBS 0.327f
C11 a_157_55# VSUBS 0.0849f
C12 a_75_305# VSUBS 0.296f
C13 a_59_207# VSUBS 0.452f
C14 w_0_269# VSUBS 0.516f
.ends

.subckt decap_3 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=0.59
C0 w_0_269# a_65_331# 0.0625f
C1 a_65_55# w_0_269# 0.0797f
C2 a_65_55# a_65_331# 0.353f
C3 a_65_331# VSUBS 0.47f
C4 a_65_55# VSUBS 0.427f
C5 w_0_269# VSUBS 0.339f
.ends

.subckt sw_top en m2_1158_361# inv_4_1/w_0_269# out vdd in m2_990_200# vss
Xdecap_8_0 vss vdd inv_4_1/w_0_269# vss decap_8
XM1_3_0 out out m2_1158_361# m2_1158_361# in m2_1158_361# m2_1158_361# m2_1158_361#
+ out in in m2_1158_361# m2_1158_361# out out m2_1158_361# m2_1158_361# in m2_1158_361#
+ vdd in in vss M1_3
XM2_2_0 m2_990_200# in m2_990_200# m2_990_200# m2_990_200# out m2_990_200# in in m2_990_200#
+ out m2_990_200# out m2_990_200# in m2_990_200# m2_990_200# vss in in out out M2_2
Xinv_4_0 inv_4_1/w_0_269# m2_1158_361# vss vdd m2_990_200# vss inv_4
Xinv_4_1 inv_4_1/w_0_269# en vss vdd m2_1158_361# vss inv_4
Xdecap_3_0 vss vdd inv_4_1/w_0_269# vss decap_3
C0 m2_1158_361# vdd 0.548f
C1 m2_1158_361# in 0.366f
C2 inv_4_1/w_0_269# en 0.00756f
C3 m2_990_200# en 0.081f
C4 out vdd 0.251f
C5 in out 3.36f
C6 m2_1158_361# en 0.0497f
C7 inv_4_1/w_0_269# m2_990_200# 0.0362f
C8 in vdd 0.441f
C9 m2_1158_361# inv_4_1/w_0_269# 0.0273f
C10 out en 0.00104f
C11 m2_1158_361# m2_990_200# 0.495f
C12 vdd en 0.0781f
C13 in en 0.0114f
C14 out m2_990_200# 0.172f
C15 inv_4_1/w_0_269# vdd -0.0142f
C16 m2_1158_361# out 0.375f
C17 inv_4_1/w_0_269# in 0.00475f
C18 m2_990_200# vdd 0.418f
C19 in m2_990_200# 0.276f
C20 en vss 0.653f
C21 vdd vss 5.79f
C22 m2_990_200# vss 2.13f
C23 out vss 0.745f
C24 in vss 1.61f
C25 m2_1158_361# vss 1.84f
C26 inv_4_1/w_0_269# vss 1.95f
.ends

.subckt C7 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt DUMMY m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C6 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt CDUM m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C4 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C2 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C5 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C3 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C1 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt C0_1 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n250_n240# m3_n450_n340# 0.503f
C1 c1_n250_n240# VSUBS 0.213f
C2 m3_n450_n340# VSUBS 0.722f
.ends

.subckt carray n2 n3 via23_4_702/m2_1_40# m3_12800_1156# m3_23200_1156# m3_28400_1156#
+ m2_800_1156# m2_19000_1156# via23_4_584/m2_1_40# via23_4_331/m2_1_40# m3_6100_1156#
+ via23_4_213/m2_1_40# m3_24500_1156# m3_29700_1156# m2_15100_1156# via23_4_347/m2_1_40#
+ via23_4_326/m2_1_40# m3_2200_1156# via23_4_459/m2_1_40# m3_7400_1156# via23_4_354/m2_1_40#
+ m3_25800_1156# m3_31000_1156# m2_11200_1156# m3_36200_1156# m2_16400_1156# via23_4_250/m2_1_40#
+ m2_27200_1156# via23_4_710/m2_1_40# m3_3500_1156# via23_4_601/m2_1_40# m3_8700_1156#
+ via23_4_709/m2_1_40# m3_32300_1156# m2_12500_1156# m3_37500_1156# m2_17700_1156#
+ via23_4_198/m2_1_40# m2_23300_1156# m2_28500_1156# m3_4800_1156# via23_4_230/m2_1_40#
+ m3_33600_1156# m2_13800_1156# m3_38800_1156# via23_4_447/m2_1_40# via23_4_598/m2_1_40#
+ via23_4_676/m2_1_40# m3_19100_1156# m2_24600_1156# m2_29800_1156# m2_35000_1156#
+ m3_34900_1156# m3_40100_1156# m2_20300_1156# m3_10000_1156# via23_4_332/m2_1_40#
+ m3_15200_1156# m2_31100_1156# m2_25900_1156# via23_4_369/m2_1_40# m2_36300_1156#
+ via23_4_590/m2_1_40# m3_41400_1156# via23_4_379/m2_1_40# via23_4_220/m2_1_40# m3_11300_1156#
+ m3_16500_1156# m2_32400_1156# m2_37600_1156# via23_4_251/m2_1_40# m3_42700_1156#
+ via23_4_711/m2_1_40# via23_4_675/m2_1_40# m3_12600_1156# via23_4_345/m2_1_40# m3_17800_1156#
+ m3_28200_1156# m2_33700_1156# m3_5000_1156# m2_38900_1156# m3_900_1156# via23_4_635/m2_1_40#
+ via23_4_455/m2_1_40# via23_4_588/m2_1_40# m3_13900_1156# via23_4_414/m2_1_40# m3_24300_1156#
+ via23_4_439/m2_1_40# m2_40200_1156# m3_1100_1156# m3_29500_1156# via23_4_460/m2_1_40#
+ via23_4_218/m2_1_40# m3_6300_1156# via23_4_704/m2_1_40# via23_4_599/m2_1_40# via23_4_677/m2_1_40#
+ via23_4_249/m2_1_40# m3_20400_1156# m3_2400_1156# m3_25600_1156# m3_36000_1156#
+ m2_41500_1156# m3_7600_1156# via23_4_333/m2_1_40# via23_4_366/m2_1_40# m3_26900_1156#
+ m3_32100_1156# via23_4_429/m2_1_40# m2_42800_1156# m3_3700_1156# m3_37300_1156#
+ m3_8900_1156# m2_6000_1156# via23_4_128/m2_1_40# via23_4_458/m2_1_40# via23_4_199/m2_1_40#
+ ndum via23_4_381/m2_1_40# m3_18000_1156# n0 via23_4_419/m2_1_40# m3_33400_1156#
+ m3_38600_1156# m2_2100_1156# m2_7300_1156# via23_4_449/m2_1_40# via23_4_200/m2_1_40#
+ via23_4_712/m2_1_40# via23_4_346/m2_1_40# m3_14100_1156# n4 m3_19300_1156# via23_4_228/m2_1_40#
+ via23_4_641/m2_1_40# via23_4_378/m2_1_40# m3_34700_1156# m3_39900_1156# n1 m2_3400_1156#
+ via23_4_589/m2_1_40# n6 m2_8600_1156# m3_10200_1156# via23_4_642/m2_1_40# via23_4_245/m2_1_40#
+ m3_15400_1156# via23_4_368/m2_1_40# via23_4_705/m2_1_40# via23_4_446/m2_1_40# m3_30800_1156#
+ via23_4_678/m2_1_40# via23_4_600/m2_1_40# m3_41200_1156# m2_4700_1156# via23_4_96/m2_1_40#
+ m2_9900_1156# n5 m3_11500_1156# m3_16700_1156# via23_4_448/m2_1_40# m3_27100_1156#
+ via23_4_334/m2_1_40# m3_42500_1156# VSUBS via23_4_380/m2_1_40# top via23_4_229/m2_1_40#
+ n7 via23_4_367/m2_1_40#
XC7_121 n7 top VSUBS C7
XC7_110 n7 top VSUBS C7
XDUMMY_80 via23_4_712/m2_1_40# top VSUBS DUMMY
XC6_20 n6 top VSUBS C6
XC6_53 n6 top VSUBS C6
XC6_31 n6 top VSUBS C6
XC6_42 n6 top VSUBS C6
XC7_122 n7 top VSUBS C7
XC7_100 n7 top VSUBS C7
XC7_111 n7 top VSUBS C7
XDUMMY_81 via23_4_709/m2_1_40# top VSUBS DUMMY
XDUMMY_70 via23_4_642/m2_1_40# top VSUBS DUMMY
XC6_21 n6 top VSUBS C6
XC6_10 n6 top VSUBS C6
XC6_54 n6 top VSUBS C6
XC6_32 n6 top VSUBS C6
XC6_43 n6 top VSUBS C6
XC6_0 n6 top VSUBS C6
XC7_123 n7 top VSUBS C7
XC7_101 n7 top VSUBS C7
XC7_112 n7 top VSUBS C7
XDUMMY_71 via23_4_641/m2_1_40# top VSUBS DUMMY
XDUMMY_82 via23_4_439/m2_1_40# top VSUBS DUMMY
XDUMMY_60 via23_4_448/m2_1_40# top VSUBS DUMMY
XC6_44 n6 top VSUBS C6
XC6_22 n6 top VSUBS C6
XC6_55 n6 top VSUBS C6
XC6_11 n6 top VSUBS C6
XC6_33 n6 top VSUBS C6
XC6_1 n6 top VSUBS C6
XC7_124 n7 top VSUBS C7
XC7_102 n7 top VSUBS C7
XC7_113 n7 top VSUBS C7
XDUMMY_72 via23_4_676/m2_1_40# top VSUBS DUMMY
XDUMMY_83 via23_4_675/m2_1_40# top VSUBS DUMMY
XDUMMY_61 via23_4_588/m2_1_40# top VSUBS DUMMY
XDUMMY_50 via23_4_429/m2_1_40# top VSUBS DUMMY
XC6_56 n6 top VSUBS C6
XC6_12 n6 top VSUBS C6
XC6_45 n6 top VSUBS C6
XC6_23 n6 top VSUBS C6
XC6_34 n6 top VSUBS C6
XC6_2 n6 top VSUBS C6
XCDUM_0 ndum top VSUBS CDUM
XC7_103 n7 top VSUBS C7
XC7_125 n7 top VSUBS C7
XC7_114 n7 top VSUBS C7
XDUMMY_73 via23_4_677/m2_1_40# top VSUBS DUMMY
XDUMMY_62 via23_4_589/m2_1_40# top VSUBS DUMMY
XDUMMY_40 via23_4_326/m2_1_40# top VSUBS DUMMY
XDUMMY_51 via23_4_414/m2_1_40# top VSUBS DUMMY
XC6_57 n6 top VSUBS C6
XC6_24 n6 top VSUBS C6
XC6_46 n6 top VSUBS C6
XC6_13 n6 top VSUBS C6
XC6_35 n6 top VSUBS C6
XDUMMY_0 via23_4_3/m2_1_40# top VSUBS DUMMY
XC6_3 n6 top VSUBS C6
XC4_0 n4 top VSUBS C4
XC7_104 n7 top VSUBS C7
XC7_115 n7 top VSUBS C7
XC7_126 n7 top VSUBS C7
XDUMMY_74 via23_4_678/m2_1_40# top VSUBS DUMMY
XDUMMY_63 via23_4_590/m2_1_40# top VSUBS DUMMY
XDUMMY_30 via23_4_251/m2_1_40# top VSUBS DUMMY
XDUMMY_52 via23_4_381/m2_1_40# top VSUBS DUMMY
XDUMMY_41 via23_4_89/m2_1_40# top VSUBS DUMMY
XC6_47 n6 top VSUBS C6
XC6_14 n6 top VSUBS C6
XC6_58 n6 top VSUBS C6
XC6_25 n6 top VSUBS C6
XC6_36 n6 top VSUBS C6
XDUMMY_1 via23_4_9/m2_1_40# top VSUBS DUMMY
XC7_90 n7 top VSUBS C7
XC6_4 n6 top VSUBS C6
XC4_1 n4 top VSUBS C4
XC7_116 n7 top VSUBS C7
XC7_105 n7 top VSUBS C7
XC7_127 n7 top VSUBS C7
XDUMMY_20 via23_4_199/m2_1_40# top VSUBS DUMMY
XDUMMY_64 via23_4_584/m2_1_40# top VSUBS DUMMY
XDUMMY_31 via23_4_245/m2_1_40# top VSUBS DUMMY
XDUMMY_75 via23_4_704/m2_1_40# top VSUBS DUMMY
XDUMMY_42 via23_4_366/m2_1_40# top VSUBS DUMMY
XDUMMY_53 via23_4_449/m2_1_40# top VSUBS DUMMY
XC6_26 n6 top VSUBS C6
XC6_15 n6 top VSUBS C6
XC6_59 n6 top VSUBS C6
XC6_48 n6 top VSUBS C6
XDUMMY_2 via23_4_1/m2_1_40# top VSUBS DUMMY
XC6_37 n6 top VSUBS C6
XC7_91 n7 top VSUBS C7
XC7_80 n7 top VSUBS C7
XC6_5 n6 top VSUBS C6
XC4_2 n4 top VSUBS C4
XC7_117 n7 top VSUBS C7
XC7_106 n7 top VSUBS C7
XDUMMY_76 via23_4_702/m2_1_40# top VSUBS DUMMY
XDUMMY_65 via23_4_600/m2_1_40# top VSUBS DUMMY
XDUMMY_32 via23_4_331/m2_1_40# top VSUBS DUMMY
XDUMMY_21 via23_4_198/m2_1_40# top VSUBS DUMMY
XDUMMY_43 via23_4_367/m2_1_40# top VSUBS DUMMY
XDUMMY_54 via23_4_446/m2_1_40# top VSUBS DUMMY
XDUMMY_10 via23_4_90/m2_1_40# top VSUBS DUMMY
XC6_27 n6 top VSUBS C6
XC6_16 n6 top VSUBS C6
XC6_49 n6 top VSUBS C6
XC6_38 n6 top VSUBS C6
XDUMMY_3 via23_4_2/m2_1_40# top VSUBS DUMMY
XC7_92 n7 top VSUBS C7
XC7_81 n7 top VSUBS C7
XC7_70 n7 top VSUBS C7
XC6_6 n6 top VSUBS C6
XC4_3 n4 top VSUBS C4
XC7_118 n7 top VSUBS C7
XC7_107 n7 top VSUBS C7
XC2_0 n2 top VSUBS C2
XDUMMY_66 via23_4_601/m2_1_40# top VSUBS DUMMY
XDUMMY_33 via23_4_332/m2_1_40# top VSUBS DUMMY
XDUMMY_22 via23_4_220/m2_1_40# top VSUBS DUMMY
XDUMMY_77 via23_4_705/m2_1_40# top VSUBS DUMMY
XDUMMY_44 via23_4_368/m2_1_40# top VSUBS DUMMY
XDUMMY_55 via23_4_447/m2_1_40# top VSUBS DUMMY
XDUMMY_11 via23_4_96/m2_1_40# top VSUBS DUMMY
XC6_28 n6 top VSUBS C6
XC6_17 n6 top VSUBS C6
XC6_39 n6 top VSUBS C6
XDUMMY_4 via23_4_20/m2_1_40# top VSUBS DUMMY
XC7_60 n7 top VSUBS C7
XC7_93 n7 top VSUBS C7
XC7_82 n7 top VSUBS C7
XC7_71 n7 top VSUBS C7
XC6_7 n6 top VSUBS C6
XC4_4 n4 top VSUBS C4
XC7_119 n7 top VSUBS C7
XC7_108 n7 top VSUBS C7
XC2_1 n2 top VSUBS C2
XDUMMY_78 via23_4_710/m2_1_40# top VSUBS DUMMY
XDUMMY_67 via23_4_599/m2_1_40# top VSUBS DUMMY
XDUMMY_34 via23_4_333/m2_1_40# top VSUBS DUMMY
XDUMMY_23 via23_4_213/m2_1_40# top VSUBS DUMMY
XDUMMY_45 via23_4_369/m2_1_40# top VSUBS DUMMY
XDUMMY_56 via23_4_458/m2_1_40# top VSUBS DUMMY
XDUMMY_12 via23_4_103/m2_1_40# top VSUBS DUMMY
XC6_18 n6 top VSUBS C6
XC6_29 n6 top VSUBS C6
XDUMMY_5 via23_4_21/m2_1_40# top VSUBS DUMMY
XC7_61 n7 top VSUBS C7
XC7_94 n7 top VSUBS C7
XC7_50 n7 top VSUBS C7
XC7_72 n7 top VSUBS C7
XC7_83 n7 top VSUBS C7
XC6_8 n6 top VSUBS C6
XC4_5 n4 top VSUBS C4
XC7_109 n7 top VSUBS C7
XC2_2 n2 top VSUBS C2
XDUMMY_79 via23_4_711/m2_1_40# top VSUBS DUMMY
XDUMMY_68 via23_4_598/m2_1_40# top VSUBS DUMMY
XDUMMY_35 via23_4_347/m2_1_40# top VSUBS DUMMY
XDUMMY_24 via23_4_229/m2_1_40# top VSUBS DUMMY
XDUMMY_46 via23_4_378/m2_1_40# top VSUBS DUMMY
XDUMMY_57 via23_4_455/m2_1_40# top VSUBS DUMMY
XDUMMY_13 via23_4_91/m2_1_40# top VSUBS DUMMY
XC6_19 n6 top VSUBS C6
XDUMMY_6 via23_4_22/m2_1_40# top VSUBS DUMMY
XC7_62 n7 top VSUBS C7
XC7_40 n7 top VSUBS C7
XC7_95 n7 top VSUBS C7
XC7_51 n7 top VSUBS C7
XC7_73 n7 top VSUBS C7
XC7_84 n7 top VSUBS C7
XC6_9 n6 top VSUBS C6
XC4_6 n4 top VSUBS C4
XC2_3 n2 top VSUBS C2
XDUMMY_36 via23_4_354/m2_1_40# top VSUBS DUMMY
XDUMMY_25 via23_4_228/m2_1_40# top VSUBS DUMMY
XDUMMY_14 via23_4_94/m2_1_40# top VSUBS DUMMY
XDUMMY_69 via23_4_635/m2_1_40# top VSUBS DUMMY
XDUMMY_47 via23_4_379/m2_1_40# top VSUBS DUMMY
XDUMMY_58 via23_4_459/m2_1_40# top VSUBS DUMMY
XDUMMY_7 via23_4_23/m2_1_40# top VSUBS DUMMY
XC7_41 n7 top VSUBS C7
XC7_63 n7 top VSUBS C7
XC7_96 n7 top VSUBS C7
XC7_52 n7 top VSUBS C7
XC7_30 n7 top VSUBS C7
XC7_74 n7 top VSUBS C7
XC7_85 n7 top VSUBS C7
XC4_7 n4 top VSUBS C4
XDUMMY_37 via23_4_345/m2_1_40# top VSUBS DUMMY
XDUMMY_26 via23_4_230/m2_1_40# top VSUBS DUMMY
XDUMMY_48 via23_4_380/m2_1_40# top VSUBS DUMMY
XDUMMY_59 via23_4_460/m2_1_40# top VSUBS DUMMY
XDUMMY_15 via23_4_117/m2_1_40# top VSUBS DUMMY
XDUMMY_8 via23_4_87/m2_1_40# top VSUBS DUMMY
XC7_97 n7 top VSUBS C7
XC7_42 n7 top VSUBS C7
XC7_53 n7 top VSUBS C7
XC7_31 n7 top VSUBS C7
XC7_86 n7 top VSUBS C7
XC7_20 n7 top VSUBS C7
XC7_64 n7 top VSUBS C7
XC7_75 n7 top VSUBS C7
XC4_10 n4 top VSUBS C4
XC4_8 n4 top VSUBS C4
XDUMMY_38 via23_4_346/m2_1_40# top VSUBS DUMMY
XDUMMY_27 via23_4_218/m2_1_40# top VSUBS DUMMY
XDUMMY_16 via23_4_111/m2_1_40# top VSUBS DUMMY
XDUMMY_49 via23_4_419/m2_1_40# top VSUBS DUMMY
XDUMMY_9 via23_4_88/m2_1_40# top VSUBS DUMMY
XC7_98 n7 top VSUBS C7
XC7_43 n7 top VSUBS C7
XC7_54 n7 top VSUBS C7
XC7_32 n7 top VSUBS C7
XC7_87 n7 top VSUBS C7
XC7_65 n7 top VSUBS C7
XC7_10 n7 top VSUBS C7
XC7_21 n7 top VSUBS C7
XC7_76 n7 top VSUBS C7
XC4_11 n4 top VSUBS C4
XC4_9 n4 top VSUBS C4
XDUMMY_39 via23_4_334/m2_1_40# top VSUBS DUMMY
XDUMMY_28 via23_4_249/m2_1_40# top VSUBS DUMMY
XDUMMY_17 via23_4_128/m2_1_40# top VSUBS DUMMY
XC7_99 n7 top VSUBS C7
XC7_33 n7 top VSUBS C7
XC7_88 n7 top VSUBS C7
XC7_55 n7 top VSUBS C7
XC7_44 n7 top VSUBS C7
XC7_66 n7 top VSUBS C7
XC7_11 n7 top VSUBS C7
XC7_77 n7 top VSUBS C7
XC7_22 n7 top VSUBS C7
XC4_12 n4 top VSUBS C4
XDUMMY_29 via23_4_250/m2_1_40# top VSUBS DUMMY
XDUMMY_18 via23_4_95/m2_1_40# top VSUBS DUMMY
XC7_45 n7 top VSUBS C7
XC7_56 n7 top VSUBS C7
XC7_34 n7 top VSUBS C7
XC7_89 n7 top VSUBS C7
XC7_12 n7 top VSUBS C7
XC7_23 n7 top VSUBS C7
XC7_78 n7 top VSUBS C7
XC7_67 n7 top VSUBS C7
XC4_13 n4 top VSUBS C4
XDUMMY_19 via23_4_200/m2_1_40# top VSUBS DUMMY
XC7_46 n7 top VSUBS C7
XC7_57 n7 top VSUBS C7
XC7_24 n7 top VSUBS C7
XC7_35 n7 top VSUBS C7
XC7_13 n7 top VSUBS C7
XC7_79 n7 top VSUBS C7
XC7_68 n7 top VSUBS C7
XC4_14 n4 top VSUBS C4
XC7_36 n7 top VSUBS C7
XC7_58 n7 top VSUBS C7
XC7_47 n7 top VSUBS C7
XC7_25 n7 top VSUBS C7
XC7_14 n7 top VSUBS C7
XC7_69 n7 top VSUBS C7
XC4_15 n4 top VSUBS C4
XC7_0 n7 top VSUBS C7
XC7_37 n7 top VSUBS C7
XC7_59 n7 top VSUBS C7
XC7_26 n7 top VSUBS C7
XC7_48 n7 top VSUBS C7
XC7_15 n7 top VSUBS C7
XC7_1 n7 top VSUBS C7
XC7_38 n7 top VSUBS C7
XC7_27 n7 top VSUBS C7
XC7_49 n7 top VSUBS C7
XC7_16 n7 top VSUBS C7
XC7_2 n7 top VSUBS C7
XC7_39 n7 top VSUBS C7
XC7_28 n7 top VSUBS C7
XC7_17 n7 top VSUBS C7
XC7_3 n7 top VSUBS C7
XC5_0 n5 top VSUBS C5
XC7_29 n7 top VSUBS C7
XC7_18 n7 top VSUBS C7
XC7_4 n7 top VSUBS C7
XC5_1 n5 top VSUBS C5
XC7_19 n7 top VSUBS C7
XC5_30 n5 top VSUBS C5
XC7_5 n7 top VSUBS C7
XC5_2 n5 top VSUBS C5
XC5_31 n5 top VSUBS C5
XC5_20 n5 top VSUBS C5
XC7_6 n7 top VSUBS C7
XC5_3 n5 top VSUBS C5
XC3_0 n3 top VSUBS C3
XC5_10 n5 top VSUBS C5
XC5_21 n5 top VSUBS C5
XC7_7 n7 top VSUBS C7
XC5_4 n5 top VSUBS C5
XC3_1 n3 top VSUBS C3
XC5_22 n5 top VSUBS C5
XC5_11 n5 top VSUBS C5
XC7_8 n7 top VSUBS C7
XC5_5 n5 top VSUBS C5
XC3_2 n3 top VSUBS C3
XC5_23 n5 top VSUBS C5
XC7_9 n7 top VSUBS C7
XC5_12 n5 top VSUBS C5
XC5_6 n5 top VSUBS C5
XC3_3 n3 top VSUBS C3
XC1_0 n1 top VSUBS C1
XC5_24 n5 top VSUBS C5
XC5_13 n5 top VSUBS C5
XC5_7 n5 top VSUBS C5
XC3_4 n3 top VSUBS C3
XC1_1 n1 top VSUBS C1
XC5_25 n5 top VSUBS C5
XC5_14 n5 top VSUBS C5
XC5_8 n5 top VSUBS C5
XC3_5 n3 top VSUBS C3
XC5_15 n5 top VSUBS C5
XC5_26 n5 top VSUBS C5
XC5_9 n5 top VSUBS C5
XC3_6 n3 top VSUBS C3
XC5_16 n5 top VSUBS C5
XC5_27 n5 top VSUBS C5
XC3_7 n3 top VSUBS C3
XC0_1_0 n0 top VSUBS C0_1
XC5_28 n5 top VSUBS C5
XC5_17 n5 top VSUBS C5
XC6_60 n6 top VSUBS C6
XC5_29 n5 top VSUBS C5
XC5_18 n5 top VSUBS C5
XC6_61 n6 top VSUBS C6
XC6_50 n6 top VSUBS C6
XC5_19 n5 top VSUBS C5
XC6_51 n6 top VSUBS C6
XC6_62 n6 top VSUBS C6
XC6_40 n6 top VSUBS C6
XC7_120 n7 top VSUBS C7
XC6_63 n6 top VSUBS C6
XC6_52 n6 top VSUBS C6
XC6_30 n6 top VSUBS C6
XC6_41 n6 top VSUBS C6
C0 m2_7300_1156# m3_7600_1156# 0.181f
C1 n2 m2_23300_1156# 0.249f
C2 m3_25600_1156# n5 0.00889f
C3 n6 m3_16500_1156# 0.181f
C4 top via23_4_641/m2_1_40# 0.216f
C5 m2_7300_1156# n1 8.05e-20
C6 via23_4_22/m2_1_40# m3_15200_1156# 0.247f
C7 top m3_19100_1156# 0.187f
C8 via23_4_218/m2_1_40# m2_4700_1156# 0.251f
C9 via23_4_600/m2_1_40# top 0.347f
C10 via23_4_711/m2_1_40# m3_40100_1156# 0.247f
C11 n7 m2_25900_1156# 1.13f
C12 m2_20300_1156# n5 2.05e-19
C13 m2_13800_1156# n3 5.59e-19
C14 via23_4_705/m2_1_40# m2_42800_1156# 0.251f
C15 m3_3700_1156# m3_4800_1156# 0.148f
C16 top m2_7300_1156# 0.267f
C17 m2_25900_1156# m3_25800_1156# 2.11f
C18 n2 m3_10000_1156# 0.021f
C19 m3_42500_1156# m3_42700_1156# 3.35f
C20 n2 via23_4_103/m2_1_40# 0.169f
C21 via23_4_23/m2_1_40# m3_16500_1156# 0.247f
C22 top m3_900_1156# 0.187f
C23 m2_40200_1156# m3_40100_1156# 2.11f
C24 ndum m2_4700_1156# 3.15e-20
C25 top via23_4_709/m2_1_40# 0.347f
C26 via23_4_96/m2_1_40# n3 4.28e-19
C27 via23_4_90/m2_1_40# m3_8900_1156# 0.247f
C28 n7 via23_4_21/m2_1_40# 0.452f
C29 via23_4_22/m2_1_40# n7 0.452f
C30 n7 m3_41200_1156# 0.00642f
C31 via23_4_367/m2_1_40# m3_42700_1156# 0.247f
C32 m2_16400_1156# m3_15400_1156# 0.0061f
C33 n6 m3_27100_1156# 0.181f
C34 via23_4_2/m2_1_40# n4 2.21e-19
C35 top via23_4_326/m2_1_40# 0.347f
C36 via23_4_220/m2_1_40# m2_800_1156# 0.251f
C37 via23_4_249/m2_1_40# m3_6300_1156# 0.247f
C38 top m3_29700_1156# 0.187f
C39 m2_12500_1156# n4 3.19e-19
C40 m3_33400_1156# m3_33600_1156# 3.35f
C41 via23_4_1/m2_1_40# n5 2.03e-19
C42 m2_4700_1156# n5 2.05e-19
C43 n7 m2_36300_1156# 1.13f
C44 via23_4_250/m2_1_40# m2_8600_1156# 0.251f
C45 m2_23300_1156# n3 1.09f
C46 m2_31100_1156# m3_31000_1156# 2.11f
C47 n2 m3_19300_1156# 0.0215f
C48 top via23_4_111/m2_1_40# 0.216f
C49 via23_4_94/m2_1_40# m3_3700_1156# 0.247f
C50 via23_4_599/m2_1_40# top 0.347f
C51 ndum m2_11200_1156# 3.15e-20
C52 n2 n4 0.147f
C53 via23_4_89/m2_1_40# m3_10200_1156# 0.247f
C54 via23_4_2/m2_1_40# n0 0.381f
C55 via23_4_449/m2_1_40# m3_28400_1156# 0.247f
C56 via23_4_381/m2_1_40# n6 0.0598f
C57 via23_4_704/m2_1_40# m3_42700_1156# 0.247f
C58 n0 m2_12500_1156# 6.36e-20
C59 n2 m2_15100_1156# 0.00855f
C60 m3_15400_1156# n5 4.08f
C61 n6 n1 0.0843f
C62 top m3_10200_1156# 0.187f
C63 m3_24300_1156# m3_24500_1156# 3.35f
C64 via23_4_103/m2_1_40# n3 4.28e-19
C65 n7 m2_17700_1156# 1.13f
C66 n6 via23_4_89/m2_1_40# 1.52e-19
C67 m2_11200_1156# n5 0.636f
C68 n2 m3_1100_1156# 0.021f
C69 via23_4_369/m2_1_40# m2_40200_1156# 0.251f
C70 n2 n0 1.42f
C71 top n6 16.4f
C72 n6 m3_37300_1156# 4.09f
C73 via23_4_710/m2_1_40# m2_38900_1156# 0.251f
C74 top m3_39900_1156# 0.187f
C75 via23_4_677/m2_1_40# m2_35000_1156# 0.251f
C76 via23_4_23/m2_1_40# n1 9.38e-20
C77 via23_4_3/m2_1_40# m3_16700_1156# 0.123f
C78 via23_4_220/m2_1_40# m3_900_1156# 0.247f
C79 n7 m3_3500_1156# 0.181f
C80 via23_4_590/m2_1_40# m3_25800_1156# 0.247f
C81 n6 m2_32400_1156# 1.13f
C82 via23_4_213/m2_1_40# top 0.216f
C83 n6 via23_4_446/m2_1_40# 0.452f
C84 top m2_35000_1156# 0.267f
C85 m3_13900_1156# m3_14100_1156# 3.35f
C86 m2_36300_1156# m3_36000_1156# 0.181f
C87 via23_4_414/m2_1_40# m2_42800_1156# 0.251f
C88 via23_4_378/m2_1_40# m3_33600_1156# 0.247f
C89 top via23_4_23/m2_1_40# 0.14f
C90 n2 m2_24600_1156# 1.37e-19
C91 m3_26900_1156# n5 0.00889f
C92 n6 m3_17800_1156# 1.98f
C93 top m3_20400_1156# 0.187f
C94 n7 m2_27200_1156# 1.05e-19
C95 n2 via23_4_3/m2_1_40# 0.169f
C96 n3 n4 10.8f
C97 top via23_4_347/m2_1_40# 0.347f
C98 top via23_4_460/m2_1_40# 0.14f
C99 n6 m2_6000_1156# 1.13f
C100 m2_15100_1156# n3 5.59e-19
C101 via23_4_20/m2_1_40# n1 9.38e-20
C102 m3_4800_1156# m3_5000_1156# 3.35f
C103 n2 m3_11300_1156# 0.021f
C104 via23_4_599/m2_1_40# m3_28400_1156# 0.247f
C105 top via23_4_20/m2_1_40# 0.14f
C106 n7 m3_12800_1156# 4.08f
C107 via23_4_675/m2_1_40# m3_32300_1156# 0.247f
C108 via23_4_601/m2_1_40# m2_31100_1156# 0.251f
C109 top m3_2200_1156# 0.187f
C110 n0 n3 1.36f
C111 via23_4_709/m2_1_40# m3_38600_1156# 0.247f
C112 m2_4700_1156# m3_3700_1156# 0.0061f
C113 via23_4_439/m2_1_40# m3_32300_1156# 0.247f
C114 m2_800_1156# m3_900_1156# 2.11f
C115 top via23_4_128/m2_1_40# 0.216f
C116 m2_16400_1156# m3_16700_1156# 0.181f
C117 n7 m3_42500_1156# 4.08f
C118 n6 via23_4_458/m2_1_40# 0.452f
C119 top via23_4_200/m2_1_40# 0.216f
C120 top m3_31000_1156# 0.187f
C121 m2_13800_1156# n4 3.19e-19
C122 via23_4_213/m2_1_40# via23_4_220/m2_1_40# 0.199f
C123 m3_33600_1156# m3_34700_1156# 0.148f
C124 via23_4_90/m2_1_40# n6 1.52e-19
C125 via23_4_332/m2_1_40# m3_12800_1156# 0.247f
C126 n7 m2_37600_1156# 2.39f
C127 top m2_25900_1156# 0.267f
C128 via23_4_446/m2_1_40# m3_31000_1156# 0.247f
C129 via23_4_88/m2_1_40# n7 0.452f
C130 via23_4_249/m2_1_40# top 0.347f
C131 ndum m2_12500_1156# 3.15e-20
C132 via23_4_3/m2_1_40# n3 4.28e-19
C133 via23_4_111/m2_1_40# m2_800_1156# 0.251f
C134 n0 m2_13800_1156# 6.36e-20
C135 via23_4_96/m2_1_40# n4 2.85e-19
C136 n2 m2_16400_1156# 0.00855f
C137 n2 m2_2100_1156# 0.00855f
C138 via23_4_21/m2_1_40# n1 9.38e-20
C139 top m3_11500_1156# 0.187f
C140 via23_4_22/m2_1_40# n1 9.38e-20
C141 m3_24500_1156# m3_25600_1156# 0.148f
C142 n7 m2_19000_1156# 2.42f
C143 via23_4_600/m2_1_40# m3_29700_1156# 0.247f
C144 via23_4_2/m2_1_40# n5 1.57e-19
C145 m2_12500_1156# n5 2.05e-19
C146 via23_4_642/m2_1_40# m3_42700_1156# 0.247f
C147 via23_4_712/m2_1_40# m2_41500_1156# 0.251f
C148 ndum n2 1.42f
C149 top via23_4_21/m2_1_40# 0.14f
C150 n2 m3_2400_1156# 0.021f
C151 via23_4_702/m2_1_40# m2_42800_1156# 0.251f
C152 n6 m3_38600_1156# 0.00746f
C153 top via23_4_22/m2_1_40# 0.14f
C154 top m3_41200_1156# 0.187f
C155 m2_23300_1156# n4 2.39f
C156 n6 m2_800_1156# 1.43e-19
C157 n7 m3_4800_1156# 2.16f
C158 n6 m2_33700_1156# 0.00135f
C159 via23_4_429/m2_1_40# via23_4_367/m2_1_40# 0.199f
C160 n2 n5 0.196f
C161 top m2_36300_1156# 0.316f
C162 m3_14100_1156# m3_15200_1156# 0.148f
C163 m2_36300_1156# m3_37300_1156# 0.0061f
C164 n2 m2_8600_1156# 0.00855f
C165 via23_4_213/m2_1_40# m2_800_1156# 0.251f
C166 via23_4_449/m2_1_40# n6 1.52e-19
C167 m2_12500_1156# m3_12600_1156# 2.11f
C168 n7 m3_33600_1156# 1.98f
C169 via23_4_103/m2_1_40# n4 2.85e-19
C170 n0 m2_23300_1156# 6.84e-20
C171 top via23_4_635/m2_1_40# 0.216f
C172 via23_4_598/m2_1_40# m3_28200_1156# 0.247f
C173 m2_17700_1156# n1 8.05e-20
C174 m3_28200_1156# n5 4.09f
C175 via23_4_111/m2_1_40# m3_900_1156# 0.247f
C176 n6 m2_7300_1156# 2.39f
C177 m2_16400_1156# n3 5.59e-19
C178 top m2_17700_1156# 0.267f
C179 n2 m3_12600_1156# 0.021f
C180 via23_4_458/m2_1_40# m2_25900_1156# 0.251f
C181 m3_5000_1156# m3_6100_1156# 0.148f
C182 m2_27200_1156# m3_27100_1156# 2.11f
C183 top via23_4_601/m2_1_40# 0.347f
C184 m2_2100_1156# n3 5.59e-19
C185 via23_4_345/m2_1_40# m3_16700_1156# 0.123f
C186 via23_4_103/m2_1_40# m3_1100_1156# 0.247f
C187 via23_4_590/m2_1_40# top 0.347f
C188 n7 m3_14100_1156# 4.08f
C189 ndum n3 1.36f
C190 via23_4_94/m2_1_40# n7 0.452f
C191 top m3_3500_1156# 0.187f
C192 via23_4_326/m2_1_40# m3_10200_1156# 0.247f
C193 m2_41500_1156# m3_41400_1156# 2.11f
C194 via23_4_459/m2_1_40# m2_23300_1156# 0.251f
C195 m2_8600_1156# m3_8700_1156# 2.11f
C196 m2_4700_1156# m3_5000_1156# 0.181f
C197 n7 m2_9900_1156# 2.39f
C198 m3_19300_1156# n4 4.08f
C199 n7 via23_4_9/m2_1_40# 0.227f
C200 via23_4_213/m2_1_40# m3_900_1156# 0.247f
C201 m2_17700_1156# m3_17800_1156# 2.11f
C202 via23_4_87/m2_1_40# m3_7400_1156# 0.247f
C203 n3 n5 0.161f
C204 m2_15100_1156# n4 3.19e-19
C205 via23_4_128/m2_1_40# m2_800_1156# 0.251f
C206 top m3_32300_1156# 0.187f
C207 m2_8600_1156# n3 5.59e-19
C208 m3_34700_1156# m3_34900_1156# 3.35f
C209 n7 m2_38900_1156# 3.52f
C210 n7 via23_4_346/m2_1_40# 0.227f
C211 via23_4_200/m2_1_40# m2_800_1156# 0.251f
C212 top m2_27200_1156# 0.267f
C213 m2_32400_1156# m3_32300_1156# 2.11f
C214 via23_4_448/m2_1_40# m3_28200_1156# 0.247f
C215 n2 m3_23200_1156# 3.41f
C216 n0 n4 0.0773f
C217 via23_4_588/m2_1_40# m3_24300_1156# 0.247f
C218 ndum m2_13800_1156# 3.15e-20
C219 n0 m2_15100_1156# 6.36e-20
C220 n7 m3_25600_1156# 4.08f
C221 n2 m2_3400_1156# 0.00855f
C222 top m3_12800_1156# 0.187f
C223 m3_25600_1156# m3_25800_1156# 3.35f
C224 n7 m2_20300_1156# 1.05e-19
C225 via23_4_95/m2_1_40# m3_6100_1156# 0.247f
C226 m2_13800_1156# n5 2.05e-19
C227 via23_4_381/m2_1_40# m2_37600_1156# 0.251f
C228 n2 m3_3700_1156# 0.021f
C229 n6 m3_39900_1156# 0.00746f
C230 via23_4_331/m2_1_40# m3_12600_1156# 0.123f
C231 top m3_42500_1156# 0.187f
C232 m2_24600_1156# n4 1.13f
C233 via23_4_88/m2_1_40# m3_7600_1156# 0.247f
C234 via23_4_128/m2_1_40# m3_900_1156# 0.247f
C235 n7 m3_6100_1156# 1.98f
C236 n6 m2_35000_1156# 0.00135f
C237 via23_4_88/m2_1_40# n1 9.38e-20
C238 via23_4_459/m2_1_40# n4 0.541f
C239 via23_4_676/m2_1_40# m3_34700_1156# 0.247f
C240 via23_4_3/m2_1_40# n4 2.85e-19
C241 top via23_4_198/m2_1_40# 0.216f
C242 via23_4_333/m2_1_40# m2_15100_1156# 0.251f
C243 top m2_37600_1156# 0.267f
C244 m3_15200_1156# m3_15400_1156# 3.35f
C245 m2_37600_1156# m3_37300_1156# 0.181f
C246 via23_4_96/m2_1_40# n5 2.03e-19
C247 via23_4_200/m2_1_40# m3_900_1156# 0.247f
C248 via23_4_249/m2_1_40# m2_7300_1156# 0.251f
C249 n6 via23_4_23/m2_1_40# 1.52e-19
C250 ndum m2_23300_1156# 1.36e-19
C251 top via23_4_88/m2_1_40# 0.14f
C252 top via23_4_367/m2_1_40# 0.136f
C253 n7 m3_34900_1156# 1.19f
C254 m3_29500_1156# n5 0.00889f
C255 m2_19000_1156# n1 8.05e-20
C256 n2 via23_4_87/m2_1_40# 0.169f
C257 n7 via23_4_1/m2_1_40# 1.18e-19
C258 n7 via23_4_250/m2_1_40# 0.452f
C259 m3_23200_1156# n3 0.174f
C260 n7 m2_4700_1156# 3.52f
C261 via23_4_251/m2_1_40# m3_10000_1156# 0.247f
C262 top m3_24300_1156# 0.187f
C263 via23_4_229/m2_1_40# m3_1100_1156# 0.247f
C264 via23_4_334/m2_1_40# m2_16400_1156# 0.251f
C265 via23_4_103/m2_1_40# m2_2100_1156# 0.251f
C266 n6 via23_4_460/m2_1_40# 1.52e-19
C267 m2_23300_1156# n5 2.05e-19
C268 via23_4_368/m2_1_40# m3_38800_1156# 0.247f
C269 top m2_19000_1156# 0.267f
C270 m3_6100_1156# m3_6300_1156# 3.35f
C271 n2 m3_13900_1156# 0.021f
C272 m2_28500_1156# m3_28200_1156# 0.181f
C273 m2_3400_1156# n3 5.59e-19
C274 n2 via23_4_91/m2_1_40# 0.169f
C275 n6 via23_4_20/m2_1_40# 0.452f
C276 top via23_4_704/m2_1_40# 0.222f
C277 n6 m3_2200_1156# 0.181f
C278 m3_10000_1156# n5 0.181f
C279 top m3_4800_1156# 0.187f
C280 via23_4_103/m2_1_40# n5 2.03e-19
C281 via23_4_334/m2_1_40# n5 0.452f
C282 n7 m2_11200_1156# 1.05e-19
C283 via23_4_347/m2_1_40# m3_20400_1156# 0.247f
C284 n6 m3_31000_1156# 1.98f
C285 m2_16400_1156# n4 3.19e-19
C286 top m3_33600_1156# 0.187f
C287 m3_34900_1156# m3_36000_1156# 0.354f
C288 m2_2100_1156# n4 3.19e-19
C289 n7 via23_4_676/m2_1_40# 0.452f
C290 n7 m2_40200_1156# 1.13f
C291 n7 via23_4_379/m2_1_40# 0.452f
C292 via23_4_245/m2_1_40# m3_6100_1156# 0.247f
C293 n6 m2_25900_1156# 2.39f
C294 via23_4_87/m2_1_40# n3 4.28e-19
C295 n2 m3_24500_1156# 3.24e-19
C296 via23_4_249/m2_1_40# n6 0.452f
C297 ndum n4 0.0771f
C298 ndum m2_15100_1156# 3.15e-20
C299 via23_4_94/m2_1_40# n1 9.38e-20
C300 n0 m2_16400_1156# 6.36e-20
C301 m2_9900_1156# n1 8.05e-20
C302 n6 m3_11500_1156# 4.08f
C303 n0 m2_2100_1156# 6.36e-20
C304 m2_2100_1156# m3_1100_1156# 0.0061f
C305 via23_4_9/m2_1_40# n1 9.38e-20
C306 via23_4_705/m2_1_40# m3_42700_1156# 0.247f
C307 top m3_14100_1156# 0.187f
C308 via23_4_91/m2_1_40# n3 4.28e-19
C309 m3_25800_1156# m3_26900_1156# 0.148f
C310 n4 n5 11.4f
C311 top via23_4_94/m2_1_40# 0.14f
C312 m2_15100_1156# n5 1.13f
C313 ndum n0 13.4f
C314 m2_8600_1156# n4 3.19e-19
C315 n6 via23_4_21/m2_1_40# 1.52e-19
C316 top m2_9900_1156# 0.267f
C317 n6 via23_4_22/m2_1_40# 1.52e-19
C318 m2_23300_1156# m3_23200_1156# 2.11f
C319 n2 m3_5000_1156# 0.021f
C320 top via23_4_9/m2_1_40# 0.14f
C321 n6 m3_41200_1156# 4.08f
C322 n2 via23_4_354/m2_1_40# 0.247f
C323 n7 m3_7400_1156# 0.181f
C324 n6 m2_36300_1156# 0.637f
C325 n0 n5 0.0772f
C326 top m2_38900_1156# 0.267f
C327 via23_4_379/m2_1_40# m3_36000_1156# 0.247f
C328 m3_15400_1156# m3_16500_1156# 0.148f
C329 m2_37600_1156# m3_38600_1156# 0.0061f
C330 top via23_4_346/m2_1_40# 0.347f
C331 via23_4_229/m2_1_40# m2_2100_1156# 0.251f
C332 n0 m2_8600_1156# 6.36e-20
C333 via23_4_366/m2_1_40# m3_42500_1156# 0.247f
C334 via23_4_198/m2_1_40# m2_800_1156# 0.251f
C335 n7 m3_36200_1156# 0.181f
C336 m2_13800_1156# m3_13900_1156# 2.11f
C337 m3_30800_1156# n5 0.00889f
C338 m2_20300_1156# n1 8.05e-20
C339 top m3_25600_1156# 0.187f
C340 via23_4_589/m2_1_40# m3_25600_1156# 0.247f
C341 via23_4_20/m2_1_40# m3_11500_1156# 0.247f
C342 n6 m2_17700_1156# 2.39f
C343 m2_24600_1156# n5 0.002f
C344 top m2_20300_1156# 0.267f
C345 via23_4_601/m2_1_40# n6 0.452f
C346 n2 m3_15200_1156# 0.021f
C347 m3_6300_1156# m3_7400_1156# 0.148f
C348 m2_28500_1156# m3_29500_1156# 0.0061f
C349 via23_4_459/m2_1_40# n5 2.03e-19
C350 via23_4_3/m2_1_40# n5 2.03e-19
C351 via23_4_590/m2_1_40# n6 0.452f
C352 via23_4_419/m2_1_40# m2_42800_1156# 0.251f
C353 n6 m3_3500_1156# 1.98f
C354 m3_11300_1156# n5 0.993f
C355 top m3_6100_1156# 0.187f
C356 m2_42800_1156# m3_42700_1156# 2.11f
C357 via23_4_2/m2_1_40# n7 9.11e-20
C358 via23_4_369/m2_1_40# m3_40100_1156# 0.247f
C359 n7 m2_12500_1156# 1.13f
C360 via23_4_250/m2_1_40# m3_7600_1156# 0.247f
C361 top via23_4_642/m2_1_40# 0.216f
C362 via23_4_677/m2_1_40# m3_34900_1156# 0.123f
C363 via23_4_710/m2_1_40# m3_38800_1156# 0.247f
C364 via23_4_1/m2_1_40# n1 9.38e-20
C365 m3_23200_1156# n4 1.99f
C366 m2_4700_1156# n1 8.05e-20
C367 n2 via23_4_95/m2_1_40# 0.169f
C368 via23_4_354/m2_1_40# n3 0.452f
C369 via23_4_419/m2_1_40# via23_4_414/m2_1_40# 0.199f
C370 via23_4_198/m2_1_40# m3_900_1156# 0.247f
C371 m2_19000_1156# m3_19100_1156# 2.11f
C372 n6 m3_32300_1156# 0.181f
C373 via23_4_709/m2_1_40# m2_37600_1156# 0.251f
C374 via23_4_90/m2_1_40# m2_9900_1156# 0.251f
C375 top m3_34900_1156# 0.221f
C376 m3_36000_1156# m3_36200_1156# 3.35f
C377 top via23_4_1/m2_1_40# 0.14f
C378 via23_4_414/m2_1_40# m3_42700_1156# 0.247f
C379 m2_3400_1156# n4 3.19e-19
C380 top m2_4700_1156# 0.267f
C381 top via23_4_250/m2_1_40# 0.347f
C382 n7 m2_41500_1156# 2.39f
C383 n2 n7 0.78f
C384 n6 m2_27200_1156# 1.13f
C385 n0 m3_23200_1156# 1.62e-19
C386 m2_33700_1156# m3_33600_1156# 2.11f
C387 ndum m2_16400_1156# 3.15e-20
C388 ndum m2_2100_1156# 3.15e-20
C389 m2_9900_1156# m3_8900_1156# 0.0061f
C390 m2_11200_1156# n1 8.05e-20
C391 m2_6000_1156# m3_6100_1156# 2.11f
C392 n0 m2_3400_1156# 6.36e-20
C393 m2_2100_1156# m3_2400_1156# 0.181f
C394 top m3_15400_1156# 0.187f
C395 m3_26900_1156# m3_27100_1156# 3.35f
C396 top via23_4_711/m2_1_40# 0.347f
C397 via23_4_89/m2_1_40# m2_11200_1156# 0.0256f
C398 m2_16400_1156# n5 2.39f
C399 top m2_11200_1156# 0.316f
C400 m2_2100_1156# n5 2.05e-19
C401 n2 m3_6300_1156# 0.021f
C402 via23_4_601/m2_1_40# m3_31000_1156# 0.247f
C403 via23_4_459/m2_1_40# m3_23200_1156# 0.247f
C404 via23_4_87/m2_1_40# n4 2.85e-19
C405 ndum n5 0.0767f
C406 n7 m3_8700_1156# 2.16f
C407 via23_4_95/m2_1_40# n3 4.28e-19
C408 n6 m2_37600_1156# 1.13f
C409 top via23_4_676/m2_1_40# 0.347f
C410 top via23_4_379/m2_1_40# 0.14f
C411 ndum m2_8600_1156# 3.15e-20
C412 top m2_40200_1156# 0.267f
C413 m2_38900_1156# m3_38600_1156# 0.181f
C414 m3_16500_1156# m3_16700_1156# 3.35f
C415 via23_4_380/m2_1_40# n7 1.18e-19
C416 via23_4_590/m2_1_40# m2_25900_1156# 0.251f
C417 via23_4_88/m2_1_40# n6 1.52e-19
C418 via23_4_91/m2_1_40# n4 2.85e-19
C419 n7 n3 0.623f
C420 via23_4_213/m2_1_40# via23_4_198/m2_1_40# 0.199f
C421 via23_4_598/m2_1_40# n5 0.452f
C422 n7 m3_37500_1156# 1.98f
C423 m3_32100_1156# n5 0.00889f
C424 via23_4_9/m2_1_40# m3_19100_1156# 0.247f
C425 top m3_26900_1156# 0.187f
C426 m2_8600_1156# n5 2.05e-19
C427 n2 via23_4_455/m2_1_40# 0.352f
C428 n6 m2_19000_1156# 1.43e-19
C429 m3_7400_1156# m3_7600_1156# 3.35f
C430 n2 m3_16500_1156# 0.021f
C431 m2_29800_1156# m3_29500_1156# 0.181f
C432 via23_4_346/m2_1_40# m3_19100_1156# 0.247f
C433 n7 m3_18000_1156# 3.1f
C434 via23_4_712/m2_1_40# m3_41400_1156# 0.247f
C435 top m3_7400_1156# 0.187f
C436 via23_4_702/m2_1_40# m3_42700_1156# 0.247f
C437 n7 m2_13800_1156# 3.52f
C438 m3_24500_1156# n4 0.181f
C439 n6 m3_33600_1156# 0.00746f
C440 top m3_36200_1156# 0.187f
C441 m3_36200_1156# m3_37300_1156# 0.148f
C442 n7 m2_42800_1156# 1.13f
C443 via23_4_218/m2_1_40# m3_3700_1156# 0.247f
C444 via23_4_584/m2_1_40# n2 0.247f
C445 via23_4_96/m2_1_40# n7 1.18e-19
C446 ndum m3_23200_1156# 3.28e-19
C447 via23_4_448/m2_1_40# n5 0.523f
C448 via23_4_200/m2_1_40# via23_4_198/m2_1_40# 0.199f
C449 via23_4_332/m2_1_40# m2_13800_1156# 0.251f
C450 via23_4_642/m2_1_40# via23_4_641/m2_1_40# 0.199f
C451 via23_4_455/m2_1_40# n3 0.453f
C452 ndum m2_3400_1156# 3.15e-20
C453 m2_9900_1156# m3_10200_1156# 0.181f
C454 n7 m3_29500_1156# 3.1f
C455 via23_4_2/m2_1_40# n1 0.251f
C456 m2_12500_1156# n1 8.05e-20
C457 via23_4_21/m2_1_40# m3_12800_1156# 0.247f
C458 m2_3400_1156# m3_2400_1156# 0.0061f
C459 top m3_16700_1156# 0.221f
C460 via23_4_230/m2_1_40# m3_2400_1156# 0.247f
C461 m3_27100_1156# m3_28200_1156# 0.148f
C462 via23_4_94/m2_1_40# n6 1.52e-19
C463 via23_4_458/m2_1_40# m3_26900_1156# 0.247f
C464 n7 m2_23300_1156# 1.05e-19
C465 n6 m2_9900_1156# 1.43e-19
C466 top via23_4_2/m2_1_40# 0.14f
C467 top m2_12500_1156# 0.267f
C468 m2_3400_1156# n5 2.05e-19
C469 n6 via23_4_9/m2_1_40# 1.52e-19
C470 m2_24600_1156# m3_24500_1156# 2.11f
C471 n2 m3_7600_1156# 0.021f
C472 via23_4_429/m2_1_40# m2_42800_1156# 0.251f
C473 n2 n1 2.02f
C474 n2 via23_4_89/m2_1_40# 0.169f
C475 n7 m3_10000_1156# 1.98f
C476 via23_4_354/m2_1_40# n0 0.247f
C477 n6 m2_38900_1156# 0.00135f
C478 top m2_41500_1156# 0.267f
C479 n7 via23_4_103/m2_1_40# 0.452f
C480 m3_16700_1156# m3_17800_1156# 0.354f
C481 top n2 1.32f
C482 m2_38900_1156# m3_39900_1156# 0.0061f
C483 via23_4_429/m2_1_40# via23_4_414/m2_1_40# 0.199f
C484 via23_4_676/m2_1_40# m2_33700_1156# 0.251f
C485 via23_4_584/m2_1_40# n3 0.452f
C486 m2_15100_1156# m3_15200_1156# 2.11f
C487 n7 m3_38800_1156# 2.16f
C488 m3_33400_1156# n5 4.08f
C489 top m3_28200_1156# 0.187f
C490 m2_28500_1156# n5 1.14f
C491 n6 m2_20300_1156# 1.43e-19
C492 m2_29800_1156# m3_30800_1156# 0.023f
C493 via23_4_87/m2_1_40# n5 2.03e-19
C494 m3_7600_1156# m3_8700_1156# 0.148f
C495 n2 m3_17800_1156# 0.021f
C496 via23_4_91/m2_1_40# m3_2400_1156# 0.247f
C497 via23_4_95/m2_1_40# n4 2.85e-19
C498 via23_4_381/m2_1_40# m3_37500_1156# 0.247f
C499 n2 m2_6000_1156# 0.00855f
C500 n6 m3_6100_1156# 0.181f
C501 via23_4_91/m2_1_40# n5 2.03e-19
C502 top m3_8700_1156# 0.187f
C503 top via23_4_705/m2_1_40# 0.216f
C504 n7 n4 0.678f
C505 n3 n1 3.36f
C506 n7 m2_15100_1156# 2.39f
C507 via23_4_89/m2_1_40# n3 4.28e-19
C508 via23_4_460/m2_1_40# m3_25600_1156# 0.247f
C509 via23_4_380/m2_1_40# top 0.14f
C510 via23_4_380/m2_1_40# m3_37300_1156# 0.247f
C511 via23_4_326/m2_1_40# m2_11200_1156# 0.0256f
C512 m2_20300_1156# m3_20400_1156# 2.11f
C513 n6 m3_34900_1156# 0.00746f
C514 top n3 2.35f
C515 via23_4_333/m2_1_40# m3_15200_1156# 0.247f
C516 top m3_37500_1156# 0.187f
C517 m3_37300_1156# m3_37500_1156# 3.35f
C518 n6 via23_4_1/m2_1_40# 1.52e-19
C519 via23_4_347/m2_1_40# m2_20300_1156# 0.251f
C520 n6 m2_4700_1156# 1.43e-19
C521 n7 n0 0.0951f
C522 via23_4_447/m2_1_40# m3_30800_1156# 0.123f
C523 n7 m3_1100_1156# 4.08f
C524 m2_35000_1156# m3_34900_1156# 2.11f
C525 via23_4_230/m2_1_40# m2_3400_1156# 0.251f
C526 top via23_4_331/m2_1_40# 0.347f
C527 via23_4_334/m2_1_40# m3_16500_1156# 0.247f
C528 via23_4_90/m2_1_40# n2 0.169f
C529 m2_11200_1156# m3_10200_1156# 0.0061f
C530 n7 m3_30800_1156# 3.14f
C531 m2_7300_1156# m3_7400_1156# 2.11f
C532 m2_13800_1156# n1 8.05e-20
C533 m3_24500_1156# n5 0.00889f
C534 m2_3400_1156# m3_3700_1156# 0.181f
C535 via23_4_22/m2_1_40# m3_14100_1156# 0.247f
C536 top m3_18000_1156# 0.187f
C537 n6 via23_4_711/m2_1_40# 0.452f
C538 m3_28200_1156# m3_28400_1156# 3.35f
C539 via23_4_588/m2_1_40# m2_23300_1156# 0.251f
C540 via23_4_1/m2_1_40# m3_20400_1156# 0.247f
C541 n7 m2_24600_1156# 2.39f
C542 n6 m2_11200_1156# 1.13f
C543 via23_4_229/m2_1_40# n7 0.452f
C544 top m2_13800_1156# 0.267f
C545 n7 via23_4_333/m2_1_40# 0.452f
C546 m2_25900_1156# m3_25600_1156# 0.181f
C547 m2_6000_1156# n3 5.59e-19
C548 n7 via23_4_459/m2_1_40# 1.18e-19
C549 top via23_4_678/m2_1_40# 0.347f
C550 n2 m3_8900_1156# 0.021f
C551 n7 via23_4_3/m2_1_40# 1.18e-19
C552 via23_4_678/m2_1_40# m3_37300_1156# 0.247f
C553 via23_4_96/m2_1_40# n1 9.38e-20
C554 via23_4_23/m2_1_40# m3_15400_1156# 0.247f
C555 n6 via23_4_379/m2_1_40# 0.0598f
C556 n6 m2_40200_1156# 2.39f
C557 top m2_42800_1156# 0.267f
C558 m2_40200_1156# m3_39900_1156# 0.181f
C559 m3_17800_1156# m3_18000_1156# 3.35f
C560 via23_4_455/m2_1_40# n4 2.21e-19
C561 top via23_4_96/m2_1_40# 0.136f
C562 n2 m2_800_1156# 0.00855f
C563 via23_4_379/m2_1_40# m2_35000_1156# 0.251f
C564 n7 m3_40100_1156# 0.181f
C565 n6 m3_26900_1156# 4.08f
C566 via23_4_366/m2_1_40# m2_41500_1156# 0.251f
C567 via23_4_91/m2_1_40# m2_3400_1156# 0.251f
C568 top via23_4_414/m2_1_40# 0.216f
C569 top m3_29500_1156# 0.187f
C570 via23_4_90/m2_1_40# n3 4.28e-19
C571 m2_29800_1156# n5 0.002f
C572 top m2_23300_1156# 0.267f
C573 m3_8700_1156# m3_8900_1156# 3.35f
C574 m2_31100_1156# m3_30800_1156# 0.181f
C575 n2 m3_19100_1156# 0.0213f
C576 via23_4_218/m2_1_40# n7 0.452f
C577 via23_4_103/m2_1_40# n1 9.38e-20
C578 n6 m3_7400_1156# 1.98f
C579 via23_4_588/m2_1_40# n4 0.452f
C580 n2 m2_7300_1156# 0.00855f
C581 m3_15200_1156# n5 0.181f
C582 top m3_10000_1156# 0.187f
C583 n7 m2_16400_1156# 1.05e-19
C584 top via23_4_103/m2_1_40# 0.14f
C585 via23_4_368/m2_1_40# n7 0.452f
C586 top via23_4_334/m2_1_40# 0.347f
C587 n7 m2_2100_1156# 2.39f
C588 n7 via23_4_251/m2_1_40# 0.452f
C589 n2 m3_900_1156# 0.021f
C590 n6 m3_36200_1156# 1f
C591 top m3_38800_1156# 0.187f
C592 m3_37500_1156# m3_38600_1156# 0.148f
C593 n7 via23_4_712/m2_1_40# 0.452f
C594 ndum n7 0.177f
C595 via23_4_447/m2_1_40# n5 0.0714f
C596 m2_800_1156# n3 5.59e-19
C597 via23_4_95/m2_1_40# n5 2.03e-19
C598 via23_4_369/m2_1_40# n7 1.18e-19
C599 via23_4_642/m2_1_40# via23_4_635/m2_1_40# 0.199f
C600 n7 n5 1.06f
C601 n4 n1 0.0766f
C602 via23_4_228/m2_1_40# top 0.276f
C603 m2_11200_1156# m3_11500_1156# 0.181f
C604 m2_15100_1156# n1 8.05e-20
C605 m3_25800_1156# n5 0.00889f
C606 n7 m2_8600_1156# 3.52f
C607 n6 m3_16700_1156# 3.14f
C608 via23_4_89/m2_1_40# n4 2.85e-19
C609 top m3_19300_1156# 0.187f
C610 m3_28400_1156# m3_29500_1156# 0.148f
C611 via23_4_711/m2_1_40# m3_41200_1156# 0.247f
C612 n6 via23_4_2/m2_1_40# 1.17e-19
C613 top n4 4.11f
C614 n6 m2_12500_1156# 2.39f
C615 top m2_15100_1156# 0.267f
C616 m2_7300_1156# n3 5.59e-19
C617 via23_4_419/m2_1_40# m3_42700_1156# 0.247f
C618 m2_25900_1156# m3_26900_1156# 0.0061f
C619 n2 m3_10200_1156# 0.021f
C620 n0 n1 13.4f
C621 via23_4_675/m2_1_40# n5 0.452f
C622 n7 m3_12600_1156# 0.181f
C623 n6 m2_41500_1156# 1.13f
C624 n2 n6 0.39f
C625 top m3_1100_1156# 0.187f
C626 m3_18000_1156# m3_19100_1156# 0.148f
C627 top n0 0.418f
C628 m2_40200_1156# m3_41200_1156# 0.0061f
C629 top via23_4_702/m2_1_40# 0.341f
C630 via23_4_439/m2_1_40# n5 0.523f
C631 via23_4_709/m2_1_40# m3_37500_1156# 0.247f
C632 via23_4_90/m2_1_40# m3_10000_1156# 0.247f
C633 via23_4_96/m2_1_40# m2_800_1156# 0.251f
C634 m2_16400_1156# m3_16500_1156# 2.11f
C635 n7 m3_41400_1156# 1.99f
C636 via23_4_249/m2_1_40# m3_7400_1156# 0.247f
C637 top m3_30800_1156# 0.221f
C638 n2 via23_4_23/m2_1_40# 0.169f
C639 ndum via23_4_455/m2_1_40# 0.381f
C640 m2_6000_1156# n4 3.19e-19
C641 via23_4_3/m2_1_40# n1 9.38e-20
C642 via23_4_448/m2_1_40# n7 1.18e-19
C643 via23_4_9/m2_1_40# m2_19000_1156# 0.251f
C644 m2_31100_1156# n5 0.002f
C645 via23_4_641/m2_1_40# m2_42800_1156# 0.251f
C646 top m2_24600_1156# 0.267f
C647 m3_8900_1156# m3_10000_1156# 0.148f
C648 via23_4_589/m2_1_40# m2_24600_1156# 0.251f
C649 m2_31100_1156# m3_32100_1156# 0.0061f
C650 n2 m3_20400_1156# 3.43f
C651 via23_4_228/m2_1_40# via23_4_220/m2_1_40# 0.199f
C652 top via23_4_333/m2_1_40# 0.347f
C653 via23_4_94/m2_1_40# m3_4800_1156# 0.247f
C654 via23_4_229/m2_1_40# top 0.347f
C655 via23_4_20/m2_1_40# m2_12500_1156# 0.251f
C656 via23_4_455/m2_1_40# n5 1.57e-19
C657 top via23_4_459/m2_1_40# 0.14f
C658 top via23_4_3/m2_1_40# 0.14f
C659 via23_4_89/m2_1_40# m3_11300_1156# 0.123f
C660 via23_4_449/m2_1_40# m3_29500_1156# 0.123f
C661 n0 m2_6000_1156# 6.36e-20
C662 via23_4_346/m2_1_40# m2_19000_1156# 0.251f
C663 m3_16500_1156# n5 1.98f
C664 top m3_11300_1156# 0.187f
C665 via23_4_380/m2_1_40# n6 0.512f
C666 n2 via23_4_20/m2_1_40# 0.169f
C667 n7 m2_3400_1156# 1.13f
C668 n2 m3_2200_1156# 0.021f
C669 via23_4_90/m2_1_40# n4 2.85e-19
C670 n6 n3 0.313f
C671 n6 m3_37500_1156# 0.188f
C672 via23_4_96/m2_1_40# m3_900_1156# 0.247f
C673 top m3_40100_1156# 0.187f
C674 m3_38600_1156# m3_38800_1156# 3.35f
C675 ndum via23_4_584/m2_1_40# 0.247f
C676 via23_4_3/m2_1_40# m3_17800_1156# 0.247f
C677 n7 m3_3700_1156# 4.08f
C678 via23_4_590/m2_1_40# m3_26900_1156# 0.247f
C679 via23_4_710/m2_1_40# n7 0.452f
C680 n6 via23_4_331/m2_1_40# 0.452f
C681 m2_36300_1156# m3_36200_1156# 2.11f
C682 via23_4_378/m2_1_40# m3_34700_1156# 0.247f
C683 via23_4_23/m2_1_40# n3 4.28e-19
C684 m2_12500_1156# m3_11500_1156# 0.0061f
C685 via23_4_218/m2_1_40# top 0.347f
C686 via23_4_598/m2_1_40# m3_27100_1156# 0.247f
C687 m2_16400_1156# n1 8.05e-20
C688 m3_27100_1156# n5 1.99f
C689 m3_20400_1156# n3 0.174f
C690 via23_4_228/m2_1_40# m2_800_1156# 0.251f
C691 m2_2100_1156# n1 8.05e-20
C692 m3_29500_1156# m3_29700_1156# 3.35f
C693 n7 m2_28500_1156# 2.42f
C694 n6 m2_13800_1156# 1.43e-19
C695 via23_4_87/m2_1_40# n7 1.18e-19
C696 top via23_4_368/m2_1_40# 0.14f
C697 top m2_16400_1156# 0.267f
C698 ndum n1 3.59f
C699 n6 via23_4_678/m2_1_40# 0.452f
C700 m2_27200_1156# m3_26900_1156# 0.181f
C701 n2 m3_11500_1156# 0.021f
C702 m2_800_1156# n4 3.19e-19
C703 top m2_2100_1156# 0.267f
C704 top via23_4_251/m2_1_40# 0.347f
C705 via23_4_599/m2_1_40# m3_29500_1156# 0.123f
C706 via23_4_20/m2_1_40# n3 4.28e-19
C707 n7 m3_13900_1156# 2.16f
C708 n7 via23_4_91/m2_1_40# 1.18e-19
C709 ndum top 0.414f
C710 via23_4_675/m2_1_40# m3_33400_1156# 0.247f
C711 top via23_4_712/m2_1_40# 0.347f
C712 n2 via23_4_21/m2_1_40# 0.169f
C713 n2 via23_4_22/m2_1_40# 0.169f
C714 top m3_2400_1156# 0.187f
C715 m3_19100_1156# m3_19300_1156# 3.35f
C716 m2_41500_1156# m3_41200_1156# 0.181f
C717 n5 n1 0.0771f
C718 via23_4_96/m2_1_40# n6 1.52e-19
C719 top via23_4_369/m2_1_40# 0.14f
C720 m2_8600_1156# m3_7600_1156# 0.0061f
C721 m2_4700_1156# m3_4800_1156# 2.11f
C722 n0 m2_800_1156# 6.36e-20
C723 m2_8600_1156# n1 8.05e-20
C724 via23_4_89/m2_1_40# n5 0.452f
C725 via23_4_439/m2_1_40# m3_33400_1156# 0.247f
C726 m2_800_1156# m3_1100_1156# 0.181f
C727 m3_19100_1156# n4 0.181f
C728 via23_4_598/m2_1_40# top 0.347f
C729 m2_17700_1156# m3_16700_1156# 0.023f
C730 n7 m3_42700_1156# 0.181f
C731 via23_4_87/m2_1_40# m3_6300_1156# 0.247f
C732 top n5 8.2f
C733 top m3_32100_1156# 0.187f
C734 m2_7300_1156# n4 3.19e-19
C735 top m2_8600_1156# 0.267f
C736 via23_4_332/m2_1_40# m3_13900_1156# 0.247f
C737 via23_4_228/m2_1_40# m3_900_1156# 0.247f
C738 n7 via23_4_378/m2_1_40# 0.452f
C739 n6 m2_23300_1156# 1.43e-19
C740 m2_32400_1156# n5 2.39f
C741 via23_4_446/m2_1_40# n5 0.0714f
C742 m2_32400_1156# m3_32100_1156# 0.181f
C743 m3_10000_1156# m3_10200_1156# 3.35f
C744 via23_4_448/m2_1_40# m3_27100_1156# 0.247f
C745 via23_4_446/m2_1_40# m3_32100_1156# 0.247f
C746 via23_4_588/m2_1_40# m3_23200_1156# 0.247f
C747 ndum m2_6000_1156# 3.15e-20
C748 n2 m2_17700_1156# 0.00855f
C749 n7 m3_24500_1156# 1.98f
C750 n0 m2_7300_1156# 6.36e-20
C751 top m3_12600_1156# 0.221f
C752 n6 via23_4_103/m2_1_40# 1.52e-19
C753 via23_4_429/m2_1_40# m3_42700_1156# 0.247f
C754 via23_4_600/m2_1_40# m3_30800_1156# 0.123f
C755 via23_4_95/m2_1_40# m3_5000_1156# 0.247f
C756 m2_6000_1156# n5 2.05e-19
C757 via23_4_94/m2_1_40# m2_4700_1156# 0.251f
C758 m3_900_1156# m3_1100_1156# 3.35f
C759 via23_4_21/m2_1_40# n3 4.28e-19
C760 n2 m3_3500_1156# 0.021f
C761 n6 m3_38800_1156# 0.00746f
C762 via23_4_22/m2_1_40# n3 4.28e-19
C763 via23_4_331/m2_1_40# m3_11500_1156# 0.247f
C764 top m3_41400_1156# 0.187f
C765 m3_38800_1156# m3_39900_1156# 0.148f
C766 via23_4_380/m2_1_40# m2_36300_1156# 0.0256f
C767 n7 m3_5000_1156# 4.08f
C768 via23_4_705/m2_1_40# via23_4_635/m2_1_40# 0.199f
C769 via23_4_96/m2_1_40# via23_4_128/m2_1_40# 0.199f
C770 via23_4_676/m2_1_40# m3_33600_1156# 0.247f
C771 via23_4_448/m2_1_40# top 0.14f
C772 top via23_4_345/m2_1_40# 0.347f
C773 via23_4_447/m2_1_40# m2_29800_1156# 0.251f
C774 m2_12500_1156# m3_12800_1156# 0.181f
C775 n7 m3_34700_1156# 4.08f
C776 m3_28400_1156# n5 0.19f
C777 via23_4_458/m2_1_40# n5 0.0714f
C778 via23_4_251/m2_1_40# m3_8900_1156# 0.247f
C779 top m3_23200_1156# 0.187f
C780 m2_3400_1156# n1 8.05e-20
C781 m3_29700_1156# m3_30800_1156# 0.354f
C782 n6 n4 0.318f
C783 via23_4_90/m2_1_40# n5 2.03e-19
C784 n7 m2_29800_1156# 3.52f
C785 n6 m2_15100_1156# 1.43e-19
C786 via23_4_21/m2_1_40# m2_13800_1156# 0.251f
C787 m2_17700_1156# n3 5.59e-19
C788 n2 m3_12800_1156# 0.021f
C789 m2_27200_1156# m3_28200_1156# 0.0061f
C790 via23_4_1/m2_1_40# m2_20300_1156# 0.251f
C791 top m2_3400_1156# 0.267f
C792 via23_4_345/m2_1_40# m3_17800_1156# 0.247f
C793 via23_4_103/m2_1_40# m3_2200_1156# 0.247f
C794 via23_4_230/m2_1_40# top 0.347f
C795 n7 m3_15200_1156# 1.98f
C796 via23_4_23/m2_1_40# n4 2.85e-19
C797 n6 n0 0.0802f
C798 via23_4_678/m2_1_40# m2_36300_1156# 0.0256f
C799 top m3_3700_1156# 0.187f
C800 via23_4_326/m2_1_40# m3_11300_1156# 0.123f
C801 m3_19300_1156# m3_20400_1156# 0.148f
C802 m2_41500_1156# m3_42500_1156# 0.0061f
C803 ndum m2_800_1156# 3.15e-20
C804 m2_8600_1156# m3_8900_1156# 0.181f
C805 top via23_4_710/m2_1_40# 0.347f
C806 via23_4_347/m2_1_40# m3_19300_1156# 0.247f
C807 m3_20400_1156# n4 1.98f
C808 m2_17700_1156# m3_18000_1156# 0.181f
C809 via23_4_347/m2_1_40# n4 0.452f
C810 n7 via23_4_447/m2_1_40# 0.452f
C811 via23_4_87/m2_1_40# n1 9.38e-20
C812 top m3_33400_1156# 0.187f
C813 via23_4_95/m2_1_40# n7 0.452f
C814 m2_800_1156# n5 2.05e-19
C815 via23_4_245/m2_1_40# m3_5000_1156# 0.247f
C816 n2 via23_4_88/m2_1_40# 0.169f
C817 n6 m2_24600_1156# 1.43e-19
C818 m2_33700_1156# n5 1.13f
C819 via23_4_635/m2_1_40# m2_42800_1156# 0.251f
C820 top m2_28500_1156# 0.267f
C821 m3_10200_1156# m3_11300_1156# 0.148f
C822 m2_32400_1156# m3_33400_1156# 0.0061f
C823 top via23_4_87/m2_1_40# 0.14f
C824 via23_4_20/m2_1_40# n4 2.85e-19
C825 n0 m3_20400_1156# 3.28e-19
C826 n2 m3_24300_1156# 4.32e-19
C827 n6 via23_4_459/m2_1_40# 1.52e-19
C828 via23_4_91/m2_1_40# n1 9.38e-20
C829 n6 via23_4_3/m2_1_40# 0.452f
C830 via23_4_449/m2_1_40# n5 0.0714f
C831 ndum m2_7300_1156# 3.15e-20
C832 n2 m2_19000_1156# 0.00869f
C833 n7 m3_25800_1156# 0.181f
C834 n6 m3_11300_1156# 0.181f
C835 top m3_13900_1156# 0.187f
C836 top via23_4_91/m2_1_40# 0.14f
C837 m2_7300_1156# n5 2.05e-19
C838 via23_4_419/m2_1_40# top 0.216f
C839 m3_1100_1156# m3_2200_1156# 0.148f
C840 n2 m3_4800_1156# 0.021f
C841 via23_4_332/m2_1_40# n7 0.452f
C842 n6 m3_40100_1156# 1.99f
C843 top m3_42700_1156# 0.187f
C844 m3_39900_1156# m3_40100_1156# 3.35f
C845 via23_4_460/m2_1_40# m2_24600_1156# 0.251f
C846 via23_4_88/m2_1_40# m3_8700_1156# 0.247f
C847 via23_4_439/m2_1_40# n7 1.18e-19
C848 via23_4_379/m2_1_40# m3_34900_1156# 0.123f
C849 top via23_4_378/m2_1_40# 0.14f
C850 m2_37600_1156# m3_37500_1156# 2.11f
C851 via23_4_366/m2_1_40# m3_41400_1156# 0.247f
C852 via23_4_88/m2_1_40# n3 4.28e-19
C853 m2_13800_1156# m3_12800_1156# 0.0061f
C854 n7 m3_36000_1156# 4.08f
C855 m3_29700_1156# n5 0.00889f
C856 via23_4_326/m2_1_40# n5 0.452f
C857 top m3_24500_1156# 0.187f
C858 m3_30800_1156# m3_31000_1156# 3.35f
C859 via23_4_229/m2_1_40# m3_2200_1156# 0.247f
C860 via23_4_589/m2_1_40# m3_24500_1156# 0.247f
C861 via23_4_21/m2_1_40# n4 2.85e-19
C862 via23_4_22/m2_1_40# n4 2.85e-19
C863 via23_4_704/m2_1_40# via23_4_705/m2_1_40# 0.199f
C864 n7 m2_31100_1156# 1.13f
C865 n6 m2_16400_1156# 1.13f
C866 via23_4_368/m2_1_40# n6 0.0598f
C867 via23_4_22/m2_1_40# m2_15100_1156# 0.251f
C868 m2_19000_1156# n3 5.59e-19
C869 via23_4_368/m2_1_40# m3_39900_1156# 0.247f
C870 n6 m2_2100_1156# 1.13f
C871 n2 m3_14100_1156# 0.021f
C872 m2_28500_1156# m3_28400_1156# 2.11f
C873 n7 via23_4_455/m2_1_40# 9.11e-20
C874 via23_4_711/m2_1_40# m2_40200_1156# 0.251f
C875 via23_4_245/m2_1_40# n7 0.452f
C876 n2 via23_4_94/m2_1_40# 0.169f
C877 ndum n6 0.0782f
C878 n2 m2_9900_1156# 0.00855f
C879 via23_4_354/m2_1_40# n1 0.251f
C880 via23_4_369/m2_1_40# n6 0.512f
C881 n6 m3_2400_1156# 4.08f
C882 m3_10200_1156# n5 4.08f
C883 n2 via23_4_9/m2_1_40# 0.169f
C884 top m3_5000_1156# 0.187f
C885 m2_42800_1156# m3_42500_1156# 0.181f
C886 via23_4_23/m2_1_40# m2_16400_1156# 0.251f
C887 top via23_4_354/m2_1_40# 0.347f
C888 n6 n5 16.1f
C889 m2_19000_1156# m3_18000_1156# 0.0061f
C890 n6 m3_32100_1156# 4.08f
C891 n6 m2_8600_1156# 1.43e-19
C892 m2_17700_1156# n4 3.19e-19
C893 top m3_34700_1156# 0.187f
C894 via23_4_367/m2_1_40# m2_42800_1156# 0.251f
C895 ndum m3_20400_1156# 1.62e-19
C896 top m2_29800_1156# 0.267f
C897 m3_11300_1156# m3_11500_1156# 3.35f
C898 m2_33700_1156# m3_33400_1156# 0.181f
C899 via23_4_23/m2_1_40# n5 0.452f
C900 top via23_4_117/m2_1_40# 0.216f
C901 n0 m2_17700_1156# 6.36e-20
C902 n2 m2_20300_1156# 0.257f
C903 m2_6000_1156# m3_5000_1156# 0.0061f
C904 n6 m3_12600_1156# 1.01f
C905 m2_2100_1156# m3_2200_1156# 2.11f
C906 top m3_15200_1156# 0.187f
C907 via23_4_94/m2_1_40# n3 4.28e-19
C908 via23_4_449/m2_1_40# m2_28500_1156# 0.251f
C909 via23_4_704/m2_1_40# m2_42800_1156# 0.251f
C910 via23_4_460/m2_1_40# n5 0.0714f
C911 m2_9900_1156# n3 5.59e-19
C912 m3_2200_1156# m3_2400_1156# 3.35f
C913 via23_4_95/m2_1_40# n1 9.38e-20
C914 m2_23300_1156# m3_24300_1156# 0.0061f
C915 n2 m3_6100_1156# 0.021f
C916 via23_4_9/m2_1_40# n3 4.28e-19
C917 n6 m3_41400_1156# 0.181f
C918 via23_4_381/m2_1_40# n7 0.452f
C919 m3_40100_1156# m3_41200_1156# 0.148f
C920 via23_4_20/m2_1_40# n5 2.03e-19
C921 top via23_4_447/m2_1_40# 0.14f
C922 n7 m3_7600_1156# 4.08f
C923 n7 n1 10.3f
C924 top via23_4_95/m2_1_40# 0.14f
C925 via23_4_87/m2_1_40# m2_7300_1156# 0.251f
C926 via23_4_448/m2_1_40# n6 1.52e-19
C927 n6 via23_4_345/m2_1_40# 0.452f
C928 n7 via23_4_677/m2_1_40# 0.452f
C929 n7 via23_4_89/m2_1_40# 1.18e-19
C930 via23_4_3/m2_1_40# m2_17700_1156# 0.251f
C931 n2 via23_4_1/m2_1_40# 0.169f
C932 n2 m2_4700_1156# 0.00855f
C933 top via23_4_199/m2_1_40# 0.216f
C934 via23_4_419/m2_1_40# via23_4_641/m2_1_40# 0.199f
C935 top n7 32.8f
C936 m2_13800_1156# m3_14100_1156# 0.181f
C937 via23_4_589/m2_1_40# n7 0.452f
C938 via23_4_378/m2_1_40# m2_33700_1156# 0.251f
C939 m3_31000_1156# n5 0.00889f
C940 via23_4_9/m2_1_40# m3_18000_1156# 0.123f
C941 via23_4_641/m2_1_40# m3_42700_1156# 0.247f
C942 top m3_25800_1156# 0.187f
C943 m3_31000_1156# m3_32100_1156# 0.148f
C944 n7 m2_32400_1156# 1.05e-19
C945 n7 via23_4_446/m2_1_40# 1.18e-19
C946 via23_4_20/m2_1_40# m3_12600_1156# 0.123f
C947 m2_25900_1156# n5 0.002f
C948 m2_20300_1156# n3 1.09f
C949 n6 m2_3400_1156# 2.39f
C950 n2 m3_15400_1156# 0.021f
C951 via23_4_230/m2_1_40# n6 0.452f
C952 via23_4_346/m2_1_40# m3_18000_1156# 0.123f
C953 top via23_4_332/m2_1_40# 0.347f
C954 via23_4_95/m2_1_40# m2_6000_1156# 0.251f
C955 n7 m3_17800_1156# 0.181f
C956 top via23_4_675/m2_1_40# 0.347f
C957 n2 m2_11200_1156# 0.00855f
C958 via23_4_88/m2_1_40# n4 2.85e-19
C959 top m3_6300_1156# 0.187f
C960 via23_4_599/m2_1_40# m2_28500_1156# 0.251f
C961 via23_4_369/m2_1_40# m3_41200_1156# 0.247f
C962 via23_4_429/m2_1_40# top 0.216f
C963 via23_4_250/m2_1_40# m3_8700_1156# 0.247f
C964 via23_4_439/m2_1_40# top 0.14f
C965 n7 m2_6000_1156# 2.39f
C966 via23_4_675/m2_1_40# m2_32400_1156# 0.251f
C967 via23_4_677/m2_1_40# m3_36000_1156# 0.247f
C968 via23_4_710/m2_1_40# m3_39900_1156# 0.247f
C969 m3_24300_1156# n4 4.08f
C970 via23_4_21/m2_1_40# n5 2.03e-19
C971 via23_4_22/m2_1_40# n5 2.03e-19
C972 m2_19000_1156# m3_19300_1156# 0.181f
C973 n6 m3_33400_1156# 0.00746f
C974 via23_4_439/m2_1_40# m2_32400_1156# 0.251f
C975 m2_19000_1156# n4 1.13f
C976 top m3_36000_1156# 0.187f
C977 via23_4_1/m2_1_40# n3 4.28e-19
C978 m2_4700_1156# n3 5.59e-19
C979 via23_4_455/m2_1_40# n1 0.251f
C980 n6 m2_28500_1156# 1.43e-19
C981 n6 via23_4_87/m2_1_40# 0.452f
C982 top m2_31100_1156# 0.267f
C983 m3_11500_1156# m3_12600_1156# 0.354f
C984 m2_33700_1156# m3_34700_1156# 0.0061f
C985 ndum m2_17700_1156# 3.15e-20
C986 top via23_4_455/m2_1_40# 0.14f
C987 via23_4_245/m2_1_40# top 0.347f
C988 n7 m3_28400_1156# 1.98f
C989 n0 m2_19000_1156# 6.36e-20
C990 n7 via23_4_458/m2_1_40# 1.18e-19
C991 via23_4_446/m2_1_40# m2_31100_1156# 0.251f
C992 m2_6000_1156# m3_6300_1156# 0.181f
C993 m2_9900_1156# m3_10000_1156# 2.11f
C994 via23_4_117/m2_1_40# m2_800_1156# 0.251f
C995 n6 via23_4_91/m2_1_40# 0.452f
C996 top m3_16500_1156# 0.187f
C997 via23_4_90/m2_1_40# n7 0.452f
C998 via23_4_458/m2_1_40# m3_25800_1156# 0.247f
C999 via23_4_702/m2_1_40# via23_4_704/m2_1_40# 0.199f
C1000 m2_17700_1156# n5 2.05e-19
C1001 m2_11200_1156# n3 5.59e-19
C1002 m2_24600_1156# m3_24300_1156# 0.181f
C1003 m3_2400_1156# m3_3500_1156# 0.148f
C1004 n2 m3_7400_1156# 0.021f
C1005 via23_4_600/m2_1_40# m2_29800_1156# 0.251f
C1006 via23_4_601/m2_1_40# m3_32100_1156# 0.247f
C1007 m3_41200_1156# m3_41400_1156# 3.35f
C1008 via23_4_459/m2_1_40# m3_24300_1156# 0.247f
C1009 via23_4_642/m2_1_40# m2_42800_1156# 0.251f
C1010 n7 m3_8900_1156# 4.08f
C1011 via23_4_584/m2_1_40# n1 0.251f
C1012 n6 via23_4_378/m2_1_40# 0.0598f
C1013 m2_38900_1156# m3_38800_1156# 2.11f
C1014 via23_4_245/m2_1_40# m2_6000_1156# 0.251f
C1015 top via23_4_588/m2_1_40# 0.347f
C1016 via23_4_584/m2_1_40# top 0.347f
C1017 via23_4_94/m2_1_40# n4 2.85e-19
C1018 m2_15100_1156# m3_14100_1156# 0.0061f
C1019 n7 m3_38600_1156# 4.08f
C1020 m3_32300_1156# n5 1.99f
C1021 via23_4_199/m2_1_40# m2_800_1156# 0.251f
C1022 top m3_27100_1156# 0.187f
C1023 m2_9900_1156# n4 3.19e-19
C1024 m3_32100_1156# m3_32300_1156# 3.35f
C1025 via23_4_117/m2_1_40# m3_900_1156# 0.247f
C1026 n7 m2_800_1156# 1.13f
C1027 via23_4_9/m2_1_40# n4 2.85e-19
C1028 n7 m2_33700_1156# 2.39f
C1029 via23_4_598/m2_1_40# m2_27200_1156# 0.251f
C1030 m2_27200_1156# n5 2.39f
C1031 via23_4_366/m2_1_40# n7 0.503f
C1032 m2_29800_1156# m3_29700_1156# 2.11f
C1033 n2 m3_16700_1156# 0.021f
C1034 via23_4_449/m2_1_40# n7 0.227f
C1035 n0 m2_9900_1156# 6.36e-20
C1036 n2 via23_4_2/m2_1_40# 0.352f
C1037 via23_4_381/m2_1_40# top 0.14f
C1038 n7 m3_19100_1156# 1.98f
C1039 n2 m2_12500_1156# 0.00855f
C1040 via23_4_89/m2_1_40# n1 9.38e-20
C1041 via23_4_345/m2_1_40# m2_17700_1156# 0.251f
C1042 via23_4_600/m2_1_40# n7 0.452f
C1043 via23_4_712/m2_1_40# m3_42500_1156# 0.247f
C1044 top m3_7600_1156# 0.187f
C1045 top n1 0.983f
C1046 top via23_4_677/m2_1_40# 0.347f
C1047 via23_4_111/m2_1_40# via23_4_117/m2_1_40# 0.199f
C1048 n7 m2_7300_1156# 1.13f
C1049 top via23_4_89/m2_1_40# 0.14f
C1050 via23_4_460/m2_1_40# m3_24500_1156# 0.247f
C1051 via23_4_380/m2_1_40# m3_36200_1156# 0.123f
C1052 m2_20300_1156# m3_19300_1156# 0.0061f
C1053 n6 m3_34700_1156# 0.00746f
C1054 via23_4_333/m2_1_40# m3_14100_1156# 0.247f
C1055 top m3_37300_1156# 0.187f
C1056 top via23_4_589/m2_1_40# 0.347f
C1057 m2_20300_1156# n4 2.39f
C1058 via23_4_199/m2_1_40# m3_900_1156# 0.247f
C1059 via23_4_447/m2_1_40# m3_29700_1156# 0.247f
C1060 n7 m3_900_1156# 0.181f
C1061 via23_4_218/m2_1_40# m3_4800_1156# 0.247f
C1062 n7 via23_4_709/m2_1_40# 0.452f
C1063 n6 m2_29800_1156# 1.43e-19
C1064 top via23_4_446/m2_1_40# 0.14f
C1065 top m2_32400_1156# 0.267f
C1066 m3_12600_1156# m3_12800_1156# 3.35f
C1067 m2_35000_1156# m3_34700_1156# 0.181f
C1068 ndum m2_19000_1156# 3.15e-20
C1069 via23_4_88/m2_1_40# n5 2.03e-19
C1070 via23_4_334/m2_1_40# m3_15400_1156# 0.247f
C1071 n7 m3_29700_1156# 2.16f
C1072 via23_4_21/m2_1_40# m3_13900_1156# 0.247f
C1073 via23_4_448/m2_1_40# m2_27200_1156# 0.251f
C1074 n0 m2_20300_1156# 2e-19
C1075 m2_7300_1156# m3_6300_1156# 0.0061f
C1076 m3_24300_1156# n5 0.00889f
C1077 via23_4_88/m2_1_40# m2_8600_1156# 0.251f
C1078 m2_3400_1156# m3_3500_1156# 2.11f
C1079 m2_6000_1156# n1 8.05e-20
C1080 top m3_17800_1156# 0.187f
C1081 via23_4_230/m2_1_40# m3_3500_1156# 0.247f
C1082 via23_4_1/m2_1_40# m3_19300_1156# 0.247f
C1083 via23_4_199/m2_1_40# via23_4_111/m2_1_40# 0.199f
C1084 m2_19000_1156# n5 2.05e-19
C1085 via23_4_2/m2_1_40# n3 0.453f
C1086 m2_12500_1156# n3 5.59e-19
C1087 via23_4_1/m2_1_40# n4 0.453f
C1088 m3_3500_1156# m3_3700_1156# 3.35f
C1089 m2_4700_1156# n4 3.19e-19
C1090 top m2_6000_1156# 0.267f
C1091 m2_24600_1156# m3_25600_1156# 0.0061f
C1092 via23_4_599/m2_1_40# n7 0.227f
C1093 n2 m3_8700_1156# 0.021f
C1094 via23_4_678/m2_1_40# m3_36200_1156# 0.123f
C1095 n6 via23_4_447/m2_1_40# 1.52e-19
C1096 m3_41400_1156# m3_42500_1156# 0.148f
C1097 via23_4_95/m2_1_40# n6 1.52e-19
C1098 via23_4_331/m2_1_40# m2_12500_1156# 0.251f
C1099 n2 n3 19.6f
C1100 n0 m2_4700_1156# 6.36e-20
C1101 n6 n7 20.9f
C1102 top via23_4_220/m2_1_40# 0.219f
C1103 via23_4_90/m2_1_40# n1 9.38e-20
C1104 m2_15100_1156# m3_15400_1156# 0.181f
C1105 n7 m3_39900_1156# 4.08f
C1106 m3_33600_1156# n5 0.181f
C1107 via23_4_635/m2_1_40# m3_42700_1156# 0.247f
C1108 n6 m3_25800_1156# 1.98f
C1109 top via23_4_458/m2_1_40# 0.14f
C1110 top m3_28400_1156# 0.187f
C1111 m2_11200_1156# n4 3.19e-19
C1112 m3_32300_1156# m3_33400_1156# 0.148f
C1113 n7 m2_35000_1156# 3.52f
C1114 via23_4_90/m2_1_40# top 0.14f
C1115 via23_4_251/m2_1_40# m2_9900_1156# 0.251f
C1116 n7 via23_4_23/m2_1_40# 1.18e-19
C1117 n2 m3_18000_1156# 0.021f
C1118 via23_4_91/m2_1_40# m3_3500_1156# 0.247f
C1119 via23_4_128/m2_1_40# via23_4_117/m2_1_40# 0.199f
C1120 ndum m2_9900_1156# 3.15e-20
C1121 via23_4_368/m2_1_40# m2_38900_1156# 0.251f
C1122 n0 m2_11200_1156# 6.36e-20
C1123 n2 m2_13800_1156# 0.00855f
C1124 via23_4_381/m2_1_40# m3_38600_1156# 0.247f
C1125 n6 m3_6300_1156# 4.08f
C1126 top m3_8900_1156# 0.187f
C1127 m3_23200_1156# m3_24300_1156# 0.148f
C1128 via23_4_94/m2_1_40# n5 2.03e-19
C1129 n7 via23_4_460/m2_1_40# 0.452f
C1130 via23_4_439/m2_1_40# n6 1.52e-19
C1131 m2_9900_1156# n5 1.13f
C1132 m2_800_1156# n1 8.05e-20
C1133 via23_4_9/m2_1_40# n5 2.03e-19
C1134 n6 m3_36000_1156# 0.00746f
C1135 top m3_38600_1156# 0.187f
C1136 n2 via23_4_96/m2_1_40# 0.169f
C1137 n7 via23_4_20/m2_1_40# 1.18e-19
C1138 top m2_800_1156# 0.267f
C1139 n7 m3_2200_1156# 1.98f
C1140 n6 m2_31100_1156# 2.39f
C1141 top m2_33700_1156# 0.267f
C1142 m3_12800_1156# m3_13900_1156# 0.148f
C1143 m2_35000_1156# m3_36000_1156# 0.0061f
C1144 top via23_4_366/m2_1_40# 0.14f
C1145 n6 via23_4_455/m2_1_40# 1.17e-19
C1146 via23_4_449/m2_1_40# top 0.14f
C1147 ndum m2_20300_1156# 1e-19
C1148 n7 m3_31000_1156# 0.181f
C1149 via23_4_200/m2_1_40# via23_4_199/m2_1_40# 0.199f
C1150 m2_11200_1156# m3_11300_1156# 2.11f
C1151 n1 VSUBS 4.59f
C1152 n5 VSUBS 20.3f
C1153 n4 VSUBS 9.84f
C1154 n3 VSUBS 7.1f
C1155 m3_42700_1156# VSUBS 1.97f
C1156 m3_42500_1156# VSUBS 1.18f
C1157 m3_41400_1156# VSUBS 1.17f
C1158 m3_41200_1156# VSUBS 1.17f
C1159 m3_40100_1156# VSUBS 1.17f
C1160 m3_39900_1156# VSUBS 1.17f
C1161 m3_38800_1156# VSUBS 1.17f
C1162 m3_38600_1156# VSUBS 1.17f
C1163 m3_37500_1156# VSUBS 1.17f
C1164 m3_37300_1156# VSUBS 1.17f
C1165 m3_36200_1156# VSUBS 1.17f
C1166 m3_36000_1156# VSUBS 1.17f
C1167 m3_34900_1156# VSUBS 1.17f
C1168 m3_34700_1156# VSUBS 1.17f
C1169 m3_33600_1156# VSUBS 1.17f
C1170 m3_33400_1156# VSUBS 1.17f
C1171 m3_32300_1156# VSUBS 1.17f
C1172 m3_32100_1156# VSUBS 1.16f
C1173 m3_31000_1156# VSUBS 1.17f
C1174 m3_30800_1156# VSUBS 1.16f
C1175 m3_29700_1156# VSUBS 1.17f
C1176 m3_29500_1156# VSUBS 1.16f
C1177 m3_28400_1156# VSUBS 1.17f
C1178 m3_28200_1156# VSUBS 1.16f
C1179 m3_27100_1156# VSUBS 1.17f
C1180 m3_26900_1156# VSUBS 1.16f
C1181 m3_25800_1156# VSUBS 1.17f
C1182 m3_25600_1156# VSUBS 1.16f
C1183 m3_24500_1156# VSUBS 1.17f
C1184 m3_24300_1156# VSUBS 1.16f
C1185 m3_23200_1156# VSUBS 1.17f
C1186 m3_20400_1156# VSUBS 1.16f
C1187 m3_19300_1156# VSUBS 1.16f
C1188 m3_19100_1156# VSUBS 1.16f
C1189 m3_18000_1156# VSUBS 1.16f
C1190 m3_17800_1156# VSUBS 1.16f
C1191 m3_16700_1156# VSUBS 1.16f
C1192 m3_16500_1156# VSUBS 1.16f
C1193 m3_15400_1156# VSUBS 1.16f
C1194 m3_15200_1156# VSUBS 1.16f
C1195 m3_14100_1156# VSUBS 1.16f
C1196 m3_13900_1156# VSUBS 1.16f
C1197 m3_12800_1156# VSUBS 1.16f
C1198 m3_12600_1156# VSUBS 1.16f
C1199 m3_11500_1156# VSUBS 1.16f
C1200 m3_11300_1156# VSUBS 1.16f
C1201 m3_10200_1156# VSUBS 1.16f
C1202 m3_10000_1156# VSUBS 1.16f
C1203 m3_8900_1156# VSUBS 1.16f
C1204 m3_8700_1156# VSUBS 1.16f
C1205 m3_7600_1156# VSUBS 1.16f
C1206 m3_7400_1156# VSUBS 1.16f
C1207 m3_6300_1156# VSUBS 1.16f
C1208 m3_6100_1156# VSUBS 1.16f
C1209 m3_5000_1156# VSUBS 1.16f
C1210 m3_4800_1156# VSUBS 1.16f
C1211 m3_3700_1156# VSUBS 1.16f
C1212 m3_3500_1156# VSUBS 1.16f
C1213 m3_2400_1156# VSUBS 1.16f
C1214 m3_2200_1156# VSUBS 1.16f
C1215 m3_1100_1156# VSUBS 1.16f
C1216 m3_900_1156# VSUBS 1.95f
C1217 m2_42800_1156# VSUBS 2.41f
C1218 m2_41500_1156# VSUBS 1.8f
C1219 m2_40200_1156# VSUBS 1.8f
C1220 m2_38900_1156# VSUBS 1.8f
C1221 m2_37600_1156# VSUBS 1.8f
C1222 m2_36300_1156# VSUBS 1.8f
C1223 m2_35000_1156# VSUBS 1.8f
C1224 m2_33700_1156# VSUBS 1.8f
C1225 m2_32400_1156# VSUBS 1.8f
C1226 m2_31100_1156# VSUBS 1.8f
C1227 m2_29800_1156# VSUBS 1.8f
C1228 m2_28500_1156# VSUBS 1.8f
C1229 m2_27200_1156# VSUBS 1.8f
C1230 m2_25900_1156# VSUBS 1.8f
C1231 m2_24600_1156# VSUBS 1.8f
C1232 m2_23300_1156# VSUBS 1.79f
C1233 m2_20300_1156# VSUBS 1.79f
C1234 m2_19000_1156# VSUBS 1.8f
C1235 m2_17700_1156# VSUBS 1.8f
C1236 m2_16400_1156# VSUBS 1.8f
C1237 m2_15100_1156# VSUBS 1.8f
C1238 m2_13800_1156# VSUBS 1.8f
C1239 m2_12500_1156# VSUBS 1.8f
C1240 m2_11200_1156# VSUBS 1.8f
C1241 m2_9900_1156# VSUBS 1.8f
C1242 m2_8600_1156# VSUBS 1.8f
C1243 m2_7300_1156# VSUBS 1.8f
C1244 m2_6000_1156# VSUBS 1.8f
C1245 m2_4700_1156# VSUBS 1.8f
C1246 m2_3400_1156# VSUBS 1.8f
C1247 m2_2100_1156# VSUBS 1.8f
C1248 m2_800_1156# VSUBS 2.41f
C1249 via23_4_326/m2_1_40# VSUBS 0.548f
C1250 via23_4_414/m2_1_40# VSUBS 0.427f
C1251 via23_4_447/m2_1_40# VSUBS 0.339f
C1252 via23_4_458/m2_1_40# VSUBS 0.339f
C1253 via23_4_446/m2_1_40# VSUBS 0.339f
C1254 via23_4_460/m2_1_40# VSUBS 0.339f
C1255 via23_4_220/m2_1_40# VSUBS 0.427f
C1256 via23_4_9/m2_1_40# VSUBS 0.418f
C1257 via23_4_459/m2_1_40# VSUBS 0.327f
C1258 via23_4_641/m2_1_40# VSUBS 0.427f
C1259 via23_4_251/m2_1_40# VSUBS 0.425f
C1260 via23_4_455/m2_1_40# VSUBS 0.283f
C1261 via23_4_635/m2_1_40# VSUBS 0.427f
C1262 via23_4_250/m2_1_40# VSUBS 0.425f
C1263 n0 VSUBS 3.21f
C1264 via23_4_3/m2_1_40# VSUBS 0.295f
C1265 via23_4_642/m2_1_40# VSUBS 0.427f
C1266 via23_4_709/m2_1_40# VSUBS 0.425f
C1267 via23_4_678/m2_1_40# VSUBS 0.548f
C1268 via23_4_117/m2_1_40# VSUBS 0.427f
C1269 via23_4_128/m2_1_40# VSUBS 0.427f
C1270 via23_4_677/m2_1_40# VSUBS 0.425f
C1271 via23_4_676/m2_1_40# VSUBS 0.425f
C1272 via23_4_21/m2_1_40# VSUBS 0.295f
C1273 via23_4_198/m2_1_40# VSUBS 0.427f
C1274 via23_4_103/m2_1_40# VSUBS 0.295f
C1275 via23_4_20/m2_1_40# VSUBS 0.295f
C1276 via23_4_91/m2_1_40# VSUBS 0.295f
C1277 via23_4_111/m2_1_40# VSUBS 0.427f
C1278 via23_4_199/m2_1_40# VSUBS 0.427f
C1279 via23_4_347/m2_1_40# VSUBS 0.425f
C1280 via23_4_379/m2_1_40# VSUBS 0.349f
C1281 via23_4_346/m2_1_40# VSUBS 0.548f
C1282 via23_4_1/m2_1_40# VSUBS 0.295f
C1283 via23_4_712/m2_1_40# VSUBS 0.425f
C1284 via23_4_378/m2_1_40# VSUBS 0.349f
C1285 via23_4_334/m2_1_40# VSUBS 0.425f
C1286 via23_4_345/m2_1_40# VSUBS 0.425f
C1287 via23_4_89/m2_1_40# VSUBS 0.418f
C1288 via23_4_23/m2_1_40# VSUBS 0.295f
C1289 via23_4_711/m2_1_40# VSUBS 0.425f
C1290 via23_4_333/m2_1_40# VSUBS 0.425f
C1291 n7 VSUBS 79.1f
C1292 via23_4_22/m2_1_40# VSUBS 0.295f
C1293 via23_4_710/m2_1_40# VSUBS 0.425f
C1294 via23_4_367/m2_1_40# VSUBS 0.575f
C1295 via23_4_332/m2_1_40# VSUBS 0.425f
C1296 via23_4_2/m2_1_40# VSUBS 0.283f
C1297 via23_4_87/m2_1_40# VSUBS 0.295f
C1298 via23_4_705/m2_1_40# VSUBS 0.427f
C1299 via23_4_366/m2_1_40# VSUBS 0.357f
C1300 via23_4_331/m2_1_40# VSUBS 0.425f
C1301 via23_4_354/m2_1_40# VSUBS 0.425f
C1302 n6 VSUBS 38.4f
C1303 via23_4_88/m2_1_40# VSUBS 0.295f
C1304 via23_4_589/m2_1_40# VSUBS 0.425f
C1305 via23_4_704/m2_1_40# VSUBS 0.427f
C1306 via23_4_369/m2_1_40# VSUBS 0.349f
C1307 via23_4_96/m2_1_40# VSUBS 0.445f
C1308 via23_4_588/m2_1_40# VSUBS 0.425f
C1309 via23_4_368/m2_1_40# VSUBS 0.349f
C1310 via23_4_95/m2_1_40# VSUBS 0.295f
C1311 via23_4_702/m2_1_40# VSUBS 0.575f
C1312 via23_4_200/m2_1_40# VSUBS 0.427f
C1313 via23_4_94/m2_1_40# VSUBS 0.295f
C1314 n2 VSUBS 8.12f
C1315 via23_4_675/m2_1_40# VSUBS 0.425f
C1316 via23_4_601/m2_1_40# VSUBS 0.425f
C1317 top VSUBS 33.9f
C1318 via23_4_381/m2_1_40# VSUBS 0.349f
C1319 via23_4_600/m2_1_40# VSUBS 0.425f
C1320 via23_4_380/m2_1_40# VSUBS 0.472f
C1321 via23_4_584/m2_1_40# VSUBS 0.425f
C1322 via23_4_599/m2_1_40# VSUBS 0.548f
C1323 via23_4_245/m2_1_40# VSUBS 0.425f
C1324 via23_4_598/m2_1_40# VSUBS 0.425f
C1325 via23_4_90/m2_1_40# VSUBS 0.295f
C1326 via23_4_218/m2_1_40# VSUBS 0.425f
C1327 via23_4_228/m2_1_40# VSUBS 0.575f
C1328 via23_4_230/m2_1_40# VSUBS 0.425f
C1329 ndum VSUBS 7.47f
C1330 via23_4_249/m2_1_40# VSUBS 0.425f
C1331 via23_4_229/m2_1_40# VSUBS 0.425f
C1332 via23_4_590/m2_1_40# VSUBS 0.425f
C1333 via23_4_419/m2_1_40# VSUBS 0.427f
C1334 via23_4_439/m2_1_40# VSUBS 0.339f
C1335 via23_4_213/m2_1_40# VSUBS 0.427f
C1336 via23_4_429/m2_1_40# VSUBS 0.427f
C1337 via23_4_449/m2_1_40# VSUBS 0.462f
C1338 via23_4_448/m2_1_40# VSUBS 0.339f
.ends

.subckt DAC ctl1 ctl0 dum ctl3 ctl4 ctl5 ctl6 ctl7 ctl2 carray_0/m3_13900_1156# carray_0/via23_4_220/m2_1_40#
+ carray_0/m3_24300_1156# carray_0/m3_6100_1156# carray_0/m2_40200_1156# carray_0/m3_29500_1156#
+ carray_0/via23_4_251/m2_1_40# carray_0/m3_20400_1156# carray_0/m3_2200_1156# carray_0/via23_4_711/m2_1_40#
+ carray_0/via23_4_675/m2_1_40# carray_0/m3_25600_1156# carray_0/m3_7400_1156# carray_0/m3_36000_1156#
+ carray_0/via23_4_345/m2_1_40# carray_0/m2_41500_1156# carray_0/via23_4_588/m2_1_40#
+ carray_0/m3_3500_1156# carray_0/m3_32100_1156# carray_0/m3_26900_1156# carray_0/m3_8700_1156#
+ carray_0/m2_42800_1156# carray_0/m3_37300_1156# carray_0/via23_4_218/m2_1_40# carray_0/m3_900_1156#
+ carray_0/via23_4_599/m2_1_40# carray_0/via23_4_677/m2_1_40# carray_0/via23_4_249/m2_1_40#
+ carray_0/m3_18000_1156# carray_0/m3_4800_1156# carray_0/m3_33400_1156# carray_0/m3_38600_1156#
+ carray_0/via23_4_333/m2_1_40# carray_0/m3_14100_1156# carray_0/m3_19300_1156# vin
+ carray_0/m3_34700_1156# carray_0/m3_39900_1156# carray_0/via23_4_199/m2_1_40# carray_0/m3_10200_1156#
+ carray_0/m3_15400_1156# carray_0/m3_30800_1156# carray_0/m3_41200_1156# enb carray_0/via23_4_712/m2_1_40#
+ carray_0/via23_4_200/m2_1_40# carray_0/via23_4_346/m2_1_40# carray_0/m3_11500_1156#
+ carray_0/m3_16700_1156# carray_0/m3_27100_1156# carray_0/via23_4_228/m2_1_40# carray_0/m3_42500_1156#
+ carray_0/via23_4_589/m2_1_40# carray_0/m3_12800_1156# carray_0/m3_5000_1156# carray_0/m3_23200_1156#
+ carray_0/via23_4_245/m2_1_40# carray_0/m3_28400_1156# carray_0/m2_19000_1156# carray_0/via23_4_600/m2_1_40#
+ carray_0/via23_4_678/m2_1_40# sample carray_0/m3_1100_1156# carray_0/m3_24500_1156#
+ carray_0/m3_6300_1156# carray_0/m3_29700_1156# carray_0/m2_15100_1156# carray_0/via23_4_334/m2_1_40#
+ carray_0/via23_4_229/m2_1_40# carray_0/via23_4_702/m2_1_40# carray_0/m3_2400_1156#
+ en_buf carray_0/m3_31000_1156# carray_0/m3_25800_1156# carray_0/m2_11200_1156# carray_0/m3_7600_1156#
+ carray_0/m3_36200_1156# carray_0/m2_16400_1156# carray_0/m2_27200_1156# carray_0/via23_4_584/m2_1_40#
+ carray_0/via23_4_331/m2_1_40# carray_0/m3_3700_1156# carray_0/m3_32300_1156# carray_0/m3_8900_1156#
+ carray_0/via23_4_213/m2_1_40# carray_0/m3_37500_1156# carray_0/m2_12500_1156# carray_0/m2_6000_1156#
+ carray_0/m2_17700_1156# carray_0/m2_800_1156# carray_0/via23_4_347/m2_1_40# carray_0/m2_23300_1156#
+ carray_0/n3 carray_0/via23_4_326/m2_1_40# carray_0/m2_28500_1156# carray_0/m3_33600_1156#
+ carray_0/via23_4_354/m2_1_40# carray_0/m2_13800_1156# carray_0/m2_2100_1156# carray_0/m3_38800_1156#
+ carray_0/m2_7300_1156# carray_0/via23_4_250/m2_1_40# carray_0/m2_24600_1156# carray_0/m3_19100_1156#
+ carray_0/m2_35000_1156# carray_0/m2_29800_1156# carray_0/via23_4_710/m2_1_40# carray_0/via23_4_601/m2_1_40#
+ carray_0/m3_40100_1156# carray_0/via23_4_709/m2_1_40# carray_0/m3_34900_1156# carray_0/m2_3400_1156#
+ carray_0/m2_20300_1156# carray_0/m2_8600_1156# carray_0/m3_10000_1156# vdd carray_0/n1
+ carray_0/m3_15200_1156# carray_0/via23_4_198/m2_1_40# carray_0/m2_31100_1156# carray_0/m2_25900_1156#
+ carray_0/m2_36300_1156# carray_0/m3_41400_1156# carray_0/m2_4700_1156# carray_0/m2_9900_1156#
+ carray_0/via23_4_230/m2_1_40# carray_0/m3_11300_1156# carray_0/n5 carray_0/via23_4_598/m2_1_40#
+ carray_0/m3_16500_1156# carray_0/via23_4_676/m2_1_40# carray_0/m2_32400_1156# carray_0/m2_37600_1156#
+ carray_0/m3_42700_1156# carray_0/n2 carray_0/n4 carray_0/m3_12600_1156# carray_0/m3_17800_1156#
+ carray_0/via23_4_332/m2_1_40# carray_0/n0 carray_0/m3_28200_1156# carray_0/m2_33700_1156#
+ carray_0/m2_38900_1156# carray_0/n6 carray_0/via23_4_590/m2_1_40# carray_0/ndum
+ vss out carray_0/n7
Xinv2_0 vdd vdd ctl7 carray_0/n7 vss vss inv2
Xinv2_1 vdd vdd ctl6 carray_0/n6 vss vss inv2
Xinv2_2 vdd vdd dum carray_0/ndum vss vss inv2
Xinv2_3 vdd vdd ctl0 carray_0/n0 vss vss inv2
Xinv2_4 vdd vdd ctl1 carray_0/n1 vss vss inv2
Xinv2_5 vdd vdd ctl5 carray_0/n5 vss vss inv2
Xinv2_6 vdd vdd ctl4 carray_0/n4 vss vss inv2
Xinv2_7 vdd vdd ctl2 carray_0/n2 vss vss inv2
Xinv2_8 vdd vdd ctl3 carray_0/n3 vss vss inv2
Xsw_top_0 sample sw_top_0/m2_1158_361# vdd out vdd vin sw_top_0/m2_990_200# vss sw_top
Xcarray_0 carray_0/n2 carray_0/n3 carray_0/via23_4_702/m2_1_40# carray_0/m3_12800_1156#
+ carray_0/m3_23200_1156# carray_0/m3_28400_1156# carray_0/m2_800_1156# carray_0/m2_19000_1156#
+ carray_0/via23_4_584/m2_1_40# carray_0/via23_4_331/m2_1_40# carray_0/m3_6100_1156#
+ carray_0/via23_4_213/m2_1_40# carray_0/m3_24500_1156# carray_0/m3_29700_1156# carray_0/m2_15100_1156#
+ carray_0/via23_4_347/m2_1_40# carray_0/via23_4_326/m2_1_40# carray_0/m3_2200_1156#
+ carray_0/via23_4_459/m2_1_40# carray_0/m3_7400_1156# carray_0/via23_4_354/m2_1_40#
+ carray_0/m3_25800_1156# carray_0/m3_31000_1156# carray_0/m2_11200_1156# carray_0/m3_36200_1156#
+ carray_0/m2_16400_1156# carray_0/via23_4_250/m2_1_40# carray_0/m2_27200_1156# carray_0/via23_4_710/m2_1_40#
+ carray_0/m3_3500_1156# carray_0/via23_4_601/m2_1_40# carray_0/m3_8700_1156# carray_0/via23_4_709/m2_1_40#
+ carray_0/m3_32300_1156# carray_0/m2_12500_1156# carray_0/m3_37500_1156# carray_0/m2_17700_1156#
+ carray_0/via23_4_198/m2_1_40# carray_0/m2_23300_1156# carray_0/m2_28500_1156# carray_0/m3_4800_1156#
+ carray_0/via23_4_230/m2_1_40# carray_0/m3_33600_1156# carray_0/m2_13800_1156# carray_0/m3_38800_1156#
+ carray_0/via23_4_447/m2_1_40# carray_0/via23_4_598/m2_1_40# carray_0/via23_4_676/m2_1_40#
+ carray_0/m3_19100_1156# carray_0/m2_24600_1156# carray_0/m2_29800_1156# carray_0/m2_35000_1156#
+ carray_0/m3_34900_1156# carray_0/m3_40100_1156# carray_0/m2_20300_1156# carray_0/m3_10000_1156#
+ carray_0/via23_4_332/m2_1_40# carray_0/m3_15200_1156# carray_0/m2_31100_1156# carray_0/m2_25900_1156#
+ carray_0/via23_4_369/m2_1_40# carray_0/m2_36300_1156# carray_0/via23_4_590/m2_1_40#
+ carray_0/m3_41400_1156# carray_0/via23_4_379/m2_1_40# carray_0/via23_4_220/m2_1_40#
+ carray_0/m3_11300_1156# carray_0/m3_16500_1156# carray_0/m2_32400_1156# carray_0/m2_37600_1156#
+ carray_0/via23_4_251/m2_1_40# carray_0/m3_42700_1156# carray_0/via23_4_711/m2_1_40#
+ carray_0/via23_4_675/m2_1_40# carray_0/m3_12600_1156# carray_0/via23_4_345/m2_1_40#
+ carray_0/m3_17800_1156# carray_0/m3_28200_1156# carray_0/m2_33700_1156# carray_0/m3_5000_1156#
+ carray_0/m2_38900_1156# carray_0/m3_900_1156# carray_0/via23_4_635/m2_1_40# carray_0/via23_4_455/m2_1_40#
+ carray_0/via23_4_588/m2_1_40# carray_0/m3_13900_1156# carray_0/via23_4_414/m2_1_40#
+ carray_0/m3_24300_1156# carray_0/via23_4_439/m2_1_40# carray_0/m2_40200_1156# carray_0/m3_1100_1156#
+ carray_0/m3_29500_1156# carray_0/via23_4_460/m2_1_40# carray_0/via23_4_218/m2_1_40#
+ carray_0/m3_6300_1156# carray_0/via23_4_704/m2_1_40# carray_0/via23_4_599/m2_1_40#
+ carray_0/via23_4_677/m2_1_40# carray_0/via23_4_249/m2_1_40# carray_0/m3_20400_1156#
+ carray_0/m3_2400_1156# carray_0/m3_25600_1156# carray_0/m3_36000_1156# carray_0/m2_41500_1156#
+ carray_0/m3_7600_1156# carray_0/via23_4_333/m2_1_40# carray_0/via23_4_366/m2_1_40#
+ carray_0/m3_26900_1156# carray_0/m3_32100_1156# carray_0/via23_4_429/m2_1_40# carray_0/m2_42800_1156#
+ carray_0/m3_3700_1156# carray_0/m3_37300_1156# carray_0/m3_8900_1156# carray_0/m2_6000_1156#
+ carray_0/via23_4_128/m2_1_40# carray_0/via23_4_458/m2_1_40# carray_0/via23_4_199/m2_1_40#
+ carray_0/ndum carray_0/via23_4_381/m2_1_40# carray_0/m3_18000_1156# carray_0/n0
+ carray_0/via23_4_419/m2_1_40# carray_0/m3_33400_1156# carray_0/m3_38600_1156# carray_0/m2_2100_1156#
+ carray_0/m2_7300_1156# carray_0/via23_4_449/m2_1_40# carray_0/via23_4_200/m2_1_40#
+ carray_0/via23_4_712/m2_1_40# carray_0/via23_4_346/m2_1_40# carray_0/m3_14100_1156#
+ carray_0/n4 carray_0/m3_19300_1156# carray_0/via23_4_228/m2_1_40# carray_0/via23_4_641/m2_1_40#
+ carray_0/via23_4_378/m2_1_40# carray_0/m3_34700_1156# carray_0/m3_39900_1156# carray_0/n1
+ carray_0/m2_3400_1156# carray_0/via23_4_589/m2_1_40# carray_0/n6 carray_0/m2_8600_1156#
+ carray_0/m3_10200_1156# carray_0/via23_4_642/m2_1_40# carray_0/via23_4_245/m2_1_40#
+ carray_0/m3_15400_1156# carray_0/via23_4_368/m2_1_40# carray_0/via23_4_705/m2_1_40#
+ carray_0/via23_4_446/m2_1_40# carray_0/m3_30800_1156# carray_0/via23_4_678/m2_1_40#
+ carray_0/via23_4_600/m2_1_40# carray_0/m3_41200_1156# carray_0/m2_4700_1156# carray_0/via23_4_96/m2_1_40#
+ carray_0/m2_9900_1156# carray_0/n5 carray_0/m3_11500_1156# carray_0/m3_16700_1156#
+ carray_0/via23_4_448/m2_1_40# carray_0/m3_27100_1156# carray_0/via23_4_334/m2_1_40#
+ carray_0/m3_42500_1156# vss carray_0/via23_4_380/m2_1_40# out carray_0/via23_4_229/m2_1_40#
+ carray_0/n7 carray_0/via23_4_367/m2_1_40# carray
Xsw_top_1 sample enb vdd out vdd vin en_buf vss sw_top
Xsw_top_2 sample enb vdd out vdd vin en_buf vss sw_top
Xsw_top_3 sample sw_top_3/m2_1158_361# vdd out vdd vin sw_top_3/m2_990_200# vss sw_top
C0 vdd carray_0/via23_4_414/m2_1_40# 0.00896f
C1 ctl5 carray_0/n4 0.0189f
C2 carray_0/n2 carray_0/via23_4_96/m2_1_40# 0.163f
C3 carray_0/n6 carray_0/n4 6.52e-20
C4 sample carray_0/m2_40200_1156# 6.55e-20
C5 sample carray_0/via23_4_378/m2_1_40# 9.23e-21
C6 ctl1 carray_0/n5 3.5e-20
C7 carray_0/via23_4_366/m2_1_40# sample 9.23e-21
C8 vdd carray_0/n4 0.156f
C9 ctl7 carray_0/n4 1.79e-20
C10 ctl6 carray_0/n4 1.79e-20
C11 carray_0/n6 ctl0 1.35e-19
C12 carray_0/ndum carray_0/n1 2.07e-19
C13 ctl0 carray_0/n0 0.0223f
C14 vdd sw_top_3/m2_1158_361# 0.0395f
C15 vdd ctl0 0.0239f
C16 vin enb 0.175f
C17 ctl5 carray_0/n5 0.022f
C18 sample carray_0/m2_41500_1156# 6.55e-20
C19 carray_0/n2 ctl3 0.0189f
C20 out carray_0/via23_4_635/m2_1_40# 0.152f
C21 carray_0/n6 carray_0/n5 1.24f
C22 carray_0/n2 carray_0/n6 4.38e-20
C23 sw_top_3/m2_990_200# sample 0.122f
C24 sample carray_0/n3 3.92e-19
C25 carray_0/n0 carray_0/n5 3.34e-19
C26 carray_0/n6 dum 6.34e-20
C27 vdd carray_0/n5 0.157f
C28 out vin 0.262f
C29 ctl7 carray_0/n5 3.5e-20
C30 ctl6 carray_0/n5 0.0191f
C31 sw_top_0/m2_1158_361# sample 0.024f
C32 carray_0/n2 vdd 0.165f
C33 carray_0/n7 ctl1 0.0197f
C34 dum carray_0/n0 0.0204f
C35 vin carray_0/via23_4_642/m2_1_40# 0.0377f
C36 vdd dum 0.0303f
C37 sample carray_0/m2_42800_1156# 3.33e-19
C38 sw_top_0/m2_1158_361# carray_0/m2_42800_1156# 0.00399f
C39 sw_top_0/m2_1158_361# carray_0/via23_4_414/m2_1_40# 0.012f
C40 sample carray_0/m2_23300_1156# 6.55e-20
C41 vin en_buf 0.0702f
C42 vdd carray_0/via23_4_367/m2_1_40# 0.0215f
C43 vdd carray_0/via23_4_702/m2_1_40# 0.0228f
C44 carray_0/n2 ctl2 0.0218f
C45 carray_0/via23_4_368/m2_1_40# sample 9.23e-21
C46 out enb 0.15f
C47 carray_0/via23_4_448/m2_1_40# sample 9.23e-21
C48 carray_0/n3 carray_0/n4 1.31f
C49 vdd carray_0/via23_4_704/m2_1_40# 0.0254f
C50 sample carray_0/n4 5.55e-19
C51 carray_0/via23_4_705/m2_1_40# sw_top_3/m2_1158_361# 0.0141f
C52 carray_0/n6 carray_0/n7 1.2f
C53 vdd carray_0/via23_4_641/m2_1_40# 0.0234f
C54 vdd carray_0/m3_42700_1156# 0.00985f
C55 sample carray_0/m2_24600_1156# 6.55e-20
C56 carray_0/via23_4_429/m2_1_40# vdd 0.0121f
C57 carray_0/n7 carray_0/n0 1.45e-19
C58 sample carray_0/via23_4_459/m2_1_40# 9.23e-21
C59 vdd carray_0/n7 0.158f
C60 sample sw_top_3/m2_1158_361# 0.024f
C61 ctl7 carray_0/n7 0.0223f
C62 vin carray_0/via23_4_419/m2_1_40# 0.0405f
C63 ctl0 sample 0.00394f
C64 ctl6 carray_0/n7 0.00154f
C65 out carray_0/via23_4_642/m2_1_40# 0.045f
C66 sample carray_0/via23_4_455/m2_1_40# 4.62e-21
C67 sw_top_3/m2_1158_361# carray_0/m2_42800_1156# 0.00317f
C68 out en_buf 0.0196f
C69 sw_top_0/m2_990_200# vin 1.53e-20
C70 carray_0/n3 carray_0/n5 5.3e-20
C71 ctl1 carray_0/n1 0.0223f
C72 sample carray_0/n5 0.0017f
C73 carray_0/n2 carray_0/n3 1.34f
C74 carray_0/via23_4_419/m2_1_40# enb 0.0282f
C75 dum sample 0.00866f
C76 sw_top_0/m2_990_200# enb 1e-20
C77 carray_0/via23_4_367/m2_1_40# sample 0.0408f
C78 sw_top_0/m2_1158_361# carray_0/via23_4_367/m2_1_40# 0.0055f
C79 out carray_0/via23_4_419/m2_1_40# 0.0571f
C80 vdd carray_0/via23_4_635/m2_1_40# 0.0119f
C81 carray_0/n6 carray_0/n1 1.07e-19
C82 carray_0/via23_4_380/m2_1_40# sample 9.23e-21
C83 carray_0/n4 carray_0/n5 1.27f
C84 sample carray_0/m2_28500_1156# 6.55e-20
C85 sw_top_0/m2_990_200# out 0.00562f
C86 carray_0/n0 carray_0/n1 1.14f
C87 carray_0/n2 carray_0/n4 4.38e-20
C88 vdd vin 0.655f
C89 vdd carray_0/n1 0.159f
C90 sample carray_0/m3_42700_1156# 0.0051f
C91 sw_top_0/m2_1158_361# carray_0/m3_42700_1156# 0.00284f
C92 ctl7 carray_0/n1 0.00154f
C93 carray_0/n7 carray_0/n3 5.65e-19
C94 ctl0 carray_0/n5 5.09e-20
C95 carray_0/via23_4_429/m2_1_40# sw_top_0/m2_1158_361# 0.0233f
C96 carray_0/via23_4_641/m2_1_40# carray_0/m2_42800_1156# 2.84e-32
C97 carray_0/m2_42800_1156# carray_0/m3_42700_1156# 5.68e-32
C98 carray_0/n7 sample 4.96f
C99 carray_0/ndum carray_0/n0 1.1f
C100 vdd carray_0/ndum 0.195f
C101 sw_top_0/m2_990_200# en_buf 0.00185f
C102 ctl0 dum 0.194f
C103 sample carray_0/m2_29800_1156# 6.55e-20
C104 carray_0/n6 carray_0/m2_800_1156# 2.66e-20
C105 vdd enb 0.0404f
C106 sample carray_0/via23_4_447/m2_1_40# 9.23e-21
C107 carray_0/n2 carray_0/n5 4.38e-20
C108 ctl3 ctl4 0.194f
C109 carray_0/n7 carray_0/n4 3.37e-19
C110 ctl5 ctl4 0.194f
C111 vdd out 0.25f
C112 sw_top_3/m2_1158_361# carray_0/m3_42700_1156# 0.00285f
C113 sample carray_0/m2_31100_1156# 6.55e-20
C114 carray_0/via23_4_381/m2_1_40# sample 9.23e-21
C115 vdd carray_0/via23_4_642/m2_1_40# 0.0195f
C116 carray_0/n7 ctl0 1.7e-19
C117 carray_0/via23_4_369/m2_1_40# sample 9.23e-21
C118 carray_0/via23_4_705/m2_1_40# vin 0.0359f
C119 vdd ctl4 0.0238f
C120 vdd en_buf 0.00727f
C121 sw_top_3/m2_990_200# vin 0.0501f
C122 carray_0/via23_4_635/m2_1_40# carray_0/m2_42800_1156# 2.84e-32
C123 carray_0/n3 carray_0/n1 8.82e-20
C124 carray_0/via23_4_449/m2_1_40# sample 9.23e-21
C125 vin sample 0.304f
C126 sample carray_0/n1 0.00248f
C127 sw_top_0/m2_1158_361# vin 0.116f
C128 carray_0/n7 carray_0/n5 3.54e-19
C129 sample carray_0/m2_32400_1156# 6.55e-20
C130 sample carray_0/via23_4_446/m2_1_40# 9.23e-21
C131 vin carray_0/m2_42800_1156# 0.00127f
C132 vin carray_0/via23_4_414/m2_1_40# 0.0351f
C133 carray_0/n2 carray_0/n7 7.53e-19
C134 carray_0/ndum sample 11.1f
C135 carray_0/n7 dum 2.69e-19
C136 sw_top_3/m2_990_200# enb 0.00762f
C137 sample carray_0/via23_4_439/m2_1_40# 9.23e-21
C138 sample carray_0/via23_4_458/m2_1_40# 9.23e-21
C139 vdd carray_0/via23_4_419/m2_1_40# 0.0238f
C140 sample enb 0.024f
C141 sw_top_0/m2_1158_361# enb 0.00667f
C142 carray_0/m2_800_1156# carray_0/n3 9.73e-19
C143 sw_top_3/m2_1158_361# carray_0/via23_4_635/m2_1_40# 0.0234f
C144 carray_0/n4 carray_0/n1 6.52e-20
C145 carray_0/n6 ctl1 1.35e-19
C146 carray_0/via23_4_705/m2_1_40# out 0.0454f
C147 enb carray_0/m2_42800_1156# 0.00753f
C148 sample carray_0/m2_33700_1156# 6.55e-20
C149 out sw_top_3/m2_990_200# 0.0098f
C150 sw_top_0/m2_990_200# vdd 0.00727f
C151 out carray_0/n3 0.00516f
C152 ctl1 carray_0/n0 0.00154f
C153 vdd ctl1 0.0238f
C154 carray_0/n2 carray_0/via23_4_128/m2_1_40# 0.0993f
C155 ctl7 ctl1 0.194f
C156 out sample 0.0065f
C157 sw_top_0/m2_1158_361# out 0.0777f
C158 vin sw_top_3/m2_1158_361# 0.143f
C159 ctl0 carray_0/n1 0.02f
C160 out carray_0/m2_42800_1156# 0.0555f
C161 ctl4 carray_0/n3 0.0189f
C162 carray_0/n6 ctl5 0.00154f
C163 sw_top_3/m2_990_200# en_buf 0.00369f
C164 out carray_0/via23_4_414/m2_1_40# 0.0451f
C165 sample carray_0/via23_4_379/m2_1_40# 9.23e-21
C166 carray_0/ndum ctl0 0.00154f
C167 vdd ctl3 0.0238f
C168 sample en_buf 0.125f
C169 sample carray_0/m2_35000_1156# 6.55e-20
C170 sw_top_0/m2_1158_361# en_buf 0.00761f
C171 carray_0/m2_800_1156# carray_0/n4 5.11e-19
C172 vdd ctl5 0.0238f
C173 carray_0/n5 carray_0/n1 8.23e-20
C174 ctl6 ctl5 0.194f
C175 sample carray_0/via23_4_460/m2_1_40# 9.23e-21
C176 carray_0/n6 carray_0/n0 1.07e-19
C177 enb sw_top_3/m2_1158_361# 0.0133f
C178 carray_0/n6 vdd 0.157f
C179 carray_0/n6 ctl7 0.0194f
C180 carray_0/n6 ctl6 0.0221f
C181 out carray_0/n4 0.00281f
C182 dum carray_0/n1 2.05e-19
C183 ctl3 ctl2 0.194f
C184 sample carray_0/m2_25900_1156# 6.55e-20
C185 vdd carray_0/n0 0.159f
C186 vdd ctl7 0.0238f
C187 vdd ctl6 0.0238f
C188 carray_0/via23_4_367/m2_1_40# vin 0.0171f
C189 carray_0/via23_4_702/m2_1_40# vin 0.0294f
C190 ctl6 ctl7 0.194f
C191 carray_0/via23_4_96/m2_1_40# carray_0/n3 8.98e-19
C192 out sw_top_3/m2_1158_361# 0.0862f
C193 carray_0/ndum dum 0.0223f
C194 ctl4 carray_0/n4 0.0219f
C195 sample carray_0/m2_36300_1156# 6.55e-20
C196 carray_0/via23_4_642/m2_1_40# sw_top_3/m2_1158_361# 0.00437f
C197 vin carray_0/via23_4_704/m2_1_40# 0.0403f
C198 vdd ctl2 0.028f
C199 carray_0/m2_800_1156# carray_0/n5 1.36e-19
C200 vin carray_0/via23_4_641/m2_1_40# 0.0326f
C201 en_buf sw_top_3/m2_1158_361# 0.00762f
C202 vin carray_0/m3_42700_1156# 9.43e-20
C203 carray_0/n2 carray_0/m2_800_1156# 0.00165f
C204 sw_top_0/m2_990_200# sample 0.122f
C205 sample carray_0/m2_27200_1156# 6.55e-20
C206 carray_0/via23_4_702/m2_1_40# enb 0.0266f
C207 out carray_0/n5 0.00162f
C208 ctl1 sample 0.00262f
C209 carray_0/via23_4_429/m2_1_40# vin 0.0184f
C210 carray_0/n7 carray_0/n1 1.17f
C211 sample carray_0/m3_42500_1156# 0.0051f
C212 carray_0/n2 out 0.0119f
C213 sample carray_0/m2_37600_1156# 6.55e-20
C214 carray_0/n2 carray_0/m3_900_1156# 0.0151f
C215 enb carray_0/via23_4_704/m2_1_40# 0.0258f
C216 carray_0/via23_4_96/m2_1_40# carray_0/n4 5.45e-19
C217 ctl3 carray_0/n3 0.0218f
C218 ctl4 carray_0/n5 0.00154f
C219 carray_0/n7 carray_0/ndum 3.26e-19
C220 out carray_0/via23_4_367/m2_1_40# 9.39e-19
C221 out carray_0/via23_4_702/m2_1_40# 0.0881f
C222 enb carray_0/via23_4_641/m2_1_40# 0.0268f
C223 enb carray_0/m3_42700_1156# 0.00374f
C224 carray_0/n6 carray_0/n3 5.3e-20
C225 out carray_0/via23_4_704/m2_1_40# 0.0571f
C226 carray_0/via23_4_705/m2_1_40# vdd 0.00979f
C227 ctl1 carray_0/n4 1.79e-20
C228 carray_0/n6 sample 0.0059f
C229 vdd sw_top_3/m2_990_200# 0.00727f
C230 sample carray_0/m2_38900_1156# 6.55e-20
C231 vdd carray_0/n3 0.154f
C232 out carray_0/via23_4_641/m2_1_40# 0.0792f
C233 out carray_0/m3_42700_1156# 0.0285f
C234 sample carray_0/n0 0.00863f
C235 vdd sample 0.362f
C236 vdd sw_top_0/m2_1158_361# 0.0386f
C237 ctl7 sample 0.00172f
C238 carray_0/via23_4_429/m2_1_40# out 0.138f
C239 ctl0 ctl1 0.194f
C240 carray_0/via23_4_96/m2_1_40# carray_0/n5 0.00116f
C241 vdd carray_0/m2_42800_1156# 0.0244f
C242 ctl3 carray_0/n4 0.00154f
C243 vin carray_0/via23_4_635/m2_1_40# 0.0176f
C244 ctl2 carray_0/n3 0.00154f
C245 ctl7 vss 0.448f
C246 ctl2 vss 0.609f
C247 sw_top_3/m2_990_200# vss 1.84f
C248 sw_top_3/m2_1158_361# vss 1.74f
C249 dum vss 0.59f
C250 en_buf vss 3.51f
C251 enb vss 3.27f
C252 ctl3 vss 0.448f
C253 carray_0/n1 vss 4.87f
C254 carray_0/n5 vss 20.6f
C255 carray_0/n4 vss 10.2f
C256 carray_0/n3 vss 7.44f
C257 carray_0/m3_42700_1156# vss 1.97f
C258 carray_0/m3_42500_1156# vss 1.18f
C259 carray_0/m3_41400_1156# vss 1.17f
C260 carray_0/m3_41200_1156# vss 1.17f
C261 carray_0/m3_40100_1156# vss 1.17f
C262 carray_0/m3_39900_1156# vss 1.17f
C263 carray_0/m3_38800_1156# vss 1.17f
C264 carray_0/m3_38600_1156# vss 1.17f
C265 carray_0/m3_37500_1156# vss 1.17f
C266 carray_0/m3_37300_1156# vss 1.17f
C267 carray_0/m3_36200_1156# vss 1.17f
C268 carray_0/m3_36000_1156# vss 1.17f
C269 carray_0/m3_34900_1156# vss 1.17f
C270 carray_0/m3_34700_1156# vss 1.17f
C271 carray_0/m3_33600_1156# vss 1.17f
C272 carray_0/m3_33400_1156# vss 1.17f
C273 carray_0/m3_32300_1156# vss 1.17f
C274 carray_0/m3_32100_1156# vss 1.16f
C275 carray_0/m3_31000_1156# vss 1.17f
C276 carray_0/m3_30800_1156# vss 1.16f
C277 carray_0/m3_29700_1156# vss 1.17f
C278 carray_0/m3_29500_1156# vss 1.16f
C279 carray_0/m3_28400_1156# vss 1.17f
C280 carray_0/m3_28200_1156# vss 1.16f
C281 carray_0/m3_27100_1156# vss 1.17f
C282 carray_0/m3_26900_1156# vss 1.16f
C283 carray_0/m3_25800_1156# vss 1.17f
C284 carray_0/m3_25600_1156# vss 1.16f
C285 carray_0/m3_24500_1156# vss 1.17f
C286 carray_0/m3_24300_1156# vss 1.16f
C287 carray_0/m3_23200_1156# vss 1.17f
C288 carray_0/m3_20400_1156# vss 1.16f
C289 carray_0/m3_19300_1156# vss 1.16f
C290 carray_0/m3_19100_1156# vss 1.16f
C291 carray_0/m3_18000_1156# vss 1.16f
C292 carray_0/m3_17800_1156# vss 1.16f
C293 carray_0/m3_16700_1156# vss 1.16f
C294 carray_0/m3_16500_1156# vss 1.16f
C295 carray_0/m3_15400_1156# vss 1.16f
C296 carray_0/m3_15200_1156# vss 1.16f
C297 carray_0/m3_14100_1156# vss 1.16f
C298 carray_0/m3_13900_1156# vss 1.16f
C299 carray_0/m3_12800_1156# vss 1.16f
C300 carray_0/m3_12600_1156# vss 1.16f
C301 carray_0/m3_11500_1156# vss 1.16f
C302 carray_0/m3_11300_1156# vss 1.16f
C303 carray_0/m3_10200_1156# vss 1.16f
C304 carray_0/m3_10000_1156# vss 1.16f
C305 carray_0/m3_8900_1156# vss 1.16f
C306 carray_0/m3_8700_1156# vss 1.16f
C307 carray_0/m3_7600_1156# vss 1.16f
C308 carray_0/m3_7400_1156# vss 1.16f
C309 carray_0/m3_6300_1156# vss 1.16f
C310 carray_0/m3_6100_1156# vss 1.16f
C311 carray_0/m3_5000_1156# vss 1.16f
C312 carray_0/m3_4800_1156# vss 1.16f
C313 carray_0/m3_3700_1156# vss 1.16f
C314 carray_0/m3_3500_1156# vss 1.16f
C315 carray_0/m3_2400_1156# vss 1.16f
C316 carray_0/m3_2200_1156# vss 1.16f
C317 carray_0/m3_1100_1156# vss 1.16f
C318 carray_0/m3_900_1156# vss 1.95f
C319 carray_0/m2_42800_1156# vss 2.41f
C320 carray_0/m2_41500_1156# vss 1.8f
C321 carray_0/m2_40200_1156# vss 1.8f
C322 carray_0/m2_38900_1156# vss 1.8f
C323 carray_0/m2_37600_1156# vss 1.8f
C324 carray_0/m2_36300_1156# vss 1.8f
C325 carray_0/m2_35000_1156# vss 1.8f
C326 carray_0/m2_33700_1156# vss 1.8f
C327 carray_0/m2_32400_1156# vss 1.8f
C328 carray_0/m2_31100_1156# vss 1.8f
C329 carray_0/m2_29800_1156# vss 1.8f
C330 carray_0/m2_28500_1156# vss 1.8f
C331 carray_0/m2_27200_1156# vss 1.8f
C332 carray_0/m2_25900_1156# vss 1.8f
C333 carray_0/m2_24600_1156# vss 1.8f
C334 carray_0/m2_23300_1156# vss 1.79f
C335 carray_0/m2_20300_1156# vss 1.79f
C336 carray_0/m2_19000_1156# vss 1.8f
C337 carray_0/m2_17700_1156# vss 1.8f
C338 carray_0/m2_16400_1156# vss 1.8f
C339 carray_0/m2_15100_1156# vss 1.8f
C340 carray_0/m2_13800_1156# vss 1.8f
C341 carray_0/m2_12500_1156# vss 1.8f
C342 carray_0/m2_11200_1156# vss 1.8f
C343 carray_0/m2_9900_1156# vss 1.8f
C344 carray_0/m2_8600_1156# vss 1.8f
C345 carray_0/m2_7300_1156# vss 1.8f
C346 carray_0/m2_6000_1156# vss 1.8f
C347 carray_0/m2_4700_1156# vss 1.8f
C348 carray_0/m2_3400_1156# vss 1.8f
C349 carray_0/m2_2100_1156# vss 1.8f
C350 carray_0/m2_800_1156# vss 2.41f
C351 carray_0/via23_4_326/m2_1_40# vss 0.548f
C352 carray_0/via23_4_414/m2_1_40# vss 0.427f
C353 carray_0/via23_4_447/m2_1_40# vss 0.339f
C354 carray_0/via23_4_458/m2_1_40# vss 0.339f
C355 carray_0/via23_4_446/m2_1_40# vss 0.339f
C356 carray_0/via23_4_460/m2_1_40# vss 0.339f
C357 carray_0/via23_4_220/m2_1_40# vss 0.427f
C358 carray_0/via23_4_9/m2_1_40# vss 0.418f
C359 carray_0/via23_4_459/m2_1_40# vss 0.327f
C360 carray_0/via23_4_641/m2_1_40# vss 0.427f
C361 carray_0/via23_4_251/m2_1_40# vss 0.425f
C362 carray_0/via23_4_455/m2_1_40# vss 0.283f
C363 carray_0/via23_4_635/m2_1_40# vss 0.427f
C364 carray_0/via23_4_250/m2_1_40# vss 0.425f
C365 carray_0/n0 vss 3.48f
C366 carray_0/via23_4_3/m2_1_40# vss 0.295f
C367 carray_0/via23_4_642/m2_1_40# vss 0.427f
C368 carray_0/via23_4_709/m2_1_40# vss 0.425f
C369 carray_0/via23_4_678/m2_1_40# vss 0.548f
C370 carray_0/via23_4_117/m2_1_40# vss 0.427f
C371 carray_0/via23_4_128/m2_1_40# vss 0.427f
C372 carray_0/via23_4_677/m2_1_40# vss 0.425f
C373 carray_0/via23_4_676/m2_1_40# vss 0.425f
C374 carray_0/via23_4_21/m2_1_40# vss 0.295f
C375 carray_0/via23_4_198/m2_1_40# vss 0.427f
C376 carray_0/via23_4_103/m2_1_40# vss 0.295f
C377 carray_0/via23_4_20/m2_1_40# vss 0.295f
C378 carray_0/via23_4_91/m2_1_40# vss 0.295f
C379 carray_0/via23_4_111/m2_1_40# vss 0.427f
C380 carray_0/via23_4_199/m2_1_40# vss 0.427f
C381 carray_0/via23_4_347/m2_1_40# vss 0.425f
C382 carray_0/via23_4_379/m2_1_40# vss 0.349f
C383 carray_0/via23_4_346/m2_1_40# vss 0.548f
C384 carray_0/via23_4_1/m2_1_40# vss 0.295f
C385 carray_0/via23_4_712/m2_1_40# vss 0.425f
C386 carray_0/via23_4_378/m2_1_40# vss 0.349f
C387 carray_0/via23_4_334/m2_1_40# vss 0.425f
C388 carray_0/via23_4_345/m2_1_40# vss 0.425f
C389 carray_0/via23_4_89/m2_1_40# vss 0.418f
C390 carray_0/via23_4_23/m2_1_40# vss 0.295f
C391 carray_0/via23_4_711/m2_1_40# vss 0.425f
C392 carray_0/via23_4_333/m2_1_40# vss 0.425f
C393 carray_0/n7 vss 78.7f
C394 carray_0/via23_4_22/m2_1_40# vss 0.295f
C395 carray_0/via23_4_710/m2_1_40# vss 0.425f
C396 carray_0/via23_4_367/m2_1_40# vss 0.575f
C397 carray_0/via23_4_332/m2_1_40# vss 0.425f
C398 carray_0/via23_4_2/m2_1_40# vss 0.283f
C399 carray_0/via23_4_87/m2_1_40# vss 0.295f
C400 carray_0/via23_4_705/m2_1_40# vss 0.427f
C401 carray_0/via23_4_366/m2_1_40# vss 0.357f
C402 carray_0/via23_4_331/m2_1_40# vss 0.425f
C403 carray_0/via23_4_354/m2_1_40# vss 0.425f
C404 carray_0/n6 vss 38.7f
C405 carray_0/via23_4_88/m2_1_40# vss 0.295f
C406 carray_0/via23_4_589/m2_1_40# vss 0.425f
C407 carray_0/via23_4_704/m2_1_40# vss 0.427f
C408 carray_0/via23_4_369/m2_1_40# vss 0.349f
C409 carray_0/via23_4_96/m2_1_40# vss 0.445f
C410 carray_0/via23_4_588/m2_1_40# vss 0.425f
C411 carray_0/via23_4_368/m2_1_40# vss 0.349f
C412 carray_0/via23_4_95/m2_1_40# vss 0.295f
C413 carray_0/via23_4_702/m2_1_40# vss 0.575f
C414 carray_0/via23_4_200/m2_1_40# vss 0.427f
C415 carray_0/via23_4_94/m2_1_40# vss 0.295f
C416 carray_0/n2 vss 8.96f
C417 carray_0/via23_4_675/m2_1_40# vss 0.425f
C418 carray_0/via23_4_601/m2_1_40# vss 0.425f
C419 out vss 37.7f
C420 carray_0/via23_4_381/m2_1_40# vss 0.349f
C421 carray_0/via23_4_600/m2_1_40# vss 0.425f
C422 carray_0/via23_4_380/m2_1_40# vss 0.472f
C423 carray_0/via23_4_584/m2_1_40# vss 0.425f
C424 carray_0/via23_4_599/m2_1_40# vss 0.548f
C425 carray_0/via23_4_245/m2_1_40# vss 0.425f
C426 carray_0/via23_4_598/m2_1_40# vss 0.425f
C427 carray_0/via23_4_90/m2_1_40# vss 0.295f
C428 carray_0/via23_4_218/m2_1_40# vss 0.425f
C429 carray_0/via23_4_228/m2_1_40# vss 0.575f
C430 carray_0/via23_4_230/m2_1_40# vss 0.425f
C431 carray_0/ndum vss 7.41f
C432 carray_0/via23_4_249/m2_1_40# vss 0.425f
C433 carray_0/via23_4_229/m2_1_40# vss 0.425f
C434 carray_0/via23_4_590/m2_1_40# vss 0.425f
C435 carray_0/via23_4_419/m2_1_40# vss 0.427f
C436 carray_0/via23_4_439/m2_1_40# vss 0.339f
C437 carray_0/via23_4_213/m2_1_40# vss 0.427f
C438 carray_0/via23_4_429/m2_1_40# vss 0.427f
C439 carray_0/via23_4_449/m2_1_40# vss 0.462f
C440 carray_0/via23_4_448/m2_1_40# vss 0.339f
C441 ctl4 vss 0.448f
C442 sample vss 27.6f
C443 sw_top_0/m2_990_200# vss 1.84f
C444 vin vss 6.69f
C445 sw_top_0/m2_1158_361# vss 1.74f
C446 ctl5 vss 0.448f
C447 vdd vss 35.1f
C448 ctl1 vss 0.448f
C449 ctl0 vss 0.448f
C450 ctl6 vss 0.448f
.ends

.subckt decap_3$1 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
C0 a_65_331# w_0_269# 0.0625f
C1 a_65_55# a_65_331# 0.353f
C2 a_65_55# w_0_269# 0.0797f
C3 a_65_331# VSUBS 0.47f
C4 a_65_55# VSUBS 0.427f
C5 w_0_269# VSUBS 0.339f
.ends

.subckt M1_1 a_30_n109# a_n88_n109# a_n33_n197# VSUBS
X0 a_30_n109# a_n33_n197# a_n88_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n109# a_n33_n197# 0.0116f
C1 a_n88_n109# a_30_n109# 0.121f
C2 a_n88_n109# a_n33_n197# 0.0116f
C3 a_30_n109# VSUBS 0.121f
C4 a_n88_n109# VSUBS 0.121f
C5 a_n33_n197# VSUBS 0.227f
.ends

.subckt trim_sw d_0 d_1 d_2 d_3 d_4 m1_1462_409# m1_1771_409# m1_799_409# m1_1226_409#
+ m1_136_409# vss
XM1_1_14 vss m1_799_409# d_2 vss M1_1
XM1_1_15 m1_799_409# vss d_2 vss M1_1
XM1_1_0 vss m1_1226_409# d_0 vss M1_1
XM1_1_1 vss m1_1771_409# d_4 vss M1_1
XM1_1_2 m1_1771_409# vss d_4 vss M1_1
XM1_1_3 vss m1_1771_409# d_4 vss M1_1
XM1_1_4 m1_1771_409# vss d_4 vss M1_1
XM1_1_5 m1_1771_409# vss d_4 vss M1_1
XM1_1_6 vss m1_1771_409# d_4 vss M1_1
XM1_1_7 vss m1_1771_409# d_4 vss M1_1
XM1_1_8 m1_1771_409# vss d_4 vss M1_1
XM1_1_9 m1_1462_409# vss d_1 vss M1_1
XM1_1_10 m1_136_409# vss d_3 vss M1_1
XM1_1_11 vss m1_136_409# d_3 vss M1_1
XM1_1_12 m1_136_409# vss d_3 vss M1_1
XM1_1_13 vss m1_136_409# d_3 vss M1_1
C0 m1_799_409# m1_1226_409# 0.153f
C1 d_4 m1_1462_409# 1.67e-19
C2 d_0 m1_1226_409# 0.0329f
C3 m1_799_409# d_2 0.0168f
C4 d_0 d_2 0.0765f
C5 m1_136_409# m1_799_409# 0.153f
C6 m1_1462_409# m1_1226_409# 0.0249f
C7 d_3 d_2 0.0446f
C8 d_4 m1_1771_409# 0.165f
C9 m1_799_409# vss 0.371f
C10 m1_1462_409# m1_1771_409# 0.0191f
C11 m1_136_409# d_3 0.069f
C12 d_0 vss 0.08f
C13 m1_1226_409# d_2 1.67e-19
C14 d_3 vss 0.272f
C15 d_0 d_1 0.113f
C16 d_4 vss 0.464f
C17 d_1 d_4 0.0454f
C18 m1_1462_409# vss 0.295f
C19 d_1 m1_1462_409# 0.0329f
C20 vss m1_1226_409# 0.168f
C21 m1_136_409# d_2 1.67e-19
C22 vss m1_1771_409# 1.08f
C23 vss d_2 0.153f
C24 m1_136_409# vss 0.789f
C25 d_0 m1_799_409# 1.67e-19
C26 d_3 m1_799_409# 1.67e-19
C27 d_1 vss 0.0843f
C28 d_2 0 0.368f
C29 m1_136_409# 0 0.38f
C30 vss 0 1.11f
C31 d_3 0 0.71f
C32 m1_1462_409# 0 0.0797f
C33 d_1 0 0.246f
C34 m1_1771_409# 0 0.401f
C35 d_4 0 1.3f
C36 m1_1226_409# 0 0.0757f
C37 d_0 0 0.233f
C38 m1_799_409# 0 0.219f
.ends

.subckt trim n1 n0 trim_sw_0/d_4 trim_sw_0/d_3 trim_sw_0/d_2 trim_sw_0/d_1 trim_sw_0/d_0
+ n4 n2 VSUBS drain n3
Xtrim_sw_0 trim_sw_0/d_0 trim_sw_0/d_1 trim_sw_0/d_2 trim_sw_0/d_3 trim_sw_0/d_4 n1
+ n4 n2 n0 n3 VSUBS trim_sw
C0 n2 n1 0.105f
C1 drain n1 0.851f
C2 trim_sw_0/d_4 n3 5.01e-19
C3 n4 n2 0.611f
C4 n4 drain 6.84f
C5 n2 n0 0.121f
C6 drain n0 0.851f
C7 n3 trim_sw_0/d_0 4.93e-20
C8 trim_sw_0/d_1 n3 4.93e-20
C9 VSUBS trim_sw_0/d_3 6.85e-20
C10 n4 n1 0.173f
C11 VSUBS n3 0.15f
C12 n1 n0 0.484f
C13 n2 trim_sw_0/d_4 0.00499f
C14 drain trim_sw_0/d_4 2.69e-20
C15 n4 n0 0.166f
C16 n2 trim_sw_0/d_0 0.00217f
C17 n2 trim_sw_0/d_1 0.00217f
C18 trim_sw_0/d_2 n3 9.86e-20
C19 n2 VSUBS 0.0689f
C20 VSUBS drain 1.76f
C21 n3 trim_sw_0/d_3 2.04e-19
C22 n1 trim_sw_0/d_1 0.00745f
C23 n4 trim_sw_0/d_4 5.97e-19
C24 VSUBS n1 0.0292f
C25 n4 trim_sw_0/d_0 2.85e-20
C26 n4 trim_sw_0/d_1 2.85e-20
C27 trim_sw_0/d_2 n2 6.21e-19
C28 trim_sw_0/d_2 drain 2.69e-20
C29 n0 trim_sw_0/d_0 0.00745f
C30 drain trim_sw_0/d_3 1.13e-19
C31 n4 VSUBS 0.204f
C32 n2 n3 0.579f
C33 drain n3 3.41f
C34 VSUBS n0 0.0289f
C35 n1 n3 0.105f
C36 VSUBS trim_sw_0/d_4 1.48e-19
C37 trim_sw_0/d_2 n4 1.64e-19
C38 n4 trim_sw_0/d_3 6.16e-20
C39 n2 drain 1.7f
C40 n4 n3 1.47f
C41 n0 n3 0.105f
C42 n1 0 0.264f
C43 n0 0 0.25f
C44 drain 0 -5.51f
C45 trim_sw_0/d_2 0 0.368f
C46 n3 0 1.47f
C47 VSUBS 0 1.91f
C48 trim_sw_0/d_3 0 0.71f
C49 trim_sw_0/d_1 0 0.246f
C50 n4 0 2.09f
C51 trim_sw_0/d_4 0 1.3f
C52 trim_sw_0/d_0 0 0.233f
C53 n2 0 0.8f
.ends

.subckt Mdiff a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_n88_n171# a_n33_51# 0.0116f
C2 a_n88_n171# a_30_n171# 0.121f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml1 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_n88_n171# a_n33_51# 0.0116f
C2 a_n88_n171# a_30_n171# 0.121f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt Minp a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_n88_n171# a_n33_51# 0.0116f
C2 a_n88_n171# a_30_n171# 0.121f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M1 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Minn a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_n88_n171# a_n33_51# 0.0116f
C2 a_n88_n171# a_30_n171# 0.121f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt Ml4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt M4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml2 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_n88_n171# a_n33_51# 0.0116f
C2 a_n88_n171# a_30_n171# 0.121f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M2 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n176# w_n124_n238# 0.00827f
C1 a_n33_55# w_n124_n238# 0.0663f
C2 a_30_n176# a_n88_n176# 0.121f
C3 a_30_n176# a_n33_55# 0.0116f
C4 a_30_n176# w_n124_n238# 0.00827f
C5 a_n33_55# a_n88_n176# 0.0116f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt comparator_core clk ip in diff outp w_302_2337# vdd vn vp vss outn
XMdiff_0 clk vss diff vss Mdiff
XMdiff_1 clk diff vss vss Mdiff
XM3_0 outp clk w_302_2337# vdd vss M3
XMl1_0 outp outn in vss Ml1
XMinp_0 vp ip diff vss Minp
XM1_0 in clk w_302_2337# vdd vss M1
XMinn_0 vn diff in vss Minn
XMl4_0 vdd outn w_302_2337# outp vss Ml4
XM4_0 vdd clk w_302_2337# ip vss M4
XMl2_0 outn ip outp vss Ml2
XM2_0 vdd clk w_302_2337# outn vss M2
XMl3_0 outn outp w_302_2337# vdd vss Ml3
C0 ip vdd 0.11f
C1 clk in 0.487f
C2 outp vdd 0.214f
C3 outn vdd 0.221f
C4 vp clk 0.105f
C5 diff vn 0.00126f
C6 ip outp 0.103f
C7 outn ip 0.0137f
C8 outn outp 1.11f
C9 in w_302_2337# 0.0589f
C10 clk vdd 0.277f
C11 vp w_302_2337# 0.0844f
C12 in vn 0.0809f
C13 in diff 0.0808f
C14 ip clk 0.487f
C15 vp vn 0.202f
C16 outp clk 0.256f
C17 vp diff 0.00126f
C18 outn clk 0.26f
C19 vdd w_302_2337# 1.19f
C20 vdd vn 0.0819f
C21 ip w_302_2337# 0.0584f
C22 outp w_302_2337# 0.305f
C23 outn w_302_2337# 0.318f
C24 ip diff 0.0808f
C25 outp vn 0.265f
C26 outp diff 0.00695f
C27 outn vn 0.212f
C28 outn diff 0.00246f
C29 in vdd 0.111f
C30 clk w_302_2337# 0.222f
C31 vp vdd 0.0812f
C32 clk vn 0.103f
C33 clk diff 0.0314f
C34 outp in 0.0137f
C35 outn in 0.103f
C36 ip vp 0.081f
C37 outp vp 0.281f
C38 outn vp 0.22f
C39 w_302_2337# vn 0.0855f
C40 clk vss 3.4f
C41 vdd vss 2.15f
C42 outn vss 1.9f
C43 w_302_2337# vss 4.58f
C44 vn vss 1.8f
C45 ip vss 1.2f
C46 vp vss 1.79f
C47 in vss 1.2f
C48 outp vss 1.89f
C49 diff vss 0.233f
.ends

.subckt comparator trim_3 trim_2 trim_0 trim_1 trim_4 trimb_4 trimb_1 trimb_0 trimb_2
+ clk comparator_core_0/w_302_2337# outp trim_1/n3 trimb_3 trim_1/drain vp outn trim_0/drain
+ trim_0/n3 vn vdd vss
Xtrim_0 trim_0/n1 trim_0/n0 trim_4 trim_3 trim_2 trim_1 trim_0 trim_0/n4 trim_0/n2
+ vss trim_0/drain trim_0/n3 trim
Xtrim_1 trim_1/n1 trim_1/n0 trimb_4 trimb_3 trimb_2 trimb_1 trimb_0 trim_1/n4 trim_1/n2
+ vss trim_1/drain trim_1/n3 trim
Xcomparator_core_0 clk trim_1/drain trim_0/drain comparator_core_0/diff outp comparator_core_0/w_302_2337#
+ vdd vn vp vss outn comparator_core
C0 trimb_4 vss 0.163f
C1 trim_3 trim_4 0.00204f
C2 outn vss 0.12f
C3 trim_2 vss 0.0538f
C4 clk outp 0.00196f
C5 trim_1/n2 vdd 0.00793f
C6 trim_0 trim_1 0.821f
C7 vdd trim_1 0.0651f
C8 trim_1/n4 trim_1/n3 0.354f
C9 trim_1/drain trim_1/n0 0.851f
C10 outn comparator_core_0/diff -1.11e-34
C11 trimb_0 trim_1/n1 3.22e-19
C12 trimb_2 trimb_1 5.25e-19
C13 outp trim_0/n4 3.21e-21
C14 trim_1/n2 trim_1/drain 1.7f
C15 vdd trimb_1 0.0651f
C16 trim_0/n1 trim_0/n4 0.0442f
C17 trim_0/n2 trim_2 7.46e-19
C18 vdd comparator_core_0/w_302_2337# 0.363f
C19 trim_1/n1 trim_1/n4 0.0442f
C20 vdd outp 0.104f
C21 trim_1/n2 vss 1.87e-20
C22 trim_0/n1 trim_0 3.22e-19
C23 trim_0/drain trim_0/n0 0.851f
C24 vp trim_1/n0 9.27e-20
C25 vn outn 8.17e-32
C26 vdd trim_1/n3 0.0276f
C27 vss trim_1 0.0907f
C28 vdd trim_0/n1 0.00185f
C29 clk trim_1/n4 2.05e-19
C30 trim_1/n2 vp 0.00276f
C31 trim_1/drain comparator_core_0/w_302_2337# 0.00517f
C32 trimb_0 trimb_2 0.969f
C33 trim_1/drain outp 0.0565f
C34 clk trim_0/n4 2.05e-19
C35 trim_1/n1 vdd 0.00185f
C36 vss trimb_1 0.0907f
C37 comparator_core_0/w_302_2337# vss 6.3e-19
C38 trimb_0 vdd 0.0787f
C39 trim_1/drain trim_1/n3 3.41f
C40 outp vss 0.12f
C41 trim_0/n2 trim_1 4.81e-20
C42 clk vdd 0.14f
C43 vss trim_1/n3 2.67e-20
C44 trim_0/n1 vss 4.36e-20
C45 vdd trim_1/n4 0.0315f
C46 trim_1/drain trim_1/n1 0.851f
C47 vp outp 5.68e-32
C48 outp comparator_core_0/diff -1.11e-34
C49 vp trim_1/n3 0.00558f
C50 vdd trim_0/n4 0.0315f
C51 trim_1/n1 vss 4.36e-20
C52 clk trim_1/drain 0.0585f
C53 trimb_0 vss 0.0594f
C54 vdd trimb_2 0.12f
C55 trim_1/drain trim_1/n4 6.86f
C56 trimb_4 trimb_3 0.00204f
C57 vdd trim_0 0.0787f
C58 trim_3 trim_2 1.07f
C59 clk vss 0.116f
C60 trim_1/n4 vss 0.0917f
C61 trim_4 trim_2 0.00289f
C62 outn trim_0/drain 0.0565f
C63 vp trim_1/n4 0.0127f
C64 vss trim_0/n4 0.0917f
C65 trim_1/drain vdd 0.0323f
C66 trimb_2 vss 0.0538f
C67 trim_0 vss 0.0594f
C68 trim_1/n2 trimb_3 6.27e-19
C69 vdd vss 5.16f
C70 trim_3 trim_1 3.55e-19
C71 clk vn 2.26e-19
C72 trim_4 trim_1 0.549f
C73 trim_0/n2 trim_0/n4 0.177f
C74 vp vdd 0.221f
C75 vdd comparator_core_0/diff 0.00201f
C76 trimb_1 trimb_3 3.55e-19
C77 trim_0/n2 trim_0 3.96e-20
C78 trim_1/drain vss 1.71f
C79 vn trim_0/n4 0.0127f
C80 trim_0/n2 vdd 0.00793f
C81 trim_1/n3 trimb_3 5.12e-19
C82 trim_1/drain vp 0.0543f
C83 trim_1/drain comparator_core_0/diff -2.84e-32
C84 comparator_core_0/w_302_2337# trim_0/drain 0.00529f
C85 vdd vn 0.221f
C86 trim_0/n3 trim_0/n4 0.354f
C87 outp trim_0/drain 4.92e-20
C88 vp vss 0.00394f
C89 trim_0/n1 trim_0/drain 0.851f
C90 trimb_0 trimb_3 3.55e-19
C91 vdd trim_0/n3 0.0276f
C92 trim_0/n2 vss 1.87e-20
C93 trim_0/n1 trim_0/n0 0.0442f
C94 vn vss 0.00394f
C95 clk trim_0/drain 0.0811f
C96 trimb_2 trimb_3 1.07f
C97 vss trim_0/n3 2.67e-20
C98 trim_4 trim_0/n4 0.00384f
C99 trim_3 trim_0 3.55e-19
C100 vdd trimb_3 0.438f
C101 trim_0/n2 vn 0.00276f
C102 trim_3 vdd 0.438f
C103 trim_0/drain trim_0/n4 6.86f
C104 trim_4 trim_0 0.0044f
C105 vdd trim_4 0.107f
C106 trim_2 trim_1 5.25e-19
C107 trim_0/n0 trim_0/n4 0.0442f
C108 vdd trim_0/drain 0.0315f
C109 trim_0 trim_0/n0 3.22e-19
C110 vn trim_0/n3 0.00558f
C111 vdd trim_0/n0 0.00149f
C112 trimb_4 trimb_1 0.549f
C113 vss trimb_3 0.0703f
C114 comparator_core_0/w_302_2337# outn -5.68e-32
C115 trim_3 vss 0.0703f
C116 outp outn 0.00414f
C117 trim_4 vss 0.163f
C118 trim_0/drain vss 1.71f
C119 trim_0/n2 trim_3 6.27e-19
C120 trim_0/drain comparator_core_0/diff -2.84e-32
C121 trimb_0 trimb_4 0.0044f
C122 trim_1/n2 trimb_1 4.81e-20
C123 trim_0/n2 trim_0/drain 1.7f
C124 clk outn 0.0885f
C125 trim_1/n4 trimb_4 0.00384f
C126 outn trim_1/n4 3.21e-21
C127 trim_1/n1 trim_1/n0 0.0442f
C128 trim_3 trim_0/n3 5.12e-19
C129 vn trim_0/drain 0.0543f
C130 trimb_0 trim_1/n0 3.22e-19
C131 trimb_2 trimb_4 0.00289f
C132 trim_1/n2 trimb_0 3.96e-20
C133 vn trim_0/n0 9.27e-20
C134 trim_1/n0 trim_1/n4 0.0442f
C135 trim_2 trim_0 0.969f
C136 trim_0/drain trim_0/n3 3.41f
C137 vdd trimb_4 0.107f
C138 vdd outn 0.105f
C139 vdd trim_2 0.12f
C140 trim_1/n2 trim_1/n4 0.177f
C141 trimb_0 trimb_1 0.821f
C142 trim_1/drain outn 4.92e-20
C143 vdd trim_1/n0 0.00149f
C144 trim_1/n2 trimb_2 7.46e-19
C145 trim_0/n4 trim_1 0.00239f
C146 trim_1/n4 trimb_1 0.00239f
C147 clk 0 3.23f
C148 vdd 0 7.35f
C149 outn 0 1.44f
C150 comparator_core_0/w_302_2337# 0 4.58f
C151 vn 0 1.65f
C152 vp 0 1.64f
C153 outp 0 1.45f
C154 comparator_core_0/diff 0 0.13f
C155 trim_1/n1 0 0.264f
C156 trim_1/n0 0 0.25f
C157 trim_1/drain 0 -4.5f
C158 trimb_2 0 0.582f
C159 trim_1/n3 0 1.47f
C160 trimb_3 0 1.6f
C161 trimb_1 0 0.399f
C162 trim_1/n4 0 2.09f
C163 trimb_4 0 1.44f
C164 trimb_0 0 0.397f
C165 trim_1/n2 0 0.8f
C166 trim_0/n1 0 0.264f
C167 trim_0/n0 0 0.25f
C168 trim_0/drain 0 -4.53f
C169 trim_2 0 0.582f
C170 trim_0/n3 0 1.47f
C171 vss 0 6.43f
C172 trim_3 0 1.6f
C173 trim_1 0 0.399f
C174 trim_0/n4 0 2.09f
C175 trim_4 0 1.44f
C176 trim_0 0 0.397f
C177 trim_0/n2 0 0.8f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.05
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.05
C0 VPWR VPB 0.0787f
C1 VPWR VGND 0.546f
C2 VGND VPB 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=2.89
C0 VPWR VPB 0.105f
C1 VPWR VGND 1.27f
C2 VGND VPB 0.22f
C3 VPWR VNB 1.14f
C4 VGND VNB 0.992f
C5 VPB VNB 0.782f
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPWR Y 0.209f
C1 VPB Y 0.0061f
C2 A Y 0.0894f
C3 VPWR VPB 0.0521f
C4 VPWR A 0.0631f
C5 VGND Y 0.155f
C6 VPWR VGND 0.0423f
C7 A VPB 0.0742f
C8 VGND VPB 0.00649f
C9 VGND A 0.0638f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND VPB VNB Q SET_B D CLK a_652_n19# a_1602_7#
+ a_562_373# a_1032_373# a_1296_7# a_796_7# a_586_7# a_1056_7# a_381_7# a_193_7# a_1140_373#
+ a_27_7# a_956_373# a_476_7# a_1224_7# a_1182_221#
X0 VPWR a_1032_373# a_1602_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1 a_1032_373# a_193_7# a_1056_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR SET_B a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_476_7# a_27_7# a_381_7# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X4 a_1296_7# a_1182_221# a_1224_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_1032_373# a_27_7# a_956_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X6 a_1182_221# a_1032_373# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X7 Q a_1602_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8 a_652_n19# a_476_7# a_796_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_1140_373# a_193_7# a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 a_586_7# a_193_7# a_476_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_381_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_1224_7# a_27_7# a_1032_373# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_1182_221# a_1032_373# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X16 VGND a_1032_373# a_1602_7# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X17 a_956_373# a_476_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 Q a_1602_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X19 a_796_7# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X20 VPWR a_476_7# a_652_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND SET_B a_1296_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X22 VGND a_652_n19# a_586_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X23 a_381_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X24 a_652_n19# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X25 a_562_373# a_27_7# a_476_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 VPWR a_1182_221# a_1140_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_476_7# a_193_7# a_381_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X29 a_1056_7# a_476_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X30 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 VPWR a_652_n19# a_562_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
C0 SET_B a_1224_7# 8.75e-19
C1 VGND a_1056_7# 0.00386f
C2 VGND a_1032_373# 0.157f
C3 a_956_373# VPWR 0.00457f
C4 a_27_7# D 0.103f
C5 a_1182_221# VGND 0.0628f
C6 VPWR a_562_373# 0.0041f
C7 SET_B Q 4.58e-19
C8 a_956_373# VGND 3.4e-19
C9 a_476_7# D 1.36e-19
C10 a_27_7# VPB 0.226f
C11 Q a_1602_7# 0.0715f
C12 a_27_7# VPWR 0.438f
C13 VPB a_652_n19# 0.0992f
C14 VPB a_476_7# 0.146f
C15 VPWR a_652_n19# 0.144f
C16 VPWR a_476_7# 0.12f
C17 a_193_7# a_1032_373# 0.0573f
C18 a_27_7# VGND 0.164f
C19 SET_B VPB 0.143f
C20 a_1182_221# a_193_7# 0.0728f
C21 SET_B VPWR 0.0807f
C22 a_586_7# VGND 0.00172f
C23 SET_B a_1296_7# 0.00167f
C24 VGND a_652_n19# 0.0761f
C25 VGND a_476_7# 0.178f
C26 a_1602_7# VPB 0.0453f
C27 VPWR a_1602_7# 0.135f
C28 SET_B VGND 0.338f
C29 a_193_7# a_562_373# 4.45e-20
C30 a_381_7# a_562_373# 8.75e-19
C31 a_1602_7# VGND 0.0942f
C32 CLK VPB 0.0702f
C33 CLK VPWR 0.0194f
C34 a_27_7# a_193_7# 0.797f
C35 a_27_7# a_381_7# 0.0729f
C36 a_796_7# VGND 0.00583f
C37 a_586_7# a_193_7# 0.00206f
C38 a_193_7# a_652_n19# 0.0849f
C39 a_381_7# a_586_7# 3.7e-19
C40 Q VPB 0.0174f
C41 CLK VGND 0.0194f
C42 a_193_7# a_476_7# 0.215f
C43 a_1224_7# VGND 0.00169f
C44 a_381_7# a_652_n19# 7.79e-20
C45 a_381_7# a_476_7# 0.0356f
C46 VPWR Q 0.0704f
C47 a_1140_373# a_1032_373# 0.00523f
C48 SET_B a_193_7# 0.202f
C49 a_1056_7# a_1032_373# 0.0016f
C50 VPB D 0.0485f
C51 VPWR D 0.0158f
C52 a_1182_221# a_1032_373# 0.344f
C53 Q VGND 0.0595f
C54 a_1602_7# a_193_7# 4.3e-19
C55 a_956_373# a_1032_373# 0.00212f
C56 VGND D 0.014f
C57 VPWR VPB 0.218f
C58 CLK a_193_7# 0.00156f
C59 VPB VGND 0.0173f
C60 a_27_7# a_1056_7# 0.00248f
C61 a_27_7# a_1032_373# 0.183f
C62 VPWR VGND 0.0687f
C63 a_1296_7# VGND 0.00523f
C64 a_27_7# a_1182_221# 0.0608f
C65 Q a_193_7# 6.4e-20
C66 a_652_n19# a_1056_7# 3.94e-19
C67 a_652_n19# a_1032_373# 0.00971f
C68 a_476_7# a_1032_373# 0.00329f
C69 a_956_373# a_27_7# 0.00294f
C70 a_193_7# D 0.0606f
C71 SET_B a_1140_373# 6.31e-19
C72 SET_B a_1056_7# 0.00152f
C73 SET_B a_1032_373# 0.215f
C74 a_381_7# D 0.14f
C75 a_1182_221# SET_B 0.12f
C76 a_27_7# a_562_373# 0.0018f
C77 a_956_373# a_652_n19# 3.11e-19
C78 a_1602_7# a_1032_373# 0.111f
C79 a_652_n19# a_562_373# 9.35e-20
C80 VPB a_193_7# 0.179f
C81 a_476_7# a_562_373# 0.00972f
C82 a_1182_221# a_1602_7# 0.144f
C83 a_381_7# VPB 0.0101f
C84 VPWR a_193_7# 0.101f
C85 VPWR a_381_7# 0.0942f
C86 a_27_7# a_652_n19# 0.19f
C87 a_1224_7# a_1032_373# 0.00536f
C88 a_27_7# a_476_7# 0.223f
C89 a_193_7# VGND 0.219f
C90 a_381_7# VGND 0.0787f
C91 a_27_7# SET_B 0.0407f
C92 a_586_7# a_476_7# 0.00807f
C93 a_476_7# a_652_n19# 0.26f
C94 Q a_1032_373# 0.00365f
C95 SET_B a_652_n19# 0.157f
C96 SET_B a_476_7# 0.203f
C97 a_27_7# a_1602_7# 2.39e-19
C98 SET_B a_1602_7# 0.00213f
C99 a_27_7# CLK 0.214f
C100 a_27_7# a_1224_7# 1.63e-19
C101 a_796_7# a_652_n19# 0.00196f
C102 VPB a_1032_373# 0.177f
C103 a_381_7# a_193_7# 0.157f
C104 a_796_7# a_476_7# 0.00184f
C105 VPWR a_1140_373# 0.00334f
C106 VPWR a_1032_373# 0.257f
C107 a_1182_221# VPB 0.112f
C108 a_1224_7# a_652_n19# 1.57e-19
C109 a_1296_7# a_1032_373# 0.00384f
C110 SET_B a_796_7# 0.00149f
C111 a_1182_221# VPWR 0.123f
C112 a_1182_221# a_1296_7# 1.84e-19
C113 a_27_7# Q 1.08e-19
C114 Q VNB 0.0834f
C115 VGND VNB 1.08f
C116 VPWR VNB 0.875f
C117 SET_B VNB 0.247f
C118 D VNB 0.107f
C119 CLK VNB 0.196f
C120 VPB VNB 1.93f
C121 a_381_7# VNB 0.0203f
C122 a_1602_7# VNB 0.126f
C123 a_1032_373# VNB 0.305f
C124 a_1182_221# VNB 0.128f
C125 a_476_7# VNB 0.286f
C126 a_652_n19# VNB 0.119f
C127 a_193_7# VNB 0.322f
C128 a_27_7# VNB 0.437f
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.97
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.97
C0 VPWR VPB 0.0858f
C1 VPB VGND 0.161f
C2 VPWR VGND 0.903f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2 a_584_7# a_346_7#
+ a_256_7# a_250_257# a_93_n19#
X0 a_346_7# A2 a_256_7# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1 a_250_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2 a_93_n19# A1 a_346_7# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X3 a_93_n19# B1 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4 VGND B2 a_584_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 VPWR a_93_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X6 VGND a_93_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X7 a_250_257# B2 a_93_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_256_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X9 a_250_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X10 a_584_7# B1 a_93_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X11 VPWR A2 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
C0 VPWR VPB 0.0756f
C1 A1 B1 0.0965f
C2 B1 a_256_7# 2.07e-20
C3 X B1 3.83e-20
C4 A3 B2 9.12e-20
C5 B2 A2 1.46e-19
C6 VGND B1 0.0344f
C7 a_584_7# B1 0.00143f
C8 A3 A2 0.0788f
C9 B2 a_93_n19# 0.0147f
C10 A3 a_93_n19# 0.124f
C11 a_93_n19# A2 0.0747f
C12 VPWR a_346_7# 0.00109f
C13 B1 a_250_257# 0.0125f
C14 B2 A1 3.14e-19
C15 B1 VPB 0.0276f
C16 A3 a_256_7# 4.42e-19
C17 A3 X 2.45e-19
C18 VGND B2 0.0469f
C19 A1 A2 0.0971f
C20 A2 a_256_7# 0.00256f
C21 X A2 1.19e-19
C22 A3 VGND 0.00974f
C23 B1 VPWR 0.01f
C24 A1 a_93_n19# 0.0641f
C25 a_93_n19# a_256_7# 0.0114f
C26 VGND A2 0.0114f
C27 X a_93_n19# 0.0841f
C28 VGND a_93_n19# 0.251f
C29 a_584_7# a_93_n19# 0.00278f
C30 B2 a_250_257# 0.0344f
C31 A3 a_250_257# 0.00602f
C32 B2 VPB 0.0355f
C33 X A1 6.03e-20
C34 B1 a_346_7# 5.39e-20
C35 A3 VPB 0.0291f
C36 a_250_257# A2 0.0129f
C37 VGND A1 0.0133f
C38 VGND a_256_7# 0.00394f
C39 VGND X 0.06f
C40 A2 VPB 0.0287f
C41 B2 VPWR 0.0108f
C42 a_93_n19# a_250_257# 0.188f
C43 A3 VPWR 0.0158f
C44 VGND a_584_7# 0.00683f
C45 a_93_n19# VPB 0.0485f
C46 VPWR A2 0.0133f
C47 A1 a_250_257# 0.0129f
C48 a_93_n19# VPWR 0.0907f
C49 X a_250_257# 5.42e-19
C50 A1 VPB 0.0296f
C51 X VPB 0.0108f
C52 VGND a_250_257# 0.0072f
C53 a_584_7# a_250_257# 2.43e-19
C54 VGND VPB 0.00788f
C55 A1 VPWR 0.016f
C56 VPWR a_256_7# 9.47e-19
C57 A2 a_346_7# 0.00252f
C58 X VPWR 0.0849f
C59 B2 B1 0.0823f
C60 a_93_n19# a_346_7# 0.0119f
C61 VGND VPWR 0.076f
C62 a_584_7# VPWR 9.47e-19
C63 A3 B1 7.88e-22
C64 B1 A2 1.44e-20
C65 a_250_257# VPB 0.00616f
C66 A1 a_346_7# 0.00465f
C67 a_93_n19# B1 0.0774f
C68 a_250_257# VPWR 0.313f
C69 VGND a_346_7# 0.00514f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_257# VNB 0.0278f
C80 a_93_n19# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X10 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X13 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X14 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X16 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X17 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X19 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X20 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X21 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X22 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X24 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X25 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X27 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 VPWR a_193_7# 0.396f
C1 VGND CLK 0.0172f
C2 VPWR D 0.0812f
C3 a_193_7# a_27_7# 0.906f
C4 VGND a_543_7# 0.123f
C5 a_651_373# RESET_B 0.0122f
C6 a_27_7# D 0.133f
C7 VPB Q 0.011f
C8 a_761_249# a_1270_373# 2.6e-19
C9 a_193_7# Q 1.81e-19
C10 VPWR a_1270_373# 7.19e-19
C11 VPB VGND 0.00999f
C12 VGND a_805_7# 0.00579f
C13 VGND a_193_7# 0.0631f
C14 RESET_B a_639_7# 9.54e-19
C15 VGND D 0.0516f
C16 a_651_373# a_761_249# 0.0977f
C17 a_651_373# VPWR 0.129f
C18 a_448_7# RESET_B 2.45e-19
C19 a_651_373# a_27_7# 9.73e-19
C20 VPB CLK 0.0693f
C21 VPB a_543_7# 0.0958f
C22 a_805_7# a_543_7# 0.00171f
C23 a_193_7# CLK 7.94e-19
C24 a_761_249# a_639_7# 3.16e-19
C25 a_193_7# a_543_7# 0.23f
C26 D a_543_7# 7.35e-20
C27 a_27_7# a_639_7# 0.00188f
C28 a_448_7# VPWR 0.0681f
C29 VPB a_193_7# 0.171f
C30 RESET_B a_1108_7# 0.237f
C31 a_1217_7# a_1108_7# 0.00742f
C32 a_448_7# a_27_7# 0.0931f
C33 RESET_B a_1217_7# 6.03e-19
C34 VPB D 0.138f
C35 a_193_7# D 0.218f
C36 VGND a_639_7# 0.00863f
C37 a_651_373# a_543_7# 0.0572f
C38 a_1283_n19# a_1108_7# 0.234f
C39 a_448_7# VGND 0.0661f
C40 RESET_B a_1283_n19# 0.278f
C41 a_761_249# a_1108_7# 0.0512f
C42 VPWR a_1108_7# 0.173f
C43 RESET_B a_761_249# 0.166f
C44 a_761_249# a_1217_7# 4.2e-19
C45 a_193_7# a_1270_373# 1.46e-19
C46 RESET_B VPWR 0.0652f
C47 a_27_7# a_1108_7# 0.102f
C48 RESET_B a_27_7# 0.296f
C49 a_651_373# VPB 0.0135f
C50 a_27_7# a_1217_7# 2.56e-19
C51 a_1462_7# RESET_B 0.00288f
C52 a_651_373# a_193_7# 0.0346f
C53 a_639_7# a_543_7# 0.0138f
C54 a_1108_7# Q 9.8e-19
C55 RESET_B Q 9.12e-19
C56 a_448_7# a_543_7# 0.0498f
C57 a_1283_n19# VPWR 0.209f
C58 VPWR a_761_249# 0.105f
C59 VGND a_1108_7# 0.148f
C60 a_1283_n19# a_27_7# 0.0436f
C61 RESET_B VGND 0.288f
C62 VGND a_1217_7# 9.68e-19
C63 a_761_249# a_27_7# 0.0701f
C64 VPWR a_27_7# 0.152f
C65 a_1462_7# a_1283_n19# 0.0074f
C66 a_193_7# a_639_7# 2.28e-19
C67 a_448_7# VPB 0.0141f
C68 a_1283_n19# Q 0.0598f
C69 a_448_7# a_193_7# 0.0642f
C70 VPWR Q 0.0997f
C71 a_448_7# D 0.156f
C72 a_1283_n19# VGND 0.24f
C73 a_27_7# Q 2.63e-20
C74 RESET_B CLK 1.09e-19
C75 VGND a_761_249# 0.0734f
C76 a_1108_7# a_543_7# 7.99e-20
C77 VGND VPWR 0.0502f
C78 RESET_B a_543_7# 0.153f
C79 VGND a_27_7# 0.254f
C80 a_1462_7# VGND 0.00221f
C81 VPB a_1108_7# 0.113f
C82 RESET_B VPB 0.138f
C83 RESET_B a_805_7# 0.00316f
C84 a_193_7# a_1108_7# 0.125f
C85 VGND Q 0.0616f
C86 RESET_B a_193_7# 0.0269f
C87 a_193_7# a_1217_7# 2.36e-20
C88 VPWR CLK 0.0174f
C89 a_761_249# a_543_7# 0.21f
C90 VPWR a_543_7# 0.1f
C91 RESET_B D 4.72e-19
C92 CLK a_27_7# 0.234f
C93 a_27_7# a_543_7# 0.115f
C94 a_1283_n19# VPB 0.137f
C95 VPB a_761_249# 0.0994f
C96 VPB VPWR 0.216f
C97 a_1270_373# a_1108_7# 0.00645f
C98 a_761_249# a_805_7# 3.69e-19
C99 RESET_B a_1270_373# 2.06e-19
C100 a_1283_n19# a_193_7# 0.0424f
C101 a_448_7# a_639_7# 4.61e-19
C102 VPB a_27_7# 0.262f
C103 a_761_249# a_193_7# 0.186f
C104 Q VNB 0.0899f
C105 VGND VNB 1.02f
C106 VPWR VNB 0.831f
C107 RESET_B VNB 0.264f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.85f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.139f
C114 a_1283_n19# VNB 0.299f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.274f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X a_27_7#
X0 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 X VPWR 0.139f
C1 A a_27_7# 0.209f
C2 A X 0.0123f
C3 a_27_7# X 0.165f
C4 VGND VPB 0.00461f
C5 VGND VPWR 0.0381f
C6 VGND A 0.0453f
C7 VPB VPWR 0.0438f
C8 A VPB 0.0335f
C9 VGND a_27_7# 0.105f
C10 VGND X 0.115f
C11 A VPWR 0.022f
C12 VPB a_27_7# 0.0686f
C13 VPB X 0.00837f
C14 a_27_7# VPWR 0.167f
C15 VGND VNB 0.263f
C16 X VNB 0.0731f
C17 VPWR VNB 0.221f
C18 A VNB 0.148f
C19 VPB VNB 0.428f
C20 a_27_7# VNB 0.32f
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B a_121_257# a_39_257#
X0 a_121_257# B a_39_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VGND a_39_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A a_39_257# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR a_39_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_39_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X6 VPWR A a_121_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_39_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 A VGND 0.0509f
C1 VGND a_121_257# 4.62e-19
C2 A B 0.0751f
C3 B VGND 0.0362f
C4 A VPWR 0.00734f
C5 VPWR VGND 0.0475f
C6 VPWR a_121_257# 0.00132f
C7 A VPB 0.0318f
C8 VPWR B 0.00593f
C9 VPB VGND 0.00955f
C10 VPB B 0.0416f
C11 A X 0.014f
C12 VGND X 0.0981f
C13 a_121_257# X 4.62e-19
C14 B X 1.51e-19
C15 A a_39_257# 0.176f
C16 VGND a_39_257# 0.14f
C17 a_39_257# a_121_257# 0.00477f
C18 B a_39_257# 0.0955f
C19 VPWR VPB 0.0714f
C20 VPWR X 0.165f
C21 VPB X 0.0108f
C22 VPWR a_39_257# 0.0899f
C23 VPB a_39_257# 0.0809f
C24 a_39_257# X 0.148f
C25 VGND VNB 0.323f
C26 X VNB 0.0724f
C27 A VNB 0.112f
C28 B VNB 0.178f
C29 VPWR VNB 0.284f
C30 VPB VNB 0.516f
C31 a_39_257# VNB 0.229f
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB X A B a_68_257# a_150_257#
X0 a_68_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_150_257# B a_68_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND A a_68_257# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_68_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR A a_150_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 X a_68_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
C0 A a_68_257# 0.158f
C1 B A 0.0751f
C2 VGND a_150_257# 4.62e-19
C3 VPWR a_68_257# 0.089f
C4 X a_68_257# 0.105f
C5 VPB VGND 0.0112f
C6 B VPWR 0.00855f
C7 X B 1.65e-19
C8 A VPWR 0.00846f
C9 X A 0.0131f
C10 a_150_257# a_68_257# 0.00477f
C11 VPB a_68_257# 0.0611f
C12 VGND a_68_257# 0.118f
C13 X VPWR 0.129f
C14 VPB B 0.0462f
C15 VGND B 0.0437f
C16 VPB A 0.031f
C17 VGND A 0.0347f
C18 a_150_257# VPWR 0.00193f
C19 X a_150_257# 4.96e-19
C20 VPB VPWR 0.0805f
C21 VGND VPWR 0.0464f
C22 X VPB 0.0209f
C23 B a_68_257# 0.0984f
C24 X VGND 0.114f
C25 VGND VNB 0.32f
C26 X VNB 0.101f
C27 A VNB 0.111f
C28 B VNB 0.183f
C29 VPWR VNB 0.269f
C30 VPB VNB 0.516f
C31 a_68_257# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y a_199_7# a_113_257#
X0 VGND A2 a_199_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1 a_113_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 a_199_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4 VPWR A1 a_113_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X5 a_113_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
C0 VPWR A1 0.0154f
C1 VGND VPB 0.00548f
C2 B1 Y 0.113f
C3 a_113_257# B1 0.00758f
C4 VGND Y 0.0654f
C5 VGND a_113_257# 0.00882f
C6 a_199_7# VPWR 4.76e-19
C7 a_199_7# A1 0.00917f
C8 VPB A2 0.0373f
C9 VPWR B1 0.0134f
C10 A1 B1 0.0518f
C11 A2 Y 0.00122f
C12 VGND VPWR 0.037f
C13 a_113_257# A2 0.0476f
C14 VGND A1 0.078f
C15 VPWR A2 0.0147f
C16 VGND a_199_7# 0.00428f
C17 A1 A2 0.0912f
C18 VGND B1 0.0436f
C19 VPB Y 0.0146f
C20 a_113_257# VPB 0.0108f
C21 a_113_257# Y 0.0909f
C22 VGND A2 0.0495f
C23 VPB VPWR 0.0424f
C24 VPB A1 0.0264f
C25 VPWR Y 0.0447f
C26 a_113_257# VPWR 0.177f
C27 A1 Y 0.0813f
C28 a_113_257# A1 0.05f
C29 VPB B1 0.0389f
C30 a_199_7# Y 0.00151f
C31 a_113_257# a_199_7# 2.42e-19
C32 VGND VNB 0.286f
C33 VPWR VNB 0.211f
C34 Y VNB 0.0544f
C35 A2 VNB 0.144f
C36 A1 VNB 0.0981f
C37 B1 VNB 0.162f
C38 VPB VNB 0.428f
C39 a_113_257# VNB 0.034f
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0 a_505_n19# a_535_334#
+ a_76_159# a_218_334# a_439_7# a_218_7#
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR a_505_n19# a_535_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_505_n19# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_76_159# A1 a_218_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_505_n19# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X5 a_439_7# A0 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6 a_218_334# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X7 a_76_159# A0 a_218_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X8 a_535_334# A1 a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X9 VGND a_505_n19# a_439_7# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_218_7# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
C0 a_218_334# VPWR 0.00177f
C1 a_218_334# VGND 7.29e-19
C2 VPWR a_535_334# 8.63e-19
C3 a_535_334# VGND 6.38e-19
C4 X a_218_7# 2.88e-19
C5 a_218_334# a_76_159# 0.00557f
C6 a_535_334# a_76_159# 6.64e-19
C7 X VPB 0.012f
C8 A1 VPB 0.0721f
C9 X VPWR 0.128f
C10 X VGND 0.0586f
C11 a_218_334# S 0.00688f
C12 VPWR A1 0.0114f
C13 A1 VGND 0.0752f
C14 S a_535_334# 0.00526f
C15 a_439_7# A1 0.00498f
C16 X a_76_159# 0.0776f
C17 A1 a_76_159# 0.187f
C18 VPWR a_218_7# 4.95e-19
C19 a_218_7# VGND 0.00328f
C20 a_218_7# a_76_159# 0.00783f
C21 A0 A1 0.267f
C22 VPWR VPB 0.11f
C23 VPB VGND 0.0134f
C24 X S 0.00823f
C25 S A1 0.0872f
C26 a_505_n19# A1 0.0993f
C27 VPB a_76_159# 0.0481f
C28 VPWR VGND 0.0804f
C29 VPWR a_439_7# 4.69e-19
C30 a_439_7# VGND 0.00354f
C31 VPWR a_76_159# 0.0542f
C32 VGND a_76_159# 0.16f
C33 A0 VPB 0.107f
C34 S VPB 0.168f
C35 a_505_n19# VPB 0.0781f
C36 VPWR A0 0.00732f
C37 A0 VGND 0.0432f
C38 a_439_7# A0 0.00369f
C39 S VPWR 0.392f
C40 VPWR a_505_n19# 0.0818f
C41 S VGND 0.033f
C42 A0 a_76_159# 0.0544f
C43 a_505_n19# VGND 0.124f
C44 S a_76_159# 0.318f
C45 S A0 0.0341f
C46 A0 a_505_n19# 0.0383f
C47 S a_505_n19# 0.198f
C48 VGND VNB 0.499f
C49 A1 VNB 0.14f
C50 A0 VNB 0.134f
C51 S VNB 0.268f
C52 VPWR VNB 0.419f
C53 X VNB 0.0924f
C54 VPB VNB 0.871f
C55 a_505_n19# VNB 0.247f
C56 a_76_159# VNB 0.139f
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=4.73
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=4.73
C0 VPB VPWR 0.142f
C1 VGND VPB 0.336f
C2 VGND VPWR 2.01f
C3 VPWR VNB 1.69f
C4 VGND VNB 1.45f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 A2 X a_448_7# a_544_257#
+ a_79_159# a_222_53#
X0 VGND A2 a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_79_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X2 a_222_53# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X3 a_448_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_544_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X5 a_448_7# a_222_53# a_79_159# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_222_53# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X7 a_79_159# a_222_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X8 a_544_257# A2 a_79_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X9 VGND a_79_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A1 a_79_159# 0.00575f
C1 A1 A2 0.0793f
C2 A1 VPB 0.0384f
C3 a_222_53# X 0.00374f
C4 a_222_53# a_79_159# 0.221f
C5 a_222_53# A2 0.0562f
C6 A1 VGND 0.017f
C7 a_222_53# VPB 0.0639f
C8 a_222_53# B1_N 0.106f
C9 A1 a_448_7# 0.0574f
C10 A1 VPWR 0.0508f
C11 a_79_159# X 0.11f
C12 a_222_53# VGND 0.0731f
C13 a_79_159# A2 0.0609f
C14 X VPB 0.0132f
C15 a_544_257# a_79_159# 0.00594f
C16 a_79_159# VPB 0.0676f
C17 a_222_53# a_448_7# 0.00596f
C18 a_544_257# A2 0.0012f
C19 X B1_N 0.00114f
C20 VPB A2 0.0259f
C21 a_222_53# VPWR 0.0224f
C22 a_79_159# B1_N 0.0833f
C23 B1_N VPB 0.0419f
C24 VGND X 0.0609f
C25 a_79_159# VGND 0.0836f
C26 VGND A2 0.0157f
C27 a_544_257# VGND 0.00166f
C28 a_448_7# a_79_159# 0.0461f
C29 VPWR X 0.0729f
C30 VGND VPB 0.0116f
C31 a_79_159# VPWR 0.263f
C32 a_448_7# A2 0.0581f
C33 VPWR A2 0.0227f
C34 VGND B1_N 0.0161f
C35 a_448_7# a_544_257# 0.00203f
C36 a_448_7# VPB 6.33e-19
C37 a_544_257# VPWR 0.0132f
C38 VPWR VPB 0.11f
C39 a_448_7# B1_N 2.55e-19
C40 VPWR B1_N 0.00448f
C41 a_448_7# VGND 0.168f
C42 VPWR VGND 0.0742f
C43 a_448_7# VPWR 0.00501f
C44 VGND VNB 0.468f
C45 B1_N VNB 0.105f
C46 VPWR VNB 0.4f
C47 X VNB 0.0865f
C48 A1 VNB 0.136f
C49 A2 VNB 0.0904f
C50 VPB VNB 0.782f
C51 a_448_7# VNB 0.0324f
C52 a_222_53# VNB 0.159f
C53 a_79_159# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR VPB VNB A X a_27_7#
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 VGND VPB 0.0142f
C1 X VPB 0.0164f
C2 a_27_7# VPB 0.266f
C3 VGND A 0.0543f
C4 A X 6.16e-19
C5 VPWR VPB 0.13f
C6 a_27_7# A 0.366f
C7 VPWR A 0.0492f
C8 VGND X 0.486f
C9 VGND a_27_7# 0.355f
C10 a_27_7# X 0.63f
C11 VGND VPWR 0.13f
C12 VPWR X 0.664f
C13 A VPB 0.0995f
C14 a_27_7# VPWR 0.465f
C15 VGND VNB 0.654f
C16 X VNB 0.0597f
C17 VPWR VNB 0.556f
C18 A VNB 0.322f
C19 VPB VNB 1.14f
C20 a_27_7# VNB 0.839f
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X9 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X11 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X16 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X17 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X20 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X22 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X23 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X26 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X28 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X29 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X30 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X33 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 a_639_7# a_27_7# 0.00188f
C1 VPB D 0.138f
C2 RESET_B a_639_7# 9.54e-19
C3 a_448_7# a_639_7# 4.61e-19
C4 a_543_7# a_639_7# 0.0138f
C5 VPB a_193_7# 0.171f
C6 a_651_373# a_761_249# 0.0977f
C7 a_761_249# VPWR 0.105f
C8 a_1108_7# VPWR 0.173f
C9 CLK a_193_7# 7.94e-19
C10 a_761_249# a_27_7# 0.0701f
C11 a_1108_7# a_27_7# 0.102f
C12 VPWR VGND 0.0779f
C13 Q a_1108_7# 0.0027f
C14 RESET_B a_761_249# 0.166f
C15 RESET_B a_1108_7# 0.237f
C16 a_543_7# a_761_249# 0.21f
C17 a_543_7# a_1108_7# 7.99e-20
C18 VGND a_27_7# 0.254f
C19 Q VGND 0.296f
C20 a_639_7# a_193_7# 2.28e-19
C21 a_1108_7# a_1283_n19# 0.234f
C22 RESET_B VGND 0.288f
C23 a_448_7# VGND 0.0661f
C24 a_543_7# VGND 0.123f
C25 a_1283_n19# VGND 0.299f
C26 VPB CLK 0.0693f
C27 a_1270_373# a_761_249# 2.6e-19
C28 RESET_B a_805_7# 0.00316f
C29 a_761_249# a_193_7# 0.186f
C30 a_1108_7# a_1270_373# 0.00645f
C31 a_1108_7# a_193_7# 0.125f
C32 D VGND 0.0516f
C33 a_543_7# a_805_7# 0.00171f
C34 a_761_249# a_1217_7# 4.2e-19
C35 a_1108_7# a_1217_7# 0.00742f
C36 VGND a_193_7# 0.0631f
C37 VGND a_1217_7# 9.68e-19
C38 VPB a_761_249# 0.0994f
C39 VPB a_1108_7# 0.115f
C40 VPB VGND 0.0123f
C41 a_651_373# VPWR 0.129f
C42 a_1462_7# VGND 0.00223f
C43 a_651_373# a_27_7# 9.73e-19
C44 a_651_373# RESET_B 0.0122f
C45 a_543_7# a_651_373# 0.0572f
C46 VGND CLK 0.0172f
C47 VPWR a_27_7# 0.152f
C48 Q VPWR 0.368f
C49 a_761_249# a_639_7# 3.16e-19
C50 RESET_B VPWR 0.0652f
C51 a_448_7# VPWR 0.0681f
C52 a_543_7# VPWR 0.1f
C53 Q a_27_7# 4.52e-20
C54 VGND a_639_7# 0.00863f
C55 a_1283_n19# VPWR 0.234f
C56 RESET_B a_27_7# 0.296f
C57 Q RESET_B 0.00188f
C58 a_448_7# a_27_7# 0.0931f
C59 a_543_7# a_27_7# 0.115f
C60 a_448_7# RESET_B 2.45e-19
C61 a_1283_n19# a_27_7# 0.0436f
C62 a_543_7# RESET_B 0.153f
C63 Q a_1283_n19# 0.367f
C64 a_448_7# a_543_7# 0.0498f
C65 RESET_B a_1283_n19# 0.28f
C66 a_651_373# a_193_7# 0.0346f
C67 a_1108_7# a_761_249# 0.0512f
C68 D VPWR 0.0812f
C69 a_1270_373# VPWR 7.19e-19
C70 VPWR a_193_7# 0.396f
C71 D a_27_7# 0.133f
C72 a_761_249# VGND 0.0734f
C73 a_1108_7# VGND 0.148f
C74 RESET_B D 4.72e-19
C75 a_448_7# D 0.156f
C76 a_27_7# a_193_7# 0.906f
C77 a_543_7# D 7.35e-20
C78 Q a_193_7# 2.64e-19
C79 RESET_B a_1270_373# 2.06e-19
C80 RESET_B a_193_7# 0.0269f
C81 a_27_7# a_1217_7# 2.56e-19
C82 a_448_7# a_193_7# 0.0642f
C83 a_543_7# a_193_7# 0.23f
C84 RESET_B a_1217_7# 6.03e-19
C85 a_1283_n19# a_193_7# 0.0427f
C86 VPB a_651_373# 0.0135f
C87 a_761_249# a_805_7# 3.69e-19
C88 VGND a_805_7# 0.00579f
C89 VPB VPWR 0.242f
C90 D a_193_7# 0.218f
C91 VPB a_27_7# 0.262f
C92 Q VPB 0.0176f
C93 a_1270_373# a_193_7# 1.46e-19
C94 VPB RESET_B 0.138f
C95 a_448_7# VPB 0.0141f
C96 a_543_7# VPB 0.0958f
C97 a_1217_7# a_193_7# 2.36e-20
C98 VPWR CLK 0.0174f
C99 VPB a_1283_n19# 0.228f
C100 a_1462_7# RESET_B 0.00288f
C101 a_27_7# CLK 0.234f
C102 a_1462_7# a_1283_n19# 0.0074f
C103 RESET_B CLK 1.09e-19
C104 Q VNB 0.0615f
C105 VGND VNB 1.18f
C106 VPWR VNB 0.977f
C107 RESET_B VNB 0.26f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 2.11f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.135f
C114 a_1283_n19# VNB 0.564f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.273f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A a_27_7#
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
C0 VGND a_27_7# 0.105f
C1 VPB A 0.0524f
C2 X VPB 0.0128f
C3 VPWR A 0.0215f
C4 X VPWR 0.0897f
C5 VGND A 0.0184f
C6 X VGND 0.0546f
C7 A a_27_7# 0.181f
C8 VPWR VPB 0.0355f
C9 X a_27_7# 0.107f
C10 VGND VPB 0.00505f
C11 VPWR VGND 0.029f
C12 X A 8.48e-19
C13 VPB a_27_7# 0.0592f
C14 VPWR a_27_7# 0.135f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_7# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 a_209_7# a_209_257#
+ a_303_7# a_80_n19#
X0 VPWR A2 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1 a_80_n19# B1 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2 a_209_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 VPWR a_80_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND B1 a_80_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_209_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X6 VGND a_80_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_209_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X8 a_303_7# A2 a_209_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X9 a_80_n19# A1 a_303_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
C0 VPWR B1 0.0177f
C1 X a_80_n19# 0.0765f
C2 a_209_257# a_303_7# 1.26e-19
C3 VPB a_80_n19# 0.051f
C4 a_209_257# a_209_7# 6.96e-20
C5 A3 a_209_7# 3.56e-19
C6 X VPWR 0.117f
C7 a_209_257# A2 0.0366f
C8 A3 A2 0.109f
C9 VPB VPWR 0.0715f
C10 B1 VGND 0.0172f
C11 A1 A2 0.104f
C12 a_209_257# a_80_n19# 0.0626f
C13 A3 a_80_n19# 0.117f
C14 X VGND 0.0572f
C15 VPB VGND 0.00769f
C16 A1 a_80_n19# 0.0367f
C17 a_209_257# VPWR 0.205f
C18 A3 VPWR 0.0403f
C19 a_303_7# A2 3.38e-19
C20 A1 VPWR 0.018f
C21 VPB B1 0.0342f
C22 a_209_257# VGND 0.0043f
C23 A3 VGND 0.0169f
C24 a_303_7# a_80_n19# 0.0115f
C25 A1 VGND 0.0135f
C26 X VPB 0.0108f
C27 a_209_7# a_80_n19# 0.0101f
C28 a_303_7# VPWR 0.00105f
C29 A2 a_80_n19# 0.0357f
C30 a_209_7# VPWR 0.00102f
C31 a_209_257# B1 0.00622f
C32 A2 VPWR 0.0227f
C33 A1 B1 0.101f
C34 a_303_7# VGND 0.00661f
C35 A3 X 0.00625f
C36 a_209_257# VPB 0.00284f
C37 A3 VPB 0.0297f
C38 VPWR a_80_n19# 0.0992f
C39 a_209_7# VGND 0.00696f
C40 A2 VGND 0.0148f
C41 A1 X 1.56e-19
C42 A1 VPB 0.0287f
C43 VGND a_80_n19# 0.216f
C44 A3 a_209_257# 0.0268f
C45 X a_303_7# 6.01e-19
C46 VPWR VGND 0.0662f
C47 A1 a_209_257# 0.0378f
C48 X a_209_7# 9.76e-19
C49 X A2 3.42e-19
C50 B1 a_80_n19# 0.111f
C51 VPB A2 0.0285f
C52 VGND VNB 0.41f
C53 VPWR VNB 0.332f
C54 X VNB 0.0895f
C55 B1 VNB 0.115f
C56 A1 VNB 0.0897f
C57 A2 VNB 0.0896f
C58 A3 VNB 0.0899f
C59 VPB VNB 0.693f
C60 a_209_257# VNB 0.00621f
C61 a_80_n19# VNB 0.211f
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X14 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X15 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X17 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X18 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X20 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X21 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X24 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X26 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X27 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X29 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 VGND VPWR 0.0719f
C1 a_448_7# a_543_7# 0.0498f
C2 VGND Q 0.11f
C3 a_543_7# VPB 0.0958f
C4 VPWR a_27_7# 0.152f
C5 a_27_7# Q 2.57e-20
C6 CLK VPWR 0.0174f
C7 a_193_7# VGND 0.0631f
C8 VGND RESET_B 0.288f
C9 a_761_249# a_1108_7# 0.0512f
C10 a_651_373# a_27_7# 9.73e-19
C11 a_448_7# VPWR 0.0681f
C12 VGND a_639_7# 0.00863f
C13 VPB VPWR 0.234f
C14 a_193_7# a_27_7# 0.906f
C15 VPB Q 0.00555f
C16 a_27_7# RESET_B 0.296f
C17 a_193_7# CLK 7.94e-19
C18 CLK RESET_B 1.09e-19
C19 a_639_7# a_27_7# 0.00188f
C20 a_543_7# a_1108_7# 7.99e-20
C21 VPWR a_1283_n19# 0.23f
C22 a_1283_n19# Q 0.0963f
C23 a_1108_7# a_1217_7# 0.00742f
C24 a_651_373# VPB 0.0135f
C25 a_193_7# a_448_7# 0.0642f
C26 a_448_7# RESET_B 2.45e-19
C27 a_193_7# VPB 0.171f
C28 VPB RESET_B 0.138f
C29 a_543_7# D 7.35e-20
C30 a_448_7# a_639_7# 4.61e-19
C31 a_193_7# a_1283_n19# 0.0425f
C32 a_805_7# a_761_249# 3.69e-19
C33 a_1283_n19# RESET_B 0.279f
C34 VGND a_27_7# 0.254f
C35 VPWR a_1108_7# 0.174f
C36 a_1108_7# Q 9.64e-19
C37 CLK VGND 0.0172f
C38 a_543_7# a_761_249# 0.21f
C39 a_761_249# a_1217_7# 4.2e-19
C40 a_1270_373# a_1108_7# 0.00645f
C41 a_543_7# a_805_7# 0.00171f
C42 CLK a_27_7# 0.234f
C43 VPWR D 0.0812f
C44 a_448_7# VGND 0.0661f
C45 VPB VGND 0.0122f
C46 a_193_7# a_1108_7# 0.125f
C47 a_1108_7# RESET_B 0.237f
C48 a_448_7# a_27_7# 0.0931f
C49 VPB a_27_7# 0.262f
C50 VPWR a_761_249# 0.105f
C51 VGND a_1283_n19# 0.259f
C52 CLK VPB 0.0693f
C53 a_193_7# D 0.218f
C54 D RESET_B 4.72e-19
C55 a_1270_373# a_761_249# 2.6e-19
C56 a_1462_7# RESET_B 0.00288f
C57 a_27_7# a_1283_n19# 0.0436f
C58 a_651_373# a_761_249# 0.0977f
C59 a_448_7# VPB 0.0141f
C60 a_543_7# VPWR 0.1f
C61 a_193_7# a_761_249# 0.186f
C62 a_761_249# RESET_B 0.166f
C63 VGND a_1108_7# 0.148f
C64 a_805_7# RESET_B 0.00316f
C65 a_639_7# a_761_249# 3.16e-19
C66 VPB a_1283_n19# 0.168f
C67 a_651_373# a_543_7# 0.0572f
C68 a_27_7# a_1108_7# 0.102f
C69 a_193_7# a_543_7# 0.23f
C70 a_193_7# a_1217_7# 2.36e-20
C71 a_543_7# RESET_B 0.153f
C72 RESET_B a_1217_7# 6.03e-19
C73 VGND D 0.0516f
C74 VPWR Q 0.169f
C75 a_1462_7# VGND 0.00221f
C76 a_543_7# a_639_7# 0.0138f
C77 D a_27_7# 0.133f
C78 a_1270_373# VPWR 7.19e-19
C79 VPB a_1108_7# 0.115f
C80 VGND a_761_249# 0.0734f
C81 a_651_373# VPWR 0.129f
C82 a_193_7# VPWR 0.396f
C83 a_193_7# Q 1.79e-19
C84 VGND a_805_7# 0.00579f
C85 VPWR RESET_B 0.0652f
C86 RESET_B Q 8.96e-19
C87 a_27_7# a_761_249# 0.0701f
C88 a_448_7# D 0.156f
C89 a_1283_n19# a_1108_7# 0.234f
C90 VPB D 0.138f
C91 a_193_7# a_1270_373# 1.46e-19
C92 a_1270_373# RESET_B 2.06e-19
C93 a_543_7# VGND 0.123f
C94 VGND a_1217_7# 9.68e-19
C95 a_193_7# a_651_373# 0.0346f
C96 a_651_373# RESET_B 0.0122f
C97 a_543_7# a_27_7# 0.115f
C98 a_193_7# RESET_B 0.0269f
C99 a_27_7# a_1217_7# 2.56e-19
C100 VPB a_761_249# 0.0994f
C101 a_1462_7# a_1283_n19# 0.0074f
C102 a_193_7# a_639_7# 2.28e-19
C103 a_639_7# RESET_B 9.54e-19
C104 Q VNB 0.0296f
C105 VGND VNB 1.1f
C106 VPWR VNB 0.902f
C107 RESET_B VNB 0.263f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.93f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.137f
C114 a_1283_n19# VNB 0.389f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.273f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X a_184_257# a_112_257# a_30_13#
X0 VPWR A a_184_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_184_257# B a_112_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_30_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X3 VPWR a_30_13# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND a_30_13# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_30_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X6 a_112_257# C a_30_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_30_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR VPB 0.0818f
C1 VPWR X 0.176f
C2 a_30_13# A 0.244f
C3 a_30_13# VPB 0.0791f
C4 a_30_13# X 0.137f
C5 B VGND 0.0151f
C6 VPWR a_184_257# 7.72e-19
C7 VPWR C 0.00459f
C8 a_30_13# a_184_257# 0.00863f
C9 B A 0.0788f
C10 B VPB 0.0972f
C11 B X 6.52e-19
C12 a_30_13# C 0.0862f
C13 a_112_257# VGND 3.96e-19
C14 a_30_13# VPWR 0.101f
C15 B C 0.0802f
C16 A a_112_257# 0.00223f
C17 B VPWR 0.148f
C18 a_30_13# B 0.121f
C19 A VGND 0.0192f
C20 VPB VGND 0.00844f
C21 X VGND 0.0786f
C22 A VPB 0.0382f
C23 a_112_257# VPWR 5.94e-19
C24 a_184_257# VGND 5.47e-19
C25 A X 0.00129f
C26 X VPB 0.00385f
C27 a_30_13# a_112_257# 0.00501f
C28 C VGND 0.0163f
C29 A a_184_257# 0.00228f
C30 A C 0.0343f
C31 VPWR VGND 0.0712f
C32 C VPB 0.0399f
C33 a_30_13# VGND 0.236f
C34 A VPWR 0.00982f
C35 VGND VNB 0.38f
C36 X VNB 0.0245f
C37 A VNB 0.117f
C38 C VNB 0.161f
C39 B VNB 0.116f
C40 VPWR VNB 0.33f
C41 VPB VNB 0.605f
C42 a_30_13# VNB 0.267f
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB A1 A2 B1 X a_382_257# a_79_n19#
+ a_297_7#
X0 a_297_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X2 a_382_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3 VPWR A1 a_382_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4 a_297_7# B1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_297_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
C0 a_382_257# VGND 8.23e-19
C1 VGND a_297_7# 0.125f
C2 VPWR a_79_n19# 0.201f
C3 B1 a_297_7# 0.00637f
C4 VPWR A2 0.0835f
C5 a_79_n19# A2 0.0889f
C6 A1 VPB 0.0412f
C7 VPWR VGND 0.0588f
C8 VPWR B1 0.0213f
C9 VGND a_79_n19# 0.129f
C10 a_382_257# A1 2.25e-19
C11 a_79_n19# B1 0.134f
C12 VGND A2 0.0171f
C13 B1 A2 0.0665f
C14 A1 a_297_7# 0.0492f
C15 VGND B1 0.0182f
C16 VPB X 0.011f
C17 VPWR A1 0.0449f
C18 A1 a_79_n19# 7.71e-19
C19 A1 A2 0.102f
C20 A1 VGND 0.0157f
C21 VPWR X 0.0958f
C22 a_79_n19# X 0.104f
C23 VPB a_297_7# 7.6e-19
C24 a_382_257# a_297_7# 8.13e-19
C25 VGND X 0.0736f
C26 B1 X 3.56e-19
C27 VPWR VPB 0.0624f
C28 VPB a_79_n19# 0.0489f
C29 VPB A2 0.0334f
C30 VPWR a_382_257# 0.00566f
C31 a_382_257# a_79_n19# 0.00145f
C32 a_382_257# A2 0.0145f
C33 VPWR a_297_7# 0.0056f
C34 VPB VGND 0.0049f
C35 VPB B1 0.0328f
C36 a_79_n19# a_297_7# 0.0326f
C37 a_297_7# A2 0.048f
C38 VGND VNB 0.352f
C39 VPWR VNB 0.304f
C40 X VNB 0.0935f
C41 A1 VNB 0.152f
C42 A2 VNB 0.0981f
C43 B1 VNB 0.101f
C44 VPB VNB 0.605f
C45 a_297_7# VNB 0.0348f
C46 a_79_n19# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=0.59
C0 VPB VGND 0.0797f
C1 VPWR VPB 0.0625f
C2 VPWR VGND 0.353f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB A B Y a_109_257#
X0 a_109_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 B VGND 0.0451f
C1 A VPB 0.0415f
C2 a_109_257# VGND 0.00128f
C3 VGND Y 0.154f
C4 B A 0.0584f
C5 VGND VPWR 0.0314f
C6 A Y 0.0471f
C7 A VPWR 0.0528f
C8 B VPB 0.0367f
C9 Y VPB 0.0139f
C10 A VGND 0.0486f
C11 VPB VPWR 0.0449f
C12 B Y 0.0877f
C13 a_109_257# Y 0.0113f
C14 B VPWR 0.0148f
C15 a_109_257# VPWR 0.00638f
C16 VGND VPB 0.00456f
C17 Y VPWR 0.0995f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_1 VGND VPWR VPB VNB Y A2_N A1_N B2 B1 a_109_257#
+ a_397_257# a_109_7# a_481_7#
X0 a_109_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A2_N a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.283 pd=1.52 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_109_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.283 ps=1.52 w=0.65 l=0.15
X3 a_109_7# A2_N a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 a_397_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_481_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B1 a_481_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B2 a_397_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_257# a_109_7# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.34 ps=2.68 w=1 l=0.15
X9 a_109_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y a_109_7# 0.192f
C1 B1 VPWR 0.018f
C2 B1 a_397_257# 0.0427f
C3 VPWR B2 0.0184f
C4 a_397_257# B2 0.0458f
C5 a_109_7# B2 0.0577f
C6 a_481_7# VPWR 6.39e-19
C7 a_481_7# a_397_257# 4.76e-19
C8 A2_N VPB 0.0308f
C9 VPWR VPB 0.0778f
C10 a_397_257# VPB 0.00776f
C11 A1_N VGND 0.0492f
C12 A2_N a_109_257# 5.93e-19
C13 a_109_7# VPB 0.0663f
C14 VPWR a_109_257# 0.00889f
C15 a_109_7# a_109_257# 0.00765f
C16 Y VGND 0.0978f
C17 A2_N VPWR 0.0192f
C18 VPWR a_397_257# 0.174f
C19 B1 VGND 0.0479f
C20 VGND B2 0.0678f
C21 A2_N a_109_7# 0.147f
C22 VPWR a_109_7# 0.0963f
C23 a_109_7# a_397_257# 0.00647f
C24 a_481_7# VGND 0.00561f
C25 A1_N VPB 0.0331f
C26 VGND VPB 0.00833f
C27 A1_N a_109_257# 8.3e-19
C28 B1 Y 0.00112f
C29 Y B2 0.0778f
C30 VGND a_109_257# 0.00196f
C31 a_481_7# Y 0.00154f
C32 B1 B2 0.118f
C33 a_481_7# B2 0.00732f
C34 Y VPB 0.0105f
C35 A2_N A1_N 0.0842f
C36 A2_N VGND 0.0187f
C37 B1 VPB 0.035f
C38 VPWR A1_N 0.0498f
C39 B2 VPB 0.0272f
C40 VPWR VGND 0.0681f
C41 VGND a_397_257# 0.00847f
C42 A1_N a_109_7# 0.0213f
C43 VGND a_109_7# 0.185f
C44 A2_N Y 5.53e-19
C45 VPWR Y 0.0595f
C46 Y a_397_257# 0.0601f
C47 VGND VNB 0.438f
C48 Y VNB 0.0102f
C49 VPWR VNB 0.354f
C50 B1 VNB 0.145f
C51 B2 VNB 0.0969f
C52 A2_N VNB 0.0969f
C53 A1_N VNB 0.141f
C54 VPB VNB 0.693f
C55 a_397_257# VNB 0.0287f
C56 a_109_7# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A a_75_172#
X0 a_75_172# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR a_75_172# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND a_75_172# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 a_75_172# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
C0 a_75_172# VPWR 0.134f
C1 VPB VPWR 0.0355f
C2 VGND X 0.0545f
C3 A X 8.48e-19
C4 a_75_172# VPB 0.0571f
C5 VGND A 0.0184f
C6 X VPWR 0.0896f
C7 VGND VPWR 0.0289f
C8 a_75_172# X 0.107f
C9 A VPWR 0.0217f
C10 VPB X 0.0128f
C11 VGND a_75_172# 0.105f
C12 VGND VPB 0.00507f
C13 a_75_172# A 0.178f
C14 VPB A 0.0525f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_172# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2 a_27_257# a_109_257#
+ a_373_7# a_109_7#
X0 VGND A2 a_373_7# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1 a_109_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3 X a_27_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 X a_27_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_27_257# B1 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_27_257# B1 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X9 a_373_7# A1 a_27_257# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_109_257# A2 0.00625f
C1 X a_373_7# 1.97e-19
C2 a_109_257# VGND 0.00426f
C3 VPWR A2 0.0178f
C4 VGND VPWR 0.0641f
C5 a_109_7# B2 4.58e-19
C6 B1 A2 1.81e-19
C7 VGND B1 0.0267f
C8 a_27_257# B2 0.0567f
C9 VGND a_109_7# 0.00792f
C10 A1 A2 0.0738f
C11 VGND A1 0.0137f
C12 a_109_257# VPB 0.00882f
C13 VPB VPWR 0.0714f
C14 a_27_257# A2 0.161f
C15 a_27_257# VGND 0.257f
C16 VPB B1 0.0317f
C17 a_109_257# X 0.00169f
C18 X VPWR 0.0914f
C19 a_373_7# VPWR 7.36e-19
C20 B2 A2 8.94e-20
C21 VPB A1 0.0387f
C22 VGND B2 0.0538f
C23 X B1 8.38e-20
C24 a_27_257# VPB 0.0591f
C25 VGND A2 0.0162f
C26 X A1 2.98e-19
C27 a_373_7# A1 0.00122f
C28 VPB B2 0.0299f
C29 a_27_257# X 0.108f
C30 a_27_257# a_373_7# 0.0134f
C31 a_109_257# VPWR 0.187f
C32 VPB A2 0.0284f
C33 VGND VPB 0.00746f
C34 X B2 3.26e-20
C35 a_109_257# B1 0.0106f
C36 VPWR B1 0.0139f
C37 a_109_7# VPWR 0.00104f
C38 X A2 0.0011f
C39 VGND X 0.0543f
C40 a_373_7# A2 6.81e-19
C41 VGND a_373_7# 0.00344f
C42 a_109_257# A1 0.0105f
C43 A1 VPWR 0.0168f
C44 a_109_257# a_27_257# 0.171f
C45 a_109_7# B1 0.00145f
C46 a_27_257# VPWR 0.13f
C47 A1 B1 0.0657f
C48 a_27_257# B1 0.0838f
C49 VPB X 0.011f
C50 a_109_257# B2 0.0015f
C51 VPWR B2 0.0126f
C52 a_27_257# a_109_7# 0.00393f
C53 a_27_257# A1 0.0839f
C54 B1 B2 0.0739f
C55 VGND VNB 0.421f
C56 X VNB 0.0917f
C57 VPWR VNB 0.328f
C58 A2 VNB 0.0927f
C59 A1 VNB 0.112f
C60 B1 VNB 0.112f
C61 B2 VNB 0.126f
C62 VPB VNB 0.693f
C63 a_109_257# VNB 0.00274f
C64 a_27_257# VNB 0.19f
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR VPB VNB A X a_110_7#
X0 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X25 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X26 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X27 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 VPWR VPB 0.184f
C1 A VGND 0.115f
C2 VPWR a_110_7# 0.67f
C3 A X 0.00292f
C4 VGND X 0.977f
C5 A VPB 0.133f
C6 VPB VGND 0.0114f
C7 A a_110_7# 0.307f
C8 a_110_7# VGND 0.512f
C9 VPB X 0.0315f
C10 a_110_7# X 1.62f
C11 VPB a_110_7# 0.528f
C12 VPWR A 0.112f
C13 VPWR VGND 0.187f
C14 VPWR X 1.36f
C15 VGND VNB 1.01f
C16 X VNB 0.111f
C17 VPWR VNB 0.835f
C18 A VNB 0.495f
C19 VPB VNB 1.85f
C20 a_110_7# VNB 1.73f
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 B1 Y A1 a_109_257# a_27_7#
X0 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 Y A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3 VGND A1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_27_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPB A2 0.0305f
C1 VPB A1 0.0327f
C2 VPB a_27_7# 8.4e-19
C3 a_109_257# VPWR 0.00401f
C4 Y VPB 0.00672f
C5 A2 VGND 0.0183f
C6 VGND A1 0.0163f
C7 a_27_7# VGND 0.142f
C8 VPB VPWR 0.056f
C9 Y VGND 0.0289f
C10 A2 A1 0.0986f
C11 A2 a_27_7# 0.0388f
C12 a_27_7# A1 0.037f
C13 Y A2 0.124f
C14 Y A1 8.9e-19
C15 Y a_27_7# 0.0517f
C16 VGND VPWR 0.0381f
C17 A2 VPWR 0.109f
C18 VPB B1 0.0741f
C19 VPWR A1 0.0497f
C20 a_27_7# VPWR 0.00663f
C21 Y VPWR 0.105f
C22 VGND B1 0.016f
C23 A2 B1 0.0472f
C24 a_27_7# B1 0.00471f
C25 Y B1 0.0811f
C26 VPWR B1 0.0433f
C27 a_109_257# VGND 4.56e-19
C28 A2 a_109_257# 0.00993f
C29 a_109_257# a_27_7# 5.37e-19
C30 VPB VGND 0.00462f
C31 Y a_109_257# 5.24e-19
C32 VGND VNB 0.254f
C33 Y VNB 0.0545f
C34 VPWR VNB 0.271f
C35 B1 VNB 0.152f
C36 A2 VNB 0.0962f
C37 A1 VNB 0.138f
C38 VPB VNB 0.428f
C39 a_27_7# VNB 0.0311f
.ends

.subckt sky130_fd_sc_hd__o221ai_4 VGND VPWR VPB VNB B2 Y A2 A1 B1 C1 a_553_257# a_1241_257#
+ a_471_7# a_27_7#
X0 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X16 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X23 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X30 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X36 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 B2 A2 5.76e-19
C1 B1 Y 0.36f
C2 VPWR a_27_7# 0.00762f
C3 VPWR a_471_7# 0.0133f
C4 VPB Y 0.0189f
C5 B1 a_1241_257# 9.99e-19
C6 a_1241_257# VPB 0.00652f
C7 Y VGND 0.0339f
C8 a_1241_257# VGND 0.00647f
C9 a_471_7# a_27_7# 0.33f
C10 VPWR Y 0.498f
C11 B1 A1 0.093f
C12 VPB A1 0.133f
C13 B1 a_553_257# 0.0481f
C14 VPWR a_1241_257# 0.465f
C15 VPB a_553_257# 0.00497f
C16 VGND A1 0.0628f
C17 Y a_27_7# 0.176f
C18 VGND a_553_257# 0.00615f
C19 a_471_7# Y 0.0206f
C20 VPWR A1 0.111f
C21 VPWR a_553_257# 0.409f
C22 a_471_7# A1 0.214f
C23 B1 C1 0.0183f
C24 B2 B1 0.254f
C25 a_1241_257# Y 0.172f
C26 a_471_7# a_553_257# 7.04e-20
C27 C1 VPB 0.131f
C28 B2 VPB 0.114f
C29 C1 VGND 0.0373f
C30 B2 VGND 0.0278f
C31 B1 A2 3.11e-19
C32 A2 VPB 0.115f
C33 A2 VGND 0.0584f
C34 Y A1 0.161f
C35 Y a_553_257# 0.286f
C36 VPWR C1 0.112f
C37 B2 VPWR 0.0281f
C38 a_1241_257# A1 0.154f
C39 a_1241_257# a_553_257# 6.98e-19
C40 VPWR A2 0.0341f
C41 C1 a_27_7# 0.0594f
C42 B2 a_27_7# 0.0264f
C43 a_471_7# C1 8.47e-20
C44 B2 a_471_7# 0.0835f
C45 a_553_257# A1 2.35e-20
C46 a_471_7# A2 0.182f
C47 C1 Y 0.324f
C48 B2 Y 0.0466f
C49 B2 a_1241_257# 1.52e-19
C50 A2 Y 0.0321f
C51 a_1241_257# A2 0.0414f
C52 B1 VPB 0.129f
C53 B2 A1 5.11e-19
C54 C1 a_553_257# 3.36e-19
C55 B2 a_553_257# 0.035f
C56 B1 VGND 0.0414f
C57 VPB VGND 0.0124f
C58 A2 A1 0.291f
C59 A2 a_553_257# 3e-20
C60 VPWR B1 0.0731f
C61 VPWR VPB 0.196f
C62 VPWR VGND 0.188f
C63 B1 a_27_7# 0.0242f
C64 B1 a_471_7# 0.215f
C65 VPB a_27_7# 3.53e-19
C66 a_471_7# VPB 0.00266f
C67 VGND a_27_7# 0.598f
C68 a_471_7# VGND 0.591f
C69 VGND VNB 1.03f
C70 Y VNB 0.0292f
C71 VPWR VNB 0.917f
C72 A2 VNB 0.352f
C73 A1 VNB 0.403f
C74 B2 VNB 0.351f
C75 B1 VNB 0.373f
C76 C1 VNB 0.41f
C77 VPB VNB 1.93f
C78 a_471_7# VNB 0.0538f
C79 a_27_7# VNB 0.0485f
C80 a_553_257# VNB 0.00146f
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X a_257_159# a_306_329#
+ a_79_n19# a_578_7# a_591_329# a_288_7#
X0 a_288_7# a_257_159# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X1 X a_79_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_257_159# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VPWR S a_591_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 a_591_329# A0 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND S a_578_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X7 a_257_159# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_79_n19# A1 a_306_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X9 a_578_7# A1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X10 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_79_n19# A0 a_288_7# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X13 a_306_329# a_257_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
C0 a_257_159# a_591_329# 0.00548f
C1 VGND a_578_7# 0.00424f
C2 a_79_n19# a_578_7# 9.96e-19
C3 VPB A1 0.0585f
C4 a_257_159# A0 0.159f
C5 VGND A1 0.0497f
C6 a_79_n19# A1 0.0307f
C7 VPB S 0.0987f
C8 VGND a_306_329# 0.00149f
C9 a_79_n19# a_306_329# 0.021f
C10 VGND S 0.0569f
C11 a_79_n19# S 0.00187f
C12 a_257_159# VPWR 0.149f
C13 a_257_159# X 0.00258f
C14 a_288_7# A1 3.38e-19
C15 a_591_329# VPWR 0.00489f
C16 VPWR A0 0.0177f
C17 a_257_159# VPB 0.108f
C18 a_257_159# VGND 0.0996f
C19 a_257_159# a_79_n19# 0.285f
C20 X VPWR 0.149f
C21 a_578_7# A1 0.00429f
C22 VGND a_591_329# 6.57e-19
C23 a_79_n19# a_591_329# 0.0015f
C24 VPB A0 0.0729f
C25 VGND A0 0.0185f
C26 a_79_n19# A0 0.0671f
C27 a_257_159# a_288_7# 4.59e-19
C28 VPB VPWR 0.0953f
C29 X VPB 0.00457f
C30 S A1 0.0662f
C31 VGND VPWR 0.0922f
C32 X VGND 0.109f
C33 a_79_n19# VPWR 0.25f
C34 X a_79_n19# 0.168f
C35 a_257_159# a_578_7# 4.09e-19
C36 a_288_7# VPWR 3.13e-19
C37 VGND VPB 0.011f
C38 a_79_n19# VPB 0.0731f
C39 a_257_159# A1 0.0371f
C40 VGND a_79_n19# 0.231f
C41 a_257_159# a_306_329# 0.0102f
C42 a_257_159# S 0.146f
C43 A1 A0 0.158f
C44 a_288_7# VGND 0.00186f
C45 a_578_7# VPWR 4.32e-19
C46 a_288_7# a_79_n19# 0.00727f
C47 S A0 0.0842f
C48 VPWR A1 0.00994f
C49 VPWR a_306_329# 0.00634f
C50 S VPWR 0.033f
C51 VGND VNB 0.516f
C52 X VNB 0.0244f
C53 VPWR VNB 0.441f
C54 S VNB 0.244f
C55 A0 VNB 0.129f
C56 A1 VNB 0.162f
C57 VPB VNB 0.871f
C58 a_257_159# VNB 0.216f
C59 a_79_n19# VNB 0.227f
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB X A1 A2 B1 C1 a_510_7# a_79_n19#
+ a_215_7# a_297_257#
X0 a_79_n19# C1 a_510_7# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X1 a_297_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 a_215_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND A1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_79_n19# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X6 VPWR B1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X7 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_510_7# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X9 a_79_n19# A2 a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
C0 X A2 2.44e-19
C1 a_79_n19# C1 0.0965f
C2 VGND a_79_n19# 0.126f
C3 B1 a_215_7# 0.00549f
C4 a_79_n19# a_297_257# 0.0174f
C5 VPB C1 0.0553f
C6 X VPWR 0.129f
C7 VGND VPB 0.0108f
C8 A1 a_215_7# 0.0493f
C9 a_79_n19# a_510_7# 0.00844f
C10 VGND A2 0.0159f
C11 C1 VPWR 0.0203f
C12 VGND VPWR 0.0732f
C13 VPWR a_297_257# 0.0107f
C14 a_510_7# VPWR 0.00153f
C15 a_79_n19# B1 0.0649f
C16 VPB B1 0.0298f
C17 a_79_n19# A1 0.0844f
C18 VGND X 0.0993f
C19 B1 A2 0.0611f
C20 VPB A1 0.0322f
C21 a_79_n19# a_215_7# 0.0458f
C22 VPWR B1 0.0185f
C23 A1 A2 0.0693f
C24 VGND C1 0.0133f
C25 VGND a_297_257# 0.002f
C26 VPB a_215_7# 9.29e-19
C27 A1 VPWR 0.0184f
C28 A2 a_215_7# 0.0461f
C29 VGND a_510_7# 0.00833f
C30 VPWR a_215_7# 0.00318f
C31 X B1 1.2e-19
C32 A1 X 3.68e-19
C33 C1 B1 0.0495f
C34 VGND B1 0.0186f
C35 VPB a_79_n19# 0.0755f
C36 X a_215_7# 5.57e-19
C37 VGND A1 0.017f
C38 a_79_n19# A2 0.0474f
C39 A1 a_297_257# 6.93e-20
C40 a_510_7# B1 0.00122f
C41 VPB A2 0.034f
C42 a_79_n19# VPWR 0.361f
C43 VGND a_215_7# 0.226f
C44 a_297_257# a_215_7# 1.98e-20
C45 VPB VPWR 0.0944f
C46 VPWR A2 0.0143f
C47 a_510_7# a_215_7# 0.00529f
C48 a_79_n19# X 0.0491f
C49 VPB X 0.0125f
C50 VGND VNB 0.45f
C51 VPWR VNB 0.377f
C52 X VNB 0.0951f
C53 C1 VNB 0.167f
C54 B1 VNB 0.095f
C55 A2 VNB 0.101f
C56 A1 VNB 0.0989f
C57 VPB VNB 0.782f
C58 a_215_7# VNB 0.0101f
C59 a_79_n19# VNB 0.225f
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB B2 A2 A1 B1 X a_78_159# a_493_257#
+ a_292_257# a_215_7#
X0 a_292_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X1 a_78_159# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_215_7# B2 a_78_159# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 VGND A2 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_215_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_493_257# A2 a_78_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X7 VGND a_78_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_78_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X9 a_78_159# B2 a_292_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
C0 a_215_7# a_78_159# 0.0907f
C1 VGND VPWR 0.0668f
C2 A1 VGND 0.0146f
C3 A2 VPB 0.0341f
C4 A1 VPWR 0.057f
C5 VPB X 0.0107f
C6 B1 a_78_159# 0.148f
C7 a_493_257# a_78_159# 3.15e-19
C8 VPB VGND 0.00596f
C9 B2 a_78_159# 0.0816f
C10 VPB VPWR 0.0744f
C11 A1 VPB 0.0319f
C12 B1 a_215_7# 0.00758f
C13 A2 a_78_159# 0.0707f
C14 X a_78_159# 0.105f
C15 a_493_257# a_215_7# 3.25e-19
C16 a_292_257# a_78_159# 0.013f
C17 B2 a_215_7# 0.0207f
C18 VGND a_78_159# 0.0684f
C19 a_78_159# VPWR 0.211f
C20 A1 a_78_159# 4.58e-19
C21 B1 B2 0.0815f
C22 A2 a_215_7# 0.0439f
C23 a_215_7# X 0.00228f
C24 B1 A2 3.91e-19
C25 B1 X 6.11e-19
C26 VPB a_78_159# 0.0517f
C27 A2 a_493_257# 0.0105f
C28 a_215_7# VGND 0.258f
C29 a_215_7# VPWR 0.00435f
C30 A1 a_215_7# 0.0498f
C31 B2 A2 0.0676f
C32 B2 X 1.65e-19
C33 B1 VGND 0.0119f
C34 B1 VPWR 0.0227f
C35 a_493_257# VGND 3.15e-19
C36 B2 a_292_257# 4.98e-20
C37 a_493_257# VPWR 0.00283f
C38 A1 a_493_257# 9.88e-20
C39 B2 VGND 0.0103f
C40 a_215_7# VPB 9.85e-19
C41 B2 VPWR 0.0104f
C42 A2 a_292_257# 4.41e-20
C43 a_292_257# X 4.46e-19
C44 B1 VPB 0.0388f
C45 A2 VGND 0.0153f
C46 VGND X 0.0472f
C47 A2 VPWR 0.12f
C48 X VPWR 0.0911f
C49 A1 A2 0.0879f
C50 B2 VPB 0.0281f
C51 VGND a_292_257# 0.00136f
C52 a_292_257# VPWR 0.00854f
C53 VGND VNB 0.403f
C54 VPWR VNB 0.359f
C55 X VNB 0.0884f
C56 A1 VNB 0.132f
C57 A2 VNB 0.0971f
C58 B2 VNB 0.0913f
C59 B1 VNB 0.11f
C60 VPB VNB 0.693f
C61 a_215_7# VNB 0.0357f
C62 a_78_159# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND VPB VNB X A1 A2 A3 B2 B1 a_323_257# a_227_7#
+ a_227_257# a_77_159# a_539_257#
X0 a_227_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_227_7# B1 a_77_159# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X2 a_539_257# B2 a_77_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3 VGND A2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_77_159# B2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X5 VGND a_77_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_227_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_323_257# A2 a_227_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X8 a_227_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X9 VPWR B1 a_539_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X10 VPWR a_77_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X11 a_77_159# A3 a_323_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
C0 X A1 0.00148f
C1 a_227_257# VPWR 0.00277f
C2 B2 B1 0.044f
C3 VPWR a_539_257# 0.00916f
C4 B2 VGND 0.0105f
C5 X VGND 0.103f
C6 a_323_257# a_227_7# 0.00186f
C7 B2 A3 0.102f
C8 X A3 1.25e-19
C9 VPWR a_227_7# 0.00742f
C10 a_77_159# B2 0.116f
C11 X a_77_159# 0.0928f
C12 a_323_257# VPWR 0.00357f
C13 A1 A2 0.0751f
C14 A2 VGND 0.0164f
C15 A1 VGND 0.0197f
C16 VPB B2 0.0338f
C17 X VPB 0.0157f
C18 VGND B1 0.0107f
C19 X a_227_257# 2.01e-21
C20 B2 a_539_257# 0.00242f
C21 A2 A3 0.106f
C22 a_77_159# A2 0.113f
C23 A1 a_77_159# 0.124f
C24 VGND A3 0.0131f
C25 a_77_159# B1 0.0468f
C26 a_77_159# VGND 0.0387f
C27 VPB A2 0.0335f
C28 B2 a_227_7# 0.0275f
C29 X a_227_7# 0.0071f
C30 VPB A1 0.029f
C31 VPB B1 0.0411f
C32 VPB VGND 0.00632f
C33 A2 a_227_257# 0.003f
C34 A1 a_227_257# 3.62e-20
C35 A2 a_539_257# 6.51e-19
C36 a_77_159# A3 0.0306f
C37 a_227_257# VGND 0.00113f
C38 VGND a_539_257# 0.00177f
C39 B2 VPWR 0.0122f
C40 X VPWR 0.102f
C41 VPB A3 0.033f
C42 VPB a_77_159# 0.0477f
C43 A2 a_227_7# 0.0413f
C44 A1 a_227_7# 0.0151f
C45 a_323_257# A2 0.0116f
C46 a_77_159# a_227_257# 0.0187f
C47 a_227_7# B1 0.0341f
C48 VGND a_227_7# 0.326f
C49 a_77_159# a_539_257# 0.0229f
C50 a_323_257# VGND 0.00153f
C51 A2 VPWR 0.0135f
C52 A1 VPWR 0.0187f
C53 VPWR B1 0.0467f
C54 VGND VPWR 0.0721f
C55 a_227_7# A3 0.0376f
C56 a_323_257# A3 0.00159f
C57 a_77_159# a_227_7# 0.0851f
C58 a_323_257# a_77_159# 0.0143f
C59 X B2 7.64e-20
C60 VPB a_227_7# 0.00182f
C61 VPWR A3 0.00881f
C62 a_77_159# VPWR 0.36f
C63 a_227_257# a_227_7# 0.00166f
C64 VPB VPWR 0.0832f
C65 B2 A2 4.92e-19
C66 X A2 2.33e-19
C67 VGND VNB 0.438f
C68 VPWR VNB 0.404f
C69 X VNB 0.101f
C70 B1 VNB 0.15f
C71 B2 VNB 0.0977f
C72 A3 VNB 0.0965f
C73 A2 VNB 0.0962f
C74 A1 VNB 0.0946f
C75 VPB VNB 0.782f
C76 a_227_7# VNB 0.0309f
C77 a_77_159# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X a_111_257# a_29_13# a_183_257#
X0 VGND A a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_29_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X2 a_111_257# C a_29_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_29_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_183_257# B a_111_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_29_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A a_183_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VGND C a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 A C 0.0343f
C1 a_111_257# VGND 3.96e-19
C2 VPWR VPB 0.0649f
C3 a_29_13# a_183_257# 0.00868f
C4 B a_29_13# 0.121f
C5 VGND a_29_13# 0.217f
C6 a_29_13# X 0.0991f
C7 a_111_257# VPWR 5.94e-19
C8 VPB a_29_13# 0.0491f
C9 VPWR a_29_13# 0.0833f
C10 B C 0.0802f
C11 VGND C 0.0161f
C12 a_111_257# a_29_13# 0.005f
C13 A a_183_257# 0.00239f
C14 B A 0.0787f
C15 A VGND 0.0187f
C16 VPB C 0.0396f
C17 VPWR C 0.00457f
C18 A X 0.00127f
C19 A VPB 0.0377f
C20 VPWR A 0.00936f
C21 a_29_13# C 0.0857f
C22 a_111_257# A 0.00223f
C23 VGND a_183_257# 5.75e-19
C24 B VGND 0.0152f
C25 B X 6.52e-19
C26 A a_29_13# 0.242f
C27 VGND X 0.036f
C28 VPWR a_183_257# 8.13e-19
C29 B VPB 0.0962f
C30 VPWR B 0.147f
C31 VGND VPB 0.00724f
C32 VPWR VGND 0.0459f
C33 VPB X 0.0109f
C34 VPWR X 0.0885f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_13# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB B1 B2 A2 A1 X C1 a_149_7# a_245_257#
+ a_240_7# a_51_257# a_512_257#
X0 a_245_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1 VPWR C1 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X2 a_512_257# A2 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
X3 a_149_7# B2 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_240_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A1 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_51_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_51_257# B2 a_245_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X8 a_240_7# B1 a_149_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X9 a_149_7# C1 a_51_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X10 VPWR A1 a_512_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X11 X a_51_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
C0 a_245_257# a_51_257# 0.0122f
C1 a_51_257# C1 0.102f
C2 a_240_7# VPWR 0.00289f
C3 B2 VPWR 0.0135f
C4 a_240_7# VGND 0.164f
C5 VGND B2 0.0107f
C6 VPB A2 0.0386f
C7 X VPWR 0.143f
C8 a_240_7# B1 0.0119f
C9 B2 B1 0.0797f
C10 VPB A1 0.0255f
C11 A1 A2 0.0801f
C12 a_240_7# a_149_7# 0.0687f
C13 a_149_7# B2 0.00653f
C14 VGND X 0.144f
C15 VPWR a_51_257# 0.414f
C16 X B1 8.13e-20
C17 VGND a_51_257# 0.0874f
C18 X a_512_257# 1.12e-19
C19 VPB a_240_7# 0.0014f
C20 a_240_7# A2 0.0566f
C21 VPB B2 0.0366f
C22 B2 A2 0.0746f
C23 B1 a_51_257# 0.0669f
C24 a_149_7# a_51_257# 0.0249f
C25 a_245_257# VPWR 0.00619f
C26 a_240_7# A1 0.023f
C27 VPWR C1 0.0201f
C28 a_512_257# a_51_257# 0.0116f
C29 a_245_257# VGND 0.001f
C30 VPB X 0.0262f
C31 A2 X 3.43e-19
C32 VGND C1 0.0141f
C33 A1 X 9.4e-19
C34 B1 C1 0.052f
C35 a_149_7# C1 0.00154f
C36 VPB a_51_257# 0.0632f
C37 A2 a_51_257# 0.0889f
C38 a_240_7# B2 0.0408f
C39 A1 a_51_257# 0.125f
C40 VGND VPWR 0.0799f
C41 B2 X 1.41e-19
C42 VPB C1 0.0515f
C43 B1 VPWR 0.0115f
C44 a_149_7# VPWR 0.00235f
C45 a_240_7# a_51_257# 0.0314f
C46 B2 a_51_257# 0.0773f
C47 VPWR a_512_257# 0.00729f
C48 VGND B1 0.00794f
C49 a_149_7# VGND 0.123f
C50 a_149_7# B1 0.017f
C51 VGND a_512_257# 7.75e-19
C52 X a_51_257# 0.101f
C53 VPB VPWR 0.0879f
C54 a_240_7# a_245_257# 7.75e-19
C55 A2 VPWR 0.0151f
C56 a_245_257# B2 7.41e-19
C57 a_240_7# C1 6.33e-20
C58 A1 VPWR 0.0215f
C59 VPB VGND 0.00816f
C60 VGND A2 0.0159f
C61 VPB B1 0.0251f
C62 VGND A1 0.0277f
C63 VPB a_149_7# 1.39e-19
C64 VGND VNB 0.494f
C65 X VNB 0.107f
C66 VPWR VNB 0.409f
C67 A1 VNB 0.0908f
C68 A2 VNB 0.107f
C69 B2 VNB 0.103f
C70 B1 VNB 0.0897f
C71 C1 VNB 0.164f
C72 VPB VNB 0.871f
C73 a_240_7# VNB 0.0138f
C74 a_149_7# VNB 0.00821f
C75 a_51_257# VNB 0.207f
.ends

.subckt sky130_fd_sc_hd__and3_2 VPWR VGND VPB VNB X C B A a_184_13# a_29_271# a_112_13#
X0 VGND C a_184_13# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
X1 VPWR a_29_271# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_29_271# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_29_271# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X4 VPWR A a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_184_13# B a_112_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR C a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X7 X a_29_271# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X8 a_112_13# A a_29_271# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND a_29_271# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 C VGND 0.0714f
C1 a_112_13# VPWR 1.15e-19
C2 X VPWR 0.193f
C3 B X 8.26e-19
C4 VPB a_29_271# 0.0835f
C5 C VPWR 0.00883f
C6 a_29_271# VGND 0.143f
C7 VPB VGND 0.00661f
C8 B C 0.0649f
C9 a_184_13# C 0.00415f
C10 a_29_271# A 0.134f
C11 VPB A 0.0443f
C12 A VGND 0.0127f
C13 C X 0.0158f
C14 a_29_271# VPWR 0.178f
C15 VPB VPWR 0.0929f
C16 VGND VPWR 0.0591f
C17 B a_29_271# 0.0596f
C18 B VPB 0.0923f
C19 a_29_271# a_184_13# 0.0026f
C20 B VGND 0.00756f
C21 a_112_13# a_29_271# 0.0049f
C22 A VPWR 0.0156f
C23 a_184_13# VGND 0.00302f
C24 a_29_271# X 0.125f
C25 VPB X 0.00641f
C26 a_112_13# VGND 5.13e-19
C27 B A 0.0835f
C28 X VGND 0.14f
C29 a_29_271# C 0.189f
C30 B VPWR 0.13f
C31 VPB C 0.0352f
C32 a_184_13# VPWR 4.26e-19
C33 VGND VNB 0.369f
C34 X VNB 0.04f
C35 C VNB 0.116f
C36 A VNB 0.17f
C37 VPWR VNB 0.336f
C38 B VNB 0.103f
C39 VPB VNB 0.605f
C40 a_29_271# VNB 0.271f
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND VPB VNB X D1 C1 B1 A2 A1 a_306_7# a_79_n19#
+ a_512_7# a_409_7# a_676_257#
X0 VPWR A1 a_676_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A2 a_512_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X2 a_512_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X4 a_79_n19# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X5 a_512_7# B1 a_409_7# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X6 a_676_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X7 a_306_7# D1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X8 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_409_7# C1 a_306_7# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X10 VPWR C1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X11 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
C0 VGND a_409_7# 0.00662f
C1 A2 A1 0.121f
C2 X VPWR 0.0949f
C3 A2 a_79_n19# 0.0969f
C4 a_306_7# a_512_7# 5.86e-19
C5 VGND C1 0.0342f
C6 VPB a_512_7# 9.45e-19
C7 VGND A1 0.0184f
C8 A1 a_676_257# 2.93e-19
C9 VGND a_79_n19# 0.142f
C10 a_79_n19# a_676_257# 2.93e-19
C11 A2 a_512_7# 0.0516f
C12 X a_79_n19# 0.091f
C13 B1 VPB 0.0377f
C14 VGND a_512_7# 0.17f
C15 a_676_257# a_512_7# 7.22e-19
C16 D1 VPWR 0.0233f
C17 B1 A2 0.0534f
C18 VPWR a_409_7# 0.0011f
C19 D1 C1 0.118f
C20 VGND B1 0.0325f
C21 D1 a_79_n19# 0.155f
C22 C1 VPWR 0.0217f
C23 C1 a_409_7# 0.00808f
C24 A2 VPB 0.0353f
C25 A1 VPWR 0.055f
C26 VPWR a_79_n19# 0.44f
C27 VGND a_306_7# 0.00515f
C28 a_79_n19# a_409_7# 0.00296f
C29 D1 a_512_7# 1.56e-19
C30 VGND VPB 0.00797f
C31 C1 a_79_n19# 0.0401f
C32 VPWR a_512_7# 0.00613f
C33 VGND A2 0.0191f
C34 X VPB 0.0108f
C35 A1 a_79_n19# 2.4e-19
C36 A2 a_676_257# 0.0099f
C37 a_409_7# a_512_7# 0.00102f
C38 C1 a_512_7# 3.26e-19
C39 VGND a_676_257# 4.92e-19
C40 A1 a_512_7# 0.0432f
C41 B1 VPWR 0.0218f
C42 a_79_n19# a_512_7# 0.0103f
C43 VGND X 0.0654f
C44 B1 a_409_7# 0.00322f
C45 D1 a_306_7# 0.0092f
C46 C1 B1 0.104f
C47 B1 A1 6.19e-19
C48 D1 VPB 0.0365f
C49 VPWR a_306_7# 8.85e-19
C50 B1 a_79_n19# 0.0351f
C51 D1 A2 1.08e-19
C52 VPWR VPB 0.0881f
C53 C1 a_306_7# 0.00228f
C54 A2 VPWR 0.0848f
C55 B1 a_512_7# 0.0468f
C56 VGND D1 0.0387f
C57 C1 VPB 0.0347f
C58 a_79_n19# a_306_7# 0.00291f
C59 A1 VPB 0.04f
C60 VGND VPWR 0.0865f
C61 C1 A2 2.05e-19
C62 D1 X 3.34e-19
C63 VPB a_79_n19# 0.0534f
C64 VPWR a_676_257# 0.00372f
C65 VGND VNB 0.491f
C66 VPWR VNB 0.414f
C67 X VNB 0.0907f
C68 A1 VNB 0.154f
C69 A2 VNB 0.104f
C70 B1 VNB 0.114f
C71 C1 VNB 0.0988f
C72 D1 VNB 0.112f
C73 VPB VNB 0.871f
C74 a_512_7# VNB 0.0326f
C75 a_79_n19# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VGND VPWR VPB VNB A2 A1 B1 B2 Y C1 a_27_257# a_301_257#
+ a_383_7# a_735_7#
X0 a_27_257# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_301_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X2 a_735_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X3 a_27_257# B1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X5 a_301_257# B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_301_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_257# B2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_301_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y C1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11 Y A1 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_735_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X15 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_383_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X17 Y B1 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_383_7# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND a_27_257# 0.00854f
C1 B1 VGND 0.0184f
C2 Y VGND 0.258f
C3 A2 B2 0.0926f
C4 B2 VPWR 0.0224f
C5 VGND C1 0.0632f
C6 B2 VPB 0.0679f
C7 B2 a_301_257# 0.0418f
C8 B2 a_27_257# 0.153f
C9 A2 VPWR 0.0455f
C10 A1 a_735_7# 0.0216f
C11 B1 B2 0.213f
C12 a_383_7# a_735_7# 2.58e-19
C13 A2 VPB 0.0709f
C14 VPWR VPB 0.108f
C15 B2 Y 0.118f
C16 A2 a_301_257# 0.186f
C17 A2 a_27_257# 1.13e-19
C18 VPWR a_301_257# 0.48f
C19 VPWR a_27_257# 0.164f
C20 a_301_257# VPB 0.0181f
C21 B1 VPWR 0.0152f
C22 a_27_257# VPB 0.0204f
C23 A2 Y 0.0455f
C24 Y VPWR 0.0129f
C25 B1 VPB 0.051f
C26 a_27_257# a_301_257# 0.191f
C27 VGND a_735_7# 0.206f
C28 B2 C1 0.0205f
C29 Y VPB 0.00812f
C30 B1 a_301_257# 0.0185f
C31 B1 a_27_257# 0.0195f
C32 Y a_301_257# 0.00522f
C33 Y a_27_257# 0.128f
C34 B1 Y 0.0643f
C35 VPWR C1 0.0192f
C36 A1 VGND 0.0175f
C37 VGND a_383_7# 0.165f
C38 C1 VPB 0.078f
C39 C1 a_27_257# 0.0611f
C40 B2 a_735_7# 1.28e-19
C41 Y C1 0.106f
C42 A2 a_735_7# 0.0309f
C43 VPWR a_735_7# 0.00213f
C44 B2 a_383_7# 0.00622f
C45 a_735_7# VPB 2.96e-19
C46 A2 A1 0.207f
C47 B1 a_735_7# 1.04e-19
C48 A1 VPWR 0.0298f
C49 VPWR a_383_7# 0.00192f
C50 Y a_735_7# 0.0886f
C51 A1 VPB 0.051f
C52 B2 VGND 0.0325f
C53 A1 a_301_257# 0.0293f
C54 A1 a_27_257# 1.01e-19
C55 B1 a_383_7# 0.0137f
C56 A2 VGND 0.0568f
C57 A1 Y 0.0483f
C58 C1 a_735_7# 1.39e-20
C59 Y a_383_7# 0.0983f
C60 VPWR VGND 0.106f
C61 VGND VPB 0.00991f
C62 VGND a_301_257# 0.00922f
C63 VGND VNB 0.682f
C64 VPWR VNB 0.52f
C65 Y VNB 0.0379f
C66 A1 VNB 0.166f
C67 A2 VNB 0.23f
C68 B1 VNB 0.166f
C69 B2 VNB 0.195f
C70 C1 VNB 0.255f
C71 VPB VNB 1.14f
C72 a_735_7# VNB 0.00532f
C73 a_383_7# VNB 0.00406f
C74 a_301_257# VNB 0.0376f
C75 a_27_257# VNB 0.0292f
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB A Y B a_113_7#
X0 Y A a_113_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_113_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 Y a_113_7# 0.00937f
C1 B VPWR 0.0478f
C2 Y A 0.0855f
C3 Y B 0.0481f
C4 VGND VPB 0.0044f
C5 B A 0.051f
C6 VGND VPWR 0.0322f
C7 VPB VPWR 0.0509f
C8 Y VGND 0.139f
C9 a_113_7# VGND 0.0019f
C10 Y VPB 0.00618f
C11 VGND A 0.00949f
C12 VPB A 0.0379f
C13 Y VPWR 0.211f
C14 a_113_7# VPWR 1.78e-19
C15 VGND B 0.0544f
C16 VPB B 0.0391f
C17 A VPWR 0.0444f
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR VPB VNB X C B A a_27_7# a_109_7# a_181_7#
X0 a_27_7# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_181_7# B a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5 VGND C a_181_7# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_109_7# A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
C0 a_27_7# X 0.087f
C1 VPB a_27_7# 0.0501f
C2 a_181_7# a_27_7# 0.00401f
C3 B VGND 0.00714f
C4 B VPWR 0.128f
C5 C VGND 0.0703f
C6 C VPWR 0.00464f
C7 A a_109_7# 6.45e-19
C8 A VGND 0.0154f
C9 A VPWR 0.0185f
C10 B X 0.00111f
C11 B VPB 0.0836f
C12 C X 0.0149f
C13 C VPB 0.0347f
C14 C a_181_7# 0.00151f
C15 A VPB 0.0426f
C16 B a_27_7# 0.0625f
C17 C a_27_7# 0.186f
C18 VGND a_109_7# 0.00123f
C19 A a_27_7# 0.157f
C20 VPWR a_109_7# 3.29e-19
C21 VGND VPWR 0.0475f
C22 C B 0.0746f
C23 VGND X 0.0708f
C24 VGND VPB 0.00604f
C25 A B 0.0869f
C26 a_181_7# VGND 0.00261f
C27 VPWR X 0.0766f
C28 VPWR VPB 0.0795f
C29 a_181_7# VPWR 3.97e-19
C30 a_27_7# a_109_7# 0.00517f
C31 VGND a_27_7# 0.134f
C32 VPWR a_27_7# 0.145f
C33 VPB X 0.0121f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_7# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR VPB VNB A1 A2 B1 B2 Y a_109_257# a_307_257#
+ a_27_7#
X0 Y B2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X1 a_109_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X3 a_27_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X5 VPWR A1 a_307_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X6 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_307_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
C0 Y A1 5.15e-19
C1 VPB a_27_7# 9.43e-19
C2 A2 VPB 0.0309f
C3 VGND VPWR 0.0459f
C4 Y a_27_7# 0.0527f
C5 a_307_257# VPWR 0.00219f
C6 A2 Y 0.063f
C7 VGND B1 0.0142f
C8 VGND A1 0.0147f
C9 a_109_257# VPWR 0.00394f
C10 VPB Y 0.00499f
C11 B2 VPWR 0.0114f
C12 VGND a_27_7# 0.244f
C13 VGND A2 0.0158f
C14 B2 B1 0.0576f
C15 a_307_257# a_27_7# 2.6e-19
C16 B2 A1 4.27e-19
C17 a_307_257# A2 0.0107f
C18 a_109_257# A2 3.1e-19
C19 VGND VPB 0.0047f
C20 B2 a_27_7# 0.0266f
C21 B2 A2 0.091f
C22 VGND Y 0.00968f
C23 a_307_257# Y 3.52e-19
C24 B1 VPWR 0.0451f
C25 VPWR A1 0.0569f
C26 B2 VPB 0.0302f
C27 a_109_257# Y 0.0135f
C28 B2 Y 0.12f
C29 VPWR a_27_7# 0.00678f
C30 VGND a_307_257# 2.4e-19
C31 A2 VPWR 0.119f
C32 B1 a_27_7# 0.0334f
C33 a_27_7# A1 0.0495f
C34 A2 A1 0.089f
C35 a_109_257# VGND 9.92e-19
C36 VPWR VPB 0.0612f
C37 B1 VPB 0.0427f
C38 VPB A1 0.0315f
C39 B2 VGND 0.0105f
C40 A2 a_27_7# 0.046f
C41 VPWR Y 0.102f
C42 a_109_257# B2 5.79e-19
C43 B1 Y 0.132f
C44 VGND VNB 0.298f
C45 Y VNB 0.0144f
C46 VPWR VNB 0.298f
C47 A1 VNB 0.131f
C48 A2 VNB 0.0973f
C49 B2 VNB 0.0939f
C50 B1 VNB 0.184f
C51 VPB VNB 0.516f
C52 a_27_7# VNB 0.0465f
.ends

.subckt sky130_fd_sc_hd__or3_4 VPWR VGND VPB VNB B C A X a_109_257# a_27_7# a_193_257#
X0 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_109_257# C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X4 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR A a_193_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X8 a_193_257# B a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND C a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X12 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B a_193_257# 0.00132f
C1 X VGND 0.265f
C2 VGND a_193_257# 2.86e-19
C3 B a_109_257# 0.00939f
C4 VGND a_109_257# 7.33e-19
C5 X VPB 0.0146f
C6 A a_27_7# 0.159f
C7 X VPWR 0.365f
C8 VPWR a_193_257# 8.05e-19
C9 a_27_7# B 0.19f
C10 VGND a_27_7# 0.352f
C11 VPWR a_109_257# 0.00187f
C12 a_27_7# C 0.0996f
C13 VPB a_27_7# 0.158f
C14 a_27_7# VPWR 0.363f
C15 A B 0.0783f
C16 A VGND 0.0164f
C17 VGND B 0.0163f
C18 B C 0.0864f
C19 A VPB 0.0324f
C20 VGND C 0.0149f
C21 VPB B 0.0302f
C22 A VPWR 0.0196f
C23 VPB VGND 0.00698f
C24 B VPWR 0.0132f
C25 VGND VPWR 0.0864f
C26 X a_27_7# 0.397f
C27 VPB C 0.0369f
C28 a_27_7# a_193_257# 0.015f
C29 a_27_7# a_109_257# 0.0105f
C30 C VPWR 0.00921f
C31 VPB VPWR 0.0867f
C32 A X 5.59e-19
C33 A a_193_257# 3.02e-21
C34 VGND VNB 0.493f
C35 X VNB 0.0611f
C36 VPWR VNB 0.418f
C37 A VNB 0.0987f
C38 B VNB 0.0938f
C39 C VNB 0.141f
C40 VPB VNB 0.871f
C41 a_27_7# VNB 0.499f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 B2 A2_N A1_N X a_226_257# a_76_159#
+ a_556_7# a_226_7# a_489_373#
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X1 a_226_7# A2_N a_226_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_76_159# a_226_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X3 a_556_7# B2 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_226_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X5 VGND B1 a_556_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_226_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X7 VGND A2_N a_226_7# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_489_373# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VPWR B2 a_489_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_489_373# a_226_7# a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_76_159# X 0.0995f
C1 a_76_159# A1_N 0.119f
C2 B2 a_226_7# 0.0975f
C3 VGND VPB 0.0128f
C4 a_226_257# A1_N 0.00184f
C5 VGND VPWR 0.0743f
C6 a_76_159# VGND 0.108f
C7 A2_N X 2.55e-19
C8 a_489_373# a_226_7# 0.00579f
C9 A2_N A1_N 0.11f
C10 a_226_7# X 0.0108f
C11 VGND a_226_257# 5.63e-19
C12 B2 B1 0.182f
C13 A1_N a_226_7# 0.0209f
C14 VPWR VPB 0.0951f
C15 a_556_7# B2 0.00291f
C16 a_76_159# VPB 0.0817f
C17 A2_N VGND 0.0174f
C18 a_76_159# VPWR 0.2f
C19 a_489_373# B2 0.0541f
C20 a_489_373# B1 0.0382f
C21 VGND a_226_7# 0.149f
C22 VPWR a_226_257# 8.54e-19
C23 a_76_159# a_226_257# 0.00354f
C24 A2_N VPB 0.0327f
C25 A2_N VPWR 0.00449f
C26 VPB a_226_7# 0.111f
C27 VGND B2 0.0335f
C28 VGND B1 0.0471f
C29 VPWR a_226_7# 0.0187f
C30 A1_N X 0.00211f
C31 a_76_159# A2_N 0.0125f
C32 VGND a_556_7# 0.00639f
C33 a_76_159# a_226_7# 0.188f
C34 a_489_373# VGND 0.0058f
C35 a_226_257# a_226_7# 0.00128f
C36 VGND X 0.0627f
C37 VPB B2 0.0645f
C38 VPB B1 0.0803f
C39 VGND A1_N 0.0261f
C40 VPWR B2 0.0161f
C41 VPWR B1 0.0188f
C42 a_556_7# VPWR 7.24e-19
C43 a_76_159# B2 0.0626f
C44 A2_N a_226_7# 0.141f
C45 a_76_159# B1 0.00185f
C46 a_489_373# VPB 0.015f
C47 a_76_159# a_556_7# 0.0017f
C48 VPB X 0.0113f
C49 a_489_373# VPWR 0.143f
C50 VPB A1_N 0.0339f
C51 VPWR X 0.0589f
C52 VPWR A1_N 0.00672f
C53 a_76_159# a_489_373# 0.0473f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_373# VNB 0.0254f
C63 a_226_7# VNB 0.162f
C64 a_76_159# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A a_27_257#
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_257# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VPWR A a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
C0 Y a_27_257# 0.152f
C1 B a_27_257# 0.0451f
C2 VGND VPWR 0.0467f
C3 VPWR VPB 0.05f
C4 Y A 0.0523f
C5 B A 0.0712f
C6 VGND VPB 0.00613f
C7 VPWR Y 0.0127f
C8 B VPWR 0.0174f
C9 a_27_257# A 0.0889f
C10 VGND Y 0.289f
C11 VGND B 0.0294f
C12 VPB Y 0.00961f
C13 B VPB 0.0566f
C14 VPWR a_27_257# 0.321f
C15 VGND a_27_257# 0.00726f
C16 VPWR A 0.0418f
C17 VPB a_27_257# 0.0203f
C18 B Y 0.179f
C19 VGND A 0.0597f
C20 VPB A 0.0563f
C21 VGND VNB 0.343f
C22 Y VNB 0.0641f
C23 VPWR VNB 0.249f
C24 B VNB 0.198f
C25 A VNB 0.207f
C26 VPB VNB 0.516f
C27 a_27_257# VNB 0.0647f
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X A B a_145_35# a_59_35#
X0 a_145_35# A a_59_35# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1 VPWR B a_59_35# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 X a_59_35# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3 VGND B a_145_35# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_59_35# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5 X a_59_35# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
C0 VPWR X 0.111f
C1 a_59_35# a_145_35# 0.00658f
C2 A VPWR 0.0362f
C3 a_145_35# VGND 0.00468f
C4 a_59_35# VPB 0.0563f
C5 A X 1.68e-19
C6 VGND VPB 0.008f
C7 a_59_35# VGND 0.116f
C8 B VPB 0.0629f
C9 a_59_35# B 0.143f
C10 VGND B 0.0115f
C11 VPWR a_145_35# 6.31e-19
C12 VPWR VPB 0.0729f
C13 a_145_35# X 5.76e-19
C14 a_59_35# VPWR 0.15f
C15 X VPB 0.0127f
C16 VPWR VGND 0.0461f
C17 A VPB 0.0806f
C18 a_59_35# X 0.109f
C19 a_59_35# A 0.0809f
C20 VPWR B 0.0117f
C21 VGND X 0.0993f
C22 A VGND 0.0147f
C23 B X 0.00276f
C24 A B 0.0971f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_35# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__or4b_4 VGND VPWR VPB VNB X D_N C B A a_403_257# a_215_257#
+ a_487_257# a_109_53# a_297_257#
X0 a_297_257# a_109_53# a_215_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X1 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_215_257# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.165 ps=1.82 w=0.65 l=0.15
X8 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X9 VPWR A a_487_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_487_257# B a_403_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND C a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X13 a_215_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_403_257# C a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X15 VGND A a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X17 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 a_487_257# a_215_257# 0.00167f
C1 C D_N 6.87e-19
C2 a_487_257# A 7.1e-19
C3 a_487_257# X 5.61e-19
C4 VPWR VPB 0.117f
C5 VPWR a_109_53# 0.0693f
C6 VPB a_109_53# 0.0623f
C7 B a_215_257# 0.0415f
C8 a_403_257# a_215_257# 0.00122f
C9 VPWR a_297_257# 0.00828f
C10 a_297_257# a_109_53# 3.03e-20
C11 B A 0.108f
C12 X B 0.0046f
C13 VGND VPWR 0.103f
C14 VGND VPB 0.0105f
C15 VGND a_109_53# 0.0965f
C16 D_N B 3.04e-19
C17 VGND a_297_257# 0.00213f
C18 C VPWR 0.0452f
C19 C VPB 0.0292f
C20 C a_109_53# 0.046f
C21 A a_215_257# 0.111f
C22 X a_215_257# 0.366f
C23 a_487_257# VPWR 0.0056f
C24 C a_297_257# 0.0109f
C25 a_487_257# a_109_53# 8.62e-21
C26 D_N a_215_257# 0.00255f
C27 X A 0.0157f
C28 C VGND 0.017f
C29 D_N A 7.84e-20
C30 D_N X 3.65e-19
C31 VPWR B 0.0819f
C32 a_487_257# VGND 1e-18
C33 B VPB 0.0282f
C34 VPWR a_403_257# 0.00597f
C35 B a_109_53# 4.77e-21
C36 a_403_257# a_109_53# 1.29e-20
C37 VGND B 0.0177f
C38 VGND a_403_257# 0.00131f
C39 VPWR a_215_257# 0.154f
C40 VPB a_215_257# 0.133f
C41 a_215_257# a_109_53# 0.152f
C42 C B 0.161f
C43 VPWR A 0.0526f
C44 VPWR X 0.358f
C45 VPB A 0.031f
C46 X VPB 0.0127f
C47 C a_403_257# 0.011f
C48 a_215_257# a_297_257# 0.0145f
C49 A a_109_53# 3.09e-21
C50 D_N VPWR 0.0486f
C51 D_N VPB 0.107f
C52 a_487_257# B 0.0126f
C53 D_N a_109_53# 0.119f
C54 VGND a_215_257# 0.294f
C55 VGND A 0.0184f
C56 VGND X 0.245f
C57 C a_215_257# 0.126f
C58 D_N VGND 0.0426f
C59 a_403_257# B 0.00615f
C60 VGND VNB 0.631f
C61 X VNB 0.0581f
C62 VPWR VNB 0.515f
C63 A VNB 0.0911f
C64 B VNB 0.0892f
C65 C VNB 0.0908f
C66 D_N VNB 0.186f
C67 VPB VNB 1.05f
C68 a_215_257# VNB 0.414f
C69 a_109_53# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VPWR VGND VPB VNB B1 Y A1 A2 A3 a_27_257# a_27_7#
+ a_277_7#
X0 VPWR A3 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR A1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_277_7# A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_277_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X7 a_27_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X9 a_27_7# A2 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A1 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_27_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X14 VGND A3 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 Y B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
C0 a_277_7# A2 0.0093f
C1 a_27_7# VPB 9.31e-19
C2 VGND B1 0.0344f
C3 A3 VGND 0.0355f
C4 a_27_7# a_27_257# 0.0108f
C5 A1 B1 0.0382f
C6 Y B1 0.177f
C7 a_27_7# VPWR 0.00469f
C8 Y A3 3.4e-19
C9 a_27_7# VGND 0.0907f
C10 a_27_7# A1 0.0129f
C11 a_27_7# Y 0.0142f
C12 VPB A2 0.0568f
C13 a_27_257# a_277_7# 1.45e-19
C14 a_277_7# VPWR 0.00227f
C15 a_27_257# A2 0.0837f
C16 VPWR A2 0.0396f
C17 VGND a_277_7# 0.169f
C18 VGND A2 0.0246f
C19 A1 a_277_7# 0.0176f
C20 Y a_277_7# 0.086f
C21 A1 A2 0.0965f
C22 Y A2 7.37e-19
C23 a_27_7# A3 0.0773f
C24 a_27_257# VPB 0.0116f
C25 VPB VPWR 0.0885f
C26 a_27_257# VPWR 0.558f
C27 VGND VPB 0.00575f
C28 A1 VPB 0.0971f
C29 Y VPB 0.00779f
C30 a_27_257# VGND 0.0107f
C31 VGND VPWR 0.0914f
C32 a_27_257# A1 0.0972f
C33 a_27_257# Y 0.13f
C34 A3 a_277_7# 7.39e-19
C35 A1 VPWR 0.0475f
C36 Y VPWR 0.0196f
C37 A3 A2 0.106f
C38 A1 VGND 0.0281f
C39 Y VGND 0.168f
C40 a_27_7# a_277_7# 0.0683f
C41 A1 Y 0.118f
C42 a_27_7# A2 0.074f
C43 VPB B1 0.0808f
C44 A3 VPB 0.0731f
C45 a_27_257# B1 0.045f
C46 a_27_257# A3 0.083f
C47 B1 VPWR 0.0218f
C48 A3 VPWR 0.0415f
C49 VGND VNB 0.538f
C50 Y VNB 0.06f
C51 VPWR VNB 0.436f
C52 B1 VNB 0.258f
C53 A1 VNB 0.24f
C54 A2 VNB 0.179f
C55 A3 VNB 0.246f
C56 VPB VNB 0.959f
C57 a_277_7# VNB 0.00976f
C58 a_27_7# VNB 0.0193f
C59 a_27_257# VNB 0.0672f
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR VPB VNB A1 A2 Y B2 C1 B1 a_213_83# a_295_257#
+ a_493_257# a_109_7#
X0 a_213_83# B2 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y B2 a_295_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 VGND A2 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X4 a_213_83# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_295_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X6 a_493_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X7 a_109_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X9 a_109_7# B1 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
C0 B2 a_109_7# 0.00286f
C1 VGND a_109_7# 0.115f
C2 A2 A1 0.0891f
C3 a_493_257# Y 3.47e-19
C4 B2 B1 0.0868f
C5 VGND B1 0.0106f
C6 a_295_257# B2 5.73e-20
C7 a_213_83# B2 0.0489f
C8 B2 Y 0.0569f
C9 VGND a_295_257# 0.00139f
C10 VGND a_213_83# 0.167f
C11 VGND Y 0.046f
C12 a_213_83# A1 0.0506f
C13 Y A1 3.82e-19
C14 C1 a_109_7# 0.00243f
C15 A2 VPWR 0.115f
C16 VPB B2 0.028f
C17 VGND VPB 0.0063f
C18 C1 B1 0.0209f
C19 a_109_7# VPWR 0.0018f
C20 C1 a_213_83# 1.34e-19
C21 C1 Y 0.127f
C22 B1 VPWR 0.0222f
C23 VPB A1 0.0359f
C24 a_295_257# VPWR 0.00875f
C25 a_213_83# VPWR 0.004f
C26 VGND a_493_257# 9.1e-20
C27 Y VPWR 0.293f
C28 VGND B2 0.0119f
C29 C1 VPB 0.038f
C30 B2 A1 5.58e-19
C31 VGND A1 0.0151f
C32 A2 B1 4.14e-19
C33 VPB VPWR 0.0746f
C34 a_295_257# A2 4.69e-20
C35 a_213_83# A2 0.0451f
C36 Y A2 0.0805f
C37 a_109_7# B1 0.00614f
C38 C1 VGND 0.0128f
C39 a_213_83# a_109_7# 0.0875f
C40 a_109_7# Y 0.0456f
C41 a_493_257# VPWR 8.66e-19
C42 B2 VPWR 0.00898f
C43 VGND VPWR 0.0645f
C44 a_213_83# B1 0.0383f
C45 Y B1 0.0768f
C46 VPB A2 0.0328f
C47 a_295_257# a_213_83# 1.01e-20
C48 a_295_257# Y 0.0137f
C49 a_213_83# Y 0.0301f
C50 A1 VPWR 0.0503f
C51 VPB a_109_7# 4.01e-19
C52 a_493_257# A2 0.0112f
C53 VPB B1 0.0341f
C54 B2 A2 0.0666f
C55 VGND A2 0.0162f
C56 a_213_83# VPB 0.00108f
C57 VPB Y 0.0205f
C58 C1 VPWR 0.0213f
C59 VGND VNB 0.39f
C60 VPWR VNB 0.362f
C61 Y VNB 0.0858f
C62 A1 VNB 0.14f
C63 A2 VNB 0.0967f
C64 B2 VNB 0.0933f
C65 B1 VNB 0.106f
C66 C1 VNB 0.145f
C67 VPB VNB 0.693f
C68 a_213_83# VNB 0.0371f
C69 a_109_7# VNB 0.0115f
.ends
