magic
tech sky130B
magscale 1 2
timestamp 1696628412
<< locali >>
rect -3060 974 -3014 980
rect -3060 -23 -3014 928
rect -1774 928 -1772 974
rect -1818 746 -1772 928
rect -1818 712 -1812 746
rect -1778 712 -1772 746
rect -1818 706 -1772 712
rect -730 463 -684 924
rect -730 429 -724 463
rect -690 429 -684 463
rect -730 423 -684 429
rect -211 447 -167 921
rect -211 413 -206 447
rect -172 413 -167 447
rect -211 408 -167 413
rect -3060 -57 -3054 -23
rect -3020 -57 -3014 -23
rect -3060 -63 -3014 -57
rect -554 -333 -520 -293
rect 4 -320 38 -299
rect -554 -367 -357 -333
rect 4 -354 201 -320
rect -3523 -394 -3493 -390
rect -3525 -502 -3491 -394
rect -3288 -502 -3254 -375
rect -3525 -505 -3254 -502
rect -3055 -505 -3021 -368
rect -2814 -505 -2780 -370
rect -3525 -513 -2780 -505
rect -1928 -513 -1893 -388
rect -1692 -513 -1657 -385
rect -946 -513 -911 -381
rect -554 -513 -520 -367
rect -4358 -516 -520 -513
rect 4 -516 38 -354
rect -4358 -547 38 -516
rect -554 -550 38 -547
<< viali >>
rect -3060 928 -3014 974
rect -1818 928 -1774 974
rect -1812 712 -1778 746
rect -730 924 -684 970
rect -724 429 -690 463
rect -211 921 -167 965
rect -206 413 -172 447
rect -3054 -57 -3020 -23
<< metal1 >>
rect -3060 986 -3014 1059
rect -1818 986 -1774 1054
rect -3066 974 -3008 986
rect -3066 928 -3060 974
rect -3014 928 -3008 974
rect -3066 916 -3008 928
rect -1824 974 -1768 986
rect -730 982 -684 1059
rect -1824 928 -1818 974
rect -1774 928 -1768 974
rect -1824 916 -1768 928
rect -736 970 -678 982
rect -211 971 -167 1059
rect -736 924 -730 970
rect -684 924 -678 970
rect -736 912 -678 924
rect -223 965 -155 971
rect -223 921 -211 965
rect -167 921 -155 965
rect -223 915 -155 921
rect -4166 845 267 874
rect -4166 -1453 -4137 845
rect -1818 746 -1772 758
rect -1818 712 -1812 746
rect -1778 712 -1772 746
rect -3990 52 -2145 81
rect -3060 -23 -3014 -11
rect -3060 -57 -3054 -23
rect -3020 -57 -3014 -23
rect -3060 -157 -3014 -57
rect -3596 -203 -2709 -157
rect -3640 -465 -3611 -352
rect -3405 -465 -3376 -360
rect -3171 -465 -3142 -363
rect -2931 -465 -2902 -335
rect -3640 -466 -2902 -465
rect -2698 -466 -2669 -325
rect -3640 -494 -2669 -466
rect -2310 -460 -2281 52
rect -1818 -157 -1772 712
rect -730 463 -684 475
rect -730 429 -724 463
rect -690 429 -684 463
rect -1584 46 -946 77
rect -1998 -203 -1586 -157
rect -1118 -250 -1087 46
rect -730 -156 -684 429
rect -212 447 -166 459
rect -212 413 -206 447
rect -172 413 -166 447
rect -212 401 -166 413
rect -1019 -202 -684 -156
rect -375 -225 -344 95
rect -1118 -281 -1028 -250
rect -2045 -460 -2016 -384
rect -1807 -460 -1778 -381
rect -2310 -462 -1778 -460
rect -1569 -462 -1540 -382
rect -2310 -489 -1540 -462
rect -1059 -458 -1028 -281
rect -211 -309 -167 401
rect 230 -216 261 104
rect 523 -254 573 1055
rect 350 -304 573 -254
rect -826 -458 -795 -343
rect -1059 -489 -795 -458
rect -1807 -491 -1540 -489
rect -3640 -657 -3611 -494
rect -2931 -495 -2669 -494
rect -3950 -686 315 -657
rect -4166 -1459 -3686 -1453
rect -4166 -1482 313 -1459
rect -3952 -1488 313 -1482
use sky130_fd_pr__nfet_01v8_lvt_3SNHZA  sky130_fd_pr__nfet_01v8_lvt_3SNHZA_0
timestamp 1696623266
transform 1 0 -3154 0 1 -304
box -639 -279 639 279
use sky130_fd_pr__nfet_01v8_lvt_763N5J  sky130_fd_pr__nfet_01v8_lvt_763N5J_0
timestamp 1696622261
transform 0 1 -311 -1 0 -291
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt_763N5J  sky130_fd_pr__nfet_01v8_lvt_763N5J_1
timestamp 1696622261
transform 0 1 248 -1 0 -278
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt_FS2HZA  sky130_fd_pr__nfet_01v8_lvt_FS2HZA_0
timestamp 1696623140
transform 1 0 -1792 0 1 -304
box -403 -279 403 279
use sky130_fd_pr__nfet_01v8_lvt_THUHZA  sky130_fd_pr__nfet_01v8_lvt_THUHZA_0
timestamp 1696623031
transform 1 0 -929 0 1 -304
box -285 -279 285 279
use trimcap  trimcap_0
timestamp 1696628372
transform 1 0 -4214 0 1 -374
box 0 376 480 1324
use trimcap  trimcap_1
timestamp 1696628372
transform 1 0 -3608 0 1 -378
box 0 376 480 1324
use trimcap  trimcap_2
timestamp 1696628372
transform 1 0 -3006 0 1 -372
box 0 376 480 1324
use trimcap  trimcap_3
timestamp 1696628372
transform 1 0 -2400 0 1 -376
box 0 376 480 1324
use trimcap  trimcap_4
timestamp 1696628372
transform 1 0 -1198 0 1 -371
box 0 376 480 1324
use trimcap  trimcap_5
timestamp 1696628372
transform 1 0 -1806 0 1 -372
box 0 376 480 1324
use trimcap  trimcap_6
timestamp 1696628372
transform 1 0 -598 0 1 -370
box 0 376 480 1324
use trimcap  trimcap_7
timestamp 1696628372
transform 1 0 8 0 1 -374
box 0 376 480 1324
use trimcap  trimcap_8
timestamp 1696628372
transform 1 0 -2393 0 -1 -211
box 0 376 480 1324
use trimcap  trimcap_9
timestamp 1696628372
transform 1 0 -2999 0 -1 -215
box 0 376 480 1324
use trimcap  trimcap_10
timestamp 1696628372
transform 1 0 -3601 0 -1 -209
box 0 376 480 1324
use trimcap  trimcap_11
timestamp 1696628372
transform 1 0 -4207 0 -1 -213
box 0 376 480 1324
use trimcap  trimcap_12
timestamp 1696628372
transform 1 0 -1193 0 -1 -211
box 0 376 480 1324
use trimcap  trimcap_13
timestamp 1696628372
transform 1 0 -1799 0 -1 -215
box 0 376 480 1324
use trimcap  trimcap_14
timestamp 1696628372
transform 1 0 15 0 -1 -213
box 0 376 480 1324
use trimcap  trimcap_15
timestamp 1696628372
transform 1 0 -591 0 -1 -217
box 0 376 480 1324
<< labels >>
flabel metal1 -3640 -686 -3611 -352 0 FreeSans 480 0 0 0 n4
flabel metal1 -2310 -489 -2281 81 0 FreeSans 480 0 0 0 n3
flabel metal1 -1118 -281 -1087 77 0 FreeSans 480 0 0 0 n2
flabel metal1 -375 -225 -344 95 0 FreeSans 480 0 0 0 n1
flabel metal1 230 -216 261 104 0 FreeSans 480 0 0 0 n0
flabel metal1 -4166 845 267 874 0 FreeSans 480 0 0 0 drain
port 0 nsew
flabel locali -4356 -547 -4322 -513 0 FreeSans 480 0 0 0 vss
port 6 nsew
flabel metal1 523 1005 573 1055 0 FreeSans 480 0 0 0 d_0_
port 5 nsew
flabel metal1 -211 1015 -167 1059 0 FreeSans 480 0 0 0 d_1_
port 4 nsew
flabel metal1 -730 1013 -684 1059 0 FreeSans 480 0 0 0 d_2_
port 3 nsew
flabel metal1 -1818 1010 -1774 1054 0 FreeSans 480 0 0 0 d_3_
port 2 nsew
flabel metal1 -3060 1009 -3014 1055 0 FreeSans 480 0 0 0 d_4_
port 1 nsew
<< end >>
