magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 275 117 459 163
rect 1 -19 459 117
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 91
rect 151 7 181 91
rect 223 7 253 91
rect 351 7 381 137
<< scpmoshvt >>
rect 79 260 109 344
rect 163 260 193 344
rect 256 260 286 344
rect 351 257 381 457
<< ndiff >>
rect 301 91 351 137
rect 27 53 79 91
rect 27 19 35 53
rect 69 19 79 53
rect 27 7 79 19
rect 109 7 151 91
rect 181 7 223 91
rect 253 69 351 91
rect 253 35 307 69
rect 341 35 351 69
rect 253 7 351 35
rect 381 79 433 137
rect 381 45 391 79
rect 425 45 433 79
rect 381 7 433 45
<< pdiff >>
rect 299 445 351 457
rect 299 411 307 445
rect 341 411 351 445
rect 299 398 351 411
rect 301 344 351 398
rect 27 306 79 344
rect 27 272 35 306
rect 69 272 79 306
rect 27 260 79 272
rect 109 336 163 344
rect 109 302 119 336
rect 153 302 163 336
rect 109 260 163 302
rect 193 317 256 344
rect 193 283 212 317
rect 246 283 256 317
rect 193 260 256 283
rect 286 260 351 344
rect 301 257 351 260
rect 381 431 433 457
rect 381 397 391 431
rect 425 397 433 431
rect 381 363 433 397
rect 381 329 391 363
rect 425 329 433 363
rect 381 257 433 329
<< ndiffc >>
rect 35 19 69 53
rect 307 35 341 69
rect 391 45 425 79
<< pdiffc >>
rect 307 411 341 445
rect 35 272 69 306
rect 119 302 153 336
rect 212 283 246 317
rect 391 397 425 431
rect 391 329 425 363
<< poly >>
rect 351 457 381 483
rect 163 436 217 452
rect 163 402 173 436
rect 207 402 217 436
rect 163 386 217 402
rect 79 344 109 385
rect 163 344 193 386
rect 256 344 286 370
rect 79 211 109 260
rect 163 242 193 260
rect 25 163 109 211
rect 25 129 35 163
rect 69 129 109 163
rect 25 106 109 129
rect 79 91 109 106
rect 151 217 193 242
rect 256 219 286 260
rect 351 225 381 257
rect 151 91 181 217
rect 235 203 289 219
rect 235 186 245 203
rect 223 169 245 186
rect 279 169 289 203
rect 223 153 289 169
rect 331 209 385 225
rect 331 175 341 209
rect 375 175 385 209
rect 331 159 385 175
rect 223 130 265 153
rect 351 137 381 159
rect 223 106 260 130
rect 223 91 253 106
rect 79 -19 109 7
rect 151 -19 181 7
rect 223 -19 253 7
rect 351 -19 381 7
<< polycont >>
rect 173 402 207 436
rect 35 129 69 163
rect 245 169 279 203
rect 341 175 375 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 17 376 138 487
rect 173 436 269 453
rect 207 402 269 436
rect 173 385 269 402
rect 303 445 354 487
rect 303 411 307 445
rect 341 411 354 445
rect 303 378 354 411
rect 388 431 443 453
rect 388 397 391 431
rect 425 397 443 431
rect 17 356 140 376
rect 103 351 140 356
rect 388 363 443 397
rect 103 336 169 351
rect 17 306 69 322
rect 17 272 35 306
rect 103 302 119 336
rect 153 302 169 336
rect 203 317 354 337
rect 203 287 212 317
rect 200 283 212 287
rect 246 283 354 317
rect 388 329 391 363
rect 425 329 443 363
rect 388 313 443 329
rect 200 280 354 283
rect 197 278 354 280
rect 196 275 375 278
rect 192 272 375 275
rect 17 232 69 272
rect 188 270 375 272
rect 183 268 375 270
rect 169 262 375 268
rect 165 256 375 262
rect 161 250 375 256
rect 155 245 375 250
rect 148 238 375 245
rect 142 237 375 238
rect 142 236 220 237
rect 142 234 215 236
rect 142 233 212 234
rect 142 232 209 233
rect 17 231 209 232
rect 17 229 207 231
rect 17 228 205 229
rect 17 226 203 228
rect 17 224 202 226
rect 17 223 201 224
rect 17 220 199 223
rect 17 217 198 220
rect 17 212 196 217
rect 17 198 195 212
rect 329 209 375 237
rect 17 163 127 164
rect 17 129 35 163
rect 69 129 127 163
rect 17 87 127 129
rect 161 53 195 198
rect 17 19 35 53
rect 69 19 195 53
rect 229 169 245 203
rect 279 169 295 203
rect 229 118 295 169
rect 329 175 341 209
rect 329 158 375 175
rect 229 21 273 118
rect 409 107 443 313
rect 307 69 357 85
rect 341 35 357 69
rect 307 -23 357 35
rect 391 79 443 107
rect 425 45 443 79
rect 391 11 443 45
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 and3_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 397 385 431 419 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 397 45 431 79 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 213 385 247 419 0 FreeSans 400 0 0 0 B
port 9 nsew
flabel locali s 29 113 63 147 0 FreeSans 400 0 0 0 A
port 10 nsew
flabel locali s 235 113 269 147 0 FreeSans 400 0 0 0 C
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 -1.000 11.500 -1.000 
<< end >>
