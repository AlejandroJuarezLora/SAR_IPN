magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -29 101 29 107
rect -29 67 -17 101
rect -29 61 29 67
<< pwell >>
rect -114 -197 114 55
<< nmos >>
rect -30 -171 30 29
<< ndiff >>
rect -88 14 -30 29
rect -88 -20 -76 14
rect -42 -20 -30 14
rect -88 -54 -30 -20
rect -88 -88 -76 -54
rect -42 -88 -30 -54
rect -88 -122 -30 -88
rect -88 -156 -76 -122
rect -42 -156 -30 -122
rect -88 -171 -30 -156
rect 30 14 88 29
rect 30 -20 42 14
rect 76 -20 88 14
rect 30 -54 88 -20
rect 30 -88 42 -54
rect 76 -88 88 -54
rect 30 -122 88 -88
rect 30 -156 42 -122
rect 76 -156 88 -122
rect 30 -171 88 -156
<< ndiffc >>
rect -76 -20 -42 14
rect -76 -88 -42 -54
rect -76 -156 -42 -122
rect 42 -20 76 14
rect 42 -88 76 -54
rect 42 -156 76 -122
<< poly >>
rect -33 101 33 117
rect -33 67 -17 101
rect 17 67 33 101
rect -33 51 33 67
rect -30 29 30 51
rect -30 -197 30 -171
<< polycont >>
rect -17 67 17 101
<< locali >>
rect -33 67 -17 101
rect 17 67 33 101
rect -76 14 -42 33
rect -76 -54 -42 -52
rect -76 -90 -42 -88
rect -76 -175 -42 -156
rect 42 14 76 33
rect 42 -54 76 -52
rect 42 -90 76 -88
rect 42 -175 76 -156
<< viali >>
rect -17 67 17 101
rect -76 -20 -42 -18
rect -76 -52 -42 -20
rect -76 -122 -42 -90
rect -76 -124 -42 -122
rect 42 -20 76 -18
rect 42 -52 76 -20
rect 42 -122 76 -90
rect 42 -124 76 -122
<< metal1 >>
rect -29 101 29 107
rect -29 67 -17 101
rect 17 67 29 101
rect -29 61 29 67
rect -82 -18 -36 29
rect -82 -52 -76 -18
rect -42 -52 -36 -18
rect -82 -90 -36 -52
rect -82 -124 -76 -90
rect -42 -124 -36 -90
rect -82 -171 -36 -124
rect 36 -18 82 29
rect 36 -52 42 -18
rect 76 -52 82 -18
rect 36 -90 82 -52
rect 36 -124 42 -90
rect 76 -124 82 -90
rect 36 -171 82 -124
<< end >>
