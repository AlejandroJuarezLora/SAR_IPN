magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 229 145 419 163
rect 33 -19 419 145
rect 33 -23 63 -19
rect 29 -57 63 -23
<< scnmos >>
rect 115 35 145 119
rect 199 35 229 119
rect 307 7 337 137
<< scpmoshvt >>
rect 115 331 145 415
rect 199 331 229 415
rect 307 257 337 457
<< ndiff >>
rect 255 119 307 137
rect 59 81 115 119
rect 59 47 71 81
rect 105 47 115 81
rect 59 35 115 47
rect 145 35 199 119
rect 229 53 307 119
rect 229 35 263 53
rect 255 19 263 35
rect 297 19 307 53
rect 255 7 307 19
rect 337 53 393 137
rect 337 19 347 53
rect 381 19 393 53
rect 337 7 393 19
<< pdiff >>
rect 255 445 307 457
rect 255 415 263 445
rect 59 403 115 415
rect 59 369 71 403
rect 105 369 115 403
rect 59 331 115 369
rect 145 403 199 415
rect 145 369 155 403
rect 189 369 199 403
rect 145 331 199 369
rect 229 411 263 415
rect 297 411 307 445
rect 229 377 307 411
rect 229 343 263 377
rect 297 343 307 377
rect 229 331 307 343
rect 245 257 307 331
rect 337 445 432 457
rect 337 411 367 445
rect 401 411 432 445
rect 337 377 432 411
rect 337 343 367 377
rect 401 343 432 377
rect 337 257 432 343
<< ndiffc >>
rect 71 47 105 81
rect 263 19 297 53
rect 347 19 381 53
<< pdiffc >>
rect 71 369 105 403
rect 155 369 189 403
rect 263 411 297 445
rect 263 343 297 377
rect 367 411 401 445
rect 367 343 401 377
<< poly >>
rect 307 457 337 483
rect 115 415 145 441
rect 199 415 229 441
rect 115 225 145 331
rect 58 209 145 225
rect 58 175 74 209
rect 108 175 145 209
rect 58 159 145 175
rect 115 119 145 159
rect 199 225 229 331
rect 307 225 337 257
rect 199 209 265 225
rect 199 175 215 209
rect 249 175 265 209
rect 199 159 265 175
rect 307 209 373 225
rect 307 175 323 209
rect 357 175 373 209
rect 307 159 373 175
rect 199 119 229 159
rect 307 137 337 159
rect 115 9 145 35
rect 199 9 229 35
rect 307 -19 337 7
<< polycont >>
rect 74 175 108 209
rect 215 175 249 209
rect 323 175 357 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 57 403 113 487
rect 247 445 313 487
rect 57 369 71 403
rect 105 369 113 403
rect 57 353 113 369
rect 147 403 207 419
rect 147 369 155 403
rect 189 369 207 403
rect 147 309 207 369
rect 247 411 263 445
rect 297 411 313 445
rect 247 377 313 411
rect 247 343 263 377
rect 297 343 313 377
rect 351 445 443 453
rect 351 411 367 445
rect 401 411 443 445
rect 351 377 443 411
rect 351 343 367 377
rect 401 343 443 377
rect 20 225 73 297
rect 147 275 335 309
rect 301 225 335 275
rect 20 209 155 225
rect 20 175 74 209
rect 108 175 155 209
rect 199 209 267 225
rect 199 175 215 209
rect 249 175 267 209
rect 301 209 359 225
rect 301 175 323 209
rect 357 175 359 209
rect 301 159 359 175
rect 301 141 335 159
rect 57 103 335 141
rect 57 81 123 103
rect 57 47 71 81
rect 105 47 123 81
rect 393 69 443 343
rect 57 31 123 47
rect 247 53 297 69
rect 247 19 263 53
rect 247 -23 297 19
rect 331 53 443 69
rect 331 19 347 53
rect 381 19 443 53
rect 331 11 443 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 and2_1
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 397 113 431 147 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 397 45 431 79 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 397 181 431 215 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 397 249 431 283 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 397 317 431 351 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 397 385 431 419 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 213 181 247 215 0 FreeSans 250 0 0 0 B
port 9 nsew
flabel locali s 121 181 155 215 0 FreeSans 250 0 0 0 A
port 8 nsew
flabel locali s 29 181 63 215 0 FreeSans 250 0 0 0 A
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 12.600 11.500 12.600 
<< end >>
