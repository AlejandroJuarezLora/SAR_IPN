magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 406 542
<< pwell >>
rect 1 -19 367 143
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 289 117
<< scpmoshvt >>
rect 79 283 289 457
<< ndiff >>
rect 27 79 79 117
rect 27 45 35 79
rect 69 45 79 79
rect 27 7 79 45
rect 289 79 341 117
rect 289 45 299 79
rect 333 45 341 79
rect 289 7 341 45
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 343 79 411
rect 27 309 35 343
rect 69 309 79 343
rect 27 283 79 309
rect 289 445 341 457
rect 289 411 299 445
rect 333 411 341 445
rect 289 343 341 411
rect 289 309 299 343
rect 333 309 341 343
rect 289 283 341 309
<< ndiffc >>
rect 35 45 69 79
rect 299 45 333 79
<< pdiffc >>
rect 35 411 69 445
rect 35 309 69 343
rect 299 411 333 445
rect 299 309 333 343
<< poly >>
rect 79 457 289 483
rect 79 257 289 283
rect 79 251 163 257
rect 21 235 163 251
rect 21 201 37 235
rect 71 201 163 235
rect 21 185 163 201
rect 205 199 347 215
rect 205 165 297 199
rect 331 165 347 199
rect 205 149 347 165
rect 205 143 289 149
rect 79 117 289 143
rect 79 -19 289 7
<< polycont >>
rect 37 201 71 235
rect 297 165 331 199
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 17 445 351 487
rect 17 411 35 445
rect 69 411 299 445
rect 333 411 351 445
rect 17 343 351 411
rect 17 309 35 343
rect 69 309 299 343
rect 333 309 351 343
rect 17 269 351 309
rect 17 201 37 235
rect 71 201 167 235
rect 17 131 167 201
rect 201 199 351 269
rect 201 165 297 199
rect 331 165 351 199
rect 17 79 351 131
rect 17 45 35 79
rect 69 45 299 79
rect 333 45 351 79
rect 17 -23 351 45
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
<< metal1 >>
rect 0 521 368 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 0 456 368 487
rect 0 -23 368 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
rect 0 -88 368 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 decap_4
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 368 504
string path 0.000 -1.000 9.200 -1.000 
<< end >>
