magic
tech sky130B
magscale 1 2
timestamp 1696623266
<< error_p >>
rect -442 141 -384 147
rect -324 141 -266 147
rect -206 141 -148 147
rect -88 141 -30 147
rect 30 141 88 147
rect 148 141 206 147
rect 266 141 324 147
rect 384 141 442 147
rect -442 107 -430 141
rect -324 107 -312 141
rect -206 107 -194 141
rect -88 107 -76 141
rect 30 107 42 141
rect 148 107 160 141
rect 266 107 278 141
rect 384 107 396 141
rect -442 101 -384 107
rect -324 101 -266 107
rect -206 101 -148 107
rect -88 101 -30 107
rect 30 101 88 107
rect 148 101 206 107
rect 266 101 324 107
rect 384 101 442 107
<< pwell >>
rect -639 -279 639 279
<< nmoslvt >>
rect -443 -131 -383 69
rect -325 -131 -265 69
rect -207 -131 -147 69
rect -89 -131 -29 69
rect 29 -131 89 69
rect 147 -131 207 69
rect 265 -131 325 69
rect 383 -131 443 69
<< ndiff >>
rect -501 39 -443 69
rect -501 -101 -489 39
rect -455 -101 -443 39
rect -501 -131 -443 -101
rect -383 39 -325 69
rect -383 -101 -371 39
rect -337 -101 -325 39
rect -383 -131 -325 -101
rect -265 39 -207 69
rect -265 -101 -253 39
rect -219 -101 -207 39
rect -265 -131 -207 -101
rect -147 39 -89 69
rect -147 -101 -135 39
rect -101 -101 -89 39
rect -147 -131 -89 -101
rect -29 39 29 69
rect -29 -101 -17 39
rect 17 -101 29 39
rect -29 -131 29 -101
rect 89 39 147 69
rect 89 -101 101 39
rect 135 -101 147 39
rect 89 -131 147 -101
rect 207 39 265 69
rect 207 -101 219 39
rect 253 -101 265 39
rect 207 -131 265 -101
rect 325 39 383 69
rect 325 -101 337 39
rect 371 -101 383 39
rect 325 -131 383 -101
rect 443 39 501 69
rect 443 -101 455 39
rect 489 -101 501 39
rect 443 -131 501 -101
<< ndiffc >>
rect -489 -101 -455 39
rect -371 -101 -337 39
rect -253 -101 -219 39
rect -135 -101 -101 39
rect -17 -101 17 39
rect 101 -101 135 39
rect 219 -101 253 39
rect 337 -101 371 39
rect 455 -101 489 39
<< psubdiff >>
rect -603 209 603 243
rect -603 -209 -569 209
rect 569 -209 603 209
rect -603 -243 -406 -209
rect 406 -243 603 -209
<< psubdiffcont >>
rect -406 -243 406 -209
<< poly >>
rect -446 141 -380 157
rect -446 107 -430 141
rect -396 107 -380 141
rect -446 91 -380 107
rect -328 141 -262 157
rect -328 107 -312 141
rect -278 107 -262 141
rect -328 91 -262 107
rect -210 141 -144 157
rect -210 107 -194 141
rect -160 107 -144 141
rect -210 91 -144 107
rect -92 141 -26 157
rect -92 107 -76 141
rect -42 107 -26 141
rect -92 91 -26 107
rect 26 141 92 157
rect 26 107 42 141
rect 76 107 92 141
rect 26 91 92 107
rect 144 141 210 157
rect 144 107 160 141
rect 194 107 210 141
rect 144 91 210 107
rect 262 141 328 157
rect 262 107 278 141
rect 312 107 328 141
rect 262 91 328 107
rect 380 141 446 157
rect 380 107 396 141
rect 430 107 446 141
rect 380 91 446 107
rect -443 69 -383 91
rect -325 69 -265 91
rect -207 69 -147 91
rect -89 69 -29 91
rect 29 69 89 91
rect 147 69 207 91
rect 265 69 325 91
rect 383 69 443 91
rect -443 -157 -383 -131
rect -325 -157 -265 -131
rect -207 -157 -147 -131
rect -89 -157 -29 -131
rect 29 -157 89 -131
rect 147 -157 207 -131
rect 265 -157 325 -131
rect 383 -157 443 -131
<< polycont >>
rect -430 107 -396 141
rect -312 107 -278 141
rect -194 107 -160 141
rect -76 107 -42 141
rect 42 107 76 141
rect 160 107 194 141
rect 278 107 312 141
rect 396 107 430 141
<< locali >>
rect -446 107 -430 141
rect -396 107 -380 141
rect -328 107 -312 141
rect -278 107 -262 141
rect -210 107 -194 141
rect -160 107 -144 141
rect -92 107 -76 141
rect -42 107 -26 141
rect 26 107 42 141
rect 76 107 92 141
rect 144 107 160 141
rect 194 107 210 141
rect 262 107 278 141
rect 312 107 328 141
rect 380 107 396 141
rect 430 107 446 141
rect -489 39 -455 55
rect -489 -117 -455 -101
rect -371 39 -337 55
rect -371 -117 -337 -101
rect -253 39 -219 55
rect -253 -117 -219 -101
rect -135 39 -101 55
rect -135 -117 -101 -101
rect -17 39 17 55
rect -17 -117 17 -101
rect 101 39 135 55
rect 101 -117 135 -101
rect 219 39 253 55
rect 219 -117 253 -101
rect 337 39 371 55
rect 337 -117 371 -101
rect 455 39 489 55
rect 455 -117 489 -101
rect -422 -243 -406 -209
rect 406 -243 422 -209
<< viali >>
rect -430 107 -396 141
rect -312 107 -278 141
rect -194 107 -160 141
rect -76 107 -42 141
rect 42 107 76 141
rect 160 107 194 141
rect 278 107 312 141
rect 396 107 430 141
rect -489 -101 -455 39
rect -371 -84 -337 22
rect -253 -101 -219 39
rect -135 -84 -101 22
rect -17 -101 17 39
rect 101 -84 135 22
rect 219 -101 253 39
rect 337 -84 371 22
rect 455 -101 489 39
<< metal1 >>
rect -442 141 -384 147
rect -442 107 -430 141
rect -396 107 -384 141
rect -442 101 -384 107
rect -324 141 -266 147
rect -324 107 -312 141
rect -278 107 -266 141
rect -324 101 -266 107
rect -206 141 -148 147
rect -206 107 -194 141
rect -160 107 -148 141
rect -206 101 -148 107
rect -88 141 -30 147
rect -88 107 -76 141
rect -42 107 -30 141
rect -88 101 -30 107
rect 30 141 88 147
rect 30 107 42 141
rect 76 107 88 141
rect 30 101 88 107
rect 148 141 206 147
rect 148 107 160 141
rect 194 107 206 141
rect 148 101 206 107
rect 266 141 324 147
rect 266 107 278 141
rect 312 107 324 141
rect 266 101 324 107
rect 384 141 442 147
rect 384 107 396 141
rect 430 107 442 141
rect 384 101 442 107
rect -495 39 -449 51
rect -495 -101 -489 39
rect -455 -101 -449 39
rect -259 39 -213 51
rect -377 22 -331 34
rect -377 -84 -371 22
rect -337 -84 -331 22
rect -377 -96 -331 -84
rect -495 -113 -449 -101
rect -259 -101 -253 39
rect -219 -101 -213 39
rect -23 39 23 51
rect -141 22 -95 34
rect -141 -84 -135 22
rect -101 -84 -95 22
rect -141 -96 -95 -84
rect -259 -113 -213 -101
rect -23 -101 -17 39
rect 17 -101 23 39
rect 213 39 259 51
rect 95 22 141 34
rect 95 -84 101 22
rect 135 -84 141 22
rect 95 -96 141 -84
rect -23 -113 23 -101
rect 213 -101 219 39
rect 253 -101 259 39
rect 449 39 495 51
rect 331 22 377 34
rect 331 -84 337 22
rect 371 -84 377 22
rect 331 -96 377 -84
rect 213 -113 259 -101
rect 449 -101 455 39
rect 489 -101 495 39
rect 449 -113 495 -101
<< properties >>
string FIXED_BBOX -586 -226 586 226
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.3 m 1 nf 8 diffcov 80 polycov 80 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
