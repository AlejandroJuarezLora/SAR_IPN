* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt M2_1 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
.ends

.subckt M2_inv a_n40_n201# a_40_n104# w_n236_n324# a_n98_n104#
X0 a_40_n104# a_n40_n201# a_n98_n104# w_n236_n324# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
.ends

.subckt M1_inv a_40_n171# a_n40_n197# a_n98_n171# VSUBS
X0 a_40_n171# a_n40_n197# a_n98_n171# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
.ends

.subckt inv_lvt M2_inv_0/a_n98_n104# M2_inv_0/w_n236_n324# M1_inv_0/a_n98_n171# m1_170_505#
+ m2_289_257# VSUBS
XM2_inv_0 m1_170_505# m2_289_257# M2_inv_0/w_n236_n324# M2_inv_0/a_n98_n104# M2_inv
XM1_inv_0 m2_289_257# m1_170_505# M1_inv_0/a_n98_n171# VSUBS M1_inv
.ends

.subckt M1_2 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
.ends

.subckt latch Qn S R Q vdd vss
XM2_1_0 vss m1_1673_493# Q vss M2_1
Xinv_lvt_0 vdd vdd vss R m1_1673_493# vss inv_lvt
Xinv_lvt_1 vdd vdd vss S m1_458_623# vss inv_lvt
Xinv_lvt_2 vdd vdd vss Qn Q vss inv_lvt
Xinv_lvt_3 vdd vdd vss Q Qn vss inv_lvt
XM1_2_0 Qn m1_458_623# vss vss M1_2
.ends

.subckt inv2 w_0_269# a_67_305# a_59_207# a_149_55# a_67_55# VSUBS
X0 a_67_55# a_59_207# a_149_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_149_55# a_59_207# a_67_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_67_305# a_59_207# a_149_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_149_55# a_59_207# a_67_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt decap_8 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=2.89
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=2.89
.ends

.subckt M1_3 a_207_n176# a_n29_n176# a_26_55# a_n328_55# a_89_n176# a_n446_55# a_n564_55#
+ a_n210_55# a_n501_n176# a_561_n176# a_n383_n176# a_498_55# a_144_55# a_443_n176#
+ a_n265_n176# a_262_55# a_380_55# a_n619_n176# a_n92_55# w_n757_n324# a_325_n176#
+ a_n147_n176#
X0 a_n383_n176# a_n446_55# a_n501_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n29_n176# a_n92_55# a_n147_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_325_n176# a_262_55# a_207_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_561_n176# a_498_55# a_443_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X4 a_n265_n176# a_n328_55# a_n383_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_89_n176# a_26_55# a_n29_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_207_n176# a_144_55# a_89_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_n501_n176# a_n564_55# a_n619_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X8 a_n147_n176# a_n210_55# a_n265_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_443_n176# a_380_55# a_325_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt M2_2 a_26_51# a_89_n171# a_n328_51# a_n446_51# a_n564_51# a_n501_n171# a_n210_51#
+ a_561_n171# a_n383_n171# a_498_51# a_443_n171# a_144_51# a_n265_n171# a_262_51#
+ a_n619_n171# a_380_51# a_n92_51# a_n721_n283# a_325_n171# a_n147_n171# a_207_n171#
+ a_n29_n171#
X0 a_89_n171# a_26_51# a_n29_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_207_n171# a_144_51# a_89_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n147_n171# a_n210_51# a_n265_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_n501_n171# a_n564_51# a_n619_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X4 a_443_n171# a_380_51# a_325_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n383_n171# a_n446_51# a_n501_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_n29_n171# a_n92_51# a_n147_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_325_n171# a_262_51# a_207_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_561_n171# a_498_51# a_443_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X9 a_n265_n171# a_n328_51# a_n383_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt inv_4 w_0_269# a_59_207# a_75_55# a_75_305# a_157_55# VSUBS
X0 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt decap_3 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=0.59
.ends

.subckt sw_top out en m2_1158_361# m2_990_200# inv_4_1/w_0_269# vdd in vss
Xdecap_8_0 vss vdd inv_4_1/w_0_269# vss decap_8
XM1_3_0 out out m2_1158_361# m2_1158_361# in m2_1158_361# m2_1158_361# m2_1158_361#
+ out in in m2_1158_361# m2_1158_361# out out m2_1158_361# m2_1158_361# in m2_1158_361#
+ vdd in in M1_3
XM2_2_0 m2_990_200# in m2_990_200# m2_990_200# m2_990_200# out m2_990_200# in in m2_990_200#
+ out m2_990_200# out m2_990_200# in m2_990_200# m2_990_200# vss in in out out M2_2
Xinv_4_0 inv_4_1/w_0_269# m2_1158_361# vss vdd m2_990_200# vss inv_4
Xinv_4_1 inv_4_1/w_0_269# en vss vdd m2_1158_361# vss inv_4
Xdecap_3_0 vss vdd inv_4_1/w_0_269# vss decap_3
.ends

.subckt C7 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt DUMMY m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C6 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt CDUM m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C4 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C2 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C5 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C3 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C1 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C0_1 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt carray n5 n7 n2 n3 n4 n1 n0 ndum top n6
XC7_121 n7 top C7
XC7_110 n7 top C7
XDUMMY_80 via23_4_712/m2_1_40# top DUMMY
XC6_20 n6 top C6
XC6_53 n6 top C6
XC6_31 n6 top C6
XC6_42 n6 top C6
XC7_122 n7 top C7
XC7_100 n7 top C7
XC7_111 n7 top C7
XDUMMY_81 via23_4_709/m2_1_40# top DUMMY
XDUMMY_70 via23_4_642/m2_1_40# top DUMMY
XC6_21 n6 top C6
XC6_10 n6 top C6
XC6_54 n6 top C6
XC6_32 n6 top C6
XC6_43 n6 top C6
XC6_0 n6 top C6
XC7_123 n7 top C7
XC7_101 n7 top C7
XC7_112 n7 top C7
XDUMMY_71 via23_4_641/m2_1_40# top DUMMY
XDUMMY_82 via23_4_439/m2_1_40# top DUMMY
XDUMMY_60 via23_4_448/m2_1_40# top DUMMY
XC6_44 n6 top C6
XC6_22 n6 top C6
XC6_55 n6 top C6
XC6_11 n6 top C6
XC6_33 n6 top C6
XC6_1 n6 top C6
XC7_124 n7 top C7
XC7_102 n7 top C7
XC7_113 n7 top C7
XDUMMY_72 via23_4_676/m2_1_40# top DUMMY
XDUMMY_83 via23_4_675/m2_1_40# top DUMMY
XDUMMY_61 via23_4_588/m2_1_40# top DUMMY
XDUMMY_50 via23_4_429/m2_1_40# top DUMMY
XC6_56 n6 top C6
XC6_12 n6 top C6
XC6_45 n6 top C6
XC6_23 n6 top C6
XC6_34 n6 top C6
XC6_2 n6 top C6
XCDUM_0 ndum top CDUM
XC7_103 n7 top C7
XC7_125 n7 top C7
XC7_114 n7 top C7
XDUMMY_73 via23_4_677/m2_1_40# top DUMMY
XDUMMY_62 via23_4_589/m2_1_40# top DUMMY
XDUMMY_40 via23_4_326/m2_1_40# top DUMMY
XDUMMY_51 via23_4_414/m2_1_40# top DUMMY
XC6_57 n6 top C6
XC6_24 n6 top C6
XC6_46 n6 top C6
XC6_13 n6 top C6
XC6_35 n6 top C6
XDUMMY_0 via23_4_3/m2_1_40# top DUMMY
XC6_3 n6 top C6
XC4_0 n4 top C4
XC7_104 n7 top C7
XC7_115 n7 top C7
XC7_126 n7 top C7
XDUMMY_74 via23_4_678/m2_1_40# top DUMMY
XDUMMY_63 via23_4_590/m2_1_40# top DUMMY
XDUMMY_30 via23_4_251/m2_1_40# top DUMMY
XDUMMY_52 via23_4_381/m2_1_40# top DUMMY
XDUMMY_41 via23_4_89/m2_1_40# top DUMMY
XC6_47 n6 top C6
XC6_14 n6 top C6
XC6_58 n6 top C6
XC6_25 n6 top C6
XC6_36 n6 top C6
XDUMMY_1 via23_4_9/m2_1_40# top DUMMY
XC7_90 n7 top C7
XC6_4 n6 top C6
XC4_1 n4 top C4
XC7_116 n7 top C7
XC7_105 n7 top C7
XC7_127 n7 top C7
XDUMMY_20 via23_4_199/m2_1_40# top DUMMY
XDUMMY_64 via23_4_584/m2_1_40# top DUMMY
XDUMMY_31 via23_4_245/m2_1_40# top DUMMY
XDUMMY_75 via23_4_704/m2_1_40# top DUMMY
XDUMMY_42 via23_4_366/m2_1_40# top DUMMY
XDUMMY_53 via23_4_449/m2_1_40# top DUMMY
XC6_26 n6 top C6
XC6_15 n6 top C6
XC6_59 n6 top C6
XC6_48 n6 top C6
XDUMMY_2 via23_4_1/m2_1_40# top DUMMY
XC6_37 n6 top C6
XC7_91 n7 top C7
XC7_80 n7 top C7
XC6_5 n6 top C6
XC4_2 n4 top C4
XC7_117 n7 top C7
XC7_106 n7 top C7
XDUMMY_76 via23_4_702/m2_1_40# top DUMMY
XDUMMY_65 via23_4_600/m2_1_40# top DUMMY
XDUMMY_32 via23_4_331/m2_1_40# top DUMMY
XDUMMY_21 via23_4_198/m2_1_40# top DUMMY
XDUMMY_43 via23_4_367/m2_1_40# top DUMMY
XDUMMY_54 via23_4_446/m2_1_40# top DUMMY
XDUMMY_10 via23_4_90/m2_1_40# top DUMMY
XC6_27 n6 top C6
XC6_16 n6 top C6
XC6_49 n6 top C6
XC6_38 n6 top C6
XDUMMY_3 via23_4_2/m2_1_40# top DUMMY
XC7_92 n7 top C7
XC7_81 n7 top C7
XC7_70 n7 top C7
XC6_6 n6 top C6
XC4_3 n4 top C4
XC7_118 n7 top C7
XC7_107 n7 top C7
XC2_0 n2 top C2
XDUMMY_66 via23_4_601/m2_1_40# top DUMMY
XDUMMY_33 via23_4_332/m2_1_40# top DUMMY
XDUMMY_22 via23_4_220/m2_1_40# top DUMMY
XDUMMY_77 via23_4_705/m2_1_40# top DUMMY
XDUMMY_44 via23_4_368/m2_1_40# top DUMMY
XDUMMY_55 via23_4_447/m2_1_40# top DUMMY
XDUMMY_11 via23_4_96/m2_1_40# top DUMMY
XC6_28 n6 top C6
XC6_17 n6 top C6
XC6_39 n6 top C6
XDUMMY_4 via23_4_20/m2_1_40# top DUMMY
XC7_60 n7 top C7
XC7_93 n7 top C7
XC7_82 n7 top C7
XC7_71 n7 top C7
XC6_7 n6 top C6
XC4_4 n4 top C4
XC7_119 n7 top C7
XC7_108 n7 top C7
XC2_1 n2 top C2
XDUMMY_78 via23_4_710/m2_1_40# top DUMMY
XDUMMY_67 via23_4_599/m2_1_40# top DUMMY
XDUMMY_34 via23_4_333/m2_1_40# top DUMMY
XDUMMY_23 via23_4_213/m2_1_40# top DUMMY
XDUMMY_45 via23_4_369/m2_1_40# top DUMMY
XDUMMY_56 via23_4_458/m2_1_40# top DUMMY
XDUMMY_12 via23_4_103/m2_1_40# top DUMMY
XC6_18 n6 top C6
XC6_29 n6 top C6
XDUMMY_5 via23_4_21/m2_1_40# top DUMMY
XC7_61 n7 top C7
XC7_94 n7 top C7
XC7_50 n7 top C7
XC7_72 n7 top C7
XC7_83 n7 top C7
XC6_8 n6 top C6
XC4_5 n4 top C4
XC7_109 n7 top C7
XC2_2 n2 top C2
XDUMMY_79 via23_4_711/m2_1_40# top DUMMY
XDUMMY_68 via23_4_598/m2_1_40# top DUMMY
XDUMMY_35 via23_4_347/m2_1_40# top DUMMY
XDUMMY_24 via23_4_229/m2_1_40# top DUMMY
XDUMMY_46 via23_4_378/m2_1_40# top DUMMY
XDUMMY_57 via23_4_455/m2_1_40# top DUMMY
XDUMMY_13 via23_4_91/m2_1_40# top DUMMY
XC6_19 n6 top C6
XDUMMY_6 via23_4_22/m2_1_40# top DUMMY
XC7_62 n7 top C7
XC7_40 n7 top C7
XC7_95 n7 top C7
XC7_51 n7 top C7
XC7_73 n7 top C7
XC7_84 n7 top C7
XC6_9 n6 top C6
XC4_6 n4 top C4
XC2_3 n2 top C2
XDUMMY_36 via23_4_354/m2_1_40# top DUMMY
XDUMMY_25 via23_4_228/m2_1_40# top DUMMY
XDUMMY_14 via23_4_94/m2_1_40# top DUMMY
XDUMMY_69 via23_4_635/m2_1_40# top DUMMY
XDUMMY_47 via23_4_379/m2_1_40# top DUMMY
XDUMMY_58 via23_4_459/m2_1_40# top DUMMY
XDUMMY_7 via23_4_23/m2_1_40# top DUMMY
XC7_41 n7 top C7
XC7_63 n7 top C7
XC7_96 n7 top C7
XC7_52 n7 top C7
XC7_30 n7 top C7
XC7_74 n7 top C7
XC7_85 n7 top C7
XC4_7 n4 top C4
XDUMMY_37 via23_4_345/m2_1_40# top DUMMY
XDUMMY_26 via23_4_230/m2_1_40# top DUMMY
XDUMMY_48 via23_4_380/m2_1_40# top DUMMY
XDUMMY_59 via23_4_460/m2_1_40# top DUMMY
XDUMMY_15 via23_4_117/m2_1_40# top DUMMY
XDUMMY_8 via23_4_87/m2_1_40# top DUMMY
XC7_97 n7 top C7
XC7_42 n7 top C7
XC7_53 n7 top C7
XC7_31 n7 top C7
XC7_86 n7 top C7
XC7_20 n7 top C7
XC7_64 n7 top C7
XC7_75 n7 top C7
XC4_10 n4 top C4
XC4_8 n4 top C4
XDUMMY_38 via23_4_346/m2_1_40# top DUMMY
XDUMMY_27 via23_4_218/m2_1_40# top DUMMY
XDUMMY_16 via23_4_111/m2_1_40# top DUMMY
XDUMMY_49 via23_4_419/m2_1_40# top DUMMY
XDUMMY_9 via23_4_88/m2_1_40# top DUMMY
XC7_98 n7 top C7
XC7_43 n7 top C7
XC7_54 n7 top C7
XC7_32 n7 top C7
XC7_87 n7 top C7
XC7_65 n7 top C7
XC7_10 n7 top C7
XC7_21 n7 top C7
XC7_76 n7 top C7
XC4_11 n4 top C4
XC4_9 n4 top C4
XDUMMY_39 via23_4_334/m2_1_40# top DUMMY
XDUMMY_28 via23_4_249/m2_1_40# top DUMMY
XDUMMY_17 via23_4_128/m2_1_40# top DUMMY
XC7_99 n7 top C7
XC7_33 n7 top C7
XC7_88 n7 top C7
XC7_55 n7 top C7
XC7_44 n7 top C7
XC7_66 n7 top C7
XC7_11 n7 top C7
XC7_77 n7 top C7
XC7_22 n7 top C7
XC4_12 n4 top C4
XDUMMY_29 via23_4_250/m2_1_40# top DUMMY
XDUMMY_18 via23_4_95/m2_1_40# top DUMMY
XC7_45 n7 top C7
XC7_56 n7 top C7
XC7_34 n7 top C7
XC7_89 n7 top C7
XC7_12 n7 top C7
XC7_23 n7 top C7
XC7_78 n7 top C7
XC7_67 n7 top C7
XC4_13 n4 top C4
XDUMMY_19 via23_4_200/m2_1_40# top DUMMY
XC7_46 n7 top C7
XC7_57 n7 top C7
XC7_24 n7 top C7
XC7_35 n7 top C7
XC7_13 n7 top C7
XC7_79 n7 top C7
XC7_68 n7 top C7
XC4_14 n4 top C4
XC7_36 n7 top C7
XC7_58 n7 top C7
XC7_47 n7 top C7
XC7_25 n7 top C7
XC7_14 n7 top C7
XC7_69 n7 top C7
XC4_15 n4 top C4
XC7_0 n7 top C7
XC7_37 n7 top C7
XC7_59 n7 top C7
XC7_26 n7 top C7
XC7_48 n7 top C7
XC7_15 n7 top C7
XC7_1 n7 top C7
XC7_38 n7 top C7
XC7_27 n7 top C7
XC7_49 n7 top C7
XC7_16 n7 top C7
XC7_2 n7 top C7
XC7_39 n7 top C7
XC7_28 n7 top C7
XC7_17 n7 top C7
XC7_3 n7 top C7
XC5_0 n5 top C5
XC7_29 n7 top C7
XC7_18 n7 top C7
XC7_4 n7 top C7
XC5_1 n5 top C5
XC7_19 n7 top C7
XC5_30 n5 top C5
XC7_5 n7 top C7
XC5_2 n5 top C5
XC5_31 n5 top C5
XC5_20 n5 top C5
XC7_6 n7 top C7
XC5_3 n5 top C5
XC3_0 n3 top C3
XC5_10 n5 top C5
XC5_21 n5 top C5
XC7_7 n7 top C7
XC5_4 n5 top C5
XC3_1 n3 top C3
XC5_22 n5 top C5
XC5_11 n5 top C5
XC7_8 n7 top C7
XC5_5 n5 top C5
XC3_2 n3 top C3
XC5_23 n5 top C5
XC7_9 n7 top C7
XC5_12 n5 top C5
XC5_6 n5 top C5
XC3_3 n3 top C3
XC1_0 n1 top C1
XC5_24 n5 top C5
XC5_13 n5 top C5
XC5_7 n5 top C5
XC3_4 n3 top C3
XC1_1 n1 top C1
XC5_25 n5 top C5
XC5_14 n5 top C5
XC5_8 n5 top C5
XC3_5 n3 top C3
XC5_15 n5 top C5
XC5_26 n5 top C5
XC5_9 n5 top C5
XC3_6 n3 top C3
XC5_16 n5 top C5
XC5_27 n5 top C5
XC3_7 n3 top C3
XC0_1_0 n0 top C0_1
XC5_28 n5 top C5
XC5_17 n5 top C5
XC6_60 n6 top C6
XC5_29 n5 top C5
XC5_18 n5 top C5
XC6_61 n6 top C6
XC6_50 n6 top C6
XC5_19 n5 top C5
XC6_51 n6 top C6
XC6_62 n6 top C6
XC6_40 n6 top C6
XC7_120 n7 top C7
XC6_63 n6 top C6
XC6_52 n6 top C6
XC6_30 n6 top C6
XC6_41 n6 top C6
.ends

.subckt DAC enb en_buf ctl1 ctl0 dum ctl3 ctl4 ctl5 ctl6 ctl7 ctl2 sample out vin
+ vdd_uq0 en_buf_uq0 enb_uq0 vss vdd
Xinv2_0 vdd vdd ctl7 carray_0/n7 vss vss inv2
Xinv2_1 vdd vdd ctl6 carray_0/n6 vss vss inv2
Xinv2_2 vdd vdd dum carray_0/ndum vss vss inv2
Xinv2_3 vdd vdd ctl0 carray_0/n0 vss vss inv2
Xinv2_4 vdd vdd ctl1 carray_0/n1 vss vss inv2
Xinv2_5 vdd vdd ctl5 carray_0/n5 vss vss inv2
Xinv2_6 vdd vdd ctl4 carray_0/n4 vss vss inv2
Xinv2_7 vdd vdd ctl2 carray_0/n2 vss vss inv2
Xinv2_8 vdd vdd ctl3 carray_0/n3 vss vss inv2
Xsw_top_0 out sample sw_top_0/m2_1158_361# sw_top_0/m2_990_200# vdd_uq0 vdd_uq0 vin
+ vss sw_top
Xcarray_0 carray_0/n5 carray_0/n7 carray_0/n2 carray_0/n3 carray_0/n4 carray_0/n1
+ carray_0/n0 carray_0/ndum out carray_0/n6 carray
Xsw_top_1 out sample enb_uq0 en_buf_uq0 vdd_uq0 vdd_uq0 vin vss sw_top
Xsw_top_2 out sample enb en_buf vdd_uq0 vdd_uq0 vin vss sw_top
Xsw_top_3 out sample sw_top_3/m2_1158_361# sw_top_3/m2_990_200# vdd_uq0 vdd_uq0 vin
+ vss sw_top
.ends

.subckt decap_3$1 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
.ends

.subckt M1_1 a_30_n109# a_n88_n109# a_n33_n197# VSUBS
X0 a_30_n109# a_n33_n197# a_n88_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt trim_sw d_0 d_1 d_2 d_3 d_4 m1_1462_409# m1_1771_409# m1_136_409# m1_799_409#
+ m1_1226_409# vss
XM1_1_14 vss m1_799_409# d_2 vss M1_1
XM1_1_15 m1_799_409# vss d_2 vss M1_1
XM1_1_0 vss m1_1226_409# d_0 vss M1_1
XM1_1_1 vss m1_1771_409# d_4 vss M1_1
XM1_1_2 m1_1771_409# vss d_4 vss M1_1
XM1_1_3 vss m1_1771_409# d_4 vss M1_1
XM1_1_4 m1_1771_409# vss d_4 vss M1_1
XM1_1_5 m1_1771_409# vss d_4 vss M1_1
XM1_1_6 vss m1_1771_409# d_4 vss M1_1
XM1_1_7 vss m1_1771_409# d_4 vss M1_1
XM1_1_8 m1_1771_409# vss d_4 vss M1_1
XM1_1_9 m1_1462_409# vss d_1 vss M1_1
XM1_1_10 m1_136_409# vss d_3 vss M1_1
XM1_1_11 vss m1_136_409# d_3 vss M1_1
XM1_1_12 m1_136_409# vss d_3 vss M1_1
XM1_1_13 vss m1_136_409# d_3 vss M1_1
.ends

.subckt trim n3 n4 n2 n1 n0 trim_sw_0/d_4 trim_sw_0/d_3 trim_sw_0/d_2 trim_sw_0/d_1
+ trim_sw_0/d_0 VSUBS drain
Xtrim_sw_0 trim_sw_0/d_0 trim_sw_0/d_1 trim_sw_0/d_2 trim_sw_0/d_3 trim_sw_0/d_4 n1
+ n4 n3 n2 n0 VSUBS trim_sw
.ends

.subckt Mdiff a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt M3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Ml1 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Minp a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt M1 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Minn a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Ml4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt M4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Ml2 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt M2 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt Ml3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176#
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt comparator_core vdd vss outp outn clk ip in diff vp vn
XMdiff_0 clk vss diff vss Mdiff
XMdiff_1 clk diff vss vss Mdiff
XM3_0 outp clk w_302_2337# vdd M3
XMl1_0 outp outn in vss Ml1
XMinp_0 vp ip diff vss Minp
XM1_0 in clk w_302_2337# vdd M1
XMinn_0 vn diff in vss Minn
XMl4_0 vdd outn w_302_2337# outp Ml4
XM4_0 vdd clk w_302_2337# ip M4
XMl2_0 outn ip outp vss Ml2
XM2_0 vdd clk w_302_2337# outn M2
XMl3_0 outn outp w_302_2337# vdd Ml3
.ends

.subckt comparator trim_3 trim_2 trim_0 trim_1 trim_4 trimb_4 trimb_1 trimb_0 trimb_2
+ trimb_3 outn outp clk vdd vp vn vss
Xtrim_0 trim_0/n3 trim_0/n4 trim_0/n2 trim_0/n1 trim_0/n0 trim_4 trim_3 trim_2 trim_1
+ trim_0 vss trim_0/drain trim
Xtrim_1 trim_1/n3 trim_1/n4 trim_1/n2 trim_1/n1 trim_1/n0 trimb_4 trimb_3 trimb_2
+ trimb_1 trimb_0 vss trim_1/drain trim
Xcomparator_core_0 vdd vss outp outn clk trim_1/drain trim_0/drain comparator_core_0/diff
+ vp vn comparator_core
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=1.05
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=2.89
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=2.89
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND VPB VNB Q SET_B D CLK
X0 VPWR a_1032_373# a_1602_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1 a_1032_373# a_193_7# a_1056_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR SET_B a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_476_7# a_27_7# a_381_7# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X4 a_1296_7# a_1182_221# a_1224_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_1032_373# a_27_7# a_956_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X6 a_1182_221# a_1032_373# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X7 Q a_1602_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8 a_652_n19# a_476_7# a_796_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_1140_373# a_193_7# a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 a_586_7# a_193_7# a_476_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_381_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_1224_7# a_27_7# a_1032_373# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_1182_221# a_1032_373# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X16 VGND a_1032_373# a_1602_7# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X17 a_956_373# a_476_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 Q a_1602_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X19 a_796_7# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X20 VPWR a_476_7# a_652_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND SET_B a_1296_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X22 VGND a_652_n19# a_586_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X23 a_381_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X24 a_652_n19# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X25 a_562_373# a_27_7# a_476_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 VPWR a_1182_221# a_1140_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_476_7# a_193_7# a_381_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X29 a_1056_7# a_476_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X30 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 VPWR a_652_n19# a_562_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=1.97
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=1.97
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_346_7# A2 a_256_7# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1 a_250_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2 a_93_n19# A1 a_346_7# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X3 a_93_n19# B1 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4 VGND B2 a_584_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 VPWR a_93_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X6 VGND a_93_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X7 a_250_257# B2 a_93_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_256_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X9 a_250_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X10 a_584_7# B1 a_93_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X11 VPWR A2 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X10 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X13 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X14 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X16 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X17 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X19 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X20 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X21 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X22 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X24 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X25 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X27 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X
X0 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_257# B a_39_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VGND a_39_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A a_39_257# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR a_39_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_39_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X6 VPWR A a_121_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_39_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB X A B
X0 a_68_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_150_257# B a_68_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND A a_68_257# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_68_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR A a_150_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 X a_68_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 VGND A2 a_199_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1 a_113_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 a_199_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4 VPWR A1 a_113_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X5 a_113_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR a_505_n19# a_535_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_505_n19# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_76_159# A1 a_218_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_505_n19# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X5 a_439_7# A0 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6 a_218_334# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X7 a_76_159# A0 a_218_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X8 a_535_334# A1 a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X9 VGND a_505_n19# a_439_7# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_218_7# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=4.73
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=4.73
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 A2 X
X0 VGND A2 a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_79_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X2 a_222_53# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X3 a_448_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_544_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X5 a_448_7# a_222_53# a_79_159# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_222_53# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X7 a_79_159# a_222_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X8 a_544_257# A2 a_79_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X9 VGND a_79_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR VPB VNB A X
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X9 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X11 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X16 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X17 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X20 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X22 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X23 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X26 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X28 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X29 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X30 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X33 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB X A3 A2 A1 B1
X0 VPWR A2 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1 a_80_n19# B1 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2 a_209_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 VPWR a_80_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND B1 a_80_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_209_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X6 VGND a_80_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_209_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X8 a_303_7# A2 a_209_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X9 a_80_n19# A1 a_303_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X14 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X15 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X17 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X18 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X20 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X21 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X24 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X26 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X27 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X29 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR A a_184_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_184_257# B a_112_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_30_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X3 VPWR a_30_13# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND a_30_13# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_30_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X6 a_112_257# C a_30_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_30_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB A1 A2 B1 X
X0 a_297_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X2 a_382_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3 VPWR A1 a_382_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4 a_297_7# B1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_297_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.143 ps=1.62 w=0.55 l=0.59
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.226 ps=2.26 w=0.87 l=0.59
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB A B Y
X0 a_109_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_1 VGND VPWR VPB VNB Y A2_N A1_N B2 B1
X0 a_109_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A2_N a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.283 pd=1.52 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_109_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.283 ps=1.52 w=0.65 l=0.15
X3 a_109_7# A2_N a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 a_397_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_481_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B1 a_481_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B2 a_397_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_257# a_109_7# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.34 ps=2.68 w=1 l=0.15
X9 a_109_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A
X0 a_75_172# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR a_75_172# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND a_75_172# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 a_75_172# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VGND A2 a_373_7# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1 a_109_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3 X a_27_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 X a_27_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_27_257# B1 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_27_257# B1 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X9 a_373_7# A1 a_27_257# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR VPB VNB A X
X0 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X25 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X26 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X27 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 B1 Y A1
X0 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 Y A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3 VGND A1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_27_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_4 VGND VPWR VPB VNB B2 Y A2 A1 B1 C1
X0 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X16 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X23 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X30 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X36 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 a_288_7# a_257_159# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X1 X a_79_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_257_159# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VPWR S a_591_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 a_591_329# A0 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND S a_578_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X7 a_257_159# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_79_n19# A1 a_306_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X9 a_578_7# A1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X10 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_79_n19# A0 a_288_7# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X13 a_306_329# a_257_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB X A1 A2 B1 C1
X0 a_79_n19# C1 a_510_7# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X1 a_297_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 a_215_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND A1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_79_n19# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X6 VPWR B1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X7 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_510_7# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X9 a_79_n19# A2 a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB B2 A2 A1 B1 X
X0 a_292_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X1 a_78_159# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_215_7# B2 a_78_159# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 VGND A2 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_215_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_493_257# A2 a_78_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X7 VGND a_78_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_78_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X9 a_78_159# B2 a_292_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND VPB VNB X A1 A2 A3 B2 B1
X0 a_227_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_227_7# B1 a_77_159# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X2 a_539_257# B2 a_77_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3 VGND A2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_77_159# B2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X5 VGND a_77_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_227_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_323_257# A2 a_227_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X8 a_227_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X9 VPWR B1 a_539_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X10 VPWR a_77_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X11 a_77_159# A3 a_323_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 VGND A a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_29_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X2 a_111_257# C a_29_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_29_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_183_257# B a_111_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_29_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A a_183_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VGND C a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB B1 B2 A2 A1 X C1
X0 a_245_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1 VPWR C1 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X2 a_512_257# A2 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
X3 a_149_7# B2 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_240_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A1 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_51_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_51_257# B2 a_245_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X8 a_240_7# B1 a_149_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X9 a_149_7# C1 a_51_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X10 VPWR A1 a_512_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X11 X a_51_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 VPWR VGND VPB VNB X C B A
X0 VGND C a_184_13# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
X1 VPWR a_29_271# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_29_271# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_29_271# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X4 VPWR A a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_184_13# B a_112_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR C a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X7 X a_29_271# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X8 a_112_13# A a_29_271# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND a_29_271# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND VPB VNB X D1 C1 B1 A2 A1
X0 VPWR A1 a_676_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A2 a_512_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X2 a_512_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X4 a_79_n19# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X5 a_512_7# B1 a_409_7# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X6 a_676_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X7 a_306_7# D1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X8 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_409_7# C1 a_306_7# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X10 VPWR C1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X11 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VGND VPWR VPB VNB A2 A1 B1 B2 Y C1
X0 a_27_257# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_301_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X2 a_735_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X3 a_27_257# B1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X5 a_301_257# B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_301_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_257# B2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_301_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y C1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11 Y A1 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_735_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X15 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_383_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X17 Y B1 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_383_7# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB A Y B
X0 Y A a_113_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_113_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR VPB VNB X C B A
X0 a_27_7# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_181_7# B a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5 VGND C a_181_7# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_109_7# A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR VPB VNB A1 A2 B1 B2 Y
X0 Y B2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X1 a_109_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X3 a_27_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X5 VPWR A1 a_307_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X6 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_307_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPWR VGND VPB VNB B C A X
X0 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_109_257# C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X4 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR A a_193_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X8 a_193_257# B a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND C a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X12 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 B2 A2_N A1_N X
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X1 a_226_7# A2_N a_226_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_76_159# a_226_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X3 a_556_7# B2 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_226_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X5 VGND B1 a_556_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_226_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X7 VGND A2_N a_226_7# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_489_373# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VPWR B2 a_489_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_489_373# a_226_7# a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_257# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VPWR A a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X A B
X0 a_145_35# A a_59_35# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1 VPWR B a_59_35# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 X a_59_35# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3 VGND B a_145_35# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_59_35# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5 X a_59_35# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 VGND VPWR VPB VNB X D_N C B A
X0 a_297_257# a_109_53# a_215_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X1 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_215_257# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.165 ps=1.82 w=0.65 l=0.15
X8 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X9 VPWR A a_487_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_487_257# B a_403_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND C a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X13 a_215_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_403_257# C a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X15 VGND A a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X17 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VPWR VGND VPB VNB B1 Y A1 A2 A3
X0 VPWR A3 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR A1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_277_7# A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_277_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X7 a_27_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X9 a_27_7# A2 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A1 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_27_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X14 VGND A3 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 Y B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR VPB VNB A1 A2 Y B2 C1 B1
X0 a_213_83# B2 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y B2 a_295_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 VGND A2 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X4 a_213_83# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_295_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X6 a_493_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X7 a_109_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X9 a_109_7# B1 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctlp[0]
+ ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] cal clk clkc comp en result[0]
+ result[1] result[2] result[3] result[4] result[5] result[6] result[7] rstn sample
+ trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4]
+ valid VPWR VGND
XFILLER_13_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_294_ VPWR VGND VPWR VGND _294_/Y _294_/A sky130_fd_sc_hd__inv_2
X_346_ VPWR VGND VPWR VGND _346_/Q _346_/SET_B _346_/D _297_/B sky130_fd_sc_hd__dfstp_1
X_277_ VPWR VGND VPWR VGND _277_/Y _277_/A sky130_fd_sc_hd__inv_2
XFILLER_5_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_200_ VGND VPWR VPWR VGND _337_/D _193_/Y _197_/X _338_/Q _337_/Q _194_/X sky130_fd_sc_hd__a32o_1
X_329_ VGND VPWR VPWR VGND _331_/CLK _329_/D _346_/SET_B _329_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput20 VGND VPWR VPWR VGND _281_/A ctlp[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput7 VGND VPWR VPWR VGND _271_/Y ctln[1] sky130_fd_sc_hd__clkbuf_2
Xoutput31 VGND VPWR VPWR VGND _285_/A trim[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_293_ VPWR VGND VPWR VGND _294_/A _340_/Q _313_/Q sky130_fd_sc_hd__or2_2
XFILLER_9_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_276_ VGND VPWR VPWR VGND _277_/A _328_/Q _319_/Q sky130_fd_sc_hd__or2_1
X_345_ VPWR VGND VPWR VGND _345_/Q _346_/SET_B _345_/D _297_/B sky130_fd_sc_hd__dfstp_1
X_328_ VGND VPWR VPWR VGND _297_/B _328_/D _346_/SET_B _328_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_259_ VPWR VGND VPWR VGND _258_/S _339_/Q _312_/Q _261_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput21 VGND VPWR VPWR VGND _283_/A ctlp[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput8 VGND VPWR VPWR VGND _273_/Y ctln[2] sky130_fd_sc_hd__clkbuf_2
Xoutput10 VGND VPWR VPWR VGND _277_/Y ctln[4] sky130_fd_sc_hd__clkbuf_2
Xoutput32 VGND VPWR VPWR VGND _288_/A trim[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_292_ VPWR VGND VPWR VGND _292_/Y _292_/A sky130_fd_sc_hd__inv_2
XFILLER_3_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_275_ VPWR VGND VPWR VGND _275_/Y _275_/A sky130_fd_sc_hd__inv_2
X_344_ VPWR VGND VPWR VGND _344_/Q _346_/SET_B _344_/D _297_/B sky130_fd_sc_hd__dfstp_1
XFILLER_5_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_327_ VGND VPWR VPWR VGND _331_/CLK _327_/D _346_/SET_B _327_/Q sky130_fd_sc_hd__dfrtp_1
X_189_ VGND VPWR VPWR VGND _196_/A _190_/A sky130_fd_sc_hd__clkbuf_2
X_258_ VGND VPWR VPWR VGND _313_/D _306_/X _258_/S _313_/Q sky130_fd_sc_hd__mux2_1
XFILLER_6_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput22 VGND VPWR VPWR VGND _315_/Q result[0] sky130_fd_sc_hd__clkbuf_2
Xoutput33 VGND VPWR VPWR VGND _290_/A trim[2] sky130_fd_sc_hd__clkbuf_2
Xoutput9 VGND VPWR VPWR VGND _275_/Y ctln[3] sky130_fd_sc_hd__clkbuf_2
Xoutput11 VGND VPWR VPWR VGND _279_/Y ctln[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_291_ VPWR VGND VPWR VGND _292_/A _339_/Q _312_/Q sky130_fd_sc_hd__or2_2
XFILLER_12_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_274_ VPWR VGND VPWR VGND _275_/A _327_/Q _318_/Q sky130_fd_sc_hd__or2_2
XFILLER_5_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_343_ VGND VPWR VPWR VGND _343_/CLK _343_/D repeater43/X _343_/Q sky130_fd_sc_hd__dfrtp_1
X_326_ VGND VPWR VPWR VGND _331_/CLK _326_/D repeater43/X _326_/Q sky130_fd_sc_hd__dfrtp_1
X_257_ VGND VPWR VPWR VGND _260_/B _190_/A _254_/Y _258_/S sky130_fd_sc_hd__o21ba_1
XFILLER_9_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_188_ VGND VPWR VPWR VGND _341_/D _255_/B _188_/S _307_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_309_ VGND VPWR VPWR VGND _340_/CLK _309_/D _346_/SET_B _309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput23 VGND VPWR VPWR VGND _316_/Q result[1] sky130_fd_sc_hd__clkbuf_2
Xoutput34 VGND VPWR VPWR VGND _292_/A trim[3] sky130_fd_sc_hd__clkbuf_2
Xoutput12 VGND VPWR VPWR VGND _281_/Y ctln[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_290_ VPWR VGND VPWR VGND _290_/Y _290_/A sky130_fd_sc_hd__inv_2
Xrepeater42 VGND VPWR VPWR VGND repeater43/X _346_/SET_B sky130_fd_sc_hd__buf_8
XFILLER_9_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_12_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_273_ VPWR VGND VPWR VGND _273_/Y _273_/A sky130_fd_sc_hd__inv_2
XFILLER_5_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_342_ VGND VPWR VPWR VGND _343_/CLK _342_/D repeater43/X _342_/Q sky130_fd_sc_hd__dfrtp_4
X_325_ VGND VPWR VPWR VGND _331_/CLK _325_/D repeater43/X _325_/Q sky130_fd_sc_hd__dfrtp_1
X_187_ VGND VPWR VPWR VGND _255_/B _341_/Q sky130_fd_sc_hd__buf_1
X_256_ VGND VPWR VPWR VGND _260_/B _255_/X _191_/B _196_/A _192_/B sky130_fd_sc_hd__a31o_1
X_239_ VPWR VGND VPWR VGND _232_/X _328_/Q _319_/Q _240_/B sky130_fd_sc_hd__a21oi_1
X_308_ VGND VPWR VPWR VGND _308_/X _227_/A _308_/S _192_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput24 VGND VPWR VPWR VGND _317_/Q result[2] sky130_fd_sc_hd__clkbuf_2
Xoutput13 VGND VPWR VPWR VGND _283_/Y ctln[7] sky130_fd_sc_hd__clkbuf_2
Xoutput35 VGND VPWR VPWR VGND _294_/A trim[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrepeater43 VGND VPWR VPWR VGND input4/X repeater43/X sky130_fd_sc_hd__buf_8
XFILLER_8_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_272_ VPWR VGND VPWR VGND _273_/A _326_/Q _317_/Q sky130_fd_sc_hd__or2_2
X_341_ VGND VPWR VPWR VGND _343_/CLK _341_/D repeater43/X _341_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_324_ VGND VPWR VPWR VGND _297_/B _324_/D repeater43/X _324_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_255_ VGND VPWR VPWR VGND _255_/B _298_/C _342_/Q _255_/X sky130_fd_sc_hd__or3_2
X_186_ VGND VPWR VPWR VGND _308_/X _188_/S _172_/A _342_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_238_ VGND VPWR VPWR VGND _242_/A _238_/B _320_/D sky130_fd_sc_hd__nor2_1
X_307_ VGND VPWR VPWR VGND _307_/X _145_/A _308_/S _296_/Y sky130_fd_sc_hd__mux2_1
X_169_ VGND VPWR VPWR VGND _172_/A _169_/B _169_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_8 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput14 VGND VPWR VPWR VGND _269_/A ctlp[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput36 VGND VPWR VPWR VGND _285_/Y trimb[0] sky130_fd_sc_hd__clkbuf_2
Xoutput25 VGND VPWR VPWR VGND _318_/Q result[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_271_ VPWR VGND VPWR VGND _271_/Y _271_/A sky130_fd_sc_hd__inv_2
X_340_ VGND VPWR VPWR VGND _340_/CLK _340_/D _346_/SET_B _340_/Q sky130_fd_sc_hd__dfrtp_1
X_185_ VPWR VGND VPWR VGND _343_/D _185_/A sky130_fd_sc_hd__inv_2
X_323_ VGND VPWR VPWR VGND _343_/CLK _323_/D repeater43/X _323_/Q sky130_fd_sc_hd__dfrtp_1
X_254_ VGND VPWR VPWR VGND _254_/A _254_/B _254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_237_ VPWR VGND VPWR VGND _232_/X _329_/Q _320_/Q _238_/B sky130_fd_sc_hd__a21oi_1
X_168_ VGND VPWR VPWR VGND _169_/B _167_/X _165_/X _167_/X _165_/X sky130_fd_sc_hd__a2bb2oi_1
X_306_ VGND VPWR VPWR VGND _306_/X _286_/B _306_/S _294_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput15 VGND VPWR VPWR VGND _271_/A ctlp[1] sky130_fd_sc_hd__clkbuf_2
Xoutput26 VGND VPWR VPWR VGND _319_/Q result[4] sky130_fd_sc_hd__clkbuf_2
Xoutput37 VGND VPWR VPWR VGND _288_/Y trimb[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_clk VGND VPWR VPWR VGND _297_/B clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_270_ VPWR VGND VPWR VGND _271_/A _325_/Q _316_/Q sky130_fd_sc_hd__or2_2
X_322_ VGND VPWR VPWR VGND _331_/CLK _322_/D repeater43/X _322_/Q sky130_fd_sc_hd__dfrtp_1
X_253_ VPWR VGND VPWR VGND _254_/A _347_/Q sky130_fd_sc_hd__inv_2
XFILLER_13_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_184_ VGND VPWR VPWR VGND _185_/A _150_/C _188_/S _182_/X sky130_fd_sc_hd__mux2_1
X_236_ VGND VPWR VPWR VGND _242_/A _236_/B _321_/D sky130_fd_sc_hd__nor2_1
X_167_ VPWR VGND VPWR VGND _166_/Y _346_/Q _162_/X _167_/X _160_/X sky130_fd_sc_hd__a22o_1
X_305_ VGND VPWR VPWR VGND _305_/X _286_/B _306_/S _254_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_219_ VGND VPWR VPWR VGND _329_/D _216_/X _330_/Q _212_/X _217_/X _329_/Q sky130_fd_sc_hd__a32o_1
XFILLER_19_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput16 VGND VPWR VPWR VGND _273_/A ctlp[2] sky130_fd_sc_hd__clkbuf_2
Xoutput38 VGND VPWR VPWR VGND _290_/Y trimb[2] sky130_fd_sc_hd__clkbuf_2
Xoutput27 VGND VPWR VPWR VGND _320_/Q result[5] sky130_fd_sc_hd__clkbuf_2
XPHY_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk VGND VPWR VPWR VGND clk clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_7_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_5_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk VGND VPWR VPWR VGND _340_/CLK clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_1
X_321_ VGND VPWR VPWR VGND _331_/CLK _321_/D repeater43/X _321_/Q sky130_fd_sc_hd__dfrtp_1
X_252_ VGND VPWR VPWR VGND _251_/X _228_/A _314_/D _297_/A sky130_fd_sc_hd__o21ai_1
X_183_ VGND VPWR VPWR VGND _298_/A _188_/S _181_/X _324_/Q _150_/C _157_/A sky130_fd_sc_hd__o221ai_4
X_235_ VPWR VGND VPWR VGND _232_/X _330_/Q _321_/Q _236_/B sky130_fd_sc_hd__a21oi_1
X_304_ VGND VPWR VPWR VGND _304_/S _227_/A _216_/X _304_/X sky130_fd_sc_hd__mux2_2
X_166_ VPWR VGND VPWR VGND _166_/Y _346_/Q sky130_fd_sc_hd__inv_2
X_218_ VGND VPWR VPWR VGND _330_/D _216_/X _304_/X _331_/Q _217_/X _330_/Q sky130_fd_sc_hd__a32o_1
XFILLER_19_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_149_ VGND VPWR VPWR VGND _149_/A _150_/C sky130_fd_sc_hd__clkbuf_2
Xoutput39 VGND VPWR VPWR VGND _292_/Y trimb[3] sky130_fd_sc_hd__clkbuf_2
Xoutput17 VGND VPWR VPWR VGND _275_/A ctlp[3] sky130_fd_sc_hd__clkbuf_2
Xoutput28 VGND VPWR VPWR VGND _321_/Q result[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_320_ VGND VPWR VPWR VGND _297_/B _320_/D _346_/SET_B _320_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_251_ VGND VPWR VPWR VGND _251_/X _324_/Q _181_/X _172_/A _250_/X sky130_fd_sc_hd__o211a_1
X_182_ VGND VPWR VPWR VGND _182_/X _175_/Y _286_/B _196_/A _181_/X sky130_fd_sc_hd__o211a_1
XFILLER_18_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_234_ VGND VPWR VPWR VGND _242_/A _234_/B _322_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1_0_clk VGND VPWR VPWR VGND _331_/CLK clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_1
X_165_ VGND VPWR VPWR VGND _164_/Y _160_/X _158_/Y _161_/Y _165_/X sky130_fd_sc_hd__o22a_1
X_303_ VPWR VGND VPWR VGND _347_/D _303_/A sky130_fd_sc_hd__inv_2
XFILLER_1_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_217_ VGND VPWR VPWR VGND _217_/A _217_/X sky130_fd_sc_hd__clkbuf_2
X_148_ VPWR VGND VPWR VGND _298_/B _341_/Q sky130_fd_sc_hd__inv_2
Xoutput18 VGND VPWR VPWR VGND _277_/A ctlp[4] sky130_fd_sc_hd__clkbuf_2
Xoutput29 VGND VPWR VPWR VGND _322_/Q result[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_181_ VGND VPWR VPWR VGND _215_/A _181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_250_ VGND VPWR VPWR VGND _190_/A _216_/A _260_/A _284_/A _250_/X sky130_fd_sc_hd__o22a_1
XFILLER_1_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_233_ VPWR VGND VPWR VGND _232_/X _331_/Q _322_/Q _234_/B sky130_fd_sc_hd__a21oi_1
X_302_ VPWR VGND VPWR VGND _303_/A _157_/A _300_/Y _301_/X _147_/A _254_/A sky130_fd_sc_hd__o32a_1
X_164_ VPWR VGND VPWR VGND _164_/Y _164_/A sky130_fd_sc_hd__inv_2
XFILLER_19_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_216_ VGND VPWR VPWR VGND _216_/A _216_/X sky130_fd_sc_hd__clkbuf_2
X_147_ VPWR VGND VPWR VGND _147_/Y _147_/A sky130_fd_sc_hd__inv_2
Xoutput19 VGND VPWR VPWR VGND _279_/A ctlp[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_clk VGND VPWR VPWR VGND _343_/CLK clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_180_ VPWR VGND VPWR VGND _298_/A _298_/B _298_/C _215_/A sky130_fd_sc_hd__or3_1
XFILLER_1_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_232_ VGND VPWR VPWR VGND _232_/A _232_/X sky130_fd_sc_hd__clkbuf_2
X_163_ VGND VPWR VPWR VGND _162_/X _160_/A _158_/Y _345_/Q _164_/A sky130_fd_sc_hd__o22a_1
X_301_ VGND VPWR VPWR VGND _162_/X _254_/A _347_/Q _160_/X _301_/X _299_/X sky130_fd_sc_hd__o221a_1
XFILLER_19_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_146_ VPWR VGND VPWR VGND _147_/A _146_/C _341_/Q _177_/A sky130_fd_sc_hd__and3_2
X_215_ VPWR VGND VPWR VGND _216_/A _215_/A sky130_fd_sc_hd__inv_2
XFILLER_21_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_231_ VPWR VGND VPWR VGND _232_/A _146_/C _255_/B _150_/C _162_/X _298_/A sky130_fd_sc_hd__o2111a_1
X_162_ VGND VPWR VPWR VGND _162_/A _162_/X sky130_fd_sc_hd__clkbuf_2
X_300_ VGND VPWR VPWR VGND _254_/A _160_/X _162_/X _347_/Q _300_/Y _299_/X sky130_fd_sc_hd__a221oi_2
XFILLER_1_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput1 VGND VPWR VPWR VGND input1/X cal sky130_fd_sc_hd__clkbuf_1
XFILLER_10_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_214_ VPWR VGND VPWR VGND _331_/Q _212_/X _181_/X _331_/D _217_/A sky130_fd_sc_hd__a22o_1
X_145_ VGND VPWR VPWR VGND _145_/A _146_/C _304_/S sky130_fd_sc_hd__nand2_1
XFILLER_21_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_7_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_8_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_230_ VGND VPWR VPWR VGND _248_/A _242_/A sky130_fd_sc_hd__clkbuf_2
X_161_ VPWR VGND VPWR VGND _161_/Y _344_/Q sky130_fd_sc_hd__inv_2
XFILLER_1_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput2 VGND VPWR VPWR VGND _162_/A comp sky130_fd_sc_hd__buf_1
XFILLER_10_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_213_ VPWR VGND VPWR VGND _217_/A _304_/X sky130_fd_sc_hd__inv_2
X_144_ VGND VPWR VPWR VGND _304_/S _144_/A sky130_fd_sc_hd__buf_1
XFILLER_21_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_160_ VGND VPWR VPWR VGND _160_/A _160_/X sky130_fd_sc_hd__clkbuf_2
Xinput3 VGND VPWR VPWR VGND en _227_/A sky130_fd_sc_hd__clkbuf_2
X_289_ VPWR VGND VPWR VGND _290_/A _338_/Q _311_/Q sky130_fd_sc_hd__or2_2
XFILLER_19_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_212_ VGND VPWR VPWR VGND _212_/X _304_/X sky130_fd_sc_hd__buf_1
X_143_ VGND VPWR VPWR VGND _144_/A _149_/A _341_/Q _177_/A sky130_fd_sc_hd__and3_1
XFILLER_18_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_130 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_1_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_288_ VPWR VGND VPWR VGND _288_/Y _288_/A sky130_fd_sc_hd__inv_2
Xinput4 VGND VPWR VPWR VGND input4/X rstn sky130_fd_sc_hd__buf_1
X_211_ VPWR VGND VPWR VGND _153_/B _332_/Q _206_/A _332_/D _197_/X sky130_fd_sc_hd__a22o_1
X_142_ VPWR VGND VPWR VGND _149_/A _343_/Q sky130_fd_sc_hd__inv_2
XFILLER_10_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_287_ VPWR VGND VPWR VGND _288_/A _337_/Q _310_/Q sky130_fd_sc_hd__or2_2
XFILLER_19_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_210_ VGND VPWR VPWR VGND _153_/A _207_/C _306_/S _209_/X _333_/D sky130_fd_sc_hd__o22ai_1
X_141_ VPWR VGND VPWR VGND _145_/A _227_/A sky130_fd_sc_hd__inv_2
X_339_ VGND VPWR VPWR VGND _340_/CLK _339_/D _346_/SET_B _339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_14_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_60 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_286_ VGND VPWR VPWR VGND _306_/S _286_/Y _286_/B sky130_fd_sc_hd__nand2_1
X_140_ VPWR VGND VPWR VGND _177_/A _342_/Q sky130_fd_sc_hd__inv_2
X_338_ VGND VPWR VPWR VGND _340_/CLK _338_/D _346_/SET_B _338_/Q sky130_fd_sc_hd__dfrtp_1
X_269_ VPWR VGND VPWR VGND _269_/Y _269_/A sky130_fd_sc_hd__inv_2
XFILLER_7_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_285_ VPWR VGND VPWR VGND _285_/Y _285_/A sky130_fd_sc_hd__inv_2
XFILLER_4_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk VGND VPWR VPWR VGND clkbuf_2_3_0_clk/A clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_268_ VPWR VGND VPWR VGND _269_/A _324_/Q _315_/Q sky130_fd_sc_hd__or2_2
XFILLER_2_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_337_ VGND VPWR VPWR VGND _340_/CLK _337_/D _346_/SET_B _337_/Q sky130_fd_sc_hd__dfrtp_1
X_199_ VGND VPWR VPWR VGND _338_/D _193_/Y _197_/X _339_/Q _338_/Q _194_/X sky130_fd_sc_hd__a32o_1
XFILLER_21_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_40 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_284_ VPWR VGND VPWR VGND _285_/A _284_/A _309_/Q sky130_fd_sc_hd__or2_2
XFILLER_19_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_198_ VGND VPWR VPWR VGND _339_/D _193_/Y _197_/X _340_/Q _339_/Q _194_/X sky130_fd_sc_hd__a32o_1
X_267_ VGND VPWR VPWR VGND _267_/A _267_/B _309_/D sky130_fd_sc_hd__nor2_1
X_336_ VGND VPWR VPWR VGND _340_/CLK _336_/D _346_/SET_B _336_/Q sky130_fd_sc_hd__dfrtp_1
X_319_ VGND VPWR VPWR VGND _297_/B _319_/D _346_/SET_B _319_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0_0_clk VGND VPWR VPWR VGND clkbuf_2_1_0_clk/A clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_283_ VPWR VGND VPWR VGND _283_/Y _283_/A sky130_fd_sc_hd__inv_2
XFILLER_18_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_335_ VGND VPWR VPWR VGND _343_/CLK _335_/D repeater43/X _335_/Q sky130_fd_sc_hd__dfrtp_1
X_197_ VGND VPWR VPWR VGND _260_/A _197_/X sky130_fd_sc_hd__clkbuf_2
X_266_ VPWR VGND VPWR VGND _258_/S _284_/A _309_/Q _267_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_318_ VGND VPWR VPWR VGND _331_/CLK _318_/D repeater43/X _318_/Q sky130_fd_sc_hd__dfrtp_1
X_249_ VPWR VGND VPWR VGND _297_/A _314_/Q sky130_fd_sc_hd__inv_2
XFILLER_20_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_282_ VPWR VGND VPWR VGND _283_/A _331_/Q _322_/Q sky130_fd_sc_hd__or2_2
XFILLER_18_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_334_ VGND VPWR VPWR VGND _343_/CLK _334_/D repeater43/X _334_/Q sky130_fd_sc_hd__dfrtp_1
X_196_ VPWR VGND VPWR VGND _260_/A _196_/A sky130_fd_sc_hd__inv_2
X_265_ VGND VPWR VPWR VGND _267_/A _265_/B _310_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_248_ VGND VPWR VPWR VGND _248_/A _248_/B _315_/D sky130_fd_sc_hd__nor2_1
X_317_ VGND VPWR VPWR VGND _331_/CLK _317_/D repeater43/X _317_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_179_ VGND VPWR VPWR VGND _191_/B _286_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_11_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_281_ VPWR VGND VPWR VGND _281_/Y _281_/A sky130_fd_sc_hd__inv_2
XPHY_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_195_ VPWR VGND VPWR VGND _340_/Q _306_/S _193_/Y _340_/D _194_/X sky130_fd_sc_hd__a22o_1
X_333_ VGND VPWR VPWR VGND _343_/CLK _333_/D repeater43/X _333_/Q sky130_fd_sc_hd__dfrtp_4
X_264_ VPWR VGND VPWR VGND _258_/S _337_/Q _310_/Q _265_/B sky130_fd_sc_hd__a21oi_1
X_316_ VGND VPWR VPWR VGND _331_/CLK _316_/D repeater43/X _316_/Q sky130_fd_sc_hd__dfrtp_1
X_247_ VPWR VGND VPWR VGND _232_/A _324_/Q _315_/Q _248_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_134 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_178_ VPWR VGND VPWR VGND _298_/A _341_/Q _298_/C _191_/B sky130_fd_sc_hd__or3_4
XFILLER_22_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_280_ VGND VPWR VPWR VGND _281_/A _330_/Q _321_/Q sky130_fd_sc_hd__or2_1
XFILLER_14_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_332_ VGND VPWR VPWR VGND _340_/CLK _332_/D repeater43/X _332_/Q sky130_fd_sc_hd__dfrtp_4
X_194_ VGND VPWR VPWR VGND _194_/X _194_/A sky130_fd_sc_hd__buf_1
X_263_ VGND VPWR VPWR VGND _267_/A _263_/B _311_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_246_ VGND VPWR VPWR VGND _248_/A _246_/B _316_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_315_ VGND VPWR VPWR VGND _343_/CLK _315_/D repeater43/X _315_/Q sky130_fd_sc_hd__dfrtp_1
X_177_ VGND VPWR VPWR VGND _177_/A _298_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_229_ VGND VPWR VPWR VGND input1/X _248_/A _226_/X _175_/Y _323_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_331_ VGND VPWR VPWR VGND _331_/CLK _331_/D repeater43/X _331_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_193_ VPWR VGND VPWR VGND _193_/Y _194_/A sky130_fd_sc_hd__inv_2
X_262_ VPWR VGND VPWR VGND _258_/S _338_/Q _311_/Q _263_/B sky130_fd_sc_hd__a21oi_1
XPHY_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_245_ VPWR VGND VPWR VGND _232_/A _325_/Q _316_/Q _246_/B sky130_fd_sc_hd__a21oi_1
XFILLER_14_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_314_ VGND VPWR VPWR VGND _297_/B _314_/D _346_/SET_B _314_/Q sky130_fd_sc_hd__dfrtp_1
X_176_ VGND VPWR VPWR VGND _298_/C _343_/Q sky130_fd_sc_hd__buf_1
XFILLER_22_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_159_ VPWR VGND VPWR VGND _160_/A _162_/A sky130_fd_sc_hd__inv_2
X_228_ VPWR VGND VPWR VGND _248_/A _228_/A sky130_fd_sc_hd__inv_2
XFILLER_17_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_330_ VGND VPWR VPWR VGND _331_/CLK _330_/D repeater43/X _330_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_261_ VGND VPWR VPWR VGND _261_/A _267_/A _312_/D sky130_fd_sc_hd__nor2_1
XPHY_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_192_ VGND VPWR VPWR VGND _194_/A _305_/X _192_/B sky130_fd_sc_hd__or2_1
XPHY_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_175_ VPWR VGND VPWR VGND _175_/Y _323_/Q sky130_fd_sc_hd__inv_2
X_244_ VGND VPWR VPWR VGND _248_/A _244_/B _317_/D sky130_fd_sc_hd__nor2_1
X_313_ VGND VPWR VPWR VGND _340_/CLK _313_/D _346_/SET_B _313_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_158_ VPWR VGND VPWR VGND _158_/Y _345_/Q sky130_fd_sc_hd__inv_2
X_227_ VGND VPWR VPWR VGND _227_/A _228_/A _304_/S sky130_fd_sc_hd__nand2_1
XFILLER_3_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_5_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_260_ VGND VPWR VPWR VGND _260_/B _267_/A _260_/A sky130_fd_sc_hd__nor2_2
XFILLER_2_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_191_ VGND VPWR VPWR VGND _323_/Q _191_/B _192_/B sky130_fd_sc_hd__nor2_1
X_243_ VPWR VGND VPWR VGND _232_/A _326_/Q _317_/Q _244_/B sky130_fd_sc_hd__a21oi_1
X_312_ VGND VPWR VPWR VGND _340_/CLK _312_/D _346_/SET_B _312_/Q sky130_fd_sc_hd__dfrtp_1
X_174_ VPWR VGND VPWR VGND _161_/Y _344_/Q _172_/A _344_/D _147_/A sky130_fd_sc_hd__a22o_1
XFILLER_22_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_226_ VGND VPWR VPWR VGND _150_/C _225_/X _147_/A _226_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_157_ VGND VPWR VPWR VGND _157_/A _172_/A sky130_fd_sc_hd__clkbuf_2
X_209_ VPWR VGND VPWR VGND _153_/A _333_/Q _332_/Q _209_/X _153_/B sky130_fd_sc_hd__a22o_1
XFILLER_14_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_190_ VGND VPWR VPWR VGND _190_/A _306_/S sky130_fd_sc_hd__clkbuf_2
X_242_ VGND VPWR VPWR VGND _242_/A _242_/B _318_/D sky130_fd_sc_hd__nor2_1
XFILLER_14_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_173_ VGND VPWR VPWR VGND _345_/Q _147_/Y _172_/Y _147_/Y _345_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_311_ VGND VPWR VPWR VGND _340_/CLK _311_/D _346_/SET_B _311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_156_ VPWR VGND VPWR VGND _157_/A _196_/A _225_/B sky130_fd_sc_hd__or2_2
X_225_ VPWR VGND VPWR VGND _225_/X _336_/Q _225_/B sky130_fd_sc_hd__and2_1
X_208_ VGND VPWR VPWR VGND _207_/X _204_/Y _206_/A _334_/Q _334_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_310_ VGND VPWR VPWR VGND _340_/CLK _310_/D _346_/SET_B _310_/Q sky130_fd_sc_hd__dfrtp_1
X_241_ VPWR VGND VPWR VGND _232_/X _327_/Q _318_/Q _242_/B sky130_fd_sc_hd__a21oi_1
X_172_ VGND VPWR VPWR VGND _172_/A _172_/B _172_/Y sky130_fd_sc_hd__nor2_1
X_224_ VGND VPWR VPWR VGND _324_/D _216_/A _325_/Q _304_/X _217_/A _324_/Q sky130_fd_sc_hd__a32o_1
XFILLER_6_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_155_ VPWR VGND VPWR VGND _225_/B _254_/B sky130_fd_sc_hd__inv_2
XFILLER_17_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_207_ VGND VPWR VPWR VGND _207_/X _207_/C _332_/Q _333_/Q sky130_fd_sc_hd__and3_1
XFILLER_0_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_26 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_240_ VGND VPWR VPWR VGND _242_/A _240_/B _319_/D sky130_fd_sc_hd__nor2_1
X_171_ VGND VPWR VPWR VGND _164_/A _164_/Y _161_/Y _344_/Q _172_/B sky130_fd_sc_hd__o22a_1
XFILLER_9_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_223_ VGND VPWR VPWR VGND _325_/D _216_/A _326_/Q _304_/X _217_/A _325_/Q sky130_fd_sc_hd__a32o_1
XFILLER_8_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_154_ VGND VPWR VPWR VGND _254_/B _154_/A sky130_fd_sc_hd__buf_1
X_206_ VPWR VGND VPWR VGND _207_/C _206_/A sky130_fd_sc_hd__inv_2
XFILLER_5_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_11_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_170_ VGND VPWR VPWR VGND _346_/Q _147_/Y _169_/Y _147_/Y _346_/D sky130_fd_sc_hd__a2bb2o_1
X_299_ VGND VPWR VPWR VGND _167_/X _160_/X _166_/Y _165_/X _299_/X sky130_fd_sc_hd__o22a_1
XFILLER_3_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_222_ VGND VPWR VPWR VGND _326_/D _216_/A _327_/Q _212_/X _217_/X _326_/Q sky130_fd_sc_hd__a32o_1
X_153_ VGND VPWR VPWR VGND _154_/A _334_/Q _335_/Q _153_/B _153_/A sky130_fd_sc_hd__or4b_4
XFILLER_10_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_205_ VGND VPWR VPWR VGND _206_/A _204_/Y _335_/Q _335_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_84 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_298_ VGND VPWR VPWR VGND _298_/X _298_/C _298_/B _298_/A sky130_fd_sc_hd__and3_1
XFILLER_9_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_221_ VGND VPWR VPWR VGND _327_/D _216_/X _328_/Q _212_/X _217_/X _327_/Q sky130_fd_sc_hd__a32o_1
X_152_ VPWR VGND VPWR VGND _153_/B _332_/Q sky130_fd_sc_hd__inv_2
X_204_ VPWR VGND VPWR VGND _190_/A _204_/Y _333_/Q _332_/Q _334_/Q sky130_fd_sc_hd__a31oi_2
XFILLER_3_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_297_ VGND VPWR VPWR VGND _297_/B _297_/Y _297_/A sky130_fd_sc_hd__nor2_2
X_220_ VGND VPWR VPWR VGND _328_/D _216_/X _329_/Q _212_/X _217_/X _328_/Q sky130_fd_sc_hd__a32o_1
X_151_ VPWR VGND VPWR VGND _153_/A _333_/Q sky130_fd_sc_hd__inv_2
XFILLER_6_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_203_ VGND VPWR VPWR VGND _206_/A _298_/C _225_/B _336_/Q _147_/Y sky130_fd_sc_hd__a31o_1
XFILLER_9_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_296_ VGND VPWR VPWR VGND _342_/Q _255_/B _296_/Y _306_/S _286_/B _284_/A sky130_fd_sc_hd__o221ai_1
XFILLER_3_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_150_ VPWR VGND VPWR VGND _298_/B _150_/C _342_/Q _196_/A sky130_fd_sc_hd__or3_4
X_279_ VPWR VGND VPWR VGND _279_/Y _279_/A sky130_fd_sc_hd__inv_2
XFILLER_17_7 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_202_ VGND VPWR VPWR VGND _336_/D _193_/Y _197_/X _337_/Q _284_/A _194_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_9_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xoutput40 VGND VPWR VPWR VGND _294_/Y trimb[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_15_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput5 VGND VPWR VPWR VGND clkc _297_/Y sky130_fd_sc_hd__buf_1
XFILLER_3_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_295_ VPWR VGND VPWR VGND _308_/S _181_/X _190_/A _286_/B _255_/B _342_/Q sky130_fd_sc_hd__o2111a_1
XFILLER_10_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_278_ VGND VPWR VPWR VGND _279_/A _329_/Q _320_/Q sky130_fd_sc_hd__or2_1
X_347_ VGND VPWR VPWR VGND _297_/B _347_/D _346_/SET_B _347_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_201_ VGND VPWR VPWR VGND _336_/Q _284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput6 VGND VPWR VPWR VGND _269_/Y ctln[0] sky130_fd_sc_hd__clkbuf_2
Xoutput41 VGND VPWR VPWR VGND _298_/X valid sky130_fd_sc_hd__clkbuf_2
Xoutput30 VGND VPWR VPWR VGND _286_/Y sample sky130_fd_sc_hd__clkbuf_2
.ends

.subckt SAR comp ctln1 ctln0 ctlp1 ctlp0 ctln7 ctln6 ctln5 ctln4 ctln3 ctln2 trim4
+ trim1 trim0 trim2 trim3 trimb3 trimb2 trimb0 trimb1 trimb4 ctlp2 ctlp3 ctlp4 ctlp5
+ ctlp6 ctlp7 clkc result7 result6 result5 result4 rstn result3 result2 result1 result0
+ valid cal en clk dvdd vinp vinn avdd dvss
Xlatch_0 latch_0/Qn latch_0/S latch_0/R comp avdd dvss latch
XDAC_0 DAC_0/enb DAC_0/en_buf ctlp1 ctlp0 avdd ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp2
+ sample DAC_0/out vinp avdd DAC_0/en_buf_uq0 DAC_0/enb_uq0 dvss avdd DAC
XDAC_1 DAC_1/enb DAC_1/en_buf ctln1 ctln0 dvss ctln3 ctln4 ctln5 ctln6 ctln7 ctln2
+ sample DAC_1/out vinn avdd DAC_1/en_buf_uq0 DAC_1/enb_uq0 dvss avdd DAC
Xdecap_3$1_0 dvss avdd avdd dvss decap_3$1
Xcomparator_0 trim3 trim2 trim0 trim1 trim4 trimb4 trimb1 trimb0 trimb2 trimb3 latch_0/R
+ latch_0/S clkc avdd DAC_0/out DAC_1/out dvss comparator
Xsarlogic_0 ctln0 ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctlp0 ctlp1 ctlp2 ctlp3
+ ctlp4 ctlp5 ctlp6 ctlp7 cal clk clkc comp en result0 result1 result2 result3 result4
+ result5 result6 result7 rstn sample trim0 trim1 trim2 trim3 trim4 trimb0 trimb1
+ trimb2 trimb3 trimb4 valid dvdd dvss sarlogic
.ends

.subckt user_analog_project_wrapper wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[1] wbs_adr_i[2] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[1]
+ wbs_dat_i[2] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[1] wbs_dat_o[2] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i wbs_dat_i[17] wbs_dat_i[18]
+ wbs_dat_i[19] wbs_adr_i[18] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23]
+ wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29]
+ wbs_adr_i[19] wbs_dat_i[30] wbs_dat_i[31] la_oenb[0] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] la_oenb[1] wbs_adr_i[30] wbs_adr_i[31] la_oenb[2] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] la_oenb[3] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] la_oenb[4] wbs_dat_o[30] wbs_dat_o[31] la_oenb[5] la_data_in[0] la_data_in[1]
+ la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5] la_data_out[0] la_data_out[1]
+ la_data_out[2] la_data_out[3] la_data_out[4] la_data_out[5] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] la_data_in[26] la_data_in[11]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[6] la_data_in[7] la_data_in[8]
+ la_data_in[9] la_data_in[15] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_in[16] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[10]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_data_in[20] la_oenb[10]
+ la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_data_in[21] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_data_in[22] la_data_in[39] la_oenb[45] la_data_in[40]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_in[41] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_in[42] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_oenb[46]
+ la_oenb[38] la_oenb[39] la_oenb[37] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_oenb[44] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_data_in[38] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[47] la_oenb[48]
+ la_oenb[49] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_out[47] la_data_out[48] la_data_out[49] la_data_in[64]
+ la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_in[65] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_in[66] la_data_in[67] la_data_in[72]
+ la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78]
+ la_data_in[79] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[69] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_data_out[68] la_data_out[69]
+ la_data_in[70] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_in[71] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_in[68] la_oenb[88] la_oenb[89]
+ la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96]
+ la_oenb[97] la_oenb[98] la_oenb[99] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[100] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94]
+ la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[93] la_data_out[106] la_data_out[94] la_data_out[107] la_data_out[95]
+ la_data_out[96] la_data_out[108] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[92] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_data_in[88] la_data_in[89] la_data_out[88]
+ la_data_out[89] la_data_out[90] la_data_out[91] la_data_in[119] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_in[116] la_data_in[117] la_data_out[123]
+ la_data_in[112] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_in[118] la_oenb[109] la_data_in[120] la_oenb[110] la_data_in[121] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_data_in[122] la_data_in[123] la_oenb[120] la_oenb[121] la_oenb[122]
+ la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_out[110] user_clock2 user_irq[0]
+ la_data_in[113] user_irq[1] la_data_in[114] user_irq[2] la_data_out[111] la_data_out[112]
+ la_data_out[109] la_data_in[109] la_data_out[113] la_data_in[110] la_data_out[114]
+ la_oenb[108] la_data_out[115] la_data_out[116] la_data_in[111] la_data_out[117]
+ la_data_in[115] la_data_out[118] la_data_out[119] gpio_analog[2] gpio_analog[3]
+ gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4]
+ gpio_noesd[5] gpio_noesd[6] io_analog[0] io_analog[1] io_analog[2] io_analog[3]
+ io_analog[4] io_clamp_high[0] io_clamp_low[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[9] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[9] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[9] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[9] vccd1 vdda1 io_in[16] io_in[17] gpio_analog[9] gpio_noesd[10] io_analog[5]
+ io_analog[6] io_analog[7] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17]
+ io_analog[8] io_analog[9] gpio_noesd[7] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ gpio_noesd[8] io_clamp_high[1] io_clamp_high[2] gpio_noesd[9] io_clamp_low[1] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_clamp_low[2] gpio_analog[10] io_analog[10] vccd2
+ gpio_analog[7] gpio_analog[8] io_in[14] io_in[15] vssa2 io_in_3v3[24] io_in_3v3[25]
+ io_in_3v3[26] gpio_analog[16] gpio_analog[17] gpio_analog[11] gpio_analog[12] gpio_noesd[11]
+ io_in[18] io_in[19] io_in[20] io_in[21] io_oeb[18] io_oeb[19] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15]
+ io_out[18] io_out[19] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] gpio_noesd[16] gpio_noesd[17] gpio_analog[13] gpio_analog[14] gpio_analog[15]
+ io_in_3v3[18] io_in_3v3[19] vdda2 io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ vssa1 io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in[1] io_oeb[0] gpio_noesd[0] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_out[1] io_in[6] io_in_3v3[1] io_in[7] io_in[8] gpio_analog[0]
+ io_oeb[1] io_in_3v3[0] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] gpio_analog[1] gpio_noesd[1] io_in[0] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] vssd1 io_in_3v3[5]
+ io_out[0] io_analog[6]_uq0 io_analog[6]_uq1 io_analog[6]_uq2 io_analog[6]_uq3 io_analog[6]_uq4
+ io_analog[4]_uq0 io_analog[4]_uq1 io_analog[4]_uq2 io_analog[4]_uq3 io_analog[4]_uq4
+ io_analog[5]_uq0 io_analog[5]_uq1 io_analog[5]_uq2 io_analog[5]_uq3 io_analog[5]_uq4
+ vssa1_uq0 vssa1_uq1 vssa1_uq2 vssd1_uq0 vdda1_uq0 vdda1_uq1 vdda1_uq2 vssd2_uq0
+ vdda2_uq0 vssa2_uq0 vccd1_uq0 vccd2_uq0
XSAR_0 SAR_0/comp SAR_0/ctln1 SAR_0/ctln0 SAR_0/ctlp1 SAR_0/ctlp0 SAR_0/ctln7 SAR_0/ctln6
+ SAR_0/ctln5 SAR_0/ctln4 SAR_0/ctln3 SAR_0/ctln2 SAR_0/trim4 SAR_0/trim1 SAR_0/trim0
+ SAR_0/trim2 SAR_0/trim3 SAR_0/trimb3 SAR_0/trimb2 SAR_0/trimb0 SAR_0/trimb1 SAR_0/trimb4
+ SAR_0/ctlp2 SAR_0/ctlp3 SAR_0/ctlp4 SAR_0/ctlp5 SAR_0/ctlp6 SAR_0/ctlp7 SAR_0/clkc
+ la_data_out[29] la_data_out[30] la_data_out[31] la_data_out[32] io_in[23] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] io_out[17] io_in[18] io_in[19] io_in[20]
+ vccd2 io_analog[5] io_analog[4] vdda1 vssa1 SAR
.ends

